module booth_multiplier (clk,
    done,
    rst,
    start,
    multiplicand,
    multiplier,
    product);
 input clk;
 output done;
 input rst;
 input start;
 input [7:0] multiplicand;
 input [7:0] multiplier;
 output [15:0] product;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire start_r;
 wire state;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _375_ (.I(state),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _376_ (.A1(_018_),
    .A2(_281_),
    .Z(_019_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _377_ (.I(_019_),
    .Z(_020_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _378_ (.I(_020_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _379_ (.A1(_018_),
    .A2(net19),
    .B(_021_),
    .ZN(_374_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _380_ (.A1(net9),
    .A2(net2),
    .Z(_284_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _381_ (.A1(net1),
    .A2(net10),
    .Z(_283_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _382_ (.A1(net1),
    .A2(net11),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _383_ (.A1(net9),
    .A2(net4),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _384_ (.A1(net10),
    .A2(net3),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _385_ (.A1(net2),
    .A2(net11),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _386_ (.A1(net1),
    .A2(net12),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _387_ (.A1(net9),
    .A2(net5),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _388_ (.A1(net10),
    .A2(net4),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _389_ (.A1(net3),
    .A2(net11),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _390_ (.A1(net2),
    .A2(net12),
    .Z(_294_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _391_ (.A1(net1),
    .A2(net13),
    .Z(_293_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _392_ (.A1(net9),
    .A2(net7),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _393_ (.A1(net10),
    .A2(net6),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _394_ (.A1(net11),
    .A2(net5),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _395_ (.A1(net10),
    .A2(net5),
    .Z(_116_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _396_ (.A1(net11),
    .A2(net4),
    .Z(_115_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _397_ (.A1(net4),
    .A2(net12),
    .Z(_109_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _398_ (.A1(net3),
    .A2(net13),
    .Z(_108_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _399_ (.A1(net2),
    .A2(net14),
    .Z(_107_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _400_ (.A1(net1),
    .A2(net15),
    .Z(_303_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _401_ (.A1(net10),
    .A2(net7),
    .ZN(_142_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _402_ (.A1(net11),
    .A2(net6),
    .ZN(_148_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _403_ (.A1(net12),
    .A2(net5),
    .ZN(_146_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _404_ (.A1(net4),
    .A2(net13),
    .ZN(_147_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _405_ (.A1(net3),
    .A2(net14),
    .Z(_153_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _406_ (.A1(net2),
    .A2(net15),
    .Z(_155_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _407_ (.I(net16),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _408_ (.A1(net1),
    .A2(_141_),
    .ZN(_154_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _409_ (.I(_165_),
    .ZN(_162_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _410_ (.A1(net11),
    .A2(net7),
    .Z(_319_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _411_ (.A1(net12),
    .A2(net6),
    .ZN(_168_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _412_ (.A1(net5),
    .A2(net13),
    .ZN(_167_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _413_ (.A1(net4),
    .A2(net14),
    .ZN(_166_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _414_ (.A1(net3),
    .A2(net15),
    .Z(_323_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _415_ (.A1(net2),
    .A2(_141_),
    .ZN(_324_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _416_ (.A1(net11),
    .A2(net8),
    .Z(_329_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _417_ (.A1(net9),
    .A2(net10),
    .A3(net8),
    .Z(_022_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _418_ (.A1(_321_),
    .A2(_022_),
    .ZN(_191_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _419_ (.A1(net12),
    .A2(net7),
    .ZN(_186_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _420_ (.A1(net13),
    .A2(net6),
    .ZN(_187_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _421_ (.A1(net5),
    .A2(net14),
    .ZN(_185_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _422_ (.A1(net4),
    .A2(net15),
    .Z(_333_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _423_ (.A1(net3),
    .A2(_141_),
    .ZN(_332_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _424_ (.A1(_330_),
    .A2(_022_),
    .ZN(_209_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _425_ (.A1(net12),
    .A2(net8),
    .Z(_204_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _426_ (.A1(net13),
    .A2(net7),
    .Z(_205_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _427_ (.A1(net6),
    .A2(net14),
    .Z(_206_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _428_ (.A1(net5),
    .A2(net15),
    .Z(_337_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _429_ (.A1(net4),
    .A2(_141_),
    .ZN(_338_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _430_ (.I(_314_),
    .ZN(_138_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _431_ (.A1(net13),
    .A2(net8),
    .Z(_225_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _432_ (.A1(net7),
    .A2(net14),
    .Z(_224_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _433_ (.A1(net6),
    .A2(net15),
    .Z(_344_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _434_ (.A1(net5),
    .A2(_141_),
    .ZN(_343_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _435_ (.A1(net14),
    .A2(net8),
    .Z(_241_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _436_ (.A1(net7),
    .A2(net15),
    .Z(_350_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _437_ (.A1(net6),
    .A2(_141_),
    .ZN(_351_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _438_ (.A1(net15),
    .A2(net8),
    .Z(_359_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _439_ (.A1(net7),
    .A2(_141_),
    .ZN(_360_));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 _440_ (.I(net17),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _441_ (.A1(net1),
    .A2(net14),
    .ZN(_120_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _442_ (.I(_295_),
    .ZN(_133_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _443_ (.A1(net2),
    .A2(net10),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _444_ (.A1(net2),
    .A2(net13),
    .ZN(_121_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _445_ (.A1(net9),
    .A2(net3),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _446_ (.A1(net3),
    .A2(net12),
    .ZN(_122_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _447_ (.A1(net9),
    .A2(net8),
    .ZN(_143_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _448_ (.I(_119_),
    .ZN(_131_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _449_ (.I(_129_),
    .ZN(_306_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _450_ (.I(_198_),
    .ZN(_199_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _451_ (.I(_208_),
    .ZN(_210_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _452_ (.I(_217_),
    .ZN(_218_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _453_ (.I(_227_),
    .ZN(_228_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _454_ (.I(_234_),
    .ZN(_235_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _455_ (.I(_243_),
    .ZN(_244_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _456_ (.I(_250_),
    .ZN(_251_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _457_ (.I(_260_),
    .ZN(_261_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _458_ (.I(_270_),
    .ZN(_271_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _459_ (.I(_118_),
    .ZN(_112_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _460_ (.I(_128_),
    .ZN(_161_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _461_ (.I(_156_),
    .ZN(_174_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _462_ (.I(_197_),
    .ZN(_221_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _463_ (.I(_216_),
    .ZN(_238_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _464_ (.I(_233_),
    .ZN(_254_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _465_ (.I(_249_),
    .ZN(_264_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _466_ (.I(_259_),
    .ZN(_274_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _467_ (.I(net18),
    .ZN(_277_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _468_ (.I(_092_),
    .ZN(_297_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _469_ (.I(_097_),
    .ZN(_130_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _470_ (.I(_134_),
    .ZN(_305_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _471_ (.I(_164_),
    .ZN(_316_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _472_ (.I(_179_),
    .ZN(_180_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _473_ (.I(_163_),
    .ZN(_326_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _474_ (.I(_169_),
    .ZN(_194_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _475_ (.I(_223_),
    .ZN(_339_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _476_ (.I(_240_),
    .ZN(_345_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _477_ (.I(_246_),
    .ZN(_349_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _478_ (.I(_256_),
    .ZN(_352_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _479_ (.I(_255_),
    .ZN(_361_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _480_ (.I(_276_),
    .ZN(_369_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _481_ (.I(start_r),
    .ZN(_280_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _482_ (.I(_085_),
    .ZN(_287_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _483_ (.I(_093_),
    .ZN(_290_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _484_ (.I(_101_),
    .ZN(_298_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _485_ (.A1(net9),
    .A2(net6),
    .Z(_117_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _486_ (.I(_114_),
    .ZN(_127_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _487_ (.I(_123_),
    .ZN(_304_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _488_ (.I(_135_),
    .ZN(_312_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _489_ (.I(_159_),
    .ZN(_181_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _490_ (.A1(net9),
    .A2(net10),
    .Z(_023_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _491_ (.A1(net8),
    .A2(_023_),
    .Z(_320_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _492_ (.I(_203_),
    .ZN(_334_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _493_ (.I(_188_),
    .ZN(_215_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _494_ (.I(_202_),
    .ZN(_340_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _495_ (.I(_222_),
    .ZN(_346_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _496_ (.I(_239_),
    .ZN(_353_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _497_ (.I(_245_),
    .ZN(_356_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _498_ (.I(_266_),
    .ZN(_362_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _499_ (.A1(net8),
    .A2(_141_),
    .ZN(_365_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _500_ (.I(_265_),
    .ZN(_370_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _501_ (.I(_308_),
    .ZN(_137_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _502_ (.I(_315_),
    .ZN(_158_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _503_ (.I(_322_),
    .ZN(_171_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _504_ (.I(_331_),
    .ZN(_190_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _505_ (.I(_296_),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _506_ (.I(_325_),
    .ZN(_175_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _507_ (.I(_309_),
    .ZN(_136_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _508_ (.A1(_018_),
    .A2(net19),
    .A3(_279_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _509_ (.A1(_018_),
    .A2(_278_),
    .B(_024_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _510_ (.A1(net9),
    .A2(net1),
    .Z(_025_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _511_ (.I(_020_),
    .Z(_026_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _512_ (.I0(net20),
    .I1(_025_),
    .S(_026_),
    .Z(_002_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _513_ (.A1(_311_),
    .A2(_314_),
    .B(_310_),
    .C(_317_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _514_ (.A1(_318_),
    .A2(_317_),
    .B(_328_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _515_ (.I(_327_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _516_ (.A1(_027_),
    .A2(_028_),
    .B(_029_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _517_ (.A1(_336_),
    .A2(_030_),
    .B(_335_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _518_ (.A1(_342_),
    .A2(_031_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _519_ (.I0(net21),
    .I1(_032_),
    .S(_026_),
    .Z(_003_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _520_ (.I(_139_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _521_ (.A1(_318_),
    .A2(_033_),
    .B(_317_),
    .C(_327_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _522_ (.A1(_328_),
    .A2(_327_),
    .B(_336_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _523_ (.I(_335_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _524_ (.A1(_034_),
    .A2(_035_),
    .B(_036_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _525_ (.A1(_342_),
    .A2(_037_),
    .B(_341_),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _526_ (.A1(_348_),
    .A2(_038_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _527_ (.I0(net22),
    .I1(_039_),
    .S(_026_),
    .Z(_004_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _528_ (.A1(_342_),
    .A2(_348_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _529_ (.A1(_348_),
    .A2(_341_),
    .B(_347_),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _530_ (.A1(_031_),
    .A2(_040_),
    .B(_041_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _531_ (.A1(_355_),
    .A2(_042_),
    .Z(_043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _532_ (.I0(net23),
    .I1(_043_),
    .S(_026_),
    .Z(_005_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _533_ (.I(_041_),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _534_ (.A1(_342_),
    .A2(_348_),
    .A3(_355_),
    .Z(_045_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _535_ (.A1(_355_),
    .A2(_044_),
    .B1(_045_),
    .B2(_037_),
    .C(_354_),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _536_ (.A1(_364_),
    .A2(_046_),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _537_ (.I0(net24),
    .I1(_047_),
    .S(_026_),
    .Z(_006_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _538_ (.I(_372_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _539_ (.A1(_348_),
    .A2(_355_),
    .A3(_364_),
    .Z(_049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _540_ (.A1(_342_),
    .A2(_049_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _541_ (.A1(_372_),
    .A2(_050_),
    .Z(_051_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _542_ (.A1(_355_),
    .A2(_364_),
    .Z(_052_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _543_ (.A1(_364_),
    .A2(_354_),
    .B1(_044_),
    .B2(_052_),
    .C(_363_),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _544_ (.I0(_048_),
    .I1(_051_),
    .S(_053_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _545_ (.I0(net25),
    .I1(_054_),
    .S(_020_),
    .Z(_055_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _546_ (.A1(_372_),
    .A2(_020_),
    .A3(_031_),
    .A4(_053_),
    .Z(_056_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _547_ (.A1(_372_),
    .A2(_021_),
    .A3(_031_),
    .A4(_050_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _548_ (.A1(_055_),
    .A2(_056_),
    .A3(_057_),
    .Z(_007_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _549_ (.A1(_272_),
    .A2(_275_),
    .Z(_058_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _550_ (.A1(_269_),
    .A2(_368_),
    .A3(_058_),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _551_ (.A1(_366_),
    .A2(_358_),
    .A3(_059_),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _552_ (.I(_341_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _553_ (.A1(_034_),
    .A2(_035_),
    .B(_036_),
    .C(_061_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _554_ (.A1(_342_),
    .A2(_341_),
    .Z(_063_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _555_ (.A1(_372_),
    .A2(_049_),
    .A3(_063_),
    .Z(_064_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _556_ (.A1(_355_),
    .A2(_347_),
    .Z(_065_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _557_ (.A1(_354_),
    .A2(_065_),
    .B(_364_),
    .C(_372_),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _558_ (.A1(_372_),
    .A2(_363_),
    .B(_371_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _559_ (.A1(_066_),
    .A2(_067_),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _560_ (.A1(_062_),
    .A2(_064_),
    .B(_068_),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _561_ (.A1(_060_),
    .A2(_069_),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _562_ (.I0(net26),
    .I1(_070_),
    .S(_026_),
    .Z(_008_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _563_ (.I0(net27),
    .I1(_286_),
    .S(_026_),
    .Z(_009_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _564_ (.I0(net28),
    .I1(_289_),
    .S(_026_),
    .Z(_010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _565_ (.I0(net29),
    .I1(_292_),
    .S(_026_),
    .Z(_011_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _566_ (.I0(net30),
    .I1(_302_),
    .S(_026_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _567_ (.I0(net31),
    .I1(_373_),
    .S(_020_),
    .Z(_013_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _568_ (.I(_140_),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _569_ (.I0(net32),
    .I1(_071_),
    .S(_020_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _570_ (.A1(_318_),
    .A2(_139_),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _571_ (.I0(net33),
    .I1(_072_),
    .S(_020_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _572_ (.A1(_311_),
    .A2(_314_),
    .Z(_073_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _573_ (.A1(_310_),
    .A2(_073_),
    .Z(_074_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _574_ (.A1(_318_),
    .A2(_074_),
    .B(_317_),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _575_ (.A1(_328_),
    .A2(_075_),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _576_ (.I0(net34),
    .I1(_076_),
    .S(_020_),
    .Z(_016_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _577_ (.A1(_318_),
    .A2(_033_),
    .Z(_077_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _578_ (.A1(_317_),
    .A2(_077_),
    .B(_328_),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _579_ (.A1(_029_),
    .A2(_078_),
    .Z(_079_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _580_ (.A1(_336_),
    .A2(_079_),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _581_ (.I0(net35),
    .I1(_080_),
    .S(_020_),
    .Z(_017_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _582_ (.A(_081_),
    .B(_082_),
    .CI(_083_),
    .CO(_084_),
    .S(_085_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _583_ (.A(_086_),
    .B(_087_),
    .CI(_088_),
    .CO(_089_),
    .S(_090_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _584_ (.A(_091_),
    .B(_084_),
    .CI(_090_),
    .CO(_092_),
    .S(_093_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _585_ (.A(_094_),
    .B(_095_),
    .CI(_096_),
    .CO(_097_),
    .S(_098_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _586_ (.A(_099_),
    .B(_089_),
    .CI(_098_),
    .CO(_100_),
    .S(_101_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _587_ (.A(_102_),
    .B(_103_),
    .CI(_104_),
    .CO(_105_),
    .S(_106_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _588_ (.A(_107_),
    .B(_108_),
    .CI(_109_),
    .CO(_110_),
    .S(_111_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _589_ (.A(_111_),
    .B(_112_),
    .CI(_106_),
    .CO(_113_),
    .S(_114_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _590_ (.A(_115_),
    .B(_116_),
    .CI(_117_),
    .CO(_118_),
    .S(_119_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _591_ (.A(_120_),
    .B(_121_),
    .CI(_122_),
    .CO(_123_),
    .S(_124_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _592_ (.A(_125_),
    .B(_126_),
    .CI(_127_),
    .CO(_128_),
    .S(_129_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _593_ (.A(_124_),
    .B(_130_),
    .CI(_131_),
    .CO(_125_),
    .S(_132_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _594_ (.A(_133_),
    .B(_100_),
    .CI(_132_),
    .CO(_134_),
    .S(_135_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _595_ (.A(_136_),
    .B(_137_),
    .CI(_138_),
    .CO(_139_),
    .S(_140_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _596_ (.A(_141_),
    .B(_142_),
    .CI(_143_),
    .CO(_144_),
    .S(_145_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _597_ (.A(_146_),
    .B(_147_),
    .CI(_148_),
    .CO(_149_),
    .S(_150_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _598_ (.A(_145_),
    .B(_105_),
    .CI(_150_),
    .CO(_151_),
    .S(_152_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _599_ (.A(_153_),
    .B(_154_),
    .CI(_155_),
    .CO(_156_),
    .S(_157_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _600_ (.A(_113_),
    .B(_152_),
    .CI(_158_),
    .CO(_159_),
    .S(_160_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _601_ (.A(_161_),
    .B(_162_),
    .CI(_160_),
    .CO(_163_),
    .S(_164_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _602_ (.A(_166_),
    .B(_167_),
    .CI(_168_),
    .CO(_169_),
    .S(_170_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _603_ (.A(_170_),
    .B(_171_),
    .CI(_144_),
    .CO(_172_),
    .S(_173_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _604_ (.A(_174_),
    .B(_149_),
    .CI(_175_),
    .CO(_176_),
    .S(_177_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _605_ (.A(_177_),
    .B(_151_),
    .CI(_173_),
    .CO(_178_),
    .S(_179_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _606_ (.A(_180_),
    .B(_181_),
    .CI(_182_),
    .CO(_183_),
    .S(_184_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _607_ (.A(_185_),
    .B(_186_),
    .CI(_187_),
    .CO(_188_),
    .S(_189_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _608_ (.A(_189_),
    .B(_190_),
    .CI(_191_),
    .CO(_192_),
    .S(_193_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _609_ (.A(_194_),
    .B(_195_),
    .CI(_196_),
    .CO(_197_),
    .S(_198_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _610_ (.A(_193_),
    .B(_172_),
    .CI(_199_),
    .CO(_200_),
    .S(_201_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _611_ (.A(_176_),
    .B(_178_),
    .CI(_201_),
    .CO(_202_),
    .S(_203_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _612_ (.A(_204_),
    .B(_205_),
    .CI(_206_),
    .CO(_207_),
    .S(_208_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _613_ (.A(_209_),
    .B(_210_),
    .CI(_190_),
    .CO(_211_),
    .S(_212_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _614_ (.A(_213_),
    .B(_214_),
    .CI(_215_),
    .CO(_216_),
    .S(_217_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _615_ (.A(_212_),
    .B(_192_),
    .CI(_218_),
    .CO(_219_),
    .S(_220_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _616_ (.A(_200_),
    .B(_221_),
    .CI(_220_),
    .CO(_222_),
    .S(_223_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _617_ (.A(_204_),
    .B(_224_),
    .CI(_225_),
    .CO(_226_),
    .S(_227_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _618_ (.A(_209_),
    .B(_190_),
    .CI(_228_),
    .CO(_229_),
    .S(_230_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _619_ (.A(_231_),
    .B(_207_),
    .CI(_232_),
    .CO(_233_),
    .S(_234_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _620_ (.A(_235_),
    .B(_211_),
    .CI(_230_),
    .CO(_236_),
    .S(_237_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _621_ (.A(_237_),
    .B(_219_),
    .CI(_238_),
    .CO(_239_),
    .S(_240_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _622_ (.A(_204_),
    .B(_241_),
    .CI(_225_),
    .CO(_242_),
    .S(_243_));
 gf180mcu_fd_sc_mcu9t5v0__addf_4 _623_ (.A(_209_),
    .B(_190_),
    .CI(_244_),
    .CO(_245_),
    .S(_246_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _624_ (.A(_226_),
    .B(_247_),
    .CI(_248_),
    .CO(_249_),
    .S(_250_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _625_ (.A(_246_),
    .B(_229_),
    .CI(_251_),
    .CO(_252_),
    .S(_253_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _626_ (.A(_253_),
    .B(_236_),
    .CI(_254_),
    .CO(_255_),
    .S(_256_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _627_ (.A(_242_),
    .B(_257_),
    .CI(_258_),
    .CO(_259_),
    .S(_260_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _628_ (.A(_246_),
    .B(_245_),
    .CI(_261_),
    .CO(_262_),
    .S(_263_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _629_ (.A(_263_),
    .B(_252_),
    .CI(_264_),
    .CO(_265_),
    .S(_266_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _630_ (.A(_242_),
    .B(_267_),
    .CI(_268_),
    .CO(_269_),
    .S(_270_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _631_ (.A(_246_),
    .B(_245_),
    .CI(_271_),
    .CO(_272_),
    .S(_273_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _632_ (.A(_262_),
    .B(_274_),
    .CI(_273_),
    .CO(_275_),
    .S(_276_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _633_ (.A(_277_),
    .B(start_r),
    .CO(_278_),
    .S(_279_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _634_ (.A(net18),
    .B(_280_),
    .CO(_281_),
    .S(_282_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _635_ (.A(_283_),
    .B(_284_),
    .CO(_285_),
    .S(_286_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _636_ (.A(_285_),
    .B(_287_),
    .CO(_288_),
    .S(_289_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _637_ (.A(_288_),
    .B(_290_),
    .CO(_291_),
    .S(_292_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _638_ (.A(_293_),
    .B(_294_),
    .CO(_295_),
    .S(_296_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _639_ (.A(_297_),
    .B(_298_),
    .CO(_299_),
    .S(_300_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _640_ (.A(_291_),
    .B(_300_),
    .CO(_301_),
    .S(_302_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _641_ (.A(_303_),
    .B(_304_),
    .CO(_165_),
    .S(_126_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _642_ (.A(_305_),
    .B(_306_),
    .CO(_307_),
    .S(_308_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _643_ (.A(_309_),
    .B(_308_),
    .CO(_310_),
    .S(_311_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _644_ (.A(_299_),
    .B(_312_),
    .CO(_309_),
    .S(_313_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _645_ (.A(_110_),
    .B(_157_),
    .CO(_182_),
    .S(_315_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _646_ (.A(_316_),
    .B(_307_),
    .CO(_317_),
    .S(_318_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _647_ (.A(_319_),
    .B(_320_),
    .CO(_321_),
    .S(_322_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _648_ (.A(_323_),
    .B(_324_),
    .CO(_195_),
    .S(_325_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _649_ (.A(_326_),
    .B(_184_),
    .CO(_327_),
    .S(_328_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _650_ (.A(_329_),
    .B(_320_),
    .CO(_330_),
    .S(_331_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _651_ (.A(_332_),
    .B(_333_),
    .CO(_214_),
    .S(_196_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _652_ (.A(_183_),
    .B(_334_),
    .CO(_335_),
    .S(_336_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _653_ (.A(_337_),
    .B(_338_),
    .CO(_231_),
    .S(_213_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _654_ (.A(_339_),
    .B(_340_),
    .CO(_341_),
    .S(_342_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _655_ (.A(_343_),
    .B(_344_),
    .CO(_248_),
    .S(_232_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _656_ (.A(_345_),
    .B(_346_),
    .CO(_347_),
    .S(_348_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _657_ (.A(_350_),
    .B(_351_),
    .CO(_257_),
    .S(_247_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _658_ (.A(_352_),
    .B(_353_),
    .CO(_354_),
    .S(_355_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _659_ (.A(_349_),
    .B(_356_),
    .CO(_357_),
    .S(_358_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _660_ (.A(_359_),
    .B(_360_),
    .CO(_268_),
    .S(_258_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _661_ (.A(_361_),
    .B(_362_),
    .CO(_363_),
    .S(_364_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _662_ (.A(_359_),
    .B(_365_),
    .CO(_366_),
    .S(_267_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _663_ (.A(_242_),
    .B(_267_),
    .CO(_367_),
    .S(_368_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _664_ (.A(_369_),
    .B(_370_),
    .CO(_371_),
    .S(_372_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _665_ (.A(_301_),
    .B(_313_),
    .CO(_314_),
    .S(_373_));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \done$_DFFE_PP0P_  (.D(_001_),
    .RN(_000_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \product[0]$_DFFE_PP0P_  (.D(_002_),
    .RN(_000_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \product[10]$_DFFE_PP0P_  (.D(_003_),
    .RN(_000_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \product[11]$_DFFE_PP0P_  (.D(_004_),
    .RN(_000_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \product[12]$_DFFE_PP0P_  (.D(_005_),
    .RN(_000_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \product[13]$_DFFE_PP0P_  (.D(_006_),
    .RN(_000_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \product[14]$_DFFE_PP0P_  (.D(_007_),
    .RN(_000_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \product[15]$_DFFE_PP0P_  (.D(_008_),
    .RN(_000_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \product[1]$_DFFE_PP0P_  (.D(_009_),
    .RN(_000_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \product[2]$_DFFE_PP0P_  (.D(_010_),
    .RN(_000_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \product[3]$_DFFE_PP0P_  (.D(_011_),
    .RN(_000_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \product[4]$_DFFE_PP0P_  (.D(_012_),
    .RN(_000_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \product[5]$_DFFE_PP0P_  (.D(_013_),
    .RN(_000_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \product[6]$_DFFE_PP0P_  (.D(_014_),
    .RN(_000_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \product[7]$_DFFE_PP0P_  (.D(_015_),
    .RN(_000_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \product[8]$_DFFE_PP0P_  (.D(_016_),
    .RN(_000_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net34));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \product[9]$_DFFE_PP0P_  (.D(_017_),
    .RN(_000_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net35));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \start_r$_DFF_PP0_  (.D(net18),
    .RN(_000_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(start_r));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \state$_DFF_PP0_  (.D(_374_),
    .RN(_000_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(state));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Right_145 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Right_146 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Right_147 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Right_148 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Right_149 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Right_150 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Right_151 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Right_152 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Right_153 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Right_154 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Right_155 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Right_156 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Right_157 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Right_158 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_159_Right_159 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_160_Right_160 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_161_Right_161 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_162_Right_162 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_163_Right_163 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_164_Right_164 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_165_Right_165 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_166_Right_166 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_167_Right_167 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_168_Right_168 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_169_Right_169 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_170_Right_170 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_171_Right_171 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_172_Right_172 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_173_Right_173 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_174_Right_174 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_175_Right_175 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_176_Right_176 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_177_Right_177 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_178_Right_178 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_179_Right_179 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_180_Right_180 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_181_Right_181 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_182_Right_182 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_183_Right_183 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_184_Right_184 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_185_Right_185 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_186_Right_186 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_187_Right_187 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_188_Right_188 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_189_Right_189 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_190_Right_190 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_191_Right_191 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_192_Right_192 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_193_Right_193 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_194_Right_194 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_195_Right_195 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_196_Right_196 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_197_Right_197 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_198_Right_198 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_199_Right_199 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_200_Right_200 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_201_Right_201 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_202_Right_202 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_203_Right_203 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_204_Right_204 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_205_Right_205 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_206_Right_206 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_207_Right_207 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_208_Right_208 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_209_Right_209 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_210_Right_210 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_211_Right_211 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_212_Right_212 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_213_Right_213 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_214_Right_214 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_215_Right_215 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_216_Right_216 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_217_Right_217 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_218_Right_218 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_219_Right_219 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_220_Right_220 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_221_Right_221 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_222_Right_222 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_223_Right_223 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_224_Right_224 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_225_Right_225 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_226_Right_226 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_227_Right_227 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_228_Right_228 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_229_Right_229 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_230_Right_230 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_231_Right_231 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_232_Right_232 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_233_Right_233 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_234_Right_234 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_235_Right_235 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_236_Right_236 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_237_Right_237 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_238_Right_238 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_239_Right_239 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_240_Right_240 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_241_Right_241 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_242_Right_242 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_243_Right_243 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_244_Right_244 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_245_Right_245 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_246_Right_246 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_247_Right_247 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_248_Right_248 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_249_Right_249 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_250_Right_250 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_251_Right_251 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_252_Right_252 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_253_Right_253 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_254_Right_254 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_255_Right_255 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_256_Right_256 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_257_Right_257 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_258_Right_258 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_259_Right_259 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_260_Right_260 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_261_Right_261 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_262_Right_262 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_263_Right_263 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_264_Right_264 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_265_Right_265 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_266_Right_266 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_267_Right_267 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_268_Right_268 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_269_Right_269 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_270_Right_270 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_271_Right_271 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_272_Right_272 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_273_Right_273 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_274_Right_274 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_275_Right_275 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_276_Right_276 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_277_Right_277 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_278_Right_278 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_279_Right_279 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_280_Right_280 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_281_Right_281 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_282_Right_282 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_283_Right_283 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_284_Right_284 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_285_Right_285 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_286_Right_286 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_287_Right_287 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_288_Right_288 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_289_Right_289 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_290_Right_290 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_291_Right_291 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_292_Right_292 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_293_Right_293 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_294_Right_294 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_295_Right_295 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_296_Right_296 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_297_Right_297 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_298_Right_298 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_299_Right_299 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_300_Right_300 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_301_Right_301 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_302_Right_302 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_303_Right_303 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_304_Right_304 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_305_Right_305 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_306_Right_306 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_307_Right_307 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_308_Right_308 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_309 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_310 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_311 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_312 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_313 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_314 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_315 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_316 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_317 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_318 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_319 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_320 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_321 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_322 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_323 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_324 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_325 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_326 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_327 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_328 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_329 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_330 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_331 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_332 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_333 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_334 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_335 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_336 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_337 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_338 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_339 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_340 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_341 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_342 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_343 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_344 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_345 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_346 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_347 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_348 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_349 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_350 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_351 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Left_352 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Left_353 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Left_354 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Left_355 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Left_356 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Left_357 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Left_358 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Left_359 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Left_360 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Left_361 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Left_362 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Left_363 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Left_364 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Left_365 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Left_366 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Left_367 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Left_368 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Left_369 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Left_370 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Left_371 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Left_372 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Left_373 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Left_374 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Left_375 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Left_376 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Left_377 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Left_378 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Left_379 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Left_380 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Left_381 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Left_382 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Left_383 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Left_384 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Left_385 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Left_386 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Left_387 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Left_388 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Left_389 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Left_390 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Left_391 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Left_392 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Left_393 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Left_394 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Left_395 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Left_396 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Left_397 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Left_398 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Left_399 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Left_400 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Left_401 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Left_402 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Left_403 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Left_404 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Left_405 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Left_406 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Left_407 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Left_408 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Left_409 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Left_410 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Left_411 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Left_412 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Left_413 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Left_414 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Left_415 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Left_416 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Left_417 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Left_418 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Left_419 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Left_420 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Left_421 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Left_422 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Left_423 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Left_424 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Left_425 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Left_426 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Left_427 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Left_428 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Left_429 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Left_430 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Left_431 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Left_432 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Left_433 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Left_434 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Left_435 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Left_436 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Left_437 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Left_438 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Left_439 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Left_440 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Left_441 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Left_442 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Left_443 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Left_444 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Left_445 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Left_446 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Left_447 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Left_448 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Left_449 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Left_450 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Left_451 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Left_452 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Left_453 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Left_454 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Left_455 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Left_456 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Left_457 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Left_458 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Left_459 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Left_460 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Left_461 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Left_462 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Left_463 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Left_464 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Left_465 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Left_466 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Left_467 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_159_Left_468 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_160_Left_469 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_161_Left_470 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_162_Left_471 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_163_Left_472 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_164_Left_473 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_165_Left_474 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_166_Left_475 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_167_Left_476 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_168_Left_477 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_169_Left_478 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_170_Left_479 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_171_Left_480 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_172_Left_481 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_173_Left_482 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_174_Left_483 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_175_Left_484 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_176_Left_485 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_177_Left_486 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_178_Left_487 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_179_Left_488 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_180_Left_489 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_181_Left_490 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_182_Left_491 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_183_Left_492 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_184_Left_493 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_185_Left_494 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_186_Left_495 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_187_Left_496 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_188_Left_497 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_189_Left_498 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_190_Left_499 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_191_Left_500 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_192_Left_501 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_193_Left_502 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_194_Left_503 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_195_Left_504 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_196_Left_505 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_197_Left_506 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_198_Left_507 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_199_Left_508 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_200_Left_509 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_201_Left_510 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_202_Left_511 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_203_Left_512 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_204_Left_513 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_205_Left_514 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_206_Left_515 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_207_Left_516 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_208_Left_517 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_209_Left_518 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_210_Left_519 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_211_Left_520 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_212_Left_521 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_213_Left_522 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_214_Left_523 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_215_Left_524 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_216_Left_525 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_217_Left_526 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_218_Left_527 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_219_Left_528 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_220_Left_529 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_221_Left_530 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_222_Left_531 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_223_Left_532 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_224_Left_533 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_225_Left_534 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_226_Left_535 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_227_Left_536 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_228_Left_537 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_229_Left_538 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_230_Left_539 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_231_Left_540 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_232_Left_541 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_233_Left_542 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_234_Left_543 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_235_Left_544 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_236_Left_545 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_237_Left_546 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_238_Left_547 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_239_Left_548 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_240_Left_549 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_241_Left_550 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_242_Left_551 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_243_Left_552 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_244_Left_553 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_245_Left_554 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_246_Left_555 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_247_Left_556 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_248_Left_557 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_249_Left_558 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_250_Left_559 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_251_Left_560 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_252_Left_561 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_253_Left_562 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_254_Left_563 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_255_Left_564 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_256_Left_565 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_257_Left_566 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_258_Left_567 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_259_Left_568 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_260_Left_569 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_261_Left_570 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_262_Left_571 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_263_Left_572 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_264_Left_573 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_265_Left_574 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_266_Left_575 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_267_Left_576 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_268_Left_577 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_269_Left_578 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_270_Left_579 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_271_Left_580 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_272_Left_581 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_273_Left_582 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_274_Left_583 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_275_Left_584 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_276_Left_585 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_277_Left_586 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_278_Left_587 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_279_Left_588 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_280_Left_589 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_281_Left_590 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_282_Left_591 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_283_Left_592 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_284_Left_593 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_285_Left_594 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_286_Left_595 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_287_Left_596 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_288_Left_597 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_289_Left_598 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_290_Left_599 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_291_Left_600 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_292_Left_601 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_293_Left_602 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_294_Left_603 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_295_Left_604 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_296_Left_605 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_297_Left_606 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_298_Left_607 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_299_Left_608 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_300_Left_609 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_301_Left_610 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_302_Left_611 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_303_Left_612 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_304_Left_613 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_305_Left_614 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_306_Left_615 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_307_Left_616 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_308_Left_617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_961 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_962 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_963 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_964 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_965 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_966 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_967 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_968 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_969 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_970 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_971 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_972 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_973 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_974 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_975 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_976 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_977 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_978 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_979 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_980 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_981 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_982 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_983 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_984 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_985 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_986 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_987 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_988 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_989 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_990 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_991 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_992 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_993 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_994 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_995 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_996 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_997 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_998 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_999 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1961 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1962 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1963 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1965 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1966 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1967 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1969 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1971 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1978 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1981 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1983 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1985 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1987 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1988 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1989 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1991 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1993 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1995 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1998 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_2001 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_2003 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_2004 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_2010 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_2014 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_2015 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_2017 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_2018 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_2019 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_2020 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_2023 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_2025 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_2027 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_2028 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_2029 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_2030 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_2031 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_2032 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_2033 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_2034 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_2035 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_2036 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_2037 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_2039 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_2041 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_2043 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_2044 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_2045 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_2047 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_2048 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_2051 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_2052 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_2053 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_2054 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_2059 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_2060 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_2061 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_2063 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_2065 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_2067 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_2069 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_2071 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_2072 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_2073 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_2074 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_2075 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_2076 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_2077 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_2078 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_2080 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_2082 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_2085 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_2086 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_2087 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_2089 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_2090 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_2091 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_2092 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_2093 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_2096 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_2098 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_2099 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_2100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_2107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_2112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_2121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_2123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_2125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_2127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_2128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_2136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_2137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_2139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_2140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_2141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_2142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_2143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_2144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_2145 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_2146 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_2147 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_2148 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_2149 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_2150 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_2151 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_2153 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_2155 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_2156 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_2157 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_2158 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_2159 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_2160 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_2161 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_2163 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_2164 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_2165 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_2166 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_2167 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_2168 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_2169 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_2170 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_2171 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_2172 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_2173 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_2174 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_2175 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_2176 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_2177 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_2178 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_2179 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_2180 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_2181 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_2182 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_2183 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_2184 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_2185 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_2186 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_2187 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_2188 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_2189 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_2190 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_2191 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_2192 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_2193 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_2194 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_2195 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_2196 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_2197 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_2198 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_2199 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_2200 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_2201 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_2203 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_2204 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_2205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_2206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_2207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_2208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_2209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_2210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_2211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_2212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_2213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_2217 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_2221 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_2222 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_2223 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_2224 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_2225 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_2226 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_2227 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_2228 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_2229 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_2230 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_2231 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_2232 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_2233 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_2234 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_2235 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_2236 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_2237 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_2238 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_2239 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_2240 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_2241 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_2242 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_2243 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_2244 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_2245 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_2246 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_2247 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_2248 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_2249 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_2250 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_2251 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_2252 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_2253 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_2254 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_2255 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_2256 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_2257 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_2258 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_2259 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_2260 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_2261 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_2262 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_2263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_2264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_2265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_2267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_2268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_2269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_2270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_2271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_2272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_2273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_2274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_2275 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_2276 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_2277 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_2278 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_2279 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_2281 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_2282 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_2283 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_2284 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_2285 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_2286 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_2287 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_2288 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_2289 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_2290 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_2291 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_2292 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_2293 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_2294 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_2295 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_2296 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_2297 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_2298 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_2299 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_2300 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_2301 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_2302 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_2303 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_2304 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_2305 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_2306 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_2307 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_2308 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_2309 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_2310 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_2311 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_2314 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_2315 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_2317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_2318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_2319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_2320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_2321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_2322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_2323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_2324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_2325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_2326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_2327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_2328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_2329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_2331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_2332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_2333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_2334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_2335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_2336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_2337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_2338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_2339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_2340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_2341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_2342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_2343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_2344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_2345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_2346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_2347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_2348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_2349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_2350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_2351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_2352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_2353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_2354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_2355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_2356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_2357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_2358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_2359 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_2360 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_2361 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_2362 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_2363 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_2364 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_2365 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_2366 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_2367 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_2368 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_2369 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_2370 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_2371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_2372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_2373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_2374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_2375 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_2376 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_2377 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_2378 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_2379 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_2381 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_2382 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_2383 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_2384 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_2385 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_2386 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_2387 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_2388 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_2389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_2390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_2391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_2392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_2393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_2395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_2396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_2397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_2398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_2399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_2400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_2401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_2402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_2403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_2404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_2405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_2406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_2407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_2408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_2409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_2410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_2411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_2412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_2413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_2414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_2415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_2416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_2417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_2418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_2419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_2420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_2421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_2422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_2423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_2424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_2425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_2426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_2427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_2428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_2429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_2430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_2431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_2432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_2433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_2434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_2435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_2436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_2437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_2438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_2439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_2440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_2441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_2442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_2443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_2445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_2446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_2447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_2448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_2449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_2450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_2451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_2452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_2453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_2454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_2455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_2456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_2457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_2459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_2460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_2461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_2462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_2463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_2464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_2465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_2466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_2467 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_2468 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_2469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_2470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_2471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_2472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_2473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_2474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_2475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_2476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_2477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_2478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_2479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_2480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_2481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_2482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_2483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_2484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_2485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_2486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_2487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_2488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_2489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_2492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_2493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_2495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_2496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_2497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_2498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_2499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_2500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_2501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_2502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_2503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_2504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_2505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_2506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_2507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_2509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_2510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_2511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_2512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_2513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_2514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_2515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_2516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_2517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_2518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_2519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_2520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_2521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_2522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_2523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_2524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_2525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_2526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_2527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_2528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_2529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_2530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_2531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_2532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_2533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_2534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_2535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_2536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_2537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_2538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_2539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_2540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_2541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_2542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_2543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_2544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_2545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_2546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_2547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_2548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_2549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_2550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_2551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_2552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_2553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_2554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_2555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_2556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_2557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_2559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_2560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_2561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_2562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_2563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_2564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_2565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_2566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_2567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_2568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_2569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_2570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_2571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_2573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_2574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_2575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_2576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_2577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_2578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_2579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_2580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_2581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_2582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_2583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_2584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_2585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_2586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_2587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_2588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_2589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_2590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_2591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_2592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_2593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_2594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_2595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_2596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_2597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_2598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_2599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_2600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_2601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_2602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_2603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_2604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_2605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_2606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_2607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_2608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_2609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_2610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_2611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_2612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_2613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_2614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_2615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_2616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_2617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_2618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_2619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_2620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_2621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_2623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_2624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_2625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_2626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_2627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_2628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_2629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_2630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_2631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_2632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_2633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_2634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_2635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_2637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_2639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_2640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_2641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_2642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_2643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_2644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_2645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_2647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_2648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_2649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_2651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_2652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_2653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_2654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_2655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_2656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_2657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_2658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_2659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_2660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_2661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_2662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_2663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_2664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_2665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_2666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_2667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_2669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_2670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_2671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_2673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_2674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_2675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_2676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_2677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_2678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_2679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_2680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_2681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_2682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_2683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_2684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_2685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_2687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_2688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_2689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_2690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_2691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_2692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_2693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_2694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_2695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_2696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_2697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_2698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_2699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_2700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_2701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_2702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_2703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_2704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_2705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_2706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_2707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_2708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_2709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_2710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_2711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_2712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_2713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_2714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_2715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_2716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_2717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_2718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_2719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_2720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_2721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_2722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_2723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_2724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_2725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_2726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_2727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_2728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_2729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_2730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_2731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_2732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_2733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_2734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_2735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_2737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_2738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_2739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_2740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_2741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_2742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_2743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_2744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_2745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_2746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_2747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_2748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_2749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_2751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_2752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_2753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_2754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_2755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_2756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_2757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_2758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_2759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_2760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_2761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_2762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_2763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_2764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_2765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_2766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_2767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_2769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_2770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_2771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_2772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_2773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_2774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_2775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_2776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_2777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_2778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_2779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_2780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_2781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_2783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_2785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_2786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_2787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_2789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_2791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_2792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_2793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_2794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_2795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_2796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_2797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_2798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_2799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_2801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_2802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_2803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_2804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_2805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_2806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_2807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_2808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_2809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_2810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_2811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_2812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_2813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_2815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_2816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_2817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_2818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_2819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_2820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_2821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_2822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_2823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_2824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_2825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_2826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_2827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_2828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_2829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_2830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_2831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_2832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_2833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_2834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_2835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_2836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_2837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_2838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_2839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_2840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_2841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_2842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_2843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_2844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_2845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_2847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_2848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_2849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_2851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_2852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_2853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_2854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_2855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_2856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_2857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_2858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_2859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_2860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_2861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_2862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_2863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_2865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_2866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_2867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_2868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_2869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_2870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_2871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_2872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_2873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_2874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_2875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_2876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_2877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_2878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_2879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_2880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_2881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_2882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_2883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_2884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_2885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_2886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_2887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_2888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_2889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_2890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_2891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_2892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_2893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_2894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_2895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_2896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_2897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_2898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_2899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_2900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_2901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_2902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_2903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_2904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_2905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_2906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_2907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_2908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_2909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_2910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_2911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_2912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_2913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_2915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_2916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_2917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_2918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_2919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_2920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_2921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_2922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_2923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_2924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_2925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_2926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_2927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_2929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_2930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_2931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_2932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_2933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_2934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_2935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_2936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_2937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_2938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_2939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_2940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_2941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_2942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_2943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_2944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_2945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_2946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_2947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_2948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_2949 ();
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input1 (.I(multiplicand[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input2 (.I(multiplicand[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input3 (.I(multiplicand[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input4 (.I(multiplicand[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input5 (.I(multiplicand[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input6 (.I(multiplicand[5]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input7 (.I(multiplicand[6]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input8 (.I(multiplicand[7]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input9 (.I(multiplier[0]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input10 (.I(multiplier[1]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input11 (.I(multiplier[2]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input12 (.I(multiplier[3]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input13 (.I(multiplier[4]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input14 (.I(multiplier[5]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input15 (.I(multiplier[6]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input16 (.I(multiplier[7]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input17 (.I(rst),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input18 (.I(start),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output19 (.I(net19),
    .Z(done));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output20 (.I(net20),
    .Z(product[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output21 (.I(net21),
    .Z(product[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output22 (.I(net22),
    .Z(product[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output23 (.I(net23),
    .Z(product[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output24 (.I(net24),
    .Z(product[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output25 (.I(net25),
    .Z(product[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output26 (.I(net26),
    .Z(product[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output27 (.I(net27),
    .Z(product[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output28 (.I(net28),
    .Z(product[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output29 (.I(net29),
    .Z(product[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output30 (.I(net30),
    .Z(product[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output31 (.I(net31),
    .Z(product[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output32 (.I(net32),
    .Z(product[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output33 (.I(net33),
    .Z(product[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output34 (.I(net34),
    .Z(product[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output35 (.I(net35),
    .Z(product[9]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload0 (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_1 (.I(net15));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_2 (.I(net11));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_2753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_2785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_2789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_2753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_2785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_2789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_2718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_2734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_2753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_2785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_2789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_2753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_2785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_2789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_208_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_208_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_210_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_210_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_214_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_214_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_215_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_216_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_216_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_218_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_218_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_219_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_220_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_220_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_221_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_222_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_222_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_223_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_224_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_224_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_227_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_228_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_228_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_229_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_230_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_230_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_230_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_231_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_232_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_232_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_233_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_233_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_234_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_234_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_235_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_235_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_236_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_236_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_236_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_236_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_237_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_237_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_238_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_238_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_238_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_238_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_239_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_239_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_240_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_240_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_240_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_240_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_241_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_241_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_242_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_242_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_242_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_242_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_243_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_243_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_244_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_244_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_244_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_244_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_245_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_245_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_246_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_246_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_246_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_246_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_247_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_247_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_248_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_248_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_248_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_248_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_249_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_249_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_250_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_250_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_250_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_250_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_251_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_251_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_252_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_252_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_252_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_252_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_253_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_253_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_254_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_254_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_254_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_254_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_255_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_255_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_256_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_256_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_256_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_256_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_257_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_257_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_258_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_258_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_258_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_258_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_259_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_259_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_260_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_260_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_260_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_260_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_261_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_261_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_262_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_262_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_262_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_262_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_263_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_263_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_264_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_264_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_264_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_264_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_265_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_265_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_266_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_266_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_266_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_266_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_267_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_267_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_268_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_268_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_268_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_268_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_269_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_269_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_270_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_270_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_270_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_270_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_271_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_271_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_272_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_272_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_272_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_272_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_273_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_273_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_274_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_274_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_274_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_274_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_275_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_275_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_276_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_276_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_276_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_276_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_277_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_277_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_278_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_278_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_278_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_278_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_279_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_279_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_280_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_280_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_280_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_280_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_281_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_281_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_282_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_282_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_282_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_282_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_283_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_283_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_284_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_284_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_284_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_284_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_285_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_285_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_286_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_286_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_286_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_286_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_287_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_287_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_288_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_288_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_288_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_288_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_289_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_289_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_290_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_290_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_290_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_290_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_291_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_291_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_292_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_292_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_292_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_292_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_293_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_293_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_294_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_294_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_294_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_294_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_295_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_295_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_296_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_296_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_296_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_296_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_297_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_297_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_298_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_298_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_298_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_298_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_299_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_299_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_300_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_300_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_300_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_300_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_301_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_301_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_302_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_302_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_302_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_302_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_303_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_303_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_304_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_304_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_304_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_304_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_305_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_305_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_306_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_306_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_306_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_306_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_307_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_307_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_307_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_307_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_307_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_307_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_307_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_307_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_307_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_307_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_307_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_308_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_308_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_308_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_308_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_308_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_308_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_308_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_308_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_308_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_308_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_308_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_308_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_308_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_308_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_308_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_308_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_308_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_308_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_308_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_308_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_308_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_308_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_308_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_308_2298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_308_2476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_308_2654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_308_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_308_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_308_2790 ();
endmodule
