module riscv (clk,
    memread,
    memwrite,
    reset,
    suspend,
    aluout,
    instr,
    pc,
    readdata,
    writedata);
 input clk;
 output memread;
 output memwrite;
 input reset;
 output suspend;
 output [31:0] aluout;
 input [31:0] instr;
 output [31:0] pc;
 input [31:0] readdata;
 output [31:0] writedata;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire net221;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire net275;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire net264;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire net181;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire net168;
 wire net187;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire net175;
 wire _02816_;
 wire net164;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire net167;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire \dp.ISRmux.d0[10] ;
 wire \dp.ISRmux.d0[11] ;
 wire \dp.ISRmux.d0[12] ;
 wire \dp.ISRmux.d0[13] ;
 wire \dp.ISRmux.d0[14] ;
 wire \dp.ISRmux.d0[15] ;
 wire \dp.ISRmux.d0[16] ;
 wire \dp.ISRmux.d0[17] ;
 wire \dp.ISRmux.d0[18] ;
 wire \dp.ISRmux.d0[19] ;
 wire \dp.ISRmux.d0[20] ;
 wire \dp.ISRmux.d0[21] ;
 wire \dp.ISRmux.d0[22] ;
 wire \dp.ISRmux.d0[23] ;
 wire \dp.ISRmux.d0[24] ;
 wire \dp.ISRmux.d0[25] ;
 wire \dp.ISRmux.d0[26] ;
 wire \dp.ISRmux.d0[27] ;
 wire \dp.ISRmux.d0[28] ;
 wire \dp.ISRmux.d0[29] ;
 wire \dp.ISRmux.d0[2] ;
 wire \dp.ISRmux.d0[30] ;
 wire \dp.ISRmux.d0[31] ;
 wire \dp.ISRmux.d0[3] ;
 wire \dp.ISRmux.d0[4] ;
 wire \dp.ISRmux.d0[5] ;
 wire \dp.ISRmux.d0[6] ;
 wire \dp.ISRmux.d0[7] ;
 wire \dp.ISRmux.d0[8] ;
 wire \dp.ISRmux.d0[9] ;
 wire \dp.rf.rf[0][0] ;
 wire \dp.rf.rf[0][10] ;
 wire \dp.rf.rf[0][11] ;
 wire \dp.rf.rf[0][12] ;
 wire \dp.rf.rf[0][13] ;
 wire \dp.rf.rf[0][14] ;
 wire \dp.rf.rf[0][15] ;
 wire \dp.rf.rf[0][16] ;
 wire \dp.rf.rf[0][17] ;
 wire \dp.rf.rf[0][18] ;
 wire \dp.rf.rf[0][19] ;
 wire \dp.rf.rf[0][1] ;
 wire \dp.rf.rf[0][20] ;
 wire \dp.rf.rf[0][21] ;
 wire \dp.rf.rf[0][22] ;
 wire \dp.rf.rf[0][23] ;
 wire \dp.rf.rf[0][24] ;
 wire \dp.rf.rf[0][25] ;
 wire \dp.rf.rf[0][26] ;
 wire \dp.rf.rf[0][27] ;
 wire \dp.rf.rf[0][28] ;
 wire \dp.rf.rf[0][29] ;
 wire \dp.rf.rf[0][2] ;
 wire \dp.rf.rf[0][30] ;
 wire \dp.rf.rf[0][31] ;
 wire \dp.rf.rf[0][3] ;
 wire \dp.rf.rf[0][4] ;
 wire \dp.rf.rf[0][5] ;
 wire \dp.rf.rf[0][6] ;
 wire \dp.rf.rf[0][7] ;
 wire \dp.rf.rf[0][8] ;
 wire \dp.rf.rf[0][9] ;
 wire \dp.rf.rf[10][0] ;
 wire \dp.rf.rf[10][10] ;
 wire \dp.rf.rf[10][11] ;
 wire \dp.rf.rf[10][12] ;
 wire \dp.rf.rf[10][13] ;
 wire \dp.rf.rf[10][14] ;
 wire \dp.rf.rf[10][15] ;
 wire \dp.rf.rf[10][16] ;
 wire \dp.rf.rf[10][17] ;
 wire \dp.rf.rf[10][18] ;
 wire \dp.rf.rf[10][19] ;
 wire \dp.rf.rf[10][1] ;
 wire \dp.rf.rf[10][20] ;
 wire \dp.rf.rf[10][21] ;
 wire \dp.rf.rf[10][22] ;
 wire \dp.rf.rf[10][23] ;
 wire \dp.rf.rf[10][24] ;
 wire \dp.rf.rf[10][25] ;
 wire \dp.rf.rf[10][26] ;
 wire \dp.rf.rf[10][27] ;
 wire \dp.rf.rf[10][28] ;
 wire \dp.rf.rf[10][29] ;
 wire \dp.rf.rf[10][2] ;
 wire \dp.rf.rf[10][30] ;
 wire \dp.rf.rf[10][31] ;
 wire \dp.rf.rf[10][3] ;
 wire \dp.rf.rf[10][4] ;
 wire \dp.rf.rf[10][5] ;
 wire \dp.rf.rf[10][6] ;
 wire \dp.rf.rf[10][7] ;
 wire \dp.rf.rf[10][8] ;
 wire \dp.rf.rf[10][9] ;
 wire \dp.rf.rf[11][0] ;
 wire \dp.rf.rf[11][10] ;
 wire \dp.rf.rf[11][11] ;
 wire \dp.rf.rf[11][12] ;
 wire \dp.rf.rf[11][13] ;
 wire \dp.rf.rf[11][14] ;
 wire \dp.rf.rf[11][15] ;
 wire \dp.rf.rf[11][16] ;
 wire \dp.rf.rf[11][17] ;
 wire \dp.rf.rf[11][18] ;
 wire \dp.rf.rf[11][19] ;
 wire \dp.rf.rf[11][1] ;
 wire \dp.rf.rf[11][20] ;
 wire \dp.rf.rf[11][21] ;
 wire \dp.rf.rf[11][22] ;
 wire \dp.rf.rf[11][23] ;
 wire \dp.rf.rf[11][24] ;
 wire \dp.rf.rf[11][25] ;
 wire \dp.rf.rf[11][26] ;
 wire \dp.rf.rf[11][27] ;
 wire \dp.rf.rf[11][28] ;
 wire \dp.rf.rf[11][29] ;
 wire \dp.rf.rf[11][2] ;
 wire \dp.rf.rf[11][30] ;
 wire \dp.rf.rf[11][31] ;
 wire \dp.rf.rf[11][3] ;
 wire \dp.rf.rf[11][4] ;
 wire \dp.rf.rf[11][5] ;
 wire \dp.rf.rf[11][6] ;
 wire \dp.rf.rf[11][7] ;
 wire \dp.rf.rf[11][8] ;
 wire \dp.rf.rf[11][9] ;
 wire \dp.rf.rf[12][0] ;
 wire \dp.rf.rf[12][10] ;
 wire \dp.rf.rf[12][11] ;
 wire \dp.rf.rf[12][12] ;
 wire \dp.rf.rf[12][13] ;
 wire \dp.rf.rf[12][14] ;
 wire \dp.rf.rf[12][15] ;
 wire \dp.rf.rf[12][16] ;
 wire \dp.rf.rf[12][17] ;
 wire \dp.rf.rf[12][18] ;
 wire \dp.rf.rf[12][19] ;
 wire \dp.rf.rf[12][1] ;
 wire \dp.rf.rf[12][20] ;
 wire \dp.rf.rf[12][21] ;
 wire \dp.rf.rf[12][22] ;
 wire \dp.rf.rf[12][23] ;
 wire \dp.rf.rf[12][24] ;
 wire \dp.rf.rf[12][25] ;
 wire \dp.rf.rf[12][26] ;
 wire \dp.rf.rf[12][27] ;
 wire \dp.rf.rf[12][28] ;
 wire \dp.rf.rf[12][29] ;
 wire \dp.rf.rf[12][2] ;
 wire \dp.rf.rf[12][30] ;
 wire \dp.rf.rf[12][31] ;
 wire \dp.rf.rf[12][3] ;
 wire \dp.rf.rf[12][4] ;
 wire \dp.rf.rf[12][5] ;
 wire \dp.rf.rf[12][6] ;
 wire \dp.rf.rf[12][7] ;
 wire \dp.rf.rf[12][8] ;
 wire \dp.rf.rf[12][9] ;
 wire \dp.rf.rf[13][0] ;
 wire \dp.rf.rf[13][10] ;
 wire \dp.rf.rf[13][11] ;
 wire \dp.rf.rf[13][12] ;
 wire \dp.rf.rf[13][13] ;
 wire \dp.rf.rf[13][14] ;
 wire \dp.rf.rf[13][15] ;
 wire \dp.rf.rf[13][16] ;
 wire \dp.rf.rf[13][17] ;
 wire \dp.rf.rf[13][18] ;
 wire \dp.rf.rf[13][19] ;
 wire \dp.rf.rf[13][1] ;
 wire \dp.rf.rf[13][20] ;
 wire \dp.rf.rf[13][21] ;
 wire \dp.rf.rf[13][22] ;
 wire \dp.rf.rf[13][23] ;
 wire \dp.rf.rf[13][24] ;
 wire \dp.rf.rf[13][25] ;
 wire \dp.rf.rf[13][26] ;
 wire \dp.rf.rf[13][27] ;
 wire \dp.rf.rf[13][28] ;
 wire \dp.rf.rf[13][29] ;
 wire \dp.rf.rf[13][2] ;
 wire \dp.rf.rf[13][30] ;
 wire \dp.rf.rf[13][31] ;
 wire \dp.rf.rf[13][3] ;
 wire \dp.rf.rf[13][4] ;
 wire \dp.rf.rf[13][5] ;
 wire \dp.rf.rf[13][6] ;
 wire \dp.rf.rf[13][7] ;
 wire \dp.rf.rf[13][8] ;
 wire \dp.rf.rf[13][9] ;
 wire \dp.rf.rf[14][0] ;
 wire \dp.rf.rf[14][10] ;
 wire \dp.rf.rf[14][11] ;
 wire \dp.rf.rf[14][12] ;
 wire \dp.rf.rf[14][13] ;
 wire \dp.rf.rf[14][14] ;
 wire \dp.rf.rf[14][15] ;
 wire \dp.rf.rf[14][16] ;
 wire \dp.rf.rf[14][17] ;
 wire \dp.rf.rf[14][18] ;
 wire \dp.rf.rf[14][19] ;
 wire \dp.rf.rf[14][1] ;
 wire \dp.rf.rf[14][20] ;
 wire \dp.rf.rf[14][21] ;
 wire \dp.rf.rf[14][22] ;
 wire \dp.rf.rf[14][23] ;
 wire \dp.rf.rf[14][24] ;
 wire \dp.rf.rf[14][25] ;
 wire \dp.rf.rf[14][26] ;
 wire \dp.rf.rf[14][27] ;
 wire \dp.rf.rf[14][28] ;
 wire \dp.rf.rf[14][29] ;
 wire \dp.rf.rf[14][2] ;
 wire \dp.rf.rf[14][30] ;
 wire \dp.rf.rf[14][31] ;
 wire \dp.rf.rf[14][3] ;
 wire \dp.rf.rf[14][4] ;
 wire \dp.rf.rf[14][5] ;
 wire \dp.rf.rf[14][6] ;
 wire \dp.rf.rf[14][7] ;
 wire \dp.rf.rf[14][8] ;
 wire \dp.rf.rf[14][9] ;
 wire \dp.rf.rf[15][0] ;
 wire \dp.rf.rf[15][10] ;
 wire \dp.rf.rf[15][11] ;
 wire \dp.rf.rf[15][12] ;
 wire \dp.rf.rf[15][13] ;
 wire \dp.rf.rf[15][14] ;
 wire \dp.rf.rf[15][15] ;
 wire \dp.rf.rf[15][16] ;
 wire \dp.rf.rf[15][17] ;
 wire \dp.rf.rf[15][18] ;
 wire \dp.rf.rf[15][19] ;
 wire \dp.rf.rf[15][1] ;
 wire \dp.rf.rf[15][20] ;
 wire \dp.rf.rf[15][21] ;
 wire \dp.rf.rf[15][22] ;
 wire \dp.rf.rf[15][23] ;
 wire \dp.rf.rf[15][24] ;
 wire \dp.rf.rf[15][25] ;
 wire \dp.rf.rf[15][26] ;
 wire \dp.rf.rf[15][27] ;
 wire \dp.rf.rf[15][28] ;
 wire \dp.rf.rf[15][29] ;
 wire \dp.rf.rf[15][2] ;
 wire \dp.rf.rf[15][30] ;
 wire \dp.rf.rf[15][31] ;
 wire \dp.rf.rf[15][3] ;
 wire \dp.rf.rf[15][4] ;
 wire \dp.rf.rf[15][5] ;
 wire \dp.rf.rf[15][6] ;
 wire \dp.rf.rf[15][7] ;
 wire \dp.rf.rf[15][8] ;
 wire \dp.rf.rf[15][9] ;
 wire \dp.rf.rf[16][0] ;
 wire \dp.rf.rf[16][10] ;
 wire \dp.rf.rf[16][11] ;
 wire \dp.rf.rf[16][12] ;
 wire \dp.rf.rf[16][13] ;
 wire \dp.rf.rf[16][14] ;
 wire \dp.rf.rf[16][15] ;
 wire \dp.rf.rf[16][16] ;
 wire \dp.rf.rf[16][17] ;
 wire \dp.rf.rf[16][18] ;
 wire \dp.rf.rf[16][19] ;
 wire \dp.rf.rf[16][1] ;
 wire \dp.rf.rf[16][20] ;
 wire \dp.rf.rf[16][21] ;
 wire \dp.rf.rf[16][22] ;
 wire \dp.rf.rf[16][23] ;
 wire \dp.rf.rf[16][24] ;
 wire \dp.rf.rf[16][25] ;
 wire \dp.rf.rf[16][26] ;
 wire \dp.rf.rf[16][27] ;
 wire \dp.rf.rf[16][28] ;
 wire \dp.rf.rf[16][29] ;
 wire \dp.rf.rf[16][2] ;
 wire \dp.rf.rf[16][30] ;
 wire \dp.rf.rf[16][31] ;
 wire \dp.rf.rf[16][3] ;
 wire \dp.rf.rf[16][4] ;
 wire \dp.rf.rf[16][5] ;
 wire \dp.rf.rf[16][6] ;
 wire \dp.rf.rf[16][7] ;
 wire \dp.rf.rf[16][8] ;
 wire \dp.rf.rf[16][9] ;
 wire \dp.rf.rf[17][0] ;
 wire \dp.rf.rf[17][10] ;
 wire \dp.rf.rf[17][11] ;
 wire \dp.rf.rf[17][12] ;
 wire \dp.rf.rf[17][13] ;
 wire \dp.rf.rf[17][14] ;
 wire \dp.rf.rf[17][15] ;
 wire \dp.rf.rf[17][16] ;
 wire \dp.rf.rf[17][17] ;
 wire \dp.rf.rf[17][18] ;
 wire \dp.rf.rf[17][19] ;
 wire \dp.rf.rf[17][1] ;
 wire \dp.rf.rf[17][20] ;
 wire \dp.rf.rf[17][21] ;
 wire \dp.rf.rf[17][22] ;
 wire \dp.rf.rf[17][23] ;
 wire \dp.rf.rf[17][24] ;
 wire \dp.rf.rf[17][25] ;
 wire \dp.rf.rf[17][26] ;
 wire \dp.rf.rf[17][27] ;
 wire \dp.rf.rf[17][28] ;
 wire \dp.rf.rf[17][29] ;
 wire \dp.rf.rf[17][2] ;
 wire \dp.rf.rf[17][30] ;
 wire \dp.rf.rf[17][31] ;
 wire \dp.rf.rf[17][3] ;
 wire \dp.rf.rf[17][4] ;
 wire \dp.rf.rf[17][5] ;
 wire \dp.rf.rf[17][6] ;
 wire \dp.rf.rf[17][7] ;
 wire \dp.rf.rf[17][8] ;
 wire \dp.rf.rf[17][9] ;
 wire \dp.rf.rf[18][0] ;
 wire \dp.rf.rf[18][10] ;
 wire \dp.rf.rf[18][11] ;
 wire \dp.rf.rf[18][12] ;
 wire \dp.rf.rf[18][13] ;
 wire \dp.rf.rf[18][14] ;
 wire \dp.rf.rf[18][15] ;
 wire \dp.rf.rf[18][16] ;
 wire \dp.rf.rf[18][17] ;
 wire \dp.rf.rf[18][18] ;
 wire \dp.rf.rf[18][19] ;
 wire \dp.rf.rf[18][1] ;
 wire \dp.rf.rf[18][20] ;
 wire \dp.rf.rf[18][21] ;
 wire \dp.rf.rf[18][22] ;
 wire \dp.rf.rf[18][23] ;
 wire \dp.rf.rf[18][24] ;
 wire \dp.rf.rf[18][25] ;
 wire \dp.rf.rf[18][26] ;
 wire \dp.rf.rf[18][27] ;
 wire \dp.rf.rf[18][28] ;
 wire \dp.rf.rf[18][29] ;
 wire \dp.rf.rf[18][2] ;
 wire \dp.rf.rf[18][30] ;
 wire \dp.rf.rf[18][31] ;
 wire \dp.rf.rf[18][3] ;
 wire \dp.rf.rf[18][4] ;
 wire \dp.rf.rf[18][5] ;
 wire \dp.rf.rf[18][6] ;
 wire \dp.rf.rf[18][7] ;
 wire \dp.rf.rf[18][8] ;
 wire \dp.rf.rf[18][9] ;
 wire \dp.rf.rf[19][0] ;
 wire \dp.rf.rf[19][10] ;
 wire \dp.rf.rf[19][11] ;
 wire \dp.rf.rf[19][12] ;
 wire \dp.rf.rf[19][13] ;
 wire \dp.rf.rf[19][14] ;
 wire \dp.rf.rf[19][15] ;
 wire \dp.rf.rf[19][16] ;
 wire \dp.rf.rf[19][17] ;
 wire \dp.rf.rf[19][18] ;
 wire \dp.rf.rf[19][19] ;
 wire \dp.rf.rf[19][1] ;
 wire \dp.rf.rf[19][20] ;
 wire \dp.rf.rf[19][21] ;
 wire \dp.rf.rf[19][22] ;
 wire \dp.rf.rf[19][23] ;
 wire \dp.rf.rf[19][24] ;
 wire \dp.rf.rf[19][25] ;
 wire \dp.rf.rf[19][26] ;
 wire \dp.rf.rf[19][27] ;
 wire \dp.rf.rf[19][28] ;
 wire \dp.rf.rf[19][29] ;
 wire \dp.rf.rf[19][2] ;
 wire \dp.rf.rf[19][30] ;
 wire \dp.rf.rf[19][31] ;
 wire \dp.rf.rf[19][3] ;
 wire \dp.rf.rf[19][4] ;
 wire \dp.rf.rf[19][5] ;
 wire \dp.rf.rf[19][6] ;
 wire \dp.rf.rf[19][7] ;
 wire \dp.rf.rf[19][8] ;
 wire \dp.rf.rf[19][9] ;
 wire \dp.rf.rf[1][0] ;
 wire \dp.rf.rf[1][10] ;
 wire \dp.rf.rf[1][11] ;
 wire \dp.rf.rf[1][12] ;
 wire \dp.rf.rf[1][13] ;
 wire \dp.rf.rf[1][14] ;
 wire \dp.rf.rf[1][15] ;
 wire \dp.rf.rf[1][16] ;
 wire \dp.rf.rf[1][17] ;
 wire \dp.rf.rf[1][18] ;
 wire \dp.rf.rf[1][19] ;
 wire \dp.rf.rf[1][1] ;
 wire \dp.rf.rf[1][20] ;
 wire \dp.rf.rf[1][21] ;
 wire \dp.rf.rf[1][22] ;
 wire \dp.rf.rf[1][23] ;
 wire \dp.rf.rf[1][24] ;
 wire \dp.rf.rf[1][25] ;
 wire \dp.rf.rf[1][26] ;
 wire \dp.rf.rf[1][27] ;
 wire \dp.rf.rf[1][28] ;
 wire \dp.rf.rf[1][29] ;
 wire \dp.rf.rf[1][2] ;
 wire \dp.rf.rf[1][30] ;
 wire \dp.rf.rf[1][31] ;
 wire \dp.rf.rf[1][3] ;
 wire \dp.rf.rf[1][4] ;
 wire \dp.rf.rf[1][5] ;
 wire \dp.rf.rf[1][6] ;
 wire \dp.rf.rf[1][7] ;
 wire \dp.rf.rf[1][8] ;
 wire \dp.rf.rf[1][9] ;
 wire \dp.rf.rf[20][0] ;
 wire \dp.rf.rf[20][10] ;
 wire \dp.rf.rf[20][11] ;
 wire \dp.rf.rf[20][12] ;
 wire \dp.rf.rf[20][13] ;
 wire \dp.rf.rf[20][14] ;
 wire \dp.rf.rf[20][15] ;
 wire \dp.rf.rf[20][16] ;
 wire \dp.rf.rf[20][17] ;
 wire \dp.rf.rf[20][18] ;
 wire \dp.rf.rf[20][19] ;
 wire \dp.rf.rf[20][1] ;
 wire \dp.rf.rf[20][20] ;
 wire \dp.rf.rf[20][21] ;
 wire \dp.rf.rf[20][22] ;
 wire \dp.rf.rf[20][23] ;
 wire \dp.rf.rf[20][24] ;
 wire \dp.rf.rf[20][25] ;
 wire \dp.rf.rf[20][26] ;
 wire \dp.rf.rf[20][27] ;
 wire \dp.rf.rf[20][28] ;
 wire \dp.rf.rf[20][29] ;
 wire \dp.rf.rf[20][2] ;
 wire \dp.rf.rf[20][30] ;
 wire \dp.rf.rf[20][31] ;
 wire \dp.rf.rf[20][3] ;
 wire \dp.rf.rf[20][4] ;
 wire \dp.rf.rf[20][5] ;
 wire \dp.rf.rf[20][6] ;
 wire \dp.rf.rf[20][7] ;
 wire \dp.rf.rf[20][8] ;
 wire \dp.rf.rf[20][9] ;
 wire \dp.rf.rf[21][0] ;
 wire \dp.rf.rf[21][10] ;
 wire \dp.rf.rf[21][11] ;
 wire \dp.rf.rf[21][12] ;
 wire \dp.rf.rf[21][13] ;
 wire \dp.rf.rf[21][14] ;
 wire \dp.rf.rf[21][15] ;
 wire \dp.rf.rf[21][16] ;
 wire \dp.rf.rf[21][17] ;
 wire \dp.rf.rf[21][18] ;
 wire \dp.rf.rf[21][19] ;
 wire \dp.rf.rf[21][1] ;
 wire \dp.rf.rf[21][20] ;
 wire \dp.rf.rf[21][21] ;
 wire \dp.rf.rf[21][22] ;
 wire \dp.rf.rf[21][23] ;
 wire \dp.rf.rf[21][24] ;
 wire \dp.rf.rf[21][25] ;
 wire \dp.rf.rf[21][26] ;
 wire \dp.rf.rf[21][27] ;
 wire \dp.rf.rf[21][28] ;
 wire \dp.rf.rf[21][29] ;
 wire \dp.rf.rf[21][2] ;
 wire \dp.rf.rf[21][30] ;
 wire \dp.rf.rf[21][31] ;
 wire \dp.rf.rf[21][3] ;
 wire \dp.rf.rf[21][4] ;
 wire \dp.rf.rf[21][5] ;
 wire \dp.rf.rf[21][6] ;
 wire \dp.rf.rf[21][7] ;
 wire \dp.rf.rf[21][8] ;
 wire \dp.rf.rf[21][9] ;
 wire \dp.rf.rf[22][0] ;
 wire \dp.rf.rf[22][10] ;
 wire \dp.rf.rf[22][11] ;
 wire \dp.rf.rf[22][12] ;
 wire \dp.rf.rf[22][13] ;
 wire \dp.rf.rf[22][14] ;
 wire \dp.rf.rf[22][15] ;
 wire \dp.rf.rf[22][16] ;
 wire \dp.rf.rf[22][17] ;
 wire \dp.rf.rf[22][18] ;
 wire \dp.rf.rf[22][19] ;
 wire \dp.rf.rf[22][1] ;
 wire \dp.rf.rf[22][20] ;
 wire \dp.rf.rf[22][21] ;
 wire \dp.rf.rf[22][22] ;
 wire \dp.rf.rf[22][23] ;
 wire \dp.rf.rf[22][24] ;
 wire \dp.rf.rf[22][25] ;
 wire \dp.rf.rf[22][26] ;
 wire \dp.rf.rf[22][27] ;
 wire \dp.rf.rf[22][28] ;
 wire \dp.rf.rf[22][29] ;
 wire \dp.rf.rf[22][2] ;
 wire \dp.rf.rf[22][30] ;
 wire \dp.rf.rf[22][31] ;
 wire \dp.rf.rf[22][3] ;
 wire \dp.rf.rf[22][4] ;
 wire \dp.rf.rf[22][5] ;
 wire \dp.rf.rf[22][6] ;
 wire \dp.rf.rf[22][7] ;
 wire \dp.rf.rf[22][8] ;
 wire \dp.rf.rf[22][9] ;
 wire \dp.rf.rf[23][0] ;
 wire \dp.rf.rf[23][10] ;
 wire \dp.rf.rf[23][11] ;
 wire \dp.rf.rf[23][12] ;
 wire \dp.rf.rf[23][13] ;
 wire \dp.rf.rf[23][14] ;
 wire \dp.rf.rf[23][15] ;
 wire \dp.rf.rf[23][16] ;
 wire \dp.rf.rf[23][17] ;
 wire \dp.rf.rf[23][18] ;
 wire \dp.rf.rf[23][19] ;
 wire \dp.rf.rf[23][1] ;
 wire \dp.rf.rf[23][20] ;
 wire \dp.rf.rf[23][21] ;
 wire \dp.rf.rf[23][22] ;
 wire \dp.rf.rf[23][23] ;
 wire \dp.rf.rf[23][24] ;
 wire \dp.rf.rf[23][25] ;
 wire \dp.rf.rf[23][26] ;
 wire \dp.rf.rf[23][27] ;
 wire \dp.rf.rf[23][28] ;
 wire \dp.rf.rf[23][29] ;
 wire \dp.rf.rf[23][2] ;
 wire \dp.rf.rf[23][30] ;
 wire \dp.rf.rf[23][31] ;
 wire \dp.rf.rf[23][3] ;
 wire \dp.rf.rf[23][4] ;
 wire \dp.rf.rf[23][5] ;
 wire \dp.rf.rf[23][6] ;
 wire \dp.rf.rf[23][7] ;
 wire \dp.rf.rf[23][8] ;
 wire \dp.rf.rf[23][9] ;
 wire \dp.rf.rf[24][0] ;
 wire \dp.rf.rf[24][10] ;
 wire \dp.rf.rf[24][11] ;
 wire \dp.rf.rf[24][12] ;
 wire \dp.rf.rf[24][13] ;
 wire \dp.rf.rf[24][14] ;
 wire \dp.rf.rf[24][15] ;
 wire \dp.rf.rf[24][16] ;
 wire \dp.rf.rf[24][17] ;
 wire \dp.rf.rf[24][18] ;
 wire \dp.rf.rf[24][19] ;
 wire \dp.rf.rf[24][1] ;
 wire \dp.rf.rf[24][20] ;
 wire \dp.rf.rf[24][21] ;
 wire \dp.rf.rf[24][22] ;
 wire \dp.rf.rf[24][23] ;
 wire \dp.rf.rf[24][24] ;
 wire \dp.rf.rf[24][25] ;
 wire \dp.rf.rf[24][26] ;
 wire \dp.rf.rf[24][27] ;
 wire \dp.rf.rf[24][28] ;
 wire \dp.rf.rf[24][29] ;
 wire \dp.rf.rf[24][2] ;
 wire \dp.rf.rf[24][30] ;
 wire \dp.rf.rf[24][31] ;
 wire \dp.rf.rf[24][3] ;
 wire \dp.rf.rf[24][4] ;
 wire \dp.rf.rf[24][5] ;
 wire \dp.rf.rf[24][6] ;
 wire \dp.rf.rf[24][7] ;
 wire \dp.rf.rf[24][8] ;
 wire \dp.rf.rf[24][9] ;
 wire \dp.rf.rf[25][0] ;
 wire \dp.rf.rf[25][10] ;
 wire \dp.rf.rf[25][11] ;
 wire \dp.rf.rf[25][12] ;
 wire \dp.rf.rf[25][13] ;
 wire \dp.rf.rf[25][14] ;
 wire \dp.rf.rf[25][15] ;
 wire \dp.rf.rf[25][16] ;
 wire \dp.rf.rf[25][17] ;
 wire \dp.rf.rf[25][18] ;
 wire \dp.rf.rf[25][19] ;
 wire \dp.rf.rf[25][1] ;
 wire \dp.rf.rf[25][20] ;
 wire \dp.rf.rf[25][21] ;
 wire \dp.rf.rf[25][22] ;
 wire \dp.rf.rf[25][23] ;
 wire \dp.rf.rf[25][24] ;
 wire \dp.rf.rf[25][25] ;
 wire \dp.rf.rf[25][26] ;
 wire \dp.rf.rf[25][27] ;
 wire \dp.rf.rf[25][28] ;
 wire \dp.rf.rf[25][29] ;
 wire \dp.rf.rf[25][2] ;
 wire \dp.rf.rf[25][30] ;
 wire \dp.rf.rf[25][31] ;
 wire \dp.rf.rf[25][3] ;
 wire \dp.rf.rf[25][4] ;
 wire \dp.rf.rf[25][5] ;
 wire \dp.rf.rf[25][6] ;
 wire \dp.rf.rf[25][7] ;
 wire \dp.rf.rf[25][8] ;
 wire \dp.rf.rf[25][9] ;
 wire \dp.rf.rf[26][0] ;
 wire \dp.rf.rf[26][10] ;
 wire \dp.rf.rf[26][11] ;
 wire \dp.rf.rf[26][12] ;
 wire \dp.rf.rf[26][13] ;
 wire \dp.rf.rf[26][14] ;
 wire \dp.rf.rf[26][15] ;
 wire \dp.rf.rf[26][16] ;
 wire \dp.rf.rf[26][17] ;
 wire \dp.rf.rf[26][18] ;
 wire \dp.rf.rf[26][19] ;
 wire \dp.rf.rf[26][1] ;
 wire \dp.rf.rf[26][20] ;
 wire \dp.rf.rf[26][21] ;
 wire \dp.rf.rf[26][22] ;
 wire \dp.rf.rf[26][23] ;
 wire \dp.rf.rf[26][24] ;
 wire \dp.rf.rf[26][25] ;
 wire \dp.rf.rf[26][26] ;
 wire \dp.rf.rf[26][27] ;
 wire \dp.rf.rf[26][28] ;
 wire \dp.rf.rf[26][29] ;
 wire \dp.rf.rf[26][2] ;
 wire \dp.rf.rf[26][30] ;
 wire \dp.rf.rf[26][31] ;
 wire \dp.rf.rf[26][3] ;
 wire \dp.rf.rf[26][4] ;
 wire \dp.rf.rf[26][5] ;
 wire \dp.rf.rf[26][6] ;
 wire \dp.rf.rf[26][7] ;
 wire \dp.rf.rf[26][8] ;
 wire \dp.rf.rf[26][9] ;
 wire \dp.rf.rf[27][0] ;
 wire \dp.rf.rf[27][10] ;
 wire \dp.rf.rf[27][11] ;
 wire \dp.rf.rf[27][12] ;
 wire \dp.rf.rf[27][13] ;
 wire \dp.rf.rf[27][14] ;
 wire \dp.rf.rf[27][15] ;
 wire \dp.rf.rf[27][16] ;
 wire \dp.rf.rf[27][17] ;
 wire \dp.rf.rf[27][18] ;
 wire \dp.rf.rf[27][19] ;
 wire \dp.rf.rf[27][1] ;
 wire \dp.rf.rf[27][20] ;
 wire \dp.rf.rf[27][21] ;
 wire \dp.rf.rf[27][22] ;
 wire \dp.rf.rf[27][23] ;
 wire \dp.rf.rf[27][24] ;
 wire \dp.rf.rf[27][25] ;
 wire \dp.rf.rf[27][26] ;
 wire \dp.rf.rf[27][27] ;
 wire \dp.rf.rf[27][28] ;
 wire \dp.rf.rf[27][29] ;
 wire \dp.rf.rf[27][2] ;
 wire \dp.rf.rf[27][30] ;
 wire \dp.rf.rf[27][31] ;
 wire \dp.rf.rf[27][3] ;
 wire \dp.rf.rf[27][4] ;
 wire \dp.rf.rf[27][5] ;
 wire \dp.rf.rf[27][6] ;
 wire \dp.rf.rf[27][7] ;
 wire \dp.rf.rf[27][8] ;
 wire \dp.rf.rf[27][9] ;
 wire \dp.rf.rf[28][0] ;
 wire \dp.rf.rf[28][10] ;
 wire \dp.rf.rf[28][11] ;
 wire \dp.rf.rf[28][12] ;
 wire \dp.rf.rf[28][13] ;
 wire \dp.rf.rf[28][14] ;
 wire \dp.rf.rf[28][15] ;
 wire \dp.rf.rf[28][16] ;
 wire \dp.rf.rf[28][17] ;
 wire \dp.rf.rf[28][18] ;
 wire \dp.rf.rf[28][19] ;
 wire \dp.rf.rf[28][1] ;
 wire \dp.rf.rf[28][20] ;
 wire \dp.rf.rf[28][21] ;
 wire \dp.rf.rf[28][22] ;
 wire \dp.rf.rf[28][23] ;
 wire \dp.rf.rf[28][24] ;
 wire \dp.rf.rf[28][25] ;
 wire \dp.rf.rf[28][26] ;
 wire \dp.rf.rf[28][27] ;
 wire \dp.rf.rf[28][28] ;
 wire \dp.rf.rf[28][29] ;
 wire \dp.rf.rf[28][2] ;
 wire \dp.rf.rf[28][30] ;
 wire \dp.rf.rf[28][31] ;
 wire \dp.rf.rf[28][3] ;
 wire \dp.rf.rf[28][4] ;
 wire \dp.rf.rf[28][5] ;
 wire \dp.rf.rf[28][6] ;
 wire \dp.rf.rf[28][7] ;
 wire \dp.rf.rf[28][8] ;
 wire \dp.rf.rf[28][9] ;
 wire \dp.rf.rf[29][0] ;
 wire \dp.rf.rf[29][10] ;
 wire \dp.rf.rf[29][11] ;
 wire \dp.rf.rf[29][12] ;
 wire \dp.rf.rf[29][13] ;
 wire \dp.rf.rf[29][14] ;
 wire \dp.rf.rf[29][15] ;
 wire \dp.rf.rf[29][16] ;
 wire \dp.rf.rf[29][17] ;
 wire \dp.rf.rf[29][18] ;
 wire \dp.rf.rf[29][19] ;
 wire \dp.rf.rf[29][1] ;
 wire \dp.rf.rf[29][20] ;
 wire \dp.rf.rf[29][21] ;
 wire \dp.rf.rf[29][22] ;
 wire \dp.rf.rf[29][23] ;
 wire \dp.rf.rf[29][24] ;
 wire \dp.rf.rf[29][25] ;
 wire \dp.rf.rf[29][26] ;
 wire \dp.rf.rf[29][27] ;
 wire \dp.rf.rf[29][28] ;
 wire \dp.rf.rf[29][29] ;
 wire \dp.rf.rf[29][2] ;
 wire \dp.rf.rf[29][30] ;
 wire \dp.rf.rf[29][31] ;
 wire \dp.rf.rf[29][3] ;
 wire \dp.rf.rf[29][4] ;
 wire \dp.rf.rf[29][5] ;
 wire \dp.rf.rf[29][6] ;
 wire \dp.rf.rf[29][7] ;
 wire \dp.rf.rf[29][8] ;
 wire \dp.rf.rf[29][9] ;
 wire \dp.rf.rf[2][0] ;
 wire \dp.rf.rf[2][10] ;
 wire \dp.rf.rf[2][11] ;
 wire \dp.rf.rf[2][12] ;
 wire \dp.rf.rf[2][13] ;
 wire \dp.rf.rf[2][14] ;
 wire \dp.rf.rf[2][15] ;
 wire \dp.rf.rf[2][16] ;
 wire \dp.rf.rf[2][17] ;
 wire \dp.rf.rf[2][18] ;
 wire \dp.rf.rf[2][19] ;
 wire \dp.rf.rf[2][1] ;
 wire \dp.rf.rf[2][20] ;
 wire \dp.rf.rf[2][21] ;
 wire \dp.rf.rf[2][22] ;
 wire \dp.rf.rf[2][23] ;
 wire \dp.rf.rf[2][24] ;
 wire \dp.rf.rf[2][25] ;
 wire \dp.rf.rf[2][26] ;
 wire \dp.rf.rf[2][27] ;
 wire \dp.rf.rf[2][28] ;
 wire \dp.rf.rf[2][29] ;
 wire \dp.rf.rf[2][2] ;
 wire \dp.rf.rf[2][30] ;
 wire \dp.rf.rf[2][31] ;
 wire \dp.rf.rf[2][3] ;
 wire \dp.rf.rf[2][4] ;
 wire \dp.rf.rf[2][5] ;
 wire \dp.rf.rf[2][6] ;
 wire \dp.rf.rf[2][7] ;
 wire \dp.rf.rf[2][8] ;
 wire \dp.rf.rf[2][9] ;
 wire \dp.rf.rf[30][0] ;
 wire \dp.rf.rf[30][10] ;
 wire \dp.rf.rf[30][11] ;
 wire \dp.rf.rf[30][12] ;
 wire \dp.rf.rf[30][13] ;
 wire \dp.rf.rf[30][14] ;
 wire \dp.rf.rf[30][15] ;
 wire \dp.rf.rf[30][16] ;
 wire \dp.rf.rf[30][17] ;
 wire \dp.rf.rf[30][18] ;
 wire \dp.rf.rf[30][19] ;
 wire \dp.rf.rf[30][1] ;
 wire \dp.rf.rf[30][20] ;
 wire \dp.rf.rf[30][21] ;
 wire \dp.rf.rf[30][22] ;
 wire \dp.rf.rf[30][23] ;
 wire \dp.rf.rf[30][24] ;
 wire \dp.rf.rf[30][25] ;
 wire \dp.rf.rf[30][26] ;
 wire \dp.rf.rf[30][27] ;
 wire \dp.rf.rf[30][28] ;
 wire \dp.rf.rf[30][29] ;
 wire \dp.rf.rf[30][2] ;
 wire \dp.rf.rf[30][30] ;
 wire \dp.rf.rf[30][31] ;
 wire \dp.rf.rf[30][3] ;
 wire \dp.rf.rf[30][4] ;
 wire \dp.rf.rf[30][5] ;
 wire \dp.rf.rf[30][6] ;
 wire \dp.rf.rf[30][7] ;
 wire \dp.rf.rf[30][8] ;
 wire \dp.rf.rf[30][9] ;
 wire \dp.rf.rf[31][0] ;
 wire \dp.rf.rf[31][10] ;
 wire \dp.rf.rf[31][11] ;
 wire \dp.rf.rf[31][12] ;
 wire \dp.rf.rf[31][13] ;
 wire \dp.rf.rf[31][14] ;
 wire \dp.rf.rf[31][15] ;
 wire \dp.rf.rf[31][16] ;
 wire \dp.rf.rf[31][17] ;
 wire \dp.rf.rf[31][18] ;
 wire \dp.rf.rf[31][19] ;
 wire \dp.rf.rf[31][1] ;
 wire \dp.rf.rf[31][20] ;
 wire \dp.rf.rf[31][21] ;
 wire \dp.rf.rf[31][22] ;
 wire \dp.rf.rf[31][23] ;
 wire \dp.rf.rf[31][24] ;
 wire \dp.rf.rf[31][25] ;
 wire \dp.rf.rf[31][26] ;
 wire \dp.rf.rf[31][27] ;
 wire \dp.rf.rf[31][28] ;
 wire \dp.rf.rf[31][29] ;
 wire \dp.rf.rf[31][2] ;
 wire \dp.rf.rf[31][30] ;
 wire \dp.rf.rf[31][31] ;
 wire \dp.rf.rf[31][3] ;
 wire \dp.rf.rf[31][4] ;
 wire \dp.rf.rf[31][5] ;
 wire \dp.rf.rf[31][6] ;
 wire \dp.rf.rf[31][7] ;
 wire \dp.rf.rf[31][8] ;
 wire \dp.rf.rf[31][9] ;
 wire \dp.rf.rf[3][0] ;
 wire \dp.rf.rf[3][10] ;
 wire \dp.rf.rf[3][11] ;
 wire \dp.rf.rf[3][12] ;
 wire \dp.rf.rf[3][13] ;
 wire \dp.rf.rf[3][14] ;
 wire \dp.rf.rf[3][15] ;
 wire \dp.rf.rf[3][16] ;
 wire \dp.rf.rf[3][17] ;
 wire \dp.rf.rf[3][18] ;
 wire \dp.rf.rf[3][19] ;
 wire \dp.rf.rf[3][1] ;
 wire \dp.rf.rf[3][20] ;
 wire \dp.rf.rf[3][21] ;
 wire \dp.rf.rf[3][22] ;
 wire \dp.rf.rf[3][23] ;
 wire \dp.rf.rf[3][24] ;
 wire \dp.rf.rf[3][25] ;
 wire \dp.rf.rf[3][26] ;
 wire \dp.rf.rf[3][27] ;
 wire \dp.rf.rf[3][28] ;
 wire \dp.rf.rf[3][29] ;
 wire \dp.rf.rf[3][2] ;
 wire \dp.rf.rf[3][30] ;
 wire \dp.rf.rf[3][31] ;
 wire \dp.rf.rf[3][3] ;
 wire \dp.rf.rf[3][4] ;
 wire \dp.rf.rf[3][5] ;
 wire \dp.rf.rf[3][6] ;
 wire \dp.rf.rf[3][7] ;
 wire \dp.rf.rf[3][8] ;
 wire \dp.rf.rf[3][9] ;
 wire \dp.rf.rf[4][0] ;
 wire \dp.rf.rf[4][10] ;
 wire \dp.rf.rf[4][11] ;
 wire \dp.rf.rf[4][12] ;
 wire \dp.rf.rf[4][13] ;
 wire \dp.rf.rf[4][14] ;
 wire \dp.rf.rf[4][15] ;
 wire \dp.rf.rf[4][16] ;
 wire \dp.rf.rf[4][17] ;
 wire \dp.rf.rf[4][18] ;
 wire \dp.rf.rf[4][19] ;
 wire \dp.rf.rf[4][1] ;
 wire \dp.rf.rf[4][20] ;
 wire \dp.rf.rf[4][21] ;
 wire \dp.rf.rf[4][22] ;
 wire \dp.rf.rf[4][23] ;
 wire \dp.rf.rf[4][24] ;
 wire \dp.rf.rf[4][25] ;
 wire \dp.rf.rf[4][26] ;
 wire \dp.rf.rf[4][27] ;
 wire \dp.rf.rf[4][28] ;
 wire \dp.rf.rf[4][29] ;
 wire \dp.rf.rf[4][2] ;
 wire \dp.rf.rf[4][30] ;
 wire \dp.rf.rf[4][31] ;
 wire \dp.rf.rf[4][3] ;
 wire \dp.rf.rf[4][4] ;
 wire \dp.rf.rf[4][5] ;
 wire \dp.rf.rf[4][6] ;
 wire \dp.rf.rf[4][7] ;
 wire \dp.rf.rf[4][8] ;
 wire \dp.rf.rf[4][9] ;
 wire \dp.rf.rf[5][0] ;
 wire \dp.rf.rf[5][10] ;
 wire \dp.rf.rf[5][11] ;
 wire \dp.rf.rf[5][12] ;
 wire \dp.rf.rf[5][13] ;
 wire \dp.rf.rf[5][14] ;
 wire \dp.rf.rf[5][15] ;
 wire \dp.rf.rf[5][16] ;
 wire \dp.rf.rf[5][17] ;
 wire \dp.rf.rf[5][18] ;
 wire \dp.rf.rf[5][19] ;
 wire \dp.rf.rf[5][1] ;
 wire \dp.rf.rf[5][20] ;
 wire \dp.rf.rf[5][21] ;
 wire \dp.rf.rf[5][22] ;
 wire \dp.rf.rf[5][23] ;
 wire \dp.rf.rf[5][24] ;
 wire \dp.rf.rf[5][25] ;
 wire \dp.rf.rf[5][26] ;
 wire \dp.rf.rf[5][27] ;
 wire \dp.rf.rf[5][28] ;
 wire \dp.rf.rf[5][29] ;
 wire \dp.rf.rf[5][2] ;
 wire \dp.rf.rf[5][30] ;
 wire \dp.rf.rf[5][31] ;
 wire \dp.rf.rf[5][3] ;
 wire \dp.rf.rf[5][4] ;
 wire \dp.rf.rf[5][5] ;
 wire \dp.rf.rf[5][6] ;
 wire \dp.rf.rf[5][7] ;
 wire \dp.rf.rf[5][8] ;
 wire \dp.rf.rf[5][9] ;
 wire \dp.rf.rf[6][0] ;
 wire \dp.rf.rf[6][10] ;
 wire \dp.rf.rf[6][11] ;
 wire \dp.rf.rf[6][12] ;
 wire \dp.rf.rf[6][13] ;
 wire \dp.rf.rf[6][14] ;
 wire \dp.rf.rf[6][15] ;
 wire \dp.rf.rf[6][16] ;
 wire \dp.rf.rf[6][17] ;
 wire \dp.rf.rf[6][18] ;
 wire \dp.rf.rf[6][19] ;
 wire \dp.rf.rf[6][1] ;
 wire \dp.rf.rf[6][20] ;
 wire \dp.rf.rf[6][21] ;
 wire \dp.rf.rf[6][22] ;
 wire \dp.rf.rf[6][23] ;
 wire \dp.rf.rf[6][24] ;
 wire \dp.rf.rf[6][25] ;
 wire \dp.rf.rf[6][26] ;
 wire \dp.rf.rf[6][27] ;
 wire \dp.rf.rf[6][28] ;
 wire \dp.rf.rf[6][29] ;
 wire \dp.rf.rf[6][2] ;
 wire \dp.rf.rf[6][30] ;
 wire \dp.rf.rf[6][31] ;
 wire \dp.rf.rf[6][3] ;
 wire \dp.rf.rf[6][4] ;
 wire \dp.rf.rf[6][5] ;
 wire \dp.rf.rf[6][6] ;
 wire \dp.rf.rf[6][7] ;
 wire \dp.rf.rf[6][8] ;
 wire \dp.rf.rf[6][9] ;
 wire \dp.rf.rf[7][0] ;
 wire \dp.rf.rf[7][10] ;
 wire \dp.rf.rf[7][11] ;
 wire \dp.rf.rf[7][12] ;
 wire \dp.rf.rf[7][13] ;
 wire \dp.rf.rf[7][14] ;
 wire \dp.rf.rf[7][15] ;
 wire \dp.rf.rf[7][16] ;
 wire \dp.rf.rf[7][17] ;
 wire \dp.rf.rf[7][18] ;
 wire \dp.rf.rf[7][19] ;
 wire \dp.rf.rf[7][1] ;
 wire \dp.rf.rf[7][20] ;
 wire \dp.rf.rf[7][21] ;
 wire \dp.rf.rf[7][22] ;
 wire \dp.rf.rf[7][23] ;
 wire \dp.rf.rf[7][24] ;
 wire \dp.rf.rf[7][25] ;
 wire \dp.rf.rf[7][26] ;
 wire \dp.rf.rf[7][27] ;
 wire \dp.rf.rf[7][28] ;
 wire \dp.rf.rf[7][29] ;
 wire \dp.rf.rf[7][2] ;
 wire \dp.rf.rf[7][30] ;
 wire \dp.rf.rf[7][31] ;
 wire \dp.rf.rf[7][3] ;
 wire \dp.rf.rf[7][4] ;
 wire \dp.rf.rf[7][5] ;
 wire \dp.rf.rf[7][6] ;
 wire \dp.rf.rf[7][7] ;
 wire \dp.rf.rf[7][8] ;
 wire \dp.rf.rf[7][9] ;
 wire \dp.rf.rf[8][0] ;
 wire \dp.rf.rf[8][10] ;
 wire \dp.rf.rf[8][11] ;
 wire \dp.rf.rf[8][12] ;
 wire \dp.rf.rf[8][13] ;
 wire \dp.rf.rf[8][14] ;
 wire \dp.rf.rf[8][15] ;
 wire \dp.rf.rf[8][16] ;
 wire \dp.rf.rf[8][17] ;
 wire \dp.rf.rf[8][18] ;
 wire \dp.rf.rf[8][19] ;
 wire \dp.rf.rf[8][1] ;
 wire \dp.rf.rf[8][20] ;
 wire \dp.rf.rf[8][21] ;
 wire \dp.rf.rf[8][22] ;
 wire \dp.rf.rf[8][23] ;
 wire \dp.rf.rf[8][24] ;
 wire \dp.rf.rf[8][25] ;
 wire \dp.rf.rf[8][26] ;
 wire \dp.rf.rf[8][27] ;
 wire \dp.rf.rf[8][28] ;
 wire \dp.rf.rf[8][29] ;
 wire \dp.rf.rf[8][2] ;
 wire \dp.rf.rf[8][30] ;
 wire \dp.rf.rf[8][31] ;
 wire \dp.rf.rf[8][3] ;
 wire \dp.rf.rf[8][4] ;
 wire \dp.rf.rf[8][5] ;
 wire \dp.rf.rf[8][6] ;
 wire \dp.rf.rf[8][7] ;
 wire \dp.rf.rf[8][8] ;
 wire \dp.rf.rf[8][9] ;
 wire \dp.rf.rf[9][0] ;
 wire \dp.rf.rf[9][10] ;
 wire \dp.rf.rf[9][11] ;
 wire \dp.rf.rf[9][12] ;
 wire \dp.rf.rf[9][13] ;
 wire \dp.rf.rf[9][14] ;
 wire \dp.rf.rf[9][15] ;
 wire \dp.rf.rf[9][16] ;
 wire \dp.rf.rf[9][17] ;
 wire \dp.rf.rf[9][18] ;
 wire \dp.rf.rf[9][19] ;
 wire \dp.rf.rf[9][1] ;
 wire \dp.rf.rf[9][20] ;
 wire \dp.rf.rf[9][21] ;
 wire \dp.rf.rf[9][22] ;
 wire \dp.rf.rf[9][23] ;
 wire \dp.rf.rf[9][24] ;
 wire \dp.rf.rf[9][25] ;
 wire \dp.rf.rf[9][26] ;
 wire \dp.rf.rf[9][27] ;
 wire \dp.rf.rf[9][28] ;
 wire \dp.rf.rf[9][29] ;
 wire \dp.rf.rf[9][2] ;
 wire \dp.rf.rf[9][30] ;
 wire \dp.rf.rf[9][31] ;
 wire \dp.rf.rf[9][3] ;
 wire \dp.rf.rf[9][4] ;
 wire \dp.rf.rf[9][5] ;
 wire \dp.rf.rf[9][6] ;
 wire \dp.rf.rf[9][7] ;
 wire \dp.rf.rf[9][8] ;
 wire \dp.rf.rf[9][9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net165;
 wire net166;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net222;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net237;
 wire net238;
 wire net251;
 wire net252;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net234;
 wire net235;
 wire net236;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;

 gf180mcu_fd_sc_mcu9t5v0__clkinv_16 _05201_ (.I(net22),
    .ZN(_01027_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05202_ (.I(_01027_),
    .Z(_01028_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _05203_ (.I(net23),
    .Z(_01029_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05204_ (.A1(_01028_),
    .A2(_01029_),
    .Z(_01030_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05205_ (.I(net24),
    .ZN(_01031_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05206_ (.A1(net10),
    .A2(net1),
    .Z(_01032_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05207_ (.I(instr[2]),
    .Z(_01033_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _05208_ (.I(_01033_),
    .Z(_01034_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _05209_ (.A1(net21),
    .A2(_01034_),
    .ZN(_01035_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _05210_ (.A1(_01031_),
    .A2(net230),
    .A3(_01035_),
    .Z(_01036_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05211_ (.A1(_01030_),
    .A2(_01036_),
    .Z(net94));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05212_ (.I(net13),
    .Z(_01037_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05213_ (.I(instr[20]),
    .Z(_01038_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _05214_ (.I(instr[21]),
    .Z(_01039_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05215_ (.I0(\dp.rf.rf[24][0] ),
    .I1(\dp.rf.rf[25][0] ),
    .I2(\dp.rf.rf[26][0] ),
    .I3(\dp.rf.rf[27][0] ),
    .S0(_01038_),
    .S1(_01039_),
    .Z(_01040_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05216_ (.I0(\dp.rf.rf[16][0] ),
    .I1(\dp.rf.rf[17][0] ),
    .I2(\dp.rf.rf[18][0] ),
    .I3(\dp.rf.rf[19][0] ),
    .S0(_01038_),
    .S1(_01039_),
    .Z(_01041_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _05217_ (.I(net12),
    .ZN(_01042_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05218_ (.I0(_01040_),
    .I1(_01041_),
    .S(_01042_),
    .Z(_01043_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05219_ (.I0(\dp.rf.rf[28][0] ),
    .I1(\dp.rf.rf[29][0] ),
    .I2(\dp.rf.rf[30][0] ),
    .I3(\dp.rf.rf[31][0] ),
    .S0(_01038_),
    .S1(_01039_),
    .Z(_01044_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05220_ (.I0(\dp.rf.rf[20][0] ),
    .I1(\dp.rf.rf[21][0] ),
    .I2(\dp.rf.rf[22][0] ),
    .I3(\dp.rf.rf[23][0] ),
    .S0(_01038_),
    .S1(_01039_),
    .Z(_01045_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05221_ (.I0(_01044_),
    .I1(_01045_),
    .S(_01042_),
    .Z(_01046_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05222_ (.I(net11),
    .Z(_01047_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _05223_ (.I0(_01043_),
    .I1(_01046_),
    .S(net196),
    .Z(_01048_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 _05224_ (.I(instr[20]),
    .Z(_01049_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05225_ (.I0(\dp.rf.rf[8][0] ),
    .I1(\dp.rf.rf[9][0] ),
    .I2(\dp.rf.rf[10][0] ),
    .I3(\dp.rf.rf[11][0] ),
    .S0(net264),
    .S1(_01039_),
    .Z(_01050_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05226_ (.I0(\dp.rf.rf[0][0] ),
    .I1(\dp.rf.rf[1][0] ),
    .I2(\dp.rf.rf[2][0] ),
    .I3(\dp.rf.rf[3][0] ),
    .S0(net264),
    .S1(_01039_),
    .Z(_01051_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05227_ (.I0(_01050_),
    .I1(_01051_),
    .S(_01042_),
    .Z(_01052_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05228_ (.I0(\dp.rf.rf[12][0] ),
    .I1(\dp.rf.rf[13][0] ),
    .I2(\dp.rf.rf[14][0] ),
    .I3(\dp.rf.rf[15][0] ),
    .S0(net264),
    .S1(_01039_),
    .Z(_01053_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05229_ (.I0(\dp.rf.rf[4][0] ),
    .I1(\dp.rf.rf[5][0] ),
    .I2(\dp.rf.rf[6][0] ),
    .I3(\dp.rf.rf[7][0] ),
    .S0(net264),
    .S1(_01039_),
    .Z(_01054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05230_ (.I0(_01053_),
    .I1(_01054_),
    .S(_01042_),
    .Z(_01055_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _05231_ (.I0(_01052_),
    .I1(_01055_),
    .S(net196),
    .Z(_01056_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _05232_ (.I(net13),
    .ZN(_01057_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05233_ (.I(_01057_),
    .Z(_01058_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05234_ (.I(instr[20]),
    .Z(_01059_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _05235_ (.A1(_01047_),
    .A2(_01059_),
    .A3(_01039_),
    .A4(net12),
    .Z(_01060_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05236_ (.A1(_01058_),
    .A2(_01060_),
    .Z(_01061_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _05237_ (.A1(_01037_),
    .A2(_01048_),
    .B1(_01056_),
    .B2(_01061_),
    .ZN(_01062_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05238_ (.I(net270),
    .ZN(net128));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _05239_ (.A1(net10),
    .A2(net1),
    .ZN(_01063_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _05240_ (.A1(net21),
    .A2(_01033_),
    .Z(_01064_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _05241_ (.A1(net24),
    .A2(_01063_),
    .A3(_01064_),
    .Z(_01065_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05242_ (.A1(_01029_),
    .A2(net19),
    .ZN(_01066_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _05243_ (.I(net4),
    .ZN(_01067_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _05244_ (.I(net5),
    .ZN(_01068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _05245_ (.A1(_01067_),
    .A2(_01068_),
    .ZN(_01069_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05246_ (.A1(net5),
    .A2(_01066_),
    .ZN(_01070_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _05247_ (.A1(_01065_),
    .A2(_01066_),
    .A3(_01069_),
    .B(_01070_),
    .ZN(_01071_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _05248_ (.A1(net5),
    .A2(_01065_),
    .B1(_01071_),
    .B2(net22),
    .ZN(_01072_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _05249_ (.A1(net21),
    .A2(net24),
    .Z(_01073_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 split62 (.I(_03041_),
    .Z(net221));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _05251_ (.A1(net1),
    .A2(_01033_),
    .A3(net10),
    .ZN(_01075_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _05252_ (.A1(_01073_),
    .A2(_01027_),
    .A3(_01075_),
    .Z(_01076_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 _05253_ (.I(_01076_),
    .Z(_01077_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 _05254_ (.I(_01077_),
    .Z(_01078_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05255_ (.A1(net230),
    .A2(_01035_),
    .Z(_01079_));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer102 (.I(_02427_),
    .Z(net275));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05257_ (.A1(_01029_),
    .A2(net24),
    .Z(_01081_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05258_ (.A1(_01028_),
    .A2(_01081_),
    .Z(_01082_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _05259_ (.A1(_01079_),
    .A2(_01082_),
    .ZN(_01083_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05260_ (.A1(_01078_),
    .A2(_01083_),
    .ZN(_01084_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _05261_ (.A1(_01084_),
    .A2(_01072_),
    .A3(net6),
    .Z(_01085_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _05262_ (.I(_01085_),
    .Z(_01086_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05263_ (.I0(net24),
    .I1(net22),
    .S(_01029_),
    .Z(_01087_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05264_ (.A1(net23),
    .A2(net24),
    .ZN(_01088_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05265_ (.I0(_01073_),
    .I1(_01088_),
    .S(_01027_),
    .Z(_01089_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _05266_ (.I(_01033_),
    .Z(_01090_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05267_ (.I(_01090_),
    .ZN(_01091_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _05268_ (.A1(_01064_),
    .A2(_01087_),
    .B1(_01089_),
    .B2(_01091_),
    .ZN(_01092_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05269_ (.A1(net232),
    .A2(_01092_),
    .Z(_01093_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _05270_ (.A1(net10),
    .A2(net1),
    .A3(net21),
    .A4(_01033_),
    .ZN(_01094_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _05271_ (.A1(_01063_),
    .A2(_01064_),
    .B1(_01094_),
    .B2(_01031_),
    .ZN(_01095_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _05272_ (.A1(net21),
    .A2(net24),
    .ZN(_01096_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _05273_ (.A1(_01032_),
    .A2(net22),
    .A3(_01033_),
    .A4(_01096_),
    .Z(_01097_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05274_ (.I(_01049_),
    .Z(_01098_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _05275_ (.I(_01098_),
    .ZN(_01099_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _05276_ (.A1(_01030_),
    .A2(_01095_),
    .B(_01097_),
    .C(_01099_),
    .ZN(_01100_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _05277_ (.I(net26),
    .ZN(_01101_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05278_ (.I(instr[21]),
    .Z(_01102_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _05279_ (.I(_01102_),
    .ZN(_01103_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _05280_ (.A1(_01101_),
    .A2(_01063_),
    .A3(_01064_),
    .B1(_01094_),
    .B2(_01103_),
    .ZN(_01104_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05281_ (.A1(_01082_),
    .A2(_01104_),
    .Z(_01105_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _05282_ (.A1(net25),
    .A2(_01030_),
    .A3(_01036_),
    .Z(_01106_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _05283_ (.A1(net22),
    .A2(_01063_),
    .A3(_01088_),
    .Z(_01107_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _05284_ (.A1(net21),
    .A2(_01033_),
    .Z(_01108_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _05285_ (.A1(_01107_),
    .A2(_01108_),
    .Z(_01109_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _05286_ (.A1(_01100_),
    .A2(_01105_),
    .A3(_01106_),
    .B(_01109_),
    .ZN(_01110_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05287_ (.I(_01037_),
    .Z(_01111_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 _05288_ (.I(_01061_),
    .Z(_01112_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_4 _05289_ (.A1(_01111_),
    .A2(net212),
    .B1(net197),
    .B2(_01112_),
    .C1(_01092_),
    .C2(_01032_),
    .ZN(_01113_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _05290_ (.A1(_01093_),
    .A2(_01110_),
    .B(_01113_),
    .ZN(_01114_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _05291_ (.I(_01114_),
    .Z(_01115_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _05292_ (.I(_01115_),
    .Z(_01116_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _05293_ (.A1(_01086_),
    .A2(_01116_),
    .ZN(_04825_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05294_ (.I(_04825_),
    .ZN(_04829_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05295_ (.I(net7),
    .Z(_01117_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05296_ (.I(_01117_),
    .Z(_01118_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05297_ (.I(_01118_),
    .Z(_01119_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 _05298_ (.I(instr[15]),
    .Z(_01120_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05299_ (.I(_01120_),
    .Z(_01121_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05300_ (.I(instr[17]),
    .Z(_01122_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05301_ (.I(_01122_),
    .Z(_01123_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05302_ (.I(_01123_),
    .Z(_01124_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05303_ (.I0(\dp.rf.rf[2][0] ),
    .I1(\dp.rf.rf[3][0] ),
    .I2(\dp.rf.rf[6][0] ),
    .I3(\dp.rf.rf[7][0] ),
    .S0(_01121_),
    .S1(_01124_),
    .Z(_01125_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05304_ (.A1(_01119_),
    .A2(_01125_),
    .Z(_01126_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05305_ (.I(instr[15]),
    .Z(_01127_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05306_ (.I(_01127_),
    .Z(_01128_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05307_ (.I(_01122_),
    .Z(_01129_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _05308_ (.A1(_01128_),
    .A2(_01129_),
    .ZN(_01130_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _05309_ (.I(net8),
    .ZN(_01131_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _05310_ (.A1(_01117_),
    .A2(_01130_),
    .B(_01131_),
    .ZN(_01132_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _05311_ (.I(net7),
    .ZN(_01133_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05312_ (.A1(_01133_),
    .A2(_01131_),
    .ZN(_01134_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05313_ (.I(_01127_),
    .Z(_01135_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05314_ (.I(_01135_),
    .Z(_01136_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05315_ (.I(_01122_),
    .Z(_01137_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05316_ (.I(_01137_),
    .Z(_01138_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05317_ (.I(_01138_),
    .Z(_01139_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _05318_ (.I0(\dp.rf.rf[0][0] ),
    .I1(\dp.rf.rf[1][0] ),
    .I2(\dp.rf.rf[4][0] ),
    .I3(\dp.rf.rf[5][0] ),
    .S0(_01136_),
    .S1(_01139_),
    .Z(_01140_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _05319_ (.I(net9),
    .ZN(_01141_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05320_ (.A1(_01141_),
    .A2(net186),
    .Z(_01142_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _05321_ (.A1(_01126_),
    .A2(_01132_),
    .B1(_01134_),
    .B2(_01140_),
    .C(_01142_),
    .ZN(_01143_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05322_ (.I(_01137_),
    .Z(_01144_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05323_ (.I(_01144_),
    .Z(_01145_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05324_ (.I(_01145_),
    .Z(_01146_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05325_ (.I(_01120_),
    .Z(_01147_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05326_ (.I0(\dp.rf.rf[14][0] ),
    .I1(\dp.rf.rf[15][0] ),
    .S(_01147_),
    .Z(_01148_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05327_ (.I(_01148_),
    .ZN(_01149_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _05328_ (.A1(net180),
    .A2(_01027_),
    .A3(net216),
    .B(net7),
    .ZN(_01150_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05329_ (.I(_01150_),
    .Z(_01151_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05330_ (.A1(_01146_),
    .A2(_01149_),
    .B(_01151_),
    .ZN(_01152_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _05331_ (.I(_01073_),
    .Z(_01153_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _05332_ (.I(net10),
    .Z(_01154_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _05333_ (.I(net1),
    .Z(_01155_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _05334_ (.A1(\dp.rf.rf[10][0] ),
    .A2(_01154_),
    .A3(_01155_),
    .A4(_01034_),
    .ZN(_01156_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05335_ (.I(_01135_),
    .Z(_01157_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05336_ (.I(\dp.rf.rf[10][0] ),
    .ZN(_01158_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _05337_ (.A1(_01028_),
    .A2(_01153_),
    .A3(_01156_),
    .B1(_01157_),
    .B2(_01158_),
    .ZN(_01159_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05338_ (.I(_01128_),
    .Z(_01160_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05339_ (.A1(\dp.rf.rf[11][0] ),
    .A2(_01160_),
    .Z(_01161_));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 _05340_ (.I(_01122_),
    .ZN(_01162_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _05341_ (.A1(net22),
    .A2(_01096_),
    .B(_01162_),
    .ZN(_01163_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _05342_ (.I(_01163_),
    .Z(_01164_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05343_ (.A1(_01137_),
    .A2(_01075_),
    .Z(_01165_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _05344_ (.I(_01165_),
    .Z(_01166_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _05345_ (.A1(_01159_),
    .A2(_01161_),
    .A3(_01164_),
    .A4(_01166_),
    .Z(_01167_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05346_ (.I(_01137_),
    .Z(_01168_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05347_ (.I(_01168_),
    .Z(_01169_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _05348_ (.I0(\dp.rf.rf[8][0] ),
    .I1(\dp.rf.rf[9][0] ),
    .I2(\dp.rf.rf[12][0] ),
    .I3(\dp.rf.rf[13][0] ),
    .S0(_01136_),
    .S1(_01169_),
    .Z(_01170_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05349_ (.I(_01133_),
    .Z(_01171_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05350_ (.I(_01171_),
    .Z(_01172_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05351_ (.I(_01172_),
    .Z(_01173_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05352_ (.I(_01075_),
    .Z(_01174_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _05353_ (.A1(_01027_),
    .A2(net167),
    .A3(_01174_),
    .B(net8),
    .ZN(_01175_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05354_ (.I(_01175_),
    .Z(_01176_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _05355_ (.A1(_01152_),
    .A2(_01167_),
    .B1(_01170_),
    .B2(_01173_),
    .C(_01176_),
    .ZN(_01177_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05356_ (.I(net8),
    .Z(_01178_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05357_ (.I(_01127_),
    .Z(_01179_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05358_ (.I0(\dp.rf.rf[20][0] ),
    .I1(\dp.rf.rf[21][0] ),
    .I2(\dp.rf.rf[22][0] ),
    .I3(\dp.rf.rf[23][0] ),
    .S0(_01179_),
    .S1(_01117_),
    .Z(_01180_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05359_ (.I0(\dp.rf.rf[16][0] ),
    .I1(\dp.rf.rf[17][0] ),
    .I2(\dp.rf.rf[18][0] ),
    .I3(\dp.rf.rf[19][0] ),
    .S0(_01179_),
    .S1(_01117_),
    .Z(_01181_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05360_ (.I(_01162_),
    .Z(_01182_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05361_ (.I0(_01180_),
    .I1(_01181_),
    .S(_01182_),
    .Z(_01183_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05362_ (.I(\dp.rf.rf[24][0] ),
    .ZN(_01184_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05363_ (.I(net180),
    .Z(_01185_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05364_ (.I(_01127_),
    .Z(_01186_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _05365_ (.A1(_01186_),
    .A2(_01117_),
    .Z(_01187_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _05366_ (.A1(_01028_),
    .A2(_01185_),
    .A3(_01174_),
    .B(_01187_),
    .ZN(_01188_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _05367_ (.I(_01127_),
    .ZN(_01189_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05368_ (.I(_01189_),
    .Z(_01190_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _05369_ (.A1(\dp.rf.rf[25][0] ),
    .A2(_01190_),
    .A3(_01118_),
    .ZN(_01191_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05370_ (.I(net161),
    .Z(_01192_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05371_ (.I(_01133_),
    .Z(_01193_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05372_ (.I(_01127_),
    .Z(_01194_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05373_ (.I0(\dp.rf.rf[26][0] ),
    .I1(\dp.rf.rf[27][0] ),
    .S(_01194_),
    .Z(_01195_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05374_ (.I(_01162_),
    .Z(_01196_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _05375_ (.A1(_01193_),
    .A2(_01195_),
    .B(_01196_),
    .ZN(_01197_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _05376_ (.A1(_01184_),
    .A2(_01188_),
    .B1(_01191_),
    .B2(_01192_),
    .C(_01197_),
    .ZN(_01198_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05377_ (.I(_01175_),
    .Z(_01199_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05378_ (.I(_01137_),
    .Z(_01200_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05379_ (.I(_01200_),
    .Z(_01201_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05380_ (.I(_01127_),
    .Z(_01202_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05381_ (.I0(\dp.rf.rf[28][0] ),
    .I1(\dp.rf.rf[29][0] ),
    .I2(\dp.rf.rf[30][0] ),
    .I3(\dp.rf.rf[31][0] ),
    .S0(_01202_),
    .S1(_01117_),
    .Z(_01203_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05382_ (.A1(_01201_),
    .A2(_01203_),
    .Z(_01204_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _05383_ (.A1(_01199_),
    .A2(_01204_),
    .Z(_01205_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05384_ (.A1(net9),
    .A2(net161),
    .Z(_01206_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05385_ (.I(_01206_),
    .Z(_01207_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _05386_ (.A1(_01178_),
    .A2(_01183_),
    .B1(_01198_),
    .B2(_01205_),
    .C(_01207_),
    .ZN(_01208_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _05387_ (.A1(_01143_),
    .A2(_01177_),
    .B(_01208_),
    .ZN(_04824_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05388_ (.I(net169),
    .ZN(_04828_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05389_ (.I(_01129_),
    .Z(_01209_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05390_ (.I(_01209_),
    .Z(_01210_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05391_ (.I(_01210_),
    .Z(_01211_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05392_ (.I(_01186_),
    .Z(_01212_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05393_ (.I(_01117_),
    .Z(_01213_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05394_ (.I0(\dp.rf.rf[28][31] ),
    .I1(\dp.rf.rf[29][31] ),
    .I2(\dp.rf.rf[30][31] ),
    .I3(\dp.rf.rf[31][31] ),
    .S0(_01212_),
    .S1(_01213_),
    .Z(_01214_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05395_ (.I(\dp.rf.rf[24][31] ),
    .ZN(_01215_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05396_ (.I(\dp.rf.rf[25][31] ),
    .ZN(_01216_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _05397_ (.A1(_01216_),
    .A2(_01160_),
    .A3(_01171_),
    .Z(_01217_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05398_ (.I(_01133_),
    .Z(_01218_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05399_ (.I0(\dp.rf.rf[26][31] ),
    .I1(\dp.rf.rf[27][31] ),
    .S(_01128_),
    .Z(_01219_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _05400_ (.A1(_01218_),
    .A2(_01219_),
    .B(_01196_),
    .ZN(_01220_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _05401_ (.A1(_01215_),
    .A2(_01188_),
    .B1(_01217_),
    .B2(_01192_),
    .C(_01220_),
    .ZN(_01221_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _05402_ (.A1(_01211_),
    .A2(_01214_),
    .B(_01221_),
    .C(_01176_),
    .ZN(_01222_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _05403_ (.A1(_01027_),
    .A2(net251),
    .A3(net218),
    .B(_01137_),
    .ZN(_01223_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05404_ (.I(_01223_),
    .Z(_01224_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05405_ (.I(_01120_),
    .Z(_01225_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05406_ (.I0(\dp.rf.rf[20][31] ),
    .I1(\dp.rf.rf[21][31] ),
    .I2(\dp.rf.rf[22][31] ),
    .I3(\dp.rf.rf[23][31] ),
    .S0(_01225_),
    .S1(_01118_),
    .Z(_01226_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05407_ (.I(_01226_),
    .ZN(_01227_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05408_ (.I(_01131_),
    .Z(_01228_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _05409_ (.A1(_01224_),
    .A2(_01227_),
    .B(_01228_),
    .ZN(_01229_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05410_ (.I(_01162_),
    .Z(_01230_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _05411_ (.A1(\dp.rf.rf[16][31] ),
    .A2(_01187_),
    .Z(_01231_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05412_ (.I0(\dp.rf.rf[17][31] ),
    .I1(\dp.rf.rf[19][31] ),
    .S(net7),
    .Z(_01232_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _05413_ (.A1(_01190_),
    .A2(_01232_),
    .Z(_01233_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _05414_ (.A1(\dp.rf.rf[18][31] ),
    .A2(_01160_),
    .A3(_01171_),
    .Z(_01234_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _05415_ (.A1(_01230_),
    .A2(_01231_),
    .A3(_01233_),
    .A4(_01234_),
    .Z(_01235_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _05416_ (.A1(_01229_),
    .A2(_01235_),
    .B(net177),
    .ZN(_01236_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05417_ (.I(_01175_),
    .Z(_01237_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05418_ (.I(_01127_),
    .Z(_01238_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05419_ (.I0(\dp.rf.rf[10][31] ),
    .I1(\dp.rf.rf[11][31] ),
    .I2(\dp.rf.rf[14][31] ),
    .I3(\dp.rf.rf[15][31] ),
    .S0(_01238_),
    .S1(_01209_),
    .Z(_01239_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05420_ (.I0(\dp.rf.rf[8][31] ),
    .I1(\dp.rf.rf[9][31] ),
    .I2(\dp.rf.rf[12][31] ),
    .I3(\dp.rf.rf[13][31] ),
    .S0(_01238_),
    .S1(_01209_),
    .Z(_01240_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05421_ (.I(_01133_),
    .Z(_01241_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05422_ (.I0(_01239_),
    .I1(_01240_),
    .S(_01241_),
    .Z(_01242_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05423_ (.A1(_01237_),
    .A2(_01242_),
    .ZN(_01243_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05424_ (.I(net9),
    .Z(_01244_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05425_ (.I(_01097_),
    .Z(_01245_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05426_ (.I0(\dp.rf.rf[2][31] ),
    .I1(\dp.rf.rf[3][31] ),
    .I2(\dp.rf.rf[6][31] ),
    .I3(\dp.rf.rf[7][31] ),
    .S0(_01194_),
    .S1(_01138_),
    .Z(_01246_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05427_ (.A1(_01213_),
    .A2(_01246_),
    .B(_01132_),
    .ZN(_01247_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05428_ (.I(_01122_),
    .Z(_01248_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05429_ (.A1(_01189_),
    .A2(_01248_),
    .Z(_01249_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05430_ (.I0(\dp.rf.rf[1][31] ),
    .I1(\dp.rf.rf[5][31] ),
    .S(_01248_),
    .Z(_01250_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05431_ (.I(\dp.rf.rf[0][31] ),
    .ZN(_01251_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _05432_ (.A1(_01202_),
    .A2(_01129_),
    .Z(_01252_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05433_ (.A1(_01117_),
    .A2(net8),
    .ZN(_01253_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _05434_ (.A1(_01251_),
    .A2(_01252_),
    .B(_01253_),
    .ZN(_01254_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _05435_ (.A1(\dp.rf.rf[4][31] ),
    .A2(_01249_),
    .B1(_01250_),
    .B2(_01212_),
    .C(_01254_),
    .ZN(_01255_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _05436_ (.A1(_01244_),
    .A2(_01245_),
    .A3(_01247_),
    .A4(_01255_),
    .Z(_01256_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _05437_ (.A1(_01222_),
    .A2(_01236_),
    .B1(_01243_),
    .B2(_01256_),
    .ZN(_01257_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _05438_ (.I(_01257_),
    .Z(_01258_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _05439_ (.I(_01258_),
    .ZN(_04837_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _05440_ (.A1(net232),
    .A2(_01092_),
    .ZN(_01259_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 _05441_ (.I(net262),
    .Z(_01260_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05442_ (.I(_01260_),
    .Z(_01261_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05443_ (.I(instr[21]),
    .Z(_01262_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _05444_ (.I(_01262_),
    .Z(_01263_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05445_ (.I0(\dp.rf.rf[24][31] ),
    .I1(\dp.rf.rf[25][31] ),
    .I2(\dp.rf.rf[26][31] ),
    .I3(\dp.rf.rf[27][31] ),
    .S0(_01261_),
    .S1(_01263_),
    .Z(_01264_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05446_ (.I0(\dp.rf.rf[16][31] ),
    .I1(\dp.rf.rf[17][31] ),
    .I2(\dp.rf.rf[18][31] ),
    .I3(\dp.rf.rf[19][31] ),
    .S0(_01261_),
    .S1(_01263_),
    .Z(_01265_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 _05447_ (.I(_01049_),
    .Z(_01266_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05448_ (.I(_01266_),
    .Z(_01267_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _05449_ (.I(_01262_),
    .Z(_01268_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05450_ (.I0(\dp.rf.rf[28][31] ),
    .I1(\dp.rf.rf[29][31] ),
    .I2(\dp.rf.rf[30][31] ),
    .I3(\dp.rf.rf[31][31] ),
    .S0(_01267_),
    .S1(_01268_),
    .Z(_01269_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05451_ (.I0(\dp.rf.rf[20][31] ),
    .I1(\dp.rf.rf[21][31] ),
    .I2(\dp.rf.rf[22][31] ),
    .I3(\dp.rf.rf[23][31] ),
    .S0(_01267_),
    .S1(_01263_),
    .Z(_01270_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 _05452_ (.I(_01042_),
    .Z(_01271_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05453_ (.I(_01271_),
    .Z(_01272_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 split89 (.I(_01049_),
    .Z(net264));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _05455_ (.I0(_01264_),
    .I1(_01265_),
    .I2(_01269_),
    .I3(_01270_),
    .S0(_01272_),
    .S1(net194),
    .Z(_01274_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05456_ (.I(_01266_),
    .Z(_01275_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05457_ (.I(_01262_),
    .Z(_01276_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05458_ (.I0(\dp.rf.rf[8][31] ),
    .I1(\dp.rf.rf[9][31] ),
    .I2(\dp.rf.rf[10][31] ),
    .I3(\dp.rf.rf[11][31] ),
    .S0(_01275_),
    .S1(_01276_),
    .Z(_01277_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05459_ (.I0(\dp.rf.rf[0][31] ),
    .I1(\dp.rf.rf[1][31] ),
    .I2(\dp.rf.rf[2][31] ),
    .I3(\dp.rf.rf[3][31] ),
    .S0(_01275_),
    .S1(_01268_),
    .Z(_01278_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 _05460_ (.I(_01266_),
    .Z(_01279_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05461_ (.I0(\dp.rf.rf[12][31] ),
    .I1(\dp.rf.rf[13][31] ),
    .I2(\dp.rf.rf[14][31] ),
    .I3(\dp.rf.rf[15][31] ),
    .S0(_01279_),
    .S1(_01276_),
    .Z(_01280_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05462_ (.I0(\dp.rf.rf[4][31] ),
    .I1(\dp.rf.rf[5][31] ),
    .I2(\dp.rf.rf[6][31] ),
    .I3(\dp.rf.rf[7][31] ),
    .S0(_01275_),
    .S1(_01276_),
    .Z(_01281_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05463_ (.I(_01271_),
    .Z(_01282_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05464_ (.I0(_01277_),
    .I1(_01278_),
    .I2(_01280_),
    .I3(_01281_),
    .S0(_01282_),
    .S1(net194),
    .Z(_01283_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _05465_ (.A1(_01037_),
    .A2(_01274_),
    .B1(_01283_),
    .B2(_01061_),
    .ZN(_01284_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05466_ (.I(net20),
    .ZN(_01285_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _05467_ (.A1(_01285_),
    .A2(net233),
    .A3(_01092_),
    .Z(_01286_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05468_ (.A1(_01259_),
    .A2(_01284_),
    .B(_01286_),
    .ZN(_01287_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _05469_ (.A1(_01086_),
    .A2(_01287_),
    .ZN(_04832_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05470_ (.I(_04832_),
    .ZN(_04836_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05471_ (.I(net247),
    .Z(_01288_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05472_ (.I(_01259_),
    .Z(_01289_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _05473_ (.I(_01289_),
    .Z(_01290_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05474_ (.A1(_01030_),
    .A2(_01079_),
    .Z(_01291_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _05475_ (.A1(_01030_),
    .A2(_01095_),
    .B(_01097_),
    .ZN(_01292_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _05476_ (.A1(net20),
    .A2(_01291_),
    .B(_01292_),
    .ZN(_01293_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _05477_ (.A1(net10),
    .A2(net1),
    .A3(net21),
    .A4(_01034_),
    .Z(_01294_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05478_ (.A1(_01082_),
    .A2(_01294_),
    .Z(_01295_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05479_ (.I(_01295_),
    .Z(_01296_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05480_ (.A1(net20),
    .A2(_01296_),
    .ZN(_01297_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05481_ (.A1(_01293_),
    .A2(_01297_),
    .Z(_01298_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _05482_ (.I(_01298_),
    .Z(_01299_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _05483_ (.I(_01245_),
    .Z(_01300_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _05484_ (.I(_01300_),
    .Z(_01301_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05485_ (.A1(net19),
    .A2(_01301_),
    .ZN(_01302_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05486_ (.A1(_01285_),
    .A2(_01292_),
    .Z(_01303_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _05487_ (.I(_01303_),
    .Z(_01304_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05488_ (.A1(_01299_),
    .A2(_01302_),
    .B(_01304_),
    .ZN(_05198_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05489_ (.I(_01275_),
    .Z(_01305_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05490_ (.I(_01276_),
    .Z(_01306_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05491_ (.I0(\dp.rf.rf[24][30] ),
    .I1(\dp.rf.rf[25][30] ),
    .I2(\dp.rf.rf[26][30] ),
    .I3(\dp.rf.rf[27][30] ),
    .S0(_01305_),
    .S1(_01306_),
    .Z(_01307_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05492_ (.I0(\dp.rf.rf[16][30] ),
    .I1(\dp.rf.rf[17][30] ),
    .I2(\dp.rf.rf[18][30] ),
    .I3(\dp.rf.rf[19][30] ),
    .S0(_01305_),
    .S1(_01306_),
    .Z(_01308_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05493_ (.I0(\dp.rf.rf[28][30] ),
    .I1(\dp.rf.rf[29][30] ),
    .I2(\dp.rf.rf[30][30] ),
    .I3(\dp.rf.rf[31][30] ),
    .S0(_01305_),
    .S1(_01306_),
    .Z(_01309_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05494_ (.I0(\dp.rf.rf[20][30] ),
    .I1(\dp.rf.rf[21][30] ),
    .I2(\dp.rf.rf[22][30] ),
    .I3(\dp.rf.rf[23][30] ),
    .S0(_01305_),
    .S1(_01306_),
    .Z(_01310_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05495_ (.I(_01282_),
    .Z(_01311_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05496_ (.I(net194),
    .Z(_01312_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05497_ (.I0(_01307_),
    .I1(_01308_),
    .I2(_01309_),
    .I3(_01310_),
    .S0(_01311_),
    .S1(_01312_),
    .Z(_01313_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05498_ (.I0(\dp.rf.rf[8][30] ),
    .I1(\dp.rf.rf[9][30] ),
    .I2(\dp.rf.rf[10][30] ),
    .I3(\dp.rf.rf[11][30] ),
    .S0(_01305_),
    .S1(_01306_),
    .Z(_01314_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05499_ (.I0(\dp.rf.rf[0][30] ),
    .I1(\dp.rf.rf[1][30] ),
    .I2(\dp.rf.rf[2][30] ),
    .I3(\dp.rf.rf[3][30] ),
    .S0(_01305_),
    .S1(_01306_),
    .Z(_01315_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _05500_ (.I(_01102_),
    .Z(_01316_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05501_ (.I(_01316_),
    .Z(_01317_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05502_ (.I0(\dp.rf.rf[12][30] ),
    .I1(\dp.rf.rf[13][30] ),
    .I2(\dp.rf.rf[14][30] ),
    .I3(\dp.rf.rf[15][30] ),
    .S0(_01305_),
    .S1(_01317_),
    .Z(_01318_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05503_ (.I0(\dp.rf.rf[4][30] ),
    .I1(\dp.rf.rf[5][30] ),
    .I2(\dp.rf.rf[6][30] ),
    .I3(\dp.rf.rf[7][30] ),
    .S0(_01305_),
    .S1(_01306_),
    .Z(_01319_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05504_ (.I0(_01314_),
    .I1(_01315_),
    .I2(_01318_),
    .I3(_01319_),
    .S0(_01311_),
    .S1(_01312_),
    .Z(_01320_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _05505_ (.A1(_01111_),
    .A2(_01313_),
    .B1(_01320_),
    .B2(_01112_),
    .ZN(_01321_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05506_ (.A1(_01290_),
    .A2(_01321_),
    .ZN(_01322_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _05507_ (.A1(_01290_),
    .A2(_05198_),
    .B(_01322_),
    .ZN(_01323_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _05508_ (.A1(_01288_),
    .A2(_01323_),
    .Z(_04841_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05509_ (.I(_04841_),
    .ZN(_04845_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05510_ (.I(net160),
    .Z(_01324_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05511_ (.A1(net257),
    .A2(_01252_),
    .Z(_01325_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05512_ (.I(\dp.rf.rf[28][30] ),
    .ZN(_01326_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05513_ (.I(_01249_),
    .Z(_01327_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05514_ (.I(_01189_),
    .Z(_01328_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05515_ (.I0(\dp.rf.rf[25][30] ),
    .I1(\dp.rf.rf[29][30] ),
    .S(_01248_),
    .Z(_01329_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05516_ (.A1(_01328_),
    .A2(_01329_),
    .ZN(_01330_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _05517_ (.A1(_01326_),
    .A2(_01327_),
    .B(_01330_),
    .C(_01213_),
    .ZN(_01331_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _05518_ (.A1(\dp.rf.rf[24][30] ),
    .A2(_01325_),
    .B1(_01331_),
    .B2(_01245_),
    .ZN(_01332_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05519_ (.A1(net7),
    .A2(net186),
    .Z(_01333_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05520_ (.I(_01333_),
    .Z(_01334_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05521_ (.I(_01334_),
    .Z(_01335_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05522_ (.I0(\dp.rf.rf[26][30] ),
    .I1(\dp.rf.rf[27][30] ),
    .I2(\dp.rf.rf[30][30] ),
    .I3(\dp.rf.rf[31][30] ),
    .S0(_01136_),
    .S1(_01139_),
    .Z(_01336_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05523_ (.I(_01131_),
    .Z(_01337_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05524_ (.A1(_01335_),
    .A2(_01336_),
    .B(_01337_),
    .ZN(_01338_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05525_ (.I(_01182_),
    .Z(_01339_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05526_ (.I(_01194_),
    .Z(_01340_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05527_ (.I0(\dp.rf.rf[22][30] ),
    .I1(\dp.rf.rf[23][30] ),
    .S(_01340_),
    .Z(_01341_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _05528_ (.A1(net180),
    .A2(_01027_),
    .A3(net217),
    .B(_01120_),
    .ZN(_01342_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05529_ (.A1(\dp.rf.rf[18][30] ),
    .A2(net201),
    .Z(_01343_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05530_ (.I(_01223_),
    .Z(_01344_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05531_ (.I(_01238_),
    .Z(_01345_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05532_ (.A1(\dp.rf.rf[19][30] ),
    .A2(_01345_),
    .ZN(_01346_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05533_ (.A1(_01344_),
    .A2(_01346_),
    .ZN(_01347_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _05534_ (.A1(_01339_),
    .A2(_01341_),
    .B1(_01343_),
    .B2(_01347_),
    .C(_01334_),
    .ZN(_01348_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _05535_ (.A1(_01174_),
    .A2(net167),
    .A3(_01027_),
    .B(_01131_),
    .ZN(_01349_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05536_ (.I(\dp.rf.rf[20][30] ),
    .ZN(_01350_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05537_ (.I0(\dp.rf.rf[17][30] ),
    .I1(\dp.rf.rf[21][30] ),
    .S(_01129_),
    .Z(_01351_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05538_ (.A1(_01190_),
    .A2(_01351_),
    .ZN(_01352_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05539_ (.I(_01117_),
    .Z(_01353_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _05540_ (.A1(_01350_),
    .A2(_01249_),
    .B(_01352_),
    .C(_01353_),
    .ZN(_01354_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _05541_ (.A1(_01127_),
    .A2(_01122_),
    .A3(net8),
    .Z(_01355_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05542_ (.A1(_01324_),
    .A2(_01355_),
    .Z(_01356_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _05543_ (.A1(net234),
    .A2(_01354_),
    .B1(_01356_),
    .B2(\dp.rf.rf[16][30] ),
    .ZN(_01357_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _05544_ (.A1(_01153_),
    .A2(_01028_),
    .A3(_01174_),
    .B(net9),
    .ZN(_01358_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _05545_ (.A1(_01332_),
    .A2(_01338_),
    .B1(_01348_),
    .B2(_01357_),
    .C(net208),
    .ZN(_01359_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05546_ (.A1(_01131_),
    .A2(net161),
    .Z(_01360_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05547_ (.I(_01360_),
    .Z(_01361_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05548_ (.I(_01353_),
    .Z(_01362_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 _05549_ (.I(_01202_),
    .Z(_01363_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05550_ (.I(_01123_),
    .Z(_01364_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05551_ (.I0(\dp.rf.rf[2][30] ),
    .I1(\dp.rf.rf[3][30] ),
    .I2(\dp.rf.rf[6][30] ),
    .I3(\dp.rf.rf[7][30] ),
    .S0(_01363_),
    .S1(_01364_),
    .Z(_01365_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05552_ (.A1(_01362_),
    .A2(_01365_),
    .ZN(_01366_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _05553_ (.A1(_01189_),
    .A2(_01137_),
    .ZN(_01367_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05554_ (.I(_01367_),
    .Z(_01368_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05555_ (.I(_01137_),
    .Z(_01369_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05556_ (.I0(\dp.rf.rf[1][30] ),
    .I1(\dp.rf.rf[5][30] ),
    .S(_01369_),
    .Z(_01370_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05557_ (.I(_01189_),
    .Z(_01371_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05558_ (.I(_01171_),
    .Z(_01372_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _05559_ (.A1(\dp.rf.rf[4][30] ),
    .A2(_01368_),
    .B1(_01370_),
    .B2(_01371_),
    .C(_01372_),
    .ZN(_01373_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _05560_ (.A1(_01361_),
    .A2(_01366_),
    .A3(_01373_),
    .ZN(_01374_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _05561_ (.A1(_01130_),
    .A2(_01253_),
    .B(net9),
    .C(net198),
    .ZN(_01375_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05562_ (.I(_01375_),
    .Z(_01376_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05563_ (.I(_01252_),
    .Z(_01377_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05564_ (.A1(net168),
    .A2(_01377_),
    .B(\dp.rf.rf[8][30] ),
    .ZN(_01378_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05565_ (.I0(\dp.rf.rf[9][30] ),
    .I1(\dp.rf.rf[13][30] ),
    .S(_01168_),
    .Z(_01379_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _05566_ (.A1(\dp.rf.rf[12][30] ),
    .A2(_01368_),
    .B1(_01379_),
    .B2(_01371_),
    .C(_01172_),
    .ZN(_01380_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05567_ (.I(_01123_),
    .Z(_01381_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05568_ (.I0(\dp.rf.rf[10][30] ),
    .I1(\dp.rf.rf[11][30] ),
    .I2(\dp.rf.rf[14][30] ),
    .I3(\dp.rf.rf[15][30] ),
    .S0(_01225_),
    .S1(_01381_),
    .Z(_01382_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05569_ (.A1(_01119_),
    .A2(_01382_),
    .ZN(_01383_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05570_ (.A1(net8),
    .A2(net162),
    .Z(_01384_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05571_ (.I(_01384_),
    .Z(_01385_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _05572_ (.A1(_01378_),
    .A2(_01380_),
    .B(_01383_),
    .C(_01385_),
    .ZN(_01386_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _05573_ (.A1(_01374_),
    .A2(_01376_),
    .A3(_01386_),
    .Z(_01387_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _05574_ (.A1(_01359_),
    .A2(_01387_),
    .Z(_01388_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _05575_ (.I(_01388_),
    .ZN(_04844_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05576_ (.A1(net18),
    .A2(_01301_),
    .ZN(_01389_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05577_ (.A1(_01299_),
    .A2(_01389_),
    .B(_01304_),
    .ZN(_05194_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05578_ (.I(_01038_),
    .Z(_01390_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05579_ (.I(_01102_),
    .Z(_01391_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05580_ (.I0(\dp.rf.rf[24][29] ),
    .I1(\dp.rf.rf[25][29] ),
    .I2(\dp.rf.rf[26][29] ),
    .I3(\dp.rf.rf[27][29] ),
    .S0(_01390_),
    .S1(_01391_),
    .Z(_01392_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05581_ (.I0(\dp.rf.rf[16][29] ),
    .I1(\dp.rf.rf[17][29] ),
    .I2(\dp.rf.rf[18][29] ),
    .I3(\dp.rf.rf[19][29] ),
    .S0(_01390_),
    .S1(_01391_),
    .Z(_01393_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05582_ (.I(_01271_),
    .Z(_01394_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05583_ (.I0(_01392_),
    .I1(_01393_),
    .S(_01394_),
    .Z(_01395_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05584_ (.I0(\dp.rf.rf[28][29] ),
    .I1(\dp.rf.rf[29][29] ),
    .I2(\dp.rf.rf[30][29] ),
    .I3(\dp.rf.rf[31][29] ),
    .S0(_01390_),
    .S1(_01391_),
    .Z(_01396_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05585_ (.I0(\dp.rf.rf[20][29] ),
    .I1(\dp.rf.rf[21][29] ),
    .I2(\dp.rf.rf[22][29] ),
    .I3(\dp.rf.rf[23][29] ),
    .S0(_01390_),
    .S1(_01391_),
    .Z(_01397_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05586_ (.I(_01042_),
    .Z(_01398_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05587_ (.I0(_01396_),
    .I1(_01397_),
    .S(_01398_),
    .Z(_01399_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05588_ (.I(net194),
    .Z(_01400_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05589_ (.I0(_01395_),
    .I1(_01399_),
    .S(_01400_),
    .Z(_01401_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05590_ (.I(_01038_),
    .Z(_01402_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05591_ (.I(_01102_),
    .Z(_01403_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05592_ (.I0(\dp.rf.rf[8][29] ),
    .I1(\dp.rf.rf[9][29] ),
    .I2(\dp.rf.rf[10][29] ),
    .I3(\dp.rf.rf[11][29] ),
    .S0(_01402_),
    .S1(_01403_),
    .Z(_01404_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05593_ (.I0(\dp.rf.rf[0][29] ),
    .I1(\dp.rf.rf[1][29] ),
    .I2(\dp.rf.rf[2][29] ),
    .I3(\dp.rf.rf[3][29] ),
    .S0(_01402_),
    .S1(_01403_),
    .Z(_01405_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05594_ (.I0(_01404_),
    .I1(_01405_),
    .S(_01398_),
    .Z(_01406_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05595_ (.I0(\dp.rf.rf[12][29] ),
    .I1(\dp.rf.rf[13][29] ),
    .I2(\dp.rf.rf[14][29] ),
    .I3(\dp.rf.rf[15][29] ),
    .S0(_01402_),
    .S1(_01403_),
    .Z(_01407_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05596_ (.I(_01039_),
    .Z(_01408_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05597_ (.I0(\dp.rf.rf[4][29] ),
    .I1(\dp.rf.rf[5][29] ),
    .I2(\dp.rf.rf[6][29] ),
    .I3(\dp.rf.rf[7][29] ),
    .S0(_01402_),
    .S1(_01408_),
    .Z(_01409_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05598_ (.I0(_01407_),
    .I1(_01409_),
    .S(_01398_),
    .Z(_01410_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05599_ (.I0(_01406_),
    .I1(_01410_),
    .S(_01400_),
    .Z(_01411_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _05600_ (.A1(_01111_),
    .A2(_01401_),
    .B1(_01411_),
    .B2(_01112_),
    .ZN(_01412_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05601_ (.A1(_01290_),
    .A2(_01412_),
    .ZN(_01413_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _05602_ (.A1(_01290_),
    .A2(_05194_),
    .B(_01413_),
    .ZN(_01414_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _05603_ (.A1(_01288_),
    .A2(_01414_),
    .Z(_04849_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05604_ (.I(_04849_),
    .ZN(_04853_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05605_ (.I(_01228_),
    .Z(_01415_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05606_ (.I(_01118_),
    .Z(_01416_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _05607_ (.A1(\dp.rf.rf[10][29] ),
    .A2(_01416_),
    .B(_01377_),
    .C(\dp.rf.rf[8][29] ),
    .ZN(_01417_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _05608_ (.A1(_01415_),
    .A2(_01244_),
    .A3(_01245_),
    .A4(_01417_),
    .Z(_01418_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05609_ (.I0(\dp.rf.rf[10][29] ),
    .I1(\dp.rf.rf[11][29] ),
    .I2(\dp.rf.rf[14][29] ),
    .I3(\dp.rf.rf[15][29] ),
    .S0(_01136_),
    .S1(_01169_),
    .Z(_01419_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05610_ (.I(_01419_),
    .ZN(_01420_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05611_ (.I0(\dp.rf.rf[9][29] ),
    .I1(\dp.rf.rf[13][29] ),
    .S(_01381_),
    .Z(_01421_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05612_ (.I(_01328_),
    .Z(_01422_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _05613_ (.A1(\dp.rf.rf[12][29] ),
    .A2(_01368_),
    .B1(_01421_),
    .B2(_01422_),
    .ZN(_01423_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05614_ (.I0(_01420_),
    .I1(_01423_),
    .S(_01173_),
    .Z(_01424_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05615_ (.I0(\dp.rf.rf[25][29] ),
    .I1(\dp.rf.rf[29][29] ),
    .S(_01381_),
    .Z(_01425_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05616_ (.A1(_01422_),
    .A2(_01425_),
    .ZN(_01426_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05617_ (.I(_01127_),
    .Z(_01427_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05618_ (.I(_01427_),
    .Z(_01428_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05619_ (.I(_01428_),
    .Z(_01429_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05620_ (.I(_01171_),
    .Z(_01430_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _05621_ (.A1(\dp.rf.rf[28][29] ),
    .A2(_01429_),
    .A3(_01230_),
    .B(_01430_),
    .ZN(_01431_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05622_ (.I(_01123_),
    .Z(_01432_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05623_ (.I0(\dp.rf.rf[26][29] ),
    .I1(\dp.rf.rf[27][29] ),
    .I2(\dp.rf.rf[30][29] ),
    .I3(\dp.rf.rf[31][29] ),
    .S0(_01121_),
    .S1(_01432_),
    .Z(_01433_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05624_ (.A1(_01416_),
    .A2(_01433_),
    .ZN(_01434_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05625_ (.I(_01324_),
    .Z(_01435_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _05626_ (.A1(_01426_),
    .A2(_01431_),
    .B(_01434_),
    .C(_01435_),
    .ZN(_01436_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05627_ (.I(\dp.rf.rf[24][29] ),
    .ZN(_01437_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05628_ (.I(_01028_),
    .Z(_01438_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05629_ (.A1(\dp.rf.rf[26][29] ),
    .A2(_01118_),
    .Z(_01439_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _05630_ (.A1(_01438_),
    .A2(_01185_),
    .A3(_01174_),
    .B1(_01377_),
    .B2(_01439_),
    .ZN(_01440_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05631_ (.A1(_01437_),
    .A2(_01440_),
    .B(_01337_),
    .ZN(_01441_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05632_ (.I(_01190_),
    .Z(_01442_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05633_ (.I(_01248_),
    .Z(_01443_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05634_ (.I0(\dp.rf.rf[17][29] ),
    .I1(\dp.rf.rf[21][29] ),
    .S(_01443_),
    .Z(_01444_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05635_ (.A1(_01442_),
    .A2(_01444_),
    .ZN(_01445_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _05636_ (.A1(\dp.rf.rf[20][29] ),
    .A2(_01429_),
    .A3(_01230_),
    .B(_01430_),
    .ZN(_01446_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05637_ (.I0(\dp.rf.rf[18][29] ),
    .I1(\dp.rf.rf[19][29] ),
    .I2(\dp.rf.rf[22][29] ),
    .I3(\dp.rf.rf[23][29] ),
    .S0(_01225_),
    .S1(_01381_),
    .Z(_01447_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05638_ (.A1(_01416_),
    .A2(_01447_),
    .ZN(_01448_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _05639_ (.A1(_01445_),
    .A2(_01446_),
    .B(_01448_),
    .C(_01435_),
    .ZN(_01449_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05640_ (.I(\dp.rf.rf[16][29] ),
    .ZN(_01450_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05641_ (.A1(\dp.rf.rf[18][29] ),
    .A2(_01118_),
    .Z(_01451_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _05642_ (.A1(_01438_),
    .A2(_01185_),
    .A3(_01174_),
    .B1(_01252_),
    .B2(_01451_),
    .ZN(_01452_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05643_ (.A1(_01450_),
    .A2(_01452_),
    .B(_01178_),
    .ZN(_01453_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _05644_ (.A1(_01436_),
    .A2(_01441_),
    .B1(_01449_),
    .B2(_01453_),
    .ZN(_01454_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05645_ (.I(net207),
    .Z(_01455_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05646_ (.I(_01353_),
    .Z(_01456_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05647_ (.I(_01137_),
    .Z(_01457_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05648_ (.I(_01457_),
    .Z(_01458_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05649_ (.I0(\dp.rf.rf[2][29] ),
    .I1(\dp.rf.rf[3][29] ),
    .I2(\dp.rf.rf[6][29] ),
    .I3(\dp.rf.rf[7][29] ),
    .S0(_01345_),
    .S1(_01458_),
    .Z(_01459_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05650_ (.A1(_01456_),
    .A2(_01459_),
    .Z(_01460_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05651_ (.I(\dp.rf.rf[4][29] ),
    .ZN(_01461_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05652_ (.I0(\dp.rf.rf[1][29] ),
    .I1(\dp.rf.rf[5][29] ),
    .S(_01381_),
    .Z(_01462_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05653_ (.A1(_01422_),
    .A2(_01462_),
    .ZN(_01463_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _05654_ (.A1(_01461_),
    .A2(_01327_),
    .B(_01463_),
    .C(_01456_),
    .ZN(_01464_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05655_ (.A1(\dp.rf.rf[2][29] ),
    .A2(_01362_),
    .B(\dp.rf.rf[0][29] ),
    .ZN(_01465_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _05656_ (.A1(_01119_),
    .A2(_01377_),
    .B(_01141_),
    .ZN(_01466_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _05657_ (.A1(_01130_),
    .A2(_01465_),
    .B(_01466_),
    .C(net234),
    .ZN(_01467_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _05658_ (.A1(_01460_),
    .A2(_01464_),
    .B(_01467_),
    .ZN(_01468_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _05659_ (.A1(_01418_),
    .A2(_01424_),
    .B1(_01454_),
    .B2(_01455_),
    .C(_01468_),
    .ZN(_01469_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _05660_ (.I(_01469_),
    .Z(_04848_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05661_ (.I(_04848_),
    .ZN(_04852_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05662_ (.A1(net17),
    .A2(_01301_),
    .ZN(_01470_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05663_ (.A1(_01299_),
    .A2(_01470_),
    .B(_01304_),
    .ZN(_05190_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05664_ (.I(_01059_),
    .Z(_01471_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05665_ (.I0(\dp.rf.rf[24][28] ),
    .I1(\dp.rf.rf[25][28] ),
    .I2(\dp.rf.rf[26][28] ),
    .I3(\dp.rf.rf[27][28] ),
    .S0(_01471_),
    .S1(_01316_),
    .Z(_01472_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05666_ (.I0(\dp.rf.rf[16][28] ),
    .I1(\dp.rf.rf[17][28] ),
    .I2(\dp.rf.rf[18][28] ),
    .I3(\dp.rf.rf[19][28] ),
    .S0(_01471_),
    .S1(_01316_),
    .Z(_01473_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05667_ (.I0(_01472_),
    .I1(_01473_),
    .S(_01282_),
    .Z(_01474_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05668_ (.I0(\dp.rf.rf[28][28] ),
    .I1(\dp.rf.rf[29][28] ),
    .I2(\dp.rf.rf[30][28] ),
    .I3(\dp.rf.rf[31][28] ),
    .S0(_01471_),
    .S1(_01316_),
    .Z(_01475_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05669_ (.I0(\dp.rf.rf[20][28] ),
    .I1(\dp.rf.rf[21][28] ),
    .I2(\dp.rf.rf[22][28] ),
    .I3(\dp.rf.rf[23][28] ),
    .S0(_01471_),
    .S1(_01316_),
    .Z(_01476_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05670_ (.I0(_01475_),
    .I1(_01476_),
    .S(_01394_),
    .Z(_01477_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05671_ (.I(net194),
    .Z(_01478_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05672_ (.I0(_01474_),
    .I1(_01477_),
    .S(_01478_),
    .Z(_01479_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05673_ (.I0(\dp.rf.rf[8][28] ),
    .I1(\dp.rf.rf[9][28] ),
    .I2(\dp.rf.rf[10][28] ),
    .I3(\dp.rf.rf[11][28] ),
    .S0(_01471_),
    .S1(_01316_),
    .Z(_01480_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05674_ (.I0(\dp.rf.rf[0][28] ),
    .I1(\dp.rf.rf[1][28] ),
    .I2(\dp.rf.rf[2][28] ),
    .I3(\dp.rf.rf[3][28] ),
    .S0(_01471_),
    .S1(_01316_),
    .Z(_01481_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05675_ (.I0(_01480_),
    .I1(_01481_),
    .S(_01394_),
    .Z(_01482_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05676_ (.I0(\dp.rf.rf[12][28] ),
    .I1(\dp.rf.rf[13][28] ),
    .I2(\dp.rf.rf[14][28] ),
    .I3(\dp.rf.rf[15][28] ),
    .S0(_01471_),
    .S1(_01316_),
    .Z(_01483_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 _05677_ (.I(_01059_),
    .Z(_01484_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05678_ (.I(_01102_),
    .Z(_01485_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05679_ (.I0(\dp.rf.rf[4][28] ),
    .I1(\dp.rf.rf[5][28] ),
    .I2(\dp.rf.rf[6][28] ),
    .I3(\dp.rf.rf[7][28] ),
    .S0(_01484_),
    .S1(_01485_),
    .Z(_01486_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05680_ (.I0(_01483_),
    .I1(_01486_),
    .S(_01394_),
    .Z(_01487_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05681_ (.I0(_01482_),
    .I1(_01487_),
    .S(_01478_),
    .Z(_01488_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _05682_ (.A1(_01111_),
    .A2(_01479_),
    .B1(_01488_),
    .B2(_01112_),
    .ZN(_01489_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05683_ (.A1(_01290_),
    .A2(_01489_),
    .ZN(_01490_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _05684_ (.A1(_01290_),
    .A2(_05190_),
    .B(_01490_),
    .ZN(_01491_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _05685_ (.A1(_01288_),
    .A2(_01491_),
    .Z(_04857_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05686_ (.I(_04857_),
    .ZN(_04861_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _05687_ (.A1(\dp.rf.rf[10][28] ),
    .A2(_01362_),
    .B(_01377_),
    .C(\dp.rf.rf[8][28] ),
    .ZN(_01492_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _05688_ (.A1(_01415_),
    .A2(_01244_),
    .A3(_01245_),
    .A4(_01492_),
    .Z(_01493_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05689_ (.I0(\dp.rf.rf[10][28] ),
    .I1(\dp.rf.rf[11][28] ),
    .I2(\dp.rf.rf[14][28] ),
    .I3(\dp.rf.rf[15][28] ),
    .S0(_01345_),
    .S1(_01458_),
    .Z(_01494_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05690_ (.I(_01494_),
    .ZN(_01495_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05691_ (.I(_01367_),
    .Z(_01496_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05692_ (.I(_01496_),
    .Z(_01497_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05693_ (.I0(\dp.rf.rf[9][28] ),
    .I1(\dp.rf.rf[13][28] ),
    .S(_01364_),
    .Z(_01498_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _05694_ (.A1(\dp.rf.rf[12][28] ),
    .A2(_01497_),
    .B1(_01498_),
    .B2(_01422_),
    .ZN(_01499_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05695_ (.I(_01372_),
    .Z(_01500_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05696_ (.I0(_01495_),
    .I1(_01499_),
    .S(_01500_),
    .Z(_01501_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05697_ (.I0(\dp.rf.rf[25][28] ),
    .I1(\dp.rf.rf[29][28] ),
    .S(_01364_),
    .Z(_01502_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05698_ (.A1(_01422_),
    .A2(_01502_),
    .ZN(_01503_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05699_ (.I(_01212_),
    .Z(_01504_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05700_ (.I(_01196_),
    .Z(_01505_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05701_ (.I(_01218_),
    .Z(_01506_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _05702_ (.A1(\dp.rf.rf[28][28] ),
    .A2(_01504_),
    .A3(_01505_),
    .B(_01506_),
    .ZN(_01507_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 _05703_ (.I(_01128_),
    .Z(_01508_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05704_ (.I0(\dp.rf.rf[26][28] ),
    .I1(\dp.rf.rf[27][28] ),
    .I2(\dp.rf.rf[30][28] ),
    .I3(\dp.rf.rf[31][28] ),
    .S0(_01508_),
    .S1(_01145_),
    .Z(_01509_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05705_ (.A1(_01362_),
    .A2(_01509_),
    .ZN(_01510_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05706_ (.I(_01192_),
    .Z(_01511_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _05707_ (.A1(_01503_),
    .A2(_01507_),
    .B(_01510_),
    .C(_01511_),
    .ZN(_01512_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05708_ (.I(\dp.rf.rf[24][28] ),
    .ZN(_01513_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05709_ (.A1(\dp.rf.rf[26][28] ),
    .A2(_01353_),
    .Z(_01514_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _05710_ (.A1(_01438_),
    .A2(_01185_),
    .A3(_01174_),
    .B1(_01377_),
    .B2(_01514_),
    .ZN(_01515_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05711_ (.A1(_01513_),
    .A2(_01515_),
    .B(_01337_),
    .ZN(_01516_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05712_ (.I0(\dp.rf.rf[17][28] ),
    .I1(\dp.rf.rf[21][28] ),
    .S(_01432_),
    .Z(_01517_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05713_ (.A1(_01422_),
    .A2(_01517_),
    .ZN(_01518_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _05714_ (.A1(\dp.rf.rf[20][28] ),
    .A2(_01504_),
    .A3(_01505_),
    .B(_01506_),
    .ZN(_01519_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05715_ (.I(_01128_),
    .Z(_01520_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05716_ (.I0(\dp.rf.rf[18][28] ),
    .I1(\dp.rf.rf[19][28] ),
    .I2(\dp.rf.rf[22][28] ),
    .I3(\dp.rf.rf[23][28] ),
    .S0(_01520_),
    .S1(_01201_),
    .Z(_01521_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05717_ (.A1(_01362_),
    .A2(_01521_),
    .ZN(_01522_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _05718_ (.A1(_01518_),
    .A2(_01519_),
    .B(_01522_),
    .C(_01511_),
    .ZN(_01523_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05719_ (.I(\dp.rf.rf[16][28] ),
    .ZN(_01524_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05720_ (.A1(\dp.rf.rf[18][28] ),
    .A2(_01353_),
    .Z(_01525_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _05721_ (.A1(_01438_),
    .A2(_01185_),
    .A3(_01174_),
    .B1(_01377_),
    .B2(_01525_),
    .ZN(_01526_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05722_ (.A1(_01524_),
    .A2(_01526_),
    .B(_01178_),
    .ZN(_01527_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _05723_ (.A1(_01512_),
    .A2(_01516_),
    .B1(_01523_),
    .B2(_01527_),
    .ZN(_01528_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05724_ (.I(_01117_),
    .Z(_01529_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05725_ (.I(_01529_),
    .Z(_01530_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05726_ (.I(_01120_),
    .Z(_01531_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05727_ (.I(_01531_),
    .Z(_01532_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05728_ (.I(_01209_),
    .Z(_01533_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05729_ (.I0(\dp.rf.rf[2][28] ),
    .I1(\dp.rf.rf[3][28] ),
    .I2(\dp.rf.rf[6][28] ),
    .I3(\dp.rf.rf[7][28] ),
    .S0(_01532_),
    .S1(_01533_),
    .Z(_01534_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05730_ (.A1(_01530_),
    .A2(_01534_),
    .Z(_01535_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05731_ (.I(\dp.rf.rf[4][28] ),
    .ZN(_01536_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05732_ (.I0(\dp.rf.rf[1][28] ),
    .I1(\dp.rf.rf[5][28] ),
    .S(_01124_),
    .Z(_01537_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05733_ (.A1(_01422_),
    .A2(_01537_),
    .ZN(_01538_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _05734_ (.A1(_01536_),
    .A2(_01327_),
    .B(_01538_),
    .C(_01456_),
    .ZN(_01539_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _05735_ (.A1(\dp.rf.rf[2][28] ),
    .A2(_01362_),
    .B(\dp.rf.rf[0][28] ),
    .ZN(_01540_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 _05736_ (.I(net227),
    .Z(_01541_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _05737_ (.A1(_01130_),
    .A2(_01540_),
    .B(_01466_),
    .C(_01541_),
    .ZN(_01542_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _05738_ (.A1(_01535_),
    .A2(_01539_),
    .B(_01542_),
    .ZN(_01543_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _05739_ (.A1(_01493_),
    .A2(_01501_),
    .B1(_01528_),
    .B2(_01455_),
    .C(_01543_),
    .ZN(_01544_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _05740_ (.I(_01544_),
    .Z(_04856_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05741_ (.I(_04856_),
    .ZN(_04860_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05742_ (.A1(net16),
    .A2(_01301_),
    .ZN(_01545_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05743_ (.A1(_01299_),
    .A2(_01545_),
    .B(_01304_),
    .ZN(_05186_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _05744_ (.I(_01289_),
    .Z(_01546_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 _05745_ (.I(_01049_),
    .Z(_01547_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 _05746_ (.I(_01547_),
    .Z(_01548_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05747_ (.I(instr[21]),
    .Z(_01549_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05748_ (.I(_01549_),
    .Z(_01550_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05749_ (.I0(\dp.rf.rf[24][27] ),
    .I1(\dp.rf.rf[25][27] ),
    .I2(\dp.rf.rf[26][27] ),
    .I3(\dp.rf.rf[27][27] ),
    .S0(net249),
    .S1(_01550_),
    .Z(_01551_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05750_ (.I0(\dp.rf.rf[16][27] ),
    .I1(\dp.rf.rf[17][27] ),
    .I2(\dp.rf.rf[18][27] ),
    .I3(\dp.rf.rf[19][27] ),
    .S0(net249),
    .S1(_01550_),
    .Z(_01552_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 _05751_ (.I(_01547_),
    .Z(_01553_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _05752_ (.I(instr[21]),
    .Z(_01554_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05753_ (.I(_01554_),
    .Z(_01555_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05754_ (.I0(\dp.rf.rf[28][27] ),
    .I1(\dp.rf.rf[29][27] ),
    .I2(\dp.rf.rf[30][27] ),
    .I3(\dp.rf.rf[31][27] ),
    .S0(net256),
    .S1(_01555_),
    .Z(_01556_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05755_ (.I0(\dp.rf.rf[20][27] ),
    .I1(\dp.rf.rf[21][27] ),
    .I2(\dp.rf.rf[22][27] ),
    .I3(\dp.rf.rf[23][27] ),
    .S0(net249),
    .S1(_01550_),
    .Z(_01557_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05756_ (.I0(_01551_),
    .I1(_01552_),
    .I2(_01556_),
    .I3(_01557_),
    .S0(_01272_),
    .S1(_01400_),
    .Z(_01558_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05757_ (.I0(\dp.rf.rf[8][27] ),
    .I1(\dp.rf.rf[9][27] ),
    .I2(\dp.rf.rf[10][27] ),
    .I3(\dp.rf.rf[11][27] ),
    .S0(net256),
    .S1(_01555_),
    .Z(_01559_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05758_ (.I0(\dp.rf.rf[0][27] ),
    .I1(\dp.rf.rf[1][27] ),
    .I2(\dp.rf.rf[2][27] ),
    .I3(\dp.rf.rf[3][27] ),
    .S0(net256),
    .S1(_01555_),
    .Z(_01560_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _05759_ (.I(_01554_),
    .Z(_01561_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05760_ (.I0(\dp.rf.rf[12][27] ),
    .I1(\dp.rf.rf[13][27] ),
    .I2(\dp.rf.rf[14][27] ),
    .I3(\dp.rf.rf[15][27] ),
    .S0(_01261_),
    .S1(_01561_),
    .Z(_01562_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05761_ (.I0(\dp.rf.rf[4][27] ),
    .I1(\dp.rf.rf[5][27] ),
    .I2(\dp.rf.rf[6][27] ),
    .I3(\dp.rf.rf[7][27] ),
    .S0(net256),
    .S1(_01555_),
    .Z(_01563_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05762_ (.I0(_01559_),
    .I1(_01560_),
    .I2(_01562_),
    .I3(_01563_),
    .S0(_01272_),
    .S1(_01400_),
    .Z(_01564_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _05763_ (.A1(_01037_),
    .A2(_01558_),
    .B1(_01564_),
    .B2(_01112_),
    .ZN(_01565_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05764_ (.A1(_01546_),
    .A2(_01565_),
    .ZN(_01566_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _05765_ (.A1(_01290_),
    .A2(_05186_),
    .B(_01566_),
    .ZN(_01567_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _05766_ (.A1(_01288_),
    .A2(_01567_),
    .Z(_04865_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05767_ (.I(_04865_),
    .ZN(_04869_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05768_ (.I(_01230_),
    .Z(_01568_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05769_ (.I(_01363_),
    .Z(_01569_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05770_ (.I0(\dp.rf.rf[14][27] ),
    .I1(\dp.rf.rf[15][27] ),
    .S(_01569_),
    .Z(_01570_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05771_ (.I(net202),
    .Z(_01571_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05772_ (.A1(\dp.rf.rf[10][27] ),
    .A2(_01571_),
    .Z(_01572_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05773_ (.A1(\dp.rf.rf[11][27] ),
    .A2(_01429_),
    .ZN(_01573_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05774_ (.A1(_01224_),
    .A2(_01573_),
    .ZN(_01574_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _05775_ (.A1(_01568_),
    .A2(_01570_),
    .B1(_01572_),
    .B2(_01574_),
    .C(_01335_),
    .ZN(_01575_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05776_ (.I(_01430_),
    .Z(_01576_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05777_ (.I(_01121_),
    .Z(_01577_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05778_ (.I(_01381_),
    .Z(_01578_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05779_ (.I0(\dp.rf.rf[8][27] ),
    .I1(\dp.rf.rf[9][27] ),
    .I2(\dp.rf.rf[12][27] ),
    .I3(\dp.rf.rf[13][27] ),
    .S0(_01577_),
    .S1(_01578_),
    .Z(_01579_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05780_ (.I(_01199_),
    .Z(_01580_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05781_ (.A1(_01576_),
    .A2(_01579_),
    .B(_01580_),
    .ZN(_01581_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05782_ (.I(_01202_),
    .Z(_01582_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05783_ (.I0(\dp.rf.rf[2][27] ),
    .I1(\dp.rf.rf[3][27] ),
    .I2(\dp.rf.rf[6][27] ),
    .I3(\dp.rf.rf[7][27] ),
    .S0(_01582_),
    .S1(_01124_),
    .Z(_01583_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05784_ (.I(_01583_),
    .ZN(_01584_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05785_ (.I0(\dp.rf.rf[1][27] ),
    .I1(\dp.rf.rf[5][27] ),
    .S(_01369_),
    .Z(_01585_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _05786_ (.A1(\dp.rf.rf[4][27] ),
    .A2(_01368_),
    .B1(_01585_),
    .B2(_01442_),
    .ZN(_01586_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05787_ (.I0(_01584_),
    .I1(_01586_),
    .S(_01506_),
    .Z(_01587_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _05788_ (.A1(_01252_),
    .A2(_01134_),
    .B(_01142_),
    .ZN(_01588_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05789_ (.I(_01588_),
    .Z(_01589_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _05790_ (.A1(_01575_),
    .A2(_01581_),
    .B1(_01587_),
    .B2(_01361_),
    .C(_01589_),
    .ZN(_01590_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05791_ (.I0(\dp.rf.rf[22][27] ),
    .I1(\dp.rf.rf[23][27] ),
    .S(_01569_),
    .Z(_01591_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05792_ (.I0(\dp.rf.rf[18][27] ),
    .I1(\dp.rf.rf[19][27] ),
    .S(_01577_),
    .Z(_01592_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05793_ (.A1(_01139_),
    .A2(_01324_),
    .Z(_01593_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _05794_ (.A1(_01568_),
    .A2(_01591_),
    .B1(_01592_),
    .B2(_01593_),
    .C(_01530_),
    .ZN(_01594_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05795_ (.I(\dp.rf.rf[20][27] ),
    .ZN(_01595_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05796_ (.I0(\dp.rf.rf[17][27] ),
    .I1(\dp.rf.rf[21][27] ),
    .S(_01138_),
    .Z(_01596_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05797_ (.A1(_01371_),
    .A2(_01596_),
    .ZN(_01597_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _05798_ (.A1(_01595_),
    .A2(_01327_),
    .B(_01597_),
    .C(_01416_),
    .ZN(_01598_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _05799_ (.A1(\dp.rf.rf[16][27] ),
    .A2(_01356_),
    .B1(_01598_),
    .B2(_01541_),
    .ZN(_01599_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05800_ (.I(_01179_),
    .Z(_01600_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05801_ (.I0(\dp.rf.rf[26][27] ),
    .I1(\dp.rf.rf[27][27] ),
    .I2(\dp.rf.rf[30][27] ),
    .I3(\dp.rf.rf[31][27] ),
    .S0(_01600_),
    .S1(_01210_),
    .Z(_01601_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05802_ (.I0(\dp.rf.rf[24][27] ),
    .I1(\dp.rf.rf[25][27] ),
    .I2(\dp.rf.rf[28][27] ),
    .I3(\dp.rf.rf[29][27] ),
    .S0(_01600_),
    .S1(_01210_),
    .Z(_01602_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _05803_ (.A1(_01335_),
    .A2(_01601_),
    .B1(_01602_),
    .B2(_01500_),
    .ZN(_01603_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _05804_ (.A1(_01594_),
    .A2(_01599_),
    .B1(_01603_),
    .B2(_01385_),
    .C(_01455_),
    .ZN(_01604_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _05805_ (.A1(_01590_),
    .A2(_01604_),
    .Z(_04864_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05806_ (.I(_04864_),
    .ZN(_04868_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05807_ (.I(_01093_),
    .Z(_01605_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05808_ (.A1(net15),
    .A2(_01301_),
    .ZN(_01606_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05809_ (.A1(_01299_),
    .A2(_01606_),
    .B(_01304_),
    .ZN(_05182_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _05810_ (.A1(_01037_),
    .A2(_01060_),
    .Z(_01607_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 _05811_ (.I(_01607_),
    .Z(_01608_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05812_ (.I(_01098_),
    .Z(_01609_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05813_ (.I0(\dp.rf.rf[24][26] ),
    .I1(\dp.rf.rf[25][26] ),
    .I2(\dp.rf.rf[26][26] ),
    .I3(\dp.rf.rf[27][26] ),
    .S0(_01609_),
    .S1(_01561_),
    .Z(_01610_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05814_ (.I0(\dp.rf.rf[16][26] ),
    .I1(\dp.rf.rf[17][26] ),
    .I2(\dp.rf.rf[18][26] ),
    .I3(\dp.rf.rf[19][26] ),
    .S0(_01553_),
    .S1(_01555_),
    .Z(_01611_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05815_ (.I0(\dp.rf.rf[28][26] ),
    .I1(\dp.rf.rf[29][26] ),
    .I2(\dp.rf.rf[30][26] ),
    .I3(\dp.rf.rf[31][26] ),
    .S0(_01261_),
    .S1(_01561_),
    .Z(_01612_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05816_ (.I0(\dp.rf.rf[20][26] ),
    .I1(\dp.rf.rf[21][26] ),
    .I2(\dp.rf.rf[22][26] ),
    .I3(\dp.rf.rf[23][26] ),
    .S0(_01609_),
    .S1(_01561_),
    .Z(_01613_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05817_ (.I0(_01610_),
    .I1(_01611_),
    .I2(_01612_),
    .I3(_01613_),
    .S0(_01272_),
    .S1(_01400_),
    .Z(_01614_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05818_ (.I0(\dp.rf.rf[8][26] ),
    .I1(\dp.rf.rf[9][26] ),
    .I2(\dp.rf.rf[10][26] ),
    .I3(\dp.rf.rf[11][26] ),
    .S0(_01609_),
    .S1(_01561_),
    .Z(_01615_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05819_ (.I0(\dp.rf.rf[0][26] ),
    .I1(\dp.rf.rf[1][26] ),
    .I2(\dp.rf.rf[2][26] ),
    .I3(\dp.rf.rf[3][26] ),
    .S0(_01609_),
    .S1(_01561_),
    .Z(_01616_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05820_ (.I0(\dp.rf.rf[12][26] ),
    .I1(\dp.rf.rf[13][26] ),
    .I2(\dp.rf.rf[14][26] ),
    .I3(\dp.rf.rf[15][26] ),
    .S0(_01261_),
    .S1(_01561_),
    .Z(_01617_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05821_ (.I0(\dp.rf.rf[4][26] ),
    .I1(\dp.rf.rf[5][26] ),
    .I2(\dp.rf.rf[6][26] ),
    .I3(\dp.rf.rf[7][26] ),
    .S0(_01609_),
    .S1(_01561_),
    .Z(_01618_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05822_ (.I0(_01615_),
    .I1(_01616_),
    .I2(_01617_),
    .I3(_01618_),
    .S0(_01272_),
    .S1(_01400_),
    .Z(_01619_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05823_ (.I0(_01614_),
    .I1(_01619_),
    .S(_01058_),
    .Z(_01620_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _05824_ (.A1(net192),
    .A2(_01620_),
    .ZN(_01621_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05825_ (.I(_01621_),
    .ZN(_01622_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05826_ (.A1(_01289_),
    .A2(_01622_),
    .Z(_01623_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05827_ (.A1(_01605_),
    .A2(_05182_),
    .B(_01623_),
    .ZN(_01624_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _05828_ (.A1(_01288_),
    .A2(_01624_),
    .Z(_04873_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05829_ (.I(_04873_),
    .ZN(_04877_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05830_ (.I0(\dp.rf.rf[14][26] ),
    .I1(\dp.rf.rf[15][26] ),
    .S(_01577_),
    .Z(_01625_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05831_ (.I(net202),
    .Z(_01626_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05832_ (.A1(\dp.rf.rf[10][26] ),
    .A2(_01626_),
    .Z(_01627_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05833_ (.A1(\dp.rf.rf[11][26] ),
    .A2(_01569_),
    .ZN(_01628_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05834_ (.A1(_01224_),
    .A2(_01628_),
    .ZN(_01629_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _05835_ (.A1(_01568_),
    .A2(_01625_),
    .B1(_01627_),
    .B2(_01629_),
    .C(_01335_),
    .ZN(_01630_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05836_ (.I0(\dp.rf.rf[8][26] ),
    .I1(\dp.rf.rf[9][26] ),
    .I2(\dp.rf.rf[12][26] ),
    .I3(\dp.rf.rf[13][26] ),
    .S0(_01532_),
    .S1(_01533_),
    .Z(_01631_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05837_ (.A1(_01576_),
    .A2(_01631_),
    .B(_01237_),
    .ZN(_01632_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05838_ (.I0(\dp.rf.rf[2][26] ),
    .I1(\dp.rf.rf[3][26] ),
    .I2(\dp.rf.rf[6][26] ),
    .I3(\dp.rf.rf[7][26] ),
    .S0(_01531_),
    .S1(_01443_),
    .Z(_01633_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05839_ (.A1(_01119_),
    .A2(_01633_),
    .ZN(_01634_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05840_ (.I0(\dp.rf.rf[1][26] ),
    .I1(\dp.rf.rf[5][26] ),
    .S(_01144_),
    .Z(_01635_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05841_ (.I(_01189_),
    .Z(_01636_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _05842_ (.A1(\dp.rf.rf[4][26] ),
    .A2(_01496_),
    .B1(_01635_),
    .B2(_01636_),
    .C(_01241_),
    .ZN(_01637_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _05843_ (.A1(_01337_),
    .A2(_01435_),
    .A3(_01634_),
    .A4(_01637_),
    .Z(_01638_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _05844_ (.A1(_01630_),
    .A2(_01632_),
    .B(_01638_),
    .C(_01589_),
    .ZN(_01639_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05845_ (.I0(\dp.rf.rf[26][26] ),
    .I1(\dp.rf.rf[27][26] ),
    .I2(\dp.rf.rf[30][26] ),
    .I3(\dp.rf.rf[31][26] ),
    .S0(_01212_),
    .S1(_01458_),
    .Z(_01640_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05846_ (.I0(\dp.rf.rf[24][26] ),
    .I1(\dp.rf.rf[25][26] ),
    .I2(\dp.rf.rf[28][26] ),
    .I3(\dp.rf.rf[29][26] ),
    .S0(_01212_),
    .S1(_01458_),
    .Z(_01641_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _05847_ (.A1(_01335_),
    .A2(_01640_),
    .B1(_01641_),
    .B2(_01500_),
    .ZN(_01642_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05848_ (.I0(\dp.rf.rf[22][26] ),
    .I1(\dp.rf.rf[23][26] ),
    .S(_01345_),
    .Z(_01643_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05849_ (.A1(\dp.rf.rf[18][26] ),
    .A2(_01626_),
    .Z(_01644_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05850_ (.I(_01147_),
    .Z(_01645_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05851_ (.A1(\dp.rf.rf[19][26] ),
    .A2(_01645_),
    .ZN(_01646_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05852_ (.A1(_01224_),
    .A2(_01646_),
    .ZN(_01647_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _05853_ (.A1(_01339_),
    .A2(_01643_),
    .B1(_01644_),
    .B2(_01647_),
    .C(_01335_),
    .ZN(_01648_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05854_ (.I(\dp.rf.rf[20][26] ),
    .ZN(_01649_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05855_ (.I0(\dp.rf.rf[17][26] ),
    .I1(\dp.rf.rf[21][26] ),
    .S(_01248_),
    .Z(_01650_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05856_ (.A1(_01328_),
    .A2(_01650_),
    .ZN(_01651_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _05857_ (.A1(_01649_),
    .A2(_01327_),
    .B(_01651_),
    .C(_01213_),
    .ZN(_01652_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _05858_ (.A1(\dp.rf.rf[16][26] ),
    .A2(_01356_),
    .B1(_01652_),
    .B2(net235),
    .ZN(_01653_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _05859_ (.A1(_01385_),
    .A2(_01642_),
    .B1(_01648_),
    .B2(_01653_),
    .C(_01455_),
    .ZN(_01654_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _05860_ (.A1(_01639_),
    .A2(_01654_),
    .Z(_04872_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _05861_ (.I(_04872_),
    .ZN(_04876_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05862_ (.A1(net14),
    .A2(_01301_),
    .ZN(_01655_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05863_ (.A1(_01299_),
    .A2(_01655_),
    .B(_01304_),
    .ZN(_05178_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _05864_ (.I(_01058_),
    .Z(_01656_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 _05865_ (.I(_01049_),
    .Z(_01657_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05866_ (.I(_01657_),
    .Z(_01658_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _05867_ (.I(_01408_),
    .Z(_01659_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05868_ (.I0(\dp.rf.rf[28][25] ),
    .I1(\dp.rf.rf[29][25] ),
    .I2(\dp.rf.rf[30][25] ),
    .I3(\dp.rf.rf[31][25] ),
    .S0(_01658_),
    .S1(_01659_),
    .Z(_01660_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05869_ (.I(_01038_),
    .Z(_01661_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05870_ (.I(_01661_),
    .Z(_01662_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05871_ (.I0(\dp.rf.rf[20][25] ),
    .I1(\dp.rf.rf[21][25] ),
    .I2(\dp.rf.rf[22][25] ),
    .I3(\dp.rf.rf[23][25] ),
    .S0(_01662_),
    .S1(_01659_),
    .Z(_01663_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05872_ (.I0(\dp.rf.rf[24][25] ),
    .I1(\dp.rf.rf[25][25] ),
    .I2(\dp.rf.rf[26][25] ),
    .I3(\dp.rf.rf[27][25] ),
    .S0(_01658_),
    .S1(_01659_),
    .Z(_01664_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05873_ (.I0(\dp.rf.rf[16][25] ),
    .I1(\dp.rf.rf[17][25] ),
    .I2(\dp.rf.rf[18][25] ),
    .I3(\dp.rf.rf[19][25] ),
    .S0(_01658_),
    .S1(_01659_),
    .Z(_01665_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05874_ (.I(_01398_),
    .Z(_01666_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _05875_ (.I(net11),
    .ZN(_01667_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05876_ (.I(_01667_),
    .Z(_01668_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05877_ (.I(_01668_),
    .Z(_01669_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _05878_ (.I0(_01660_),
    .I1(_01663_),
    .I2(_01664_),
    .I3(_01665_),
    .S0(_01666_),
    .S1(_01669_),
    .Z(_01670_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _05879_ (.I(net12),
    .Z(_01671_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _05880_ (.A1(_01057_),
    .A2(_01671_),
    .ZN(_01672_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05881_ (.I0(\dp.rf.rf[12][25] ),
    .I1(\dp.rf.rf[13][25] ),
    .I2(\dp.rf.rf[14][25] ),
    .I3(\dp.rf.rf[15][25] ),
    .S0(_01657_),
    .S1(_01408_),
    .Z(_01673_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05882_ (.I0(\dp.rf.rf[8][25] ),
    .I1(\dp.rf.rf[9][25] ),
    .I2(\dp.rf.rf[10][25] ),
    .I3(\dp.rf.rf[11][25] ),
    .S0(_01657_),
    .S1(_01408_),
    .Z(_01674_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05883_ (.I0(_01673_),
    .I1(_01674_),
    .S(_01668_),
    .Z(_01675_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _05884_ (.A1(_01672_),
    .A2(_01675_),
    .Z(_01676_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _05885_ (.A1(_01398_),
    .A2(_01057_),
    .ZN(_01677_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05886_ (.I0(\dp.rf.rf[4][25] ),
    .I1(\dp.rf.rf[5][25] ),
    .I2(\dp.rf.rf[6][25] ),
    .I3(\dp.rf.rf[7][25] ),
    .S0(net226),
    .S1(_01549_),
    .Z(_01678_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05887_ (.I0(\dp.rf.rf[0][25] ),
    .I1(\dp.rf.rf[1][25] ),
    .I2(\dp.rf.rf[2][25] ),
    .I3(\dp.rf.rf[3][25] ),
    .S0(net226),
    .S1(_01549_),
    .Z(_01679_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05888_ (.I0(_01678_),
    .I1(_01679_),
    .S(_01668_),
    .Z(_01680_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _05889_ (.A1(net224),
    .A2(_01680_),
    .Z(_01681_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _05890_ (.A1(net192),
    .A2(_01676_),
    .A3(_01681_),
    .Z(_01682_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _05891_ (.A1(_01656_),
    .A2(_01670_),
    .B(_01682_),
    .ZN(_01683_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05892_ (.A1(_01605_),
    .A2(_01683_),
    .ZN(_01684_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05893_ (.A1(_01605_),
    .A2(_05178_),
    .B(_01684_),
    .ZN(_01685_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _05894_ (.A1(_01288_),
    .A2(_01685_),
    .Z(_04881_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05895_ (.I(_04881_),
    .ZN(_04885_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05896_ (.I0(\dp.rf.rf[10][25] ),
    .I1(\dp.rf.rf[11][25] ),
    .I2(\dp.rf.rf[14][25] ),
    .I3(\dp.rf.rf[15][25] ),
    .S0(_01582_),
    .S1(_01124_),
    .Z(_01686_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05897_ (.I0(\dp.rf.rf[8][25] ),
    .I1(\dp.rf.rf[9][25] ),
    .I2(\dp.rf.rf[12][25] ),
    .I3(\dp.rf.rf[13][25] ),
    .S0(_01582_),
    .S1(_01124_),
    .Z(_01687_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05898_ (.I0(_01686_),
    .I1(_01687_),
    .S(_01372_),
    .Z(_01688_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _05899_ (.A1(_01580_),
    .A2(_01688_),
    .Z(_01689_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05900_ (.I0(\dp.rf.rf[2][25] ),
    .I1(\dp.rf.rf[3][25] ),
    .I2(\dp.rf.rf[6][25] ),
    .I3(\dp.rf.rf[7][25] ),
    .S0(_01532_),
    .S1(_01533_),
    .Z(_01690_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05901_ (.A1(_01530_),
    .A2(_01690_),
    .ZN(_01691_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05902_ (.I0(\dp.rf.rf[1][25] ),
    .I1(\dp.rf.rf[5][25] ),
    .S(_01145_),
    .Z(_01692_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05903_ (.I(_01636_),
    .Z(_01693_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _05904_ (.A1(\dp.rf.rf[4][25] ),
    .A2(_01497_),
    .B1(_01692_),
    .B2(_01693_),
    .C(_01173_),
    .ZN(_01694_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _05905_ (.A1(_01361_),
    .A2(_01691_),
    .A3(_01694_),
    .ZN(_01695_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _05906_ (.A1(_01376_),
    .A2(_01689_),
    .A3(_01695_),
    .Z(_01696_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _05907_ (.A1(_01141_),
    .A2(net273),
    .Z(_01697_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05908_ (.I0(\dp.rf.rf[18][25] ),
    .I1(\dp.rf.rf[19][25] ),
    .I2(\dp.rf.rf[22][25] ),
    .I3(\dp.rf.rf[23][25] ),
    .S0(_01645_),
    .S1(_01533_),
    .Z(_01698_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05909_ (.I(_01698_),
    .ZN(_01699_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05910_ (.I0(\dp.rf.rf[16][25] ),
    .I1(\dp.rf.rf[17][25] ),
    .I2(\dp.rf.rf[20][25] ),
    .I3(\dp.rf.rf[21][25] ),
    .S0(_01157_),
    .S1(_01458_),
    .Z(_01700_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05911_ (.A1(_01500_),
    .A2(_01700_),
    .B(_01178_),
    .ZN(_01701_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _05912_ (.A1(_01697_),
    .A2(_01699_),
    .B1(_01701_),
    .B2(_01455_),
    .ZN(_01702_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05913_ (.I0(\dp.rf.rf[30][25] ),
    .I1(\dp.rf.rf[31][25] ),
    .S(_01645_),
    .Z(_01703_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _05914_ (.A1(_01568_),
    .A2(_01703_),
    .B(_01511_),
    .C(_01456_),
    .ZN(_01704_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05915_ (.A1(\dp.rf.rf[27][25] ),
    .A2(_01577_),
    .Z(_01705_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _05916_ (.A1(_01146_),
    .A2(_01435_),
    .B1(_01571_),
    .B2(\dp.rf.rf[26][25] ),
    .C(_01705_),
    .ZN(_01706_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05917_ (.I0(\dp.rf.rf[24][25] ),
    .I1(\dp.rf.rf[25][25] ),
    .I2(\dp.rf.rf[28][25] ),
    .I3(\dp.rf.rf[29][25] ),
    .S0(_01345_),
    .S1(_01458_),
    .Z(_01707_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05918_ (.A1(_01500_),
    .A2(_01707_),
    .ZN(_01708_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _05919_ (.A1(_01704_),
    .A2(_01706_),
    .B(_01708_),
    .C(_01385_),
    .ZN(_01709_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05920_ (.A1(_01702_),
    .A2(_01709_),
    .Z(_01710_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _05921_ (.A1(_01696_),
    .A2(_01710_),
    .Z(_04880_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05922_ (.I(_04880_),
    .ZN(_04884_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05923_ (.I0(\dp.rf.rf[24][24] ),
    .I1(\dp.rf.rf[25][24] ),
    .I2(\dp.rf.rf[26][24] ),
    .I3(\dp.rf.rf[27][24] ),
    .S0(_01484_),
    .S1(_01485_),
    .Z(_01711_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05924_ (.I0(\dp.rf.rf[16][24] ),
    .I1(\dp.rf.rf[17][24] ),
    .I2(\dp.rf.rf[18][24] ),
    .I3(\dp.rf.rf[19][24] ),
    .S0(_01484_),
    .S1(_01485_),
    .Z(_01712_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05925_ (.I0(_01711_),
    .I1(_01712_),
    .S(_01394_),
    .Z(_01713_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05926_ (.A1(_01669_),
    .A2(_01713_),
    .ZN(_01714_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05927_ (.I0(\dp.rf.rf[28][24] ),
    .I1(\dp.rf.rf[29][24] ),
    .I2(\dp.rf.rf[30][24] ),
    .I3(\dp.rf.rf[31][24] ),
    .S0(_01390_),
    .S1(_01391_),
    .Z(_01715_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05928_ (.I0(\dp.rf.rf[20][24] ),
    .I1(\dp.rf.rf[21][24] ),
    .I2(\dp.rf.rf[22][24] ),
    .I3(\dp.rf.rf[23][24] ),
    .S0(_01390_),
    .S1(_01391_),
    .Z(_01716_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05929_ (.I0(_01715_),
    .I1(_01716_),
    .S(_01394_),
    .Z(_01717_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05930_ (.A1(_01478_),
    .A2(_01717_),
    .B(_01058_),
    .ZN(_01718_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05931_ (.I0(\dp.rf.rf[12][24] ),
    .I1(\dp.rf.rf[13][24] ),
    .I2(\dp.rf.rf[14][24] ),
    .I3(\dp.rf.rf[15][24] ),
    .S0(_01661_),
    .S1(_01391_),
    .Z(_01719_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05932_ (.I0(\dp.rf.rf[8][24] ),
    .I1(\dp.rf.rf[9][24] ),
    .I2(\dp.rf.rf[10][24] ),
    .I3(\dp.rf.rf[11][24] ),
    .S0(_01661_),
    .S1(_01391_),
    .Z(_01720_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05933_ (.I0(_01719_),
    .I1(_01720_),
    .S(_01668_),
    .Z(_01721_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05934_ (.I0(\dp.rf.rf[4][24] ),
    .I1(\dp.rf.rf[5][24] ),
    .I2(\dp.rf.rf[6][24] ),
    .I3(\dp.rf.rf[7][24] ),
    .S0(_01657_),
    .S1(_01408_),
    .Z(_01722_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05935_ (.I0(\dp.rf.rf[0][24] ),
    .I1(\dp.rf.rf[1][24] ),
    .I2(\dp.rf.rf[2][24] ),
    .I3(\dp.rf.rf[3][24] ),
    .S0(_01657_),
    .S1(_01408_),
    .Z(_01723_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05936_ (.I0(_01722_),
    .I1(_01723_),
    .S(_01668_),
    .Z(_01724_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _05937_ (.A1(_01672_),
    .A2(_01721_),
    .B1(_01724_),
    .B2(net225),
    .C(_01607_),
    .ZN(_01725_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _05938_ (.A1(_01714_),
    .A2(_01718_),
    .B(_01725_),
    .ZN(_01726_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05939_ (.A1(_01111_),
    .A2(_01301_),
    .ZN(_01727_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05940_ (.A1(_01299_),
    .A2(_01727_),
    .B(_01304_),
    .ZN(_05174_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05941_ (.A1(_01605_),
    .A2(_05174_),
    .Z(_01728_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05942_ (.A1(_01290_),
    .A2(_01726_),
    .B(_01728_),
    .ZN(_01729_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _05943_ (.A1(_01288_),
    .A2(_01729_),
    .Z(_04889_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05944_ (.I(_04889_),
    .ZN(_04893_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05945_ (.I0(\dp.rf.rf[18][24] ),
    .I1(\dp.rf.rf[19][24] ),
    .I2(\dp.rf.rf[22][24] ),
    .I3(\dp.rf.rf[23][24] ),
    .S0(_01577_),
    .S1(_01578_),
    .Z(_01730_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05946_ (.I0(\dp.rf.rf[17][24] ),
    .I1(\dp.rf.rf[21][24] ),
    .S(_01209_),
    .Z(_01731_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05947_ (.A1(_01442_),
    .A2(_01731_),
    .ZN(_01732_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _05948_ (.A1(\dp.rf.rf[20][24] ),
    .A2(_01429_),
    .A3(_01230_),
    .B(_01372_),
    .ZN(_01733_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _05949_ (.A1(_01732_),
    .A2(_01733_),
    .B(_01337_),
    .C(_01435_),
    .ZN(_01734_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05950_ (.I(\dp.rf.rf[16][24] ),
    .ZN(_01735_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _05951_ (.A1(_01027_),
    .A2(net180),
    .A3(_01174_),
    .B(_01355_),
    .ZN(_01736_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05952_ (.I(_01736_),
    .Z(_01737_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05953_ (.A1(_01735_),
    .A2(_01737_),
    .ZN(_01738_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _05954_ (.A1(_01335_),
    .A2(_01730_),
    .B1(_01734_),
    .B2(_01738_),
    .ZN(_01739_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05955_ (.I0(\dp.rf.rf[26][24] ),
    .I1(\dp.rf.rf[27][24] ),
    .I2(\dp.rf.rf[30][24] ),
    .I3(\dp.rf.rf[31][24] ),
    .S0(_01520_),
    .S1(_01364_),
    .Z(_01740_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05956_ (.I0(\dp.rf.rf[24][24] ),
    .I1(\dp.rf.rf[25][24] ),
    .I2(\dp.rf.rf[28][24] ),
    .I3(\dp.rf.rf[29][24] ),
    .S0(_01363_),
    .S1(_01364_),
    .Z(_01741_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05957_ (.I0(_01740_),
    .I1(_01741_),
    .S(_01430_),
    .Z(_01742_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _05958_ (.A1(_01415_),
    .A2(_01742_),
    .B(net205),
    .ZN(_01743_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05959_ (.I0(\dp.rf.rf[14][24] ),
    .I1(\dp.rf.rf[15][24] ),
    .S(_01508_),
    .Z(_01744_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05960_ (.I(_01744_),
    .ZN(_01745_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05961_ (.A1(_01146_),
    .A2(_01745_),
    .B(_01151_),
    .ZN(_01746_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _05962_ (.A1(_01154_),
    .A2(_01155_),
    .A3(_01090_),
    .A4(\dp.rf.rf[10][24] ),
    .ZN(_01747_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05963_ (.I(\dp.rf.rf[10][24] ),
    .ZN(_01748_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _05964_ (.A1(_01028_),
    .A2(_01185_),
    .A3(_01747_),
    .B1(_01748_),
    .B2(_01212_),
    .ZN(_01749_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05965_ (.A1(\dp.rf.rf[11][24] ),
    .A2(_01428_),
    .Z(_01750_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _05966_ (.A1(_01164_),
    .A2(_01166_),
    .A3(_01749_),
    .A4(_01750_),
    .Z(_01751_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05967_ (.I0(\dp.rf.rf[8][24] ),
    .I1(\dp.rf.rf[9][24] ),
    .I2(\dp.rf.rf[12][24] ),
    .I3(\dp.rf.rf[13][24] ),
    .S0(_01345_),
    .S1(_01458_),
    .Z(_01752_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _05968_ (.A1(_01746_),
    .A2(_01751_),
    .B1(_01752_),
    .B2(_01500_),
    .C(_01237_),
    .ZN(_01753_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05969_ (.I0(\dp.rf.rf[2][24] ),
    .I1(\dp.rf.rf[3][24] ),
    .I2(\dp.rf.rf[6][24] ),
    .I3(\dp.rf.rf[7][24] ),
    .S0(_01520_),
    .S1(_01201_),
    .Z(_01754_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05970_ (.A1(_01416_),
    .A2(_01754_),
    .Z(_01755_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05971_ (.I(\dp.rf.rf[4][24] ),
    .ZN(_01756_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05972_ (.I0(\dp.rf.rf[1][24] ),
    .I1(\dp.rf.rf[5][24] ),
    .S(_01168_),
    .Z(_01757_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05973_ (.A1(_01371_),
    .A2(_01757_),
    .ZN(_01758_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _05974_ (.A1(_01756_),
    .A2(_01327_),
    .B(_01758_),
    .C(_01416_),
    .ZN(_01759_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _05975_ (.A1(_01541_),
    .A2(_01755_),
    .A3(_01759_),
    .B(_01376_),
    .ZN(_01760_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _05976_ (.A1(_01739_),
    .A2(_01743_),
    .B1(_01753_),
    .B2(_01760_),
    .ZN(_04888_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05977_ (.I(_04888_),
    .ZN(_04892_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05978_ (.I(_01671_),
    .Z(_01761_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05979_ (.A1(_01761_),
    .A2(_01301_),
    .ZN(_01762_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05980_ (.A1(_01299_),
    .A2(_01762_),
    .B(_01304_),
    .ZN(_05170_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _05981_ (.I(_01671_),
    .Z(_01763_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05982_ (.I0(\dp.rf.rf[6][23] ),
    .I1(\dp.rf.rf[7][23] ),
    .I2(\dp.rf.rf[14][23] ),
    .I3(\dp.rf.rf[15][23] ),
    .S0(_01279_),
    .S1(_01763_),
    .Z(_01764_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05983_ (.I0(\dp.rf.rf[4][23] ),
    .I1(\dp.rf.rf[5][23] ),
    .I2(\dp.rf.rf[12][23] ),
    .I3(\dp.rf.rf[13][23] ),
    .S0(_01279_),
    .S1(_01763_),
    .Z(_01765_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05984_ (.I(_01103_),
    .Z(_01766_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05985_ (.I0(_01764_),
    .I1(_01765_),
    .S(_01766_),
    .Z(_01767_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05986_ (.I0(\dp.rf.rf[8][23] ),
    .I1(\dp.rf.rf[9][23] ),
    .I2(\dp.rf.rf[10][23] ),
    .I3(\dp.rf.rf[11][23] ),
    .S0(net226),
    .S1(_01549_),
    .Z(_01768_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05987_ (.I0(\dp.rf.rf[0][23] ),
    .I1(\dp.rf.rf[1][23] ),
    .I2(\dp.rf.rf[2][23] ),
    .I3(\dp.rf.rf[3][23] ),
    .S0(net226),
    .S1(_01549_),
    .Z(_01769_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05988_ (.I0(_01768_),
    .I1(_01769_),
    .S(_01398_),
    .Z(_01770_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05989_ (.A1(_01607_),
    .A2(_01770_),
    .Z(_01771_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05990_ (.I0(_01767_),
    .I1(_01771_),
    .S(_01669_),
    .Z(_01772_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _05991_ (.I(_01471_),
    .Z(_01773_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _05992_ (.I(_01485_),
    .Z(_01774_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05993_ (.I0(\dp.rf.rf[28][23] ),
    .I1(\dp.rf.rf[29][23] ),
    .I2(\dp.rf.rf[30][23] ),
    .I3(\dp.rf.rf[31][23] ),
    .S0(_01773_),
    .S1(_01774_),
    .Z(_01775_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05994_ (.I0(\dp.rf.rf[20][23] ),
    .I1(\dp.rf.rf[21][23] ),
    .I2(\dp.rf.rf[22][23] ),
    .I3(\dp.rf.rf[23][23] ),
    .S0(_01773_),
    .S1(_01774_),
    .Z(_01776_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05995_ (.I0(_01775_),
    .I1(_01776_),
    .S(_01311_),
    .Z(_01777_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05996_ (.A1(net13),
    .A2(net195),
    .Z(_01778_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _05997_ (.I(_01667_),
    .Z(_01779_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05998_ (.A1(_01037_),
    .A2(_01779_),
    .Z(_01780_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05999_ (.I0(\dp.rf.rf[18][23] ),
    .I1(\dp.rf.rf[19][23] ),
    .I2(\dp.rf.rf[26][23] ),
    .I3(\dp.rf.rf[27][23] ),
    .S0(_01609_),
    .S1(_01763_),
    .Z(_01781_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06000_ (.I0(\dp.rf.rf[16][23] ),
    .I1(\dp.rf.rf[17][23] ),
    .I2(\dp.rf.rf[24][23] ),
    .I3(\dp.rf.rf[25][23] ),
    .S0(_01609_),
    .S1(_01763_),
    .Z(_01782_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06001_ (.I0(_01781_),
    .I1(_01782_),
    .S(_01766_),
    .Z(_01783_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06002_ (.A1(_01780_),
    .A2(_01783_),
    .Z(_01784_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _06003_ (.A1(_01656_),
    .A2(_01772_),
    .B1(_01777_),
    .B2(net214),
    .C(_01784_),
    .ZN(_01785_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06004_ (.A1(_01546_),
    .A2(_01785_),
    .ZN(_01786_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06005_ (.A1(_01290_),
    .A2(_05170_),
    .B(_01786_),
    .ZN(_01787_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06006_ (.A1(_01288_),
    .A2(_01787_),
    .Z(_04897_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06007_ (.I(_04897_),
    .ZN(_04901_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06008_ (.I0(\dp.rf.rf[25][23] ),
    .I1(\dp.rf.rf[29][23] ),
    .S(_01533_),
    .Z(_01788_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06009_ (.A1(_01693_),
    .A2(_01788_),
    .ZN(_01789_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06010_ (.A1(_01372_),
    .A2(_01244_),
    .Z(_01790_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06011_ (.A1(\dp.rf.rf[24][23] ),
    .A2(_01377_),
    .B1(_01497_),
    .B2(\dp.rf.rf[28][23] ),
    .C(_01790_),
    .ZN(_01791_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _06012_ (.A1(_01580_),
    .A2(_01789_),
    .A3(_01791_),
    .Z(_01792_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06013_ (.I0(\dp.rf.rf[17][23] ),
    .I1(\dp.rf.rf[21][23] ),
    .S(_01533_),
    .Z(_01793_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06014_ (.A1(_01693_),
    .A2(_01793_),
    .ZN(_01794_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06015_ (.A1(\dp.rf.rf[16][23] ),
    .A2(_01377_),
    .B1(_01497_),
    .B2(\dp.rf.rf[20][23] ),
    .C(_01790_),
    .ZN(_01795_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _06016_ (.A1(_01541_),
    .A2(_01794_),
    .A3(_01795_),
    .Z(_01796_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06017_ (.I0(\dp.rf.rf[26][23] ),
    .I1(\dp.rf.rf[27][23] ),
    .I2(\dp.rf.rf[30][23] ),
    .I3(\dp.rf.rf[31][23] ),
    .S0(_01532_),
    .S1(_01210_),
    .Z(_01797_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06018_ (.I0(\dp.rf.rf[18][23] ),
    .I1(\dp.rf.rf[19][23] ),
    .I2(\dp.rf.rf[22][23] ),
    .I3(\dp.rf.rf[23][23] ),
    .S0(_01532_),
    .S1(_01210_),
    .Z(_01798_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06019_ (.I0(_01797_),
    .I1(_01798_),
    .S(_01337_),
    .Z(_01799_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _06020_ (.A1(_01244_),
    .A2(_01335_),
    .A3(_01799_),
    .ZN(_01800_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06021_ (.I0(\dp.rf.rf[1][23] ),
    .I1(\dp.rf.rf[5][23] ),
    .S(_01201_),
    .Z(_01801_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06022_ (.A1(\dp.rf.rf[4][23] ),
    .A2(_01497_),
    .B1(_01801_),
    .B2(_01693_),
    .C(_01173_),
    .ZN(_01802_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06023_ (.I0(\dp.rf.rf[2][23] ),
    .I1(\dp.rf.rf[6][23] ),
    .S(_01369_),
    .Z(_01803_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _06024_ (.A1(_01442_),
    .A2(_01529_),
    .A3(_01803_),
    .Z(_01804_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06025_ (.I0(\dp.rf.rf[3][23] ),
    .I1(\dp.rf.rf[7][23] ),
    .S(_01138_),
    .Z(_01805_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _06026_ (.A1(_01569_),
    .A2(_01213_),
    .A3(_01805_),
    .Z(_01806_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _06027_ (.A1(_01245_),
    .A2(_01804_),
    .A3(_01806_),
    .ZN(_01807_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _06028_ (.A1(\dp.rf.rf[2][23] ),
    .A2(_01213_),
    .B(_01169_),
    .C(_01645_),
    .ZN(_01808_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06029_ (.I(_01808_),
    .ZN(_01809_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06030_ (.A1(_01435_),
    .A2(_01809_),
    .B(\dp.rf.rf[0][23] ),
    .ZN(_01810_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _06031_ (.A1(_01802_),
    .A2(_01807_),
    .B(_01810_),
    .C(_01385_),
    .ZN(_01811_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06032_ (.I0(\dp.rf.rf[10][23] ),
    .I1(\dp.rf.rf[11][23] ),
    .I2(\dp.rf.rf[14][23] ),
    .I3(\dp.rf.rf[15][23] ),
    .S0(_01121_),
    .S1(_01432_),
    .Z(_01812_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06033_ (.I0(\dp.rf.rf[8][23] ),
    .I1(\dp.rf.rf[9][23] ),
    .I2(\dp.rf.rf[12][23] ),
    .I3(\dp.rf.rf[13][23] ),
    .S0(_01121_),
    .S1(_01432_),
    .Z(_01813_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06034_ (.I0(_01812_),
    .I1(_01813_),
    .S(_01372_),
    .Z(_01814_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06035_ (.A1(_01385_),
    .A2(_01814_),
    .Z(_01815_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06036_ (.A1(_01811_),
    .A2(_01815_),
    .B(_01376_),
    .ZN(_01816_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _06037_ (.A1(_01792_),
    .A2(_01796_),
    .A3(_01800_),
    .A4(_01816_),
    .ZN(_01817_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _06038_ (.I(_01817_),
    .Z(_04896_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06039_ (.I(_04896_),
    .ZN(_04900_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06040_ (.A1(_01312_),
    .A2(_01301_),
    .ZN(_01818_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06041_ (.A1(_01299_),
    .A2(_01818_),
    .B(_01304_),
    .ZN(_05166_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _06042_ (.I(_01550_),
    .Z(_01819_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _06043_ (.I(_01657_),
    .Z(_01820_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06044_ (.I0(\dp.rf.rf[16][22] ),
    .I1(\dp.rf.rf[17][22] ),
    .I2(\dp.rf.rf[24][22] ),
    .I3(\dp.rf.rf[25][22] ),
    .S0(_01820_),
    .S1(_01761_),
    .Z(_01821_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06045_ (.A1(_01819_),
    .A2(_01821_),
    .ZN(_01822_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06046_ (.A1(_01408_),
    .A2(_01671_),
    .ZN(_01823_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06047_ (.I0(\dp.rf.rf[26][22] ),
    .I1(\dp.rf.rf[27][22] ),
    .S(_01658_),
    .Z(_01824_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06048_ (.I0(\dp.rf.rf[18][22] ),
    .I1(\dp.rf.rf[19][22] ),
    .S(_01657_),
    .Z(_01825_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _06049_ (.A1(_01766_),
    .A2(_01763_),
    .A3(_01825_),
    .Z(_01826_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _06050_ (.A1(_01823_),
    .A2(_01824_),
    .B(_01826_),
    .C(_01779_),
    .ZN(_01827_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _06051_ (.A1(_01058_),
    .A2(_01822_),
    .A3(_01827_),
    .Z(_01828_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06052_ (.I0(\dp.rf.rf[6][22] ),
    .I1(\dp.rf.rf[7][22] ),
    .I2(\dp.rf.rf[14][22] ),
    .I3(\dp.rf.rf[15][22] ),
    .S0(_01609_),
    .S1(_01763_),
    .Z(_01829_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06053_ (.I0(\dp.rf.rf[4][22] ),
    .I1(\dp.rf.rf[5][22] ),
    .I2(\dp.rf.rf[12][22] ),
    .I3(\dp.rf.rf[13][22] ),
    .S0(_01609_),
    .S1(_01763_),
    .Z(_01830_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06054_ (.I0(_01829_),
    .I1(_01830_),
    .S(_01766_),
    .Z(_01831_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _06055_ (.A1(_01058_),
    .A2(_01312_),
    .A3(_01831_),
    .ZN(_01832_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06056_ (.I0(\dp.rf.rf[28][22] ),
    .I1(\dp.rf.rf[29][22] ),
    .I2(\dp.rf.rf[30][22] ),
    .I3(\dp.rf.rf[31][22] ),
    .S0(_01261_),
    .S1(_01263_),
    .Z(_01833_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06057_ (.I0(\dp.rf.rf[20][22] ),
    .I1(\dp.rf.rf[21][22] ),
    .I2(\dp.rf.rf[22][22] ),
    .I3(\dp.rf.rf[23][22] ),
    .S0(_01261_),
    .S1(_01263_),
    .Z(_01834_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06058_ (.I0(_01833_),
    .I1(_01834_),
    .S(_01272_),
    .Z(_01835_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06059_ (.A1(_01669_),
    .A2(_01061_),
    .Z(_01836_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06060_ (.I0(\dp.rf.rf[2][22] ),
    .I1(\dp.rf.rf[3][22] ),
    .I2(\dp.rf.rf[10][22] ),
    .I3(\dp.rf.rf[11][22] ),
    .S0(_01275_),
    .S1(_01763_),
    .Z(_01837_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06061_ (.I0(\dp.rf.rf[0][22] ),
    .I1(\dp.rf.rf[1][22] ),
    .I2(\dp.rf.rf[8][22] ),
    .I3(\dp.rf.rf[9][22] ),
    .S0(_01279_),
    .S1(_01763_),
    .Z(_01838_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06062_ (.I0(_01837_),
    .I1(_01838_),
    .S(_01766_),
    .Z(_01839_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06063_ (.A1(net213),
    .A2(_01835_),
    .B1(_01836_),
    .B2(_01839_),
    .ZN(_01840_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _06064_ (.A1(_01828_),
    .A2(_01832_),
    .A3(_01840_),
    .Z(_01841_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06065_ (.A1(_01546_),
    .A2(_01841_),
    .ZN(_01842_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06066_ (.A1(_01290_),
    .A2(_05166_),
    .B(_01842_),
    .ZN(_01843_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06067_ (.A1(_01288_),
    .A2(_01843_),
    .Z(_04905_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06068_ (.I(_04905_),
    .ZN(_04909_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06069_ (.I0(\dp.rf.rf[14][22] ),
    .I1(\dp.rf.rf[15][22] ),
    .S(_01186_),
    .Z(_01844_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06070_ (.I(_01844_),
    .ZN(_01845_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06071_ (.A1(_01578_),
    .A2(_01845_),
    .B(_01151_),
    .ZN(_01846_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _06072_ (.A1(_01154_),
    .A2(_01155_),
    .A3(_01034_),
    .A4(\dp.rf.rf[10][22] ),
    .ZN(_01847_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06073_ (.I(\dp.rf.rf[10][22] ),
    .ZN(_01848_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _06074_ (.A1(_01028_),
    .A2(_01153_),
    .A3(_01847_),
    .B1(_01848_),
    .B2(_01582_),
    .ZN(_01849_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06075_ (.A1(\dp.rf.rf[11][22] ),
    .A2(_01531_),
    .Z(_01850_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _06076_ (.A1(_01163_),
    .A2(_01165_),
    .A3(_01849_),
    .A4(_01850_),
    .Z(_01851_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06077_ (.I0(\dp.rf.rf[8][22] ),
    .I1(\dp.rf.rf[9][22] ),
    .I2(\dp.rf.rf[12][22] ),
    .I3(\dp.rf.rf[13][22] ),
    .S0(_01520_),
    .S1(_01364_),
    .Z(_01852_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _06078_ (.A1(_01846_),
    .A2(_01851_),
    .B1(_01852_),
    .B2(_01506_),
    .C(_01199_),
    .ZN(_01853_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _06079_ (.I(_01360_),
    .Z(_01854_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06080_ (.I0(\dp.rf.rf[2][22] ),
    .I1(\dp.rf.rf[3][22] ),
    .I2(\dp.rf.rf[6][22] ),
    .I3(\dp.rf.rf[7][22] ),
    .S0(_01238_),
    .S1(_01209_),
    .Z(_01855_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06081_ (.A1(_01529_),
    .A2(_01855_),
    .ZN(_01856_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06082_ (.I0(\dp.rf.rf[1][22] ),
    .I1(\dp.rf.rf[5][22] ),
    .S(_01123_),
    .Z(_01857_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06083_ (.A1(\dp.rf.rf[4][22] ),
    .A2(_01496_),
    .B1(_01857_),
    .B2(_01328_),
    .C(_01241_),
    .ZN(_01858_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _06084_ (.A1(_01854_),
    .A2(_01856_),
    .A3(_01858_),
    .Z(_01859_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06085_ (.I0(\dp.rf.rf[24][22] ),
    .I1(\dp.rf.rf[25][22] ),
    .I2(\dp.rf.rf[28][22] ),
    .I3(\dp.rf.rf[29][22] ),
    .S0(_01600_),
    .S1(_01210_),
    .Z(_01860_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06086_ (.I0(\dp.rf.rf[26][22] ),
    .I1(\dp.rf.rf[27][22] ),
    .S(_01147_),
    .Z(_01861_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06087_ (.I(_01861_),
    .ZN(_01862_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06088_ (.I0(\dp.rf.rf[30][22] ),
    .I1(\dp.rf.rf[31][22] ),
    .S(_01238_),
    .Z(_01863_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06089_ (.A1(_01182_),
    .A2(_01863_),
    .B(_01213_),
    .ZN(_01864_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06090_ (.A1(_01224_),
    .A2(_01862_),
    .B(_01864_),
    .ZN(_01865_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _06091_ (.A1(_01576_),
    .A2(_01860_),
    .B(_01865_),
    .C(_01237_),
    .ZN(_01866_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06092_ (.I0(\dp.rf.rf[18][22] ),
    .I1(\dp.rf.rf[19][22] ),
    .I2(\dp.rf.rf[22][22] ),
    .I3(\dp.rf.rf[23][22] ),
    .S0(_01531_),
    .S1(_01443_),
    .Z(_01867_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06093_ (.I0(\dp.rf.rf[16][22] ),
    .I1(\dp.rf.rf[17][22] ),
    .I2(\dp.rf.rf[20][22] ),
    .I3(\dp.rf.rf[21][22] ),
    .S0(_01531_),
    .S1(_01443_),
    .Z(_01868_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06094_ (.I0(_01867_),
    .I1(_01868_),
    .S(_01172_),
    .Z(_01869_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06095_ (.A1(_01178_),
    .A2(_01869_),
    .B(net205),
    .ZN(_01870_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _06096_ (.A1(_01589_),
    .A2(_01853_),
    .A3(_01859_),
    .B1(_01866_),
    .B2(_01870_),
    .ZN(_01871_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _06097_ (.I(_01871_),
    .Z(_04904_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06098_ (.I(_04904_),
    .ZN(_04908_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06099_ (.A1(_01819_),
    .A2(_01301_),
    .ZN(_01872_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06100_ (.A1(_01299_),
    .A2(_01872_),
    .B(_01304_),
    .ZN(_05162_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06101_ (.I0(\dp.rf.rf[28][21] ),
    .I1(\dp.rf.rf[29][21] ),
    .I2(\dp.rf.rf[30][21] ),
    .I3(\dp.rf.rf[31][21] ),
    .S0(_01267_),
    .S1(_01263_),
    .Z(_01873_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06102_ (.I0(\dp.rf.rf[20][21] ),
    .I1(\dp.rf.rf[21][21] ),
    .I2(\dp.rf.rf[22][21] ),
    .I3(\dp.rf.rf[23][21] ),
    .S0(_01267_),
    .S1(_01263_),
    .Z(_01874_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06103_ (.I0(\dp.rf.rf[24][21] ),
    .I1(\dp.rf.rf[25][21] ),
    .I2(\dp.rf.rf[26][21] ),
    .I3(\dp.rf.rf[27][21] ),
    .S0(_01275_),
    .S1(_01268_),
    .Z(_01875_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06104_ (.I0(\dp.rf.rf[16][21] ),
    .I1(\dp.rf.rf[17][21] ),
    .I2(\dp.rf.rf[18][21] ),
    .I3(\dp.rf.rf[19][21] ),
    .S0(_01267_),
    .S1(_01263_),
    .Z(_01876_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06105_ (.I0(_01873_),
    .I1(_01874_),
    .I2(_01875_),
    .I3(_01876_),
    .S0(_01282_),
    .S1(_01669_),
    .Z(_01877_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06106_ (.I0(\dp.rf.rf[4][21] ),
    .I1(\dp.rf.rf[5][21] ),
    .I2(\dp.rf.rf[6][21] ),
    .I3(\dp.rf.rf[7][21] ),
    .S0(_01261_),
    .S1(_01561_),
    .Z(_01878_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06107_ (.I0(\dp.rf.rf[0][21] ),
    .I1(\dp.rf.rf[1][21] ),
    .I2(\dp.rf.rf[2][21] ),
    .I3(\dp.rf.rf[3][21] ),
    .S0(_01261_),
    .S1(_01263_),
    .Z(_01879_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06108_ (.I0(_01878_),
    .I1(_01879_),
    .S(_01779_),
    .Z(_01880_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06109_ (.I0(\dp.rf.rf[12][21] ),
    .I1(\dp.rf.rf[13][21] ),
    .I2(\dp.rf.rf[14][21] ),
    .I3(\dp.rf.rf[15][21] ),
    .S0(_01059_),
    .S1(_01102_),
    .Z(_01881_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06110_ (.I0(\dp.rf.rf[8][21] ),
    .I1(\dp.rf.rf[9][21] ),
    .I2(\dp.rf.rf[10][21] ),
    .I3(\dp.rf.rf[11][21] ),
    .S0(_01059_),
    .S1(_01102_),
    .Z(_01882_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06111_ (.I0(_01881_),
    .I1(_01882_),
    .S(_01667_),
    .Z(_01883_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _06112_ (.A1(_01672_),
    .A2(_01883_),
    .Z(_01884_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06113_ (.A1(_01607_),
    .A2(_01884_),
    .Z(_01885_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _06114_ (.A1(_01656_),
    .A2(_01877_),
    .B1(_01880_),
    .B2(net223),
    .C(_01885_),
    .ZN(_01886_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06115_ (.A1(_01605_),
    .A2(_01886_),
    .ZN(_01887_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06116_ (.A1(_01605_),
    .A2(_05162_),
    .B(_01887_),
    .ZN(_01888_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06117_ (.A1(_01288_),
    .A2(_01888_),
    .Z(_04913_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06118_ (.I(_04913_),
    .ZN(_04917_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _06119_ (.I(_01193_),
    .Z(_01889_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06120_ (.I0(\dp.rf.rf[8][21] ),
    .I1(\dp.rf.rf[9][21] ),
    .I2(\dp.rf.rf[12][21] ),
    .I3(\dp.rf.rf[13][21] ),
    .S0(_01508_),
    .S1(_01201_),
    .Z(_01890_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06121_ (.I0(\dp.rf.rf[10][21] ),
    .I1(\dp.rf.rf[11][21] ),
    .S(_01427_),
    .Z(_01891_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06122_ (.I(_01891_),
    .ZN(_01892_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06123_ (.I0(\dp.rf.rf[14][21] ),
    .I1(\dp.rf.rf[15][21] ),
    .S(_01202_),
    .Z(_01893_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06124_ (.A1(_01196_),
    .A2(_01893_),
    .B(_01118_),
    .ZN(_01894_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06125_ (.A1(_01344_),
    .A2(_01892_),
    .B(_01894_),
    .ZN(_01895_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _06126_ (.A1(_01889_),
    .A2(_01890_),
    .B(_01895_),
    .C(_01199_),
    .ZN(_01896_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06127_ (.I0(\dp.rf.rf[2][21] ),
    .I1(\dp.rf.rf[3][21] ),
    .I2(\dp.rf.rf[6][21] ),
    .I3(\dp.rf.rf[7][21] ),
    .S0(_01135_),
    .S1(_01369_),
    .Z(_01897_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06128_ (.A1(_01213_),
    .A2(_01897_),
    .ZN(_01898_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06129_ (.I0(\dp.rf.rf[1][21] ),
    .I1(\dp.rf.rf[5][21] ),
    .S(_01248_),
    .Z(_01899_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06130_ (.A1(\dp.rf.rf[4][21] ),
    .A2(_01367_),
    .B1(_01899_),
    .B2(_01190_),
    .C(_01193_),
    .ZN(_01900_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _06131_ (.A1(_01854_),
    .A2(_01898_),
    .A3(_01900_),
    .Z(_01901_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06132_ (.I0(\dp.rf.rf[18][21] ),
    .I1(\dp.rf.rf[19][21] ),
    .I2(\dp.rf.rf[22][21] ),
    .I3(\dp.rf.rf[23][21] ),
    .S0(_01238_),
    .S1(_01457_),
    .Z(_01902_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06133_ (.I0(\dp.rf.rf[16][21] ),
    .I1(\dp.rf.rf[17][21] ),
    .I2(\dp.rf.rf[20][21] ),
    .I3(\dp.rf.rf[21][21] ),
    .S0(_01238_),
    .S1(_01457_),
    .Z(_01903_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06134_ (.I0(_01902_),
    .I1(_01903_),
    .S(_01241_),
    .Z(_01904_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06135_ (.A1(_01178_),
    .A2(_01904_),
    .B(_01511_),
    .ZN(_01905_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06136_ (.I0(\dp.rf.rf[30][21] ),
    .I1(\dp.rf.rf[31][21] ),
    .S(_01120_),
    .Z(_01906_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _06137_ (.A1(_01162_),
    .A2(_01906_),
    .Z(_01907_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _06138_ (.A1(_01529_),
    .A2(_01244_),
    .A3(_01192_),
    .A4(_01907_),
    .Z(_01908_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _06139_ (.A1(_01154_),
    .A2(_01155_),
    .A3(_01034_),
    .A4(\dp.rf.rf[26][21] ),
    .ZN(_01909_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06140_ (.I(\dp.rf.rf[26][21] ),
    .ZN(_01910_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _06141_ (.A1(_01028_),
    .A2(_01153_),
    .A3(_01909_),
    .B1(_01910_),
    .B2(_01428_),
    .ZN(_01911_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06142_ (.A1(\dp.rf.rf[27][21] ),
    .A2(_01520_),
    .Z(_01912_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _06143_ (.A1(_01164_),
    .A2(_01166_),
    .A3(_01911_),
    .A4(_01912_),
    .Z(_01913_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06144_ (.I0(\dp.rf.rf[24][21] ),
    .I1(\dp.rf.rf[25][21] ),
    .I2(\dp.rf.rf[28][21] ),
    .I3(\dp.rf.rf[29][21] ),
    .S0(_01120_),
    .S1(_01248_),
    .Z(_01914_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _06145_ (.A1(_01171_),
    .A2(net9),
    .A3(_01914_),
    .Z(_01915_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _06146_ (.A1(_01175_),
    .A2(_01915_),
    .Z(_01916_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06147_ (.A1(_01908_),
    .A2(_01913_),
    .B1(_01916_),
    .B2(_01244_),
    .ZN(_01917_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _06148_ (.A1(net191),
    .A2(_01896_),
    .A3(_01901_),
    .B1(_01905_),
    .B2(_01917_),
    .ZN(_01918_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _06149_ (.I(_01918_),
    .Z(_04912_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06150_ (.I(_04912_),
    .ZN(_04916_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _06151_ (.I(_01261_),
    .Z(_01919_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06152_ (.A1(_01293_),
    .A2(_01297_),
    .ZN(_01920_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06153_ (.A1(_01919_),
    .A2(_01300_),
    .B(_01920_),
    .ZN(_01921_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _06154_ (.A1(_01303_),
    .A2(_01921_),
    .Z(_01922_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06155_ (.I0(\dp.rf.rf[28][20] ),
    .I1(\dp.rf.rf[29][20] ),
    .I2(\dp.rf.rf[30][20] ),
    .I3(\dp.rf.rf[31][20] ),
    .S0(_01553_),
    .S1(_01555_),
    .Z(_01923_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06156_ (.I0(\dp.rf.rf[20][20] ),
    .I1(\dp.rf.rf[21][20] ),
    .I2(\dp.rf.rf[22][20] ),
    .I3(\dp.rf.rf[23][20] ),
    .S0(_01553_),
    .S1(_01555_),
    .Z(_01924_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06157_ (.I0(\dp.rf.rf[24][20] ),
    .I1(\dp.rf.rf[25][20] ),
    .I2(\dp.rf.rf[26][20] ),
    .I3(\dp.rf.rf[27][20] ),
    .S0(_01609_),
    .S1(_01561_),
    .Z(_01925_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06158_ (.I0(\dp.rf.rf[16][20] ),
    .I1(\dp.rf.rf[17][20] ),
    .I2(\dp.rf.rf[18][20] ),
    .I3(\dp.rf.rf[19][20] ),
    .S0(_01553_),
    .S1(_01555_),
    .Z(_01926_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06159_ (.I0(_01923_),
    .I1(_01924_),
    .I2(_01925_),
    .I3(_01926_),
    .S0(_01272_),
    .S1(_01669_),
    .Z(_01927_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _06160_ (.I(net226),
    .Z(_01928_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _06161_ (.I(_01549_),
    .Z(_01929_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06162_ (.I0(\dp.rf.rf[4][20] ),
    .I1(\dp.rf.rf[5][20] ),
    .I2(\dp.rf.rf[6][20] ),
    .I3(\dp.rf.rf[7][20] ),
    .S0(_01928_),
    .S1(_01929_),
    .Z(_01930_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06163_ (.I0(\dp.rf.rf[0][20] ),
    .I1(\dp.rf.rf[1][20] ),
    .I2(\dp.rf.rf[2][20] ),
    .I3(\dp.rf.rf[3][20] ),
    .S0(_01928_),
    .S1(_01929_),
    .Z(_01931_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06164_ (.I0(_01930_),
    .I1(_01931_),
    .S(_01779_),
    .Z(_01932_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06165_ (.I0(\dp.rf.rf[12][20] ),
    .I1(\dp.rf.rf[13][20] ),
    .I2(\dp.rf.rf[14][20] ),
    .I3(\dp.rf.rf[15][20] ),
    .S0(_01059_),
    .S1(_01262_),
    .Z(_01933_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06166_ (.I0(\dp.rf.rf[8][20] ),
    .I1(\dp.rf.rf[9][20] ),
    .I2(\dp.rf.rf[10][20] ),
    .I3(\dp.rf.rf[11][20] ),
    .S0(_01059_),
    .S1(_01262_),
    .Z(_01934_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06167_ (.I0(_01933_),
    .I1(_01934_),
    .S(_01667_),
    .Z(_01935_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _06168_ (.A1(_01672_),
    .A2(_01935_),
    .Z(_01936_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06169_ (.A1(_01607_),
    .A2(_01936_),
    .Z(_01937_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _06170_ (.A1(_01656_),
    .A2(_01927_),
    .B1(_01932_),
    .B2(net224),
    .C(_01937_),
    .ZN(_01938_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06171_ (.I0(_01922_),
    .I1(_01938_),
    .S(_01546_),
    .Z(_01939_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06172_ (.A1(_01086_),
    .A2(_01939_),
    .Z(_04921_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06173_ (.I(_04921_),
    .ZN(_04925_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06174_ (.I0(\dp.rf.rf[26][20] ),
    .I1(\dp.rf.rf[27][20] ),
    .I2(\dp.rf.rf[30][20] ),
    .I3(\dp.rf.rf[31][20] ),
    .S0(_01186_),
    .S1(_01457_),
    .Z(_01940_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06175_ (.I0(\dp.rf.rf[24][20] ),
    .I1(\dp.rf.rf[25][20] ),
    .I2(\dp.rf.rf[28][20] ),
    .I3(\dp.rf.rf[29][20] ),
    .S0(_01186_),
    .S1(_01457_),
    .Z(_01941_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06176_ (.I0(_01940_),
    .I1(_01941_),
    .S(_01193_),
    .Z(_01942_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06177_ (.A1(_01415_),
    .A2(_01942_),
    .ZN(_01943_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06178_ (.I0(\dp.rf.rf[22][20] ),
    .I1(\dp.rf.rf[23][20] ),
    .S(_01225_),
    .Z(_01944_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06179_ (.I(_01944_),
    .ZN(_01945_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06180_ (.A1(_01146_),
    .A2(_01945_),
    .B(_01151_),
    .ZN(_01946_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _06181_ (.A1(_01154_),
    .A2(_01155_),
    .A3(_01034_),
    .A4(\dp.rf.rf[18][20] ),
    .ZN(_01947_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06182_ (.I(\dp.rf.rf[18][20] ),
    .ZN(_01948_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _06183_ (.A1(_01028_),
    .A2(_01153_),
    .A3(_01947_),
    .B1(_01948_),
    .B2(_01160_),
    .ZN(_01949_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06184_ (.A1(\dp.rf.rf[19][20] ),
    .A2(_01582_),
    .Z(_01950_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _06185_ (.A1(_01164_),
    .A2(_01166_),
    .A3(_01949_),
    .A4(_01950_),
    .Z(_01951_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06186_ (.I0(\dp.rf.rf[17][20] ),
    .I1(\dp.rf.rf[21][20] ),
    .S(_01144_),
    .Z(_01952_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06187_ (.A1(_01636_),
    .A2(_01952_),
    .ZN(_01953_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06188_ (.A1(\dp.rf.rf[20][20] ),
    .A2(_01600_),
    .A3(_01196_),
    .B(_01193_),
    .ZN(_01954_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _06189_ (.A1(_01953_),
    .A2(_01954_),
    .B(_01228_),
    .C(net168),
    .ZN(_01955_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06190_ (.I(\dp.rf.rf[16][20] ),
    .ZN(_01956_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06191_ (.A1(_01956_),
    .A2(_01737_),
    .ZN(_01957_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06192_ (.A1(_01946_),
    .A2(_01951_),
    .B1(_01955_),
    .B2(_01957_),
    .ZN(_01958_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06193_ (.I0(\dp.rf.rf[14][20] ),
    .I1(\dp.rf.rf[15][20] ),
    .S(_01135_),
    .Z(_01959_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06194_ (.I(_01959_),
    .ZN(_01960_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06195_ (.A1(_01533_),
    .A2(_01960_),
    .B(net274),
    .ZN(_01961_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _06196_ (.A1(net10),
    .A2(net1),
    .A3(_01034_),
    .A4(\dp.rf.rf[10][20] ),
    .ZN(_01962_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06197_ (.I(\dp.rf.rf[10][20] ),
    .ZN(_01963_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _06198_ (.A1(_01028_),
    .A2(_01153_),
    .A3(_01962_),
    .B1(_01963_),
    .B2(_01147_),
    .ZN(_01964_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06199_ (.A1(\dp.rf.rf[11][20] ),
    .A2(_01179_),
    .Z(_01965_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _06200_ (.A1(_01163_),
    .A2(_01165_),
    .A3(_01964_),
    .A4(_01965_),
    .Z(_01966_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06201_ (.I0(\dp.rf.rf[8][20] ),
    .I1(\dp.rf.rf[9][20] ),
    .I2(\dp.rf.rf[12][20] ),
    .I3(\dp.rf.rf[13][20] ),
    .S0(_01582_),
    .S1(_01124_),
    .Z(_01967_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _06202_ (.A1(_01961_),
    .A2(_01966_),
    .B1(_01967_),
    .B2(_01506_),
    .C(_01199_),
    .ZN(_01968_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06203_ (.I0(\dp.rf.rf[2][20] ),
    .I1(\dp.rf.rf[3][20] ),
    .I2(\dp.rf.rf[6][20] ),
    .I3(\dp.rf.rf[7][20] ),
    .S0(_01186_),
    .S1(_01457_),
    .Z(_01969_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06204_ (.A1(_01529_),
    .A2(_01969_),
    .ZN(_01970_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06205_ (.I0(\dp.rf.rf[1][20] ),
    .I1(\dp.rf.rf[5][20] ),
    .S(_01248_),
    .Z(_01971_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06206_ (.A1(\dp.rf.rf[4][20] ),
    .A2(_01496_),
    .B1(_01971_),
    .B2(_01328_),
    .C(_01193_),
    .ZN(_01972_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _06207_ (.A1(_01854_),
    .A2(_01970_),
    .A3(_01972_),
    .Z(_01973_));
 gf180mcu_fd_sc_mcu9t5v0__oai33_4 _06208_ (.A1(_01455_),
    .A2(_01943_),
    .A3(_01958_),
    .B1(_01968_),
    .B2(_01973_),
    .B3(net191),
    .ZN(_01974_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _06209_ (.I(_01974_),
    .Z(_04920_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06210_ (.I(_04920_),
    .ZN(_04924_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06211_ (.A1(_01178_),
    .A2(_01300_),
    .B1(_01296_),
    .B2(_01244_),
    .ZN(_01975_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06212_ (.A1(_01293_),
    .A2(_01975_),
    .B(_01303_),
    .ZN(_01976_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06213_ (.A1(_01244_),
    .A2(_01300_),
    .ZN(_01977_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06214_ (.A1(_01298_),
    .A2(_01977_),
    .B(_01303_),
    .ZN(_01978_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06215_ (.I0(_01976_),
    .I1(_01978_),
    .S(_01109_),
    .Z(_05154_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06216_ (.I0(\dp.rf.rf[24][19] ),
    .I1(\dp.rf.rf[25][19] ),
    .I2(\dp.rf.rf[26][19] ),
    .I3(\dp.rf.rf[27][19] ),
    .S0(_01773_),
    .S1(_01774_),
    .Z(_01979_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06217_ (.I0(\dp.rf.rf[16][19] ),
    .I1(\dp.rf.rf[17][19] ),
    .I2(\dp.rf.rf[18][19] ),
    .I3(\dp.rf.rf[19][19] ),
    .S0(_01773_),
    .S1(_01774_),
    .Z(_01980_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06218_ (.I0(\dp.rf.rf[28][19] ),
    .I1(\dp.rf.rf[29][19] ),
    .I2(\dp.rf.rf[30][19] ),
    .I3(\dp.rf.rf[31][19] ),
    .S0(_01662_),
    .S1(_01659_),
    .Z(_01981_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06219_ (.I0(\dp.rf.rf[20][19] ),
    .I1(\dp.rf.rf[21][19] ),
    .I2(\dp.rf.rf[22][19] ),
    .I3(\dp.rf.rf[23][19] ),
    .S0(_01662_),
    .S1(_01774_),
    .Z(_01982_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _06220_ (.I0(_01979_),
    .I1(_01980_),
    .I2(_01981_),
    .I3(_01982_),
    .S0(_01666_),
    .S1(_01312_),
    .Z(_01983_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06221_ (.I0(\dp.rf.rf[8][19] ),
    .I1(\dp.rf.rf[9][19] ),
    .I2(\dp.rf.rf[10][19] ),
    .I3(\dp.rf.rf[11][19] ),
    .S0(_01662_),
    .S1(_01659_),
    .Z(_01984_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06222_ (.I0(\dp.rf.rf[0][19] ),
    .I1(\dp.rf.rf[1][19] ),
    .I2(\dp.rf.rf[2][19] ),
    .I3(\dp.rf.rf[3][19] ),
    .S0(_01662_),
    .S1(_01659_),
    .Z(_01985_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06223_ (.I0(\dp.rf.rf[12][19] ),
    .I1(\dp.rf.rf[13][19] ),
    .I2(\dp.rf.rf[14][19] ),
    .I3(\dp.rf.rf[15][19] ),
    .S0(_01662_),
    .S1(_01659_),
    .Z(_01986_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06224_ (.I0(\dp.rf.rf[4][19] ),
    .I1(\dp.rf.rf[5][19] ),
    .I2(\dp.rf.rf[6][19] ),
    .I3(\dp.rf.rf[7][19] ),
    .S0(_01662_),
    .S1(_01659_),
    .Z(_01987_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06225_ (.I0(_01984_),
    .I1(_01985_),
    .I2(_01986_),
    .I3(_01987_),
    .S0(_01666_),
    .S1(_01478_),
    .Z(_01988_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _06226_ (.A1(_01111_),
    .A2(_01983_),
    .B1(_01988_),
    .B2(_01112_),
    .ZN(_01989_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _06227_ (.I(_01989_),
    .ZN(_01990_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06228_ (.I0(_05154_),
    .I1(_01990_),
    .S(_01289_),
    .Z(_01991_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _06229_ (.A1(_01086_),
    .A2(_01991_),
    .ZN(_04929_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06230_ (.I(_04929_),
    .ZN(_04933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06231_ (.A1(\dp.rf.rf[26][19] ),
    .A2(_01571_),
    .ZN(_01992_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06232_ (.A1(\dp.rf.rf[27][19] ),
    .A2(_01429_),
    .B1(_01533_),
    .B2(_01192_),
    .ZN(_01993_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06233_ (.I0(\dp.rf.rf[30][19] ),
    .I1(\dp.rf.rf[31][19] ),
    .S(_01147_),
    .Z(_01994_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _06234_ (.A1(_01230_),
    .A2(_01994_),
    .B(_01192_),
    .C(_01529_),
    .ZN(_01995_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06235_ (.A1(_01992_),
    .A2(_01993_),
    .B(_01995_),
    .ZN(_01996_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06236_ (.I0(\dp.rf.rf[24][19] ),
    .I1(\dp.rf.rf[25][19] ),
    .I2(\dp.rf.rf[28][19] ),
    .I3(\dp.rf.rf[29][19] ),
    .S0(_01508_),
    .S1(_01145_),
    .Z(_01997_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06237_ (.A1(_01889_),
    .A2(_01997_),
    .Z(_01998_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _06238_ (.A1(_01580_),
    .A2(_01996_),
    .A3(_01998_),
    .ZN(_01999_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06239_ (.I0(\dp.rf.rf[22][19] ),
    .I1(\dp.rf.rf[23][19] ),
    .S(_01340_),
    .Z(_02000_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06240_ (.A1(\dp.rf.rf[18][19] ),
    .A2(net204),
    .Z(_02001_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06241_ (.A1(\dp.rf.rf[19][19] ),
    .A2(_01345_),
    .ZN(_02002_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06242_ (.A1(_01344_),
    .A2(_02002_),
    .ZN(_02003_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06243_ (.A1(_01339_),
    .A2(_02000_),
    .B1(_02001_),
    .B2(_02003_),
    .C(_01334_),
    .ZN(_02004_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06244_ (.I(\dp.rf.rf[20][19] ),
    .ZN(_02005_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06245_ (.I0(\dp.rf.rf[17][19] ),
    .I1(\dp.rf.rf[21][19] ),
    .S(_01129_),
    .Z(_02006_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06246_ (.A1(_01190_),
    .A2(_02006_),
    .ZN(_02007_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _06247_ (.A1(_02005_),
    .A2(_01249_),
    .B(_02007_),
    .C(_01353_),
    .ZN(_02008_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _06248_ (.A1(\dp.rf.rf[16][19] ),
    .A2(_01356_),
    .B1(_02008_),
    .B2(net229),
    .ZN(_02009_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06249_ (.A1(_02004_),
    .A2(_02009_),
    .Z(_02010_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06250_ (.I(\dp.rf.rf[0][19] ),
    .ZN(_02011_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _06251_ (.A1(_01438_),
    .A2(_01185_),
    .A3(_01174_),
    .B(_01252_),
    .ZN(_02012_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06252_ (.I0(\dp.rf.rf[1][19] ),
    .I1(\dp.rf.rf[5][19] ),
    .S(_01209_),
    .Z(_02013_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06253_ (.A1(\dp.rf.rf[4][19] ),
    .A2(_01368_),
    .B1(_02013_),
    .B2(_01442_),
    .C(_01506_),
    .ZN(_02014_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06254_ (.A1(_02011_),
    .A2(_02012_),
    .B1(_02014_),
    .B2(_01511_),
    .ZN(_02015_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06255_ (.I0(\dp.rf.rf[2][19] ),
    .I1(\dp.rf.rf[3][19] ),
    .I2(\dp.rf.rf[6][19] ),
    .I3(\dp.rf.rf[7][19] ),
    .S0(_01428_),
    .S1(_01169_),
    .Z(_02016_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06256_ (.A1(_01456_),
    .A2(_02016_),
    .ZN(_02017_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06257_ (.A1(_01415_),
    .A2(_02017_),
    .B(_01245_),
    .ZN(_02018_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _06258_ (.I(net272),
    .Z(_02019_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06259_ (.I0(\dp.rf.rf[14][19] ),
    .I1(\dp.rf.rf[15][19] ),
    .S(_01428_),
    .Z(_02020_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06260_ (.A1(_01339_),
    .A2(_02020_),
    .ZN(_02021_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06261_ (.A1(\dp.rf.rf[11][19] ),
    .A2(_01340_),
    .Z(_02022_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _06262_ (.A1(_01578_),
    .A2(net168),
    .B1(_01626_),
    .B2(\dp.rf.rf[10][19] ),
    .C(_02022_),
    .ZN(_02023_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06263_ (.I0(\dp.rf.rf[8][19] ),
    .I1(\dp.rf.rf[9][19] ),
    .I2(\dp.rf.rf[12][19] ),
    .I3(\dp.rf.rf[13][19] ),
    .S0(_01363_),
    .S1(_01124_),
    .Z(_02024_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06264_ (.A1(_01506_),
    .A2(_02024_),
    .B(_01199_),
    .ZN(_02025_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06265_ (.A1(_02019_),
    .A2(_02021_),
    .A3(_02023_),
    .B(_02025_),
    .ZN(_02026_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _06266_ (.A1(_02015_),
    .A2(_02018_),
    .B(_02026_),
    .C(_01376_),
    .ZN(_02027_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _06267_ (.A1(_01455_),
    .A2(_01999_),
    .A3(_02010_),
    .B(_02027_),
    .ZN(_04928_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _06268_ (.I(_04928_),
    .ZN(_04932_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06269_ (.A1(_01211_),
    .A2(_01300_),
    .B1(_01296_),
    .B2(_01178_),
    .ZN(_02028_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06270_ (.A1(_01293_),
    .A2(_02028_),
    .B(_01303_),
    .ZN(_02029_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _06271_ (.A1(_01063_),
    .A2(_01108_),
    .A3(_01088_),
    .A4(net22),
    .ZN(_02030_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06272_ (.I0(_01976_),
    .I1(_02029_),
    .S(net241),
    .Z(_05150_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06273_ (.I(_05150_),
    .ZN(_02031_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _06274_ (.I(_01279_),
    .Z(_02032_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06275_ (.I0(\dp.rf.rf[18][18] ),
    .I1(\dp.rf.rf[19][18] ),
    .S(_02032_),
    .Z(_02033_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06276_ (.I0(\dp.rf.rf[16][18] ),
    .I1(\dp.rf.rf[17][18] ),
    .S(_02032_),
    .Z(_02034_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06277_ (.I0(\dp.rf.rf[26][18] ),
    .I1(\dp.rf.rf[27][18] ),
    .S(_01773_),
    .Z(_02035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06278_ (.I0(\dp.rf.rf[24][18] ),
    .I1(\dp.rf.rf[25][18] ),
    .S(_02032_),
    .Z(_02036_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06279_ (.I0(_02033_),
    .I1(_02034_),
    .I2(_02035_),
    .I3(_02036_),
    .S0(_01766_),
    .S1(_01761_),
    .Z(_02037_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06280_ (.A1(_01780_),
    .A2(_02037_),
    .ZN(_02038_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06281_ (.I0(\dp.rf.rf[12][18] ),
    .I1(\dp.rf.rf[13][18] ),
    .I2(\dp.rf.rf[14][18] ),
    .I3(\dp.rf.rf[15][18] ),
    .S0(_01773_),
    .S1(_01317_),
    .Z(_02039_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06282_ (.I0(\dp.rf.rf[4][18] ),
    .I1(\dp.rf.rf[5][18] ),
    .I2(\dp.rf.rf[6][18] ),
    .I3(\dp.rf.rf[7][18] ),
    .S0(_01773_),
    .S1(_01317_),
    .Z(_02040_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06283_ (.I0(_02039_),
    .I1(_02040_),
    .S(_01311_),
    .Z(_02041_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _06284_ (.A1(_01656_),
    .A2(_01312_),
    .A3(_02041_),
    .ZN(_02042_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06285_ (.I0(\dp.rf.rf[28][18] ),
    .I1(\dp.rf.rf[29][18] ),
    .I2(\dp.rf.rf[30][18] ),
    .I3(\dp.rf.rf[31][18] ),
    .S0(_01773_),
    .S1(_01774_),
    .Z(_02043_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06286_ (.I0(\dp.rf.rf[20][18] ),
    .I1(\dp.rf.rf[21][18] ),
    .I2(\dp.rf.rf[22][18] ),
    .I3(\dp.rf.rf[23][18] ),
    .S0(_01773_),
    .S1(_01774_),
    .Z(_02044_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06287_ (.I0(_02043_),
    .I1(_02044_),
    .S(_01311_),
    .Z(_02045_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06288_ (.I0(\dp.rf.rf[8][18] ),
    .I1(\dp.rf.rf[9][18] ),
    .I2(\dp.rf.rf[10][18] ),
    .I3(\dp.rf.rf[11][18] ),
    .S0(_01662_),
    .S1(_01774_),
    .Z(_02046_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06289_ (.I0(\dp.rf.rf[0][18] ),
    .I1(\dp.rf.rf[1][18] ),
    .I2(\dp.rf.rf[2][18] ),
    .I3(\dp.rf.rf[3][18] ),
    .S0(_01662_),
    .S1(_01774_),
    .Z(_02047_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06290_ (.I0(_02046_),
    .I1(_02047_),
    .S(_01666_),
    .Z(_02048_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06291_ (.A1(net215),
    .A2(_02045_),
    .B1(_02048_),
    .B2(_01836_),
    .ZN(_02049_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _06292_ (.A1(_02038_),
    .A2(_02042_),
    .A3(_02049_),
    .Z(_02050_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06293_ (.I0(_02031_),
    .I1(_02050_),
    .S(_01546_),
    .Z(_02051_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06294_ (.A1(_01086_),
    .A2(_02051_),
    .Z(_04937_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06295_ (.I(_04937_),
    .ZN(_04941_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06296_ (.A1(\dp.rf.rf[2][18] ),
    .A2(_01353_),
    .Z(_02052_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _06297_ (.A1(_01355_),
    .A2(_02052_),
    .Z(_02053_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06298_ (.A1(net206),
    .A2(_02053_),
    .B(\dp.rf.rf[0][18] ),
    .ZN(_02054_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06299_ (.I0(\dp.rf.rf[10][18] ),
    .I1(\dp.rf.rf[11][18] ),
    .I2(\dp.rf.rf[14][18] ),
    .I3(\dp.rf.rf[15][18] ),
    .S0(_01531_),
    .S1(_01443_),
    .Z(_02055_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06300_ (.I0(\dp.rf.rf[8][18] ),
    .I1(\dp.rf.rf[9][18] ),
    .I2(\dp.rf.rf[12][18] ),
    .I3(\dp.rf.rf[13][18] ),
    .S0(_01531_),
    .S1(_01443_),
    .Z(_02056_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06301_ (.I0(_02055_),
    .I1(_02056_),
    .S(_01172_),
    .Z(_02057_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06302_ (.A1(_01237_),
    .A2(_02057_),
    .ZN(_02058_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06303_ (.I0(\dp.rf.rf[2][18] ),
    .I1(\dp.rf.rf[3][18] ),
    .I2(\dp.rf.rf[6][18] ),
    .I3(\dp.rf.rf[7][18] ),
    .S0(_01147_),
    .S1(_01432_),
    .Z(_02059_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06304_ (.A1(_01416_),
    .A2(_02059_),
    .ZN(_02060_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06305_ (.I0(\dp.rf.rf[1][18] ),
    .I1(\dp.rf.rf[5][18] ),
    .S(_01168_),
    .Z(_02061_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06306_ (.A1(\dp.rf.rf[4][18] ),
    .A2(_01368_),
    .B1(_02061_),
    .B2(_01371_),
    .C(_01172_),
    .ZN(_02062_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _06307_ (.A1(_01854_),
    .A2(_02060_),
    .A3(_02062_),
    .Z(_02063_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _06308_ (.A1(_01589_),
    .A2(_02054_),
    .A3(_02058_),
    .A4(_02063_),
    .Z(_02064_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06309_ (.A1(\dp.rf.rf[18][18] ),
    .A2(_01571_),
    .ZN(_02065_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06310_ (.A1(\dp.rf.rf[19][18] ),
    .A2(_01504_),
    .B1(_01211_),
    .B2(_01511_),
    .ZN(_02066_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06311_ (.I0(\dp.rf.rf[22][18] ),
    .I1(\dp.rf.rf[23][18] ),
    .S(_01645_),
    .Z(_02067_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06312_ (.A1(_01568_),
    .A2(_02067_),
    .ZN(_02068_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _06313_ (.A1(_02065_),
    .A2(_02066_),
    .B(_02019_),
    .C(_02068_),
    .ZN(_02069_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06314_ (.I(\dp.rf.rf[16][18] ),
    .ZN(_02070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06315_ (.I0(\dp.rf.rf[17][18] ),
    .I1(\dp.rf.rf[21][18] ),
    .S(_01201_),
    .Z(_02071_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06316_ (.A1(\dp.rf.rf[20][18] ),
    .A2(_01497_),
    .B1(_02071_),
    .B2(_01693_),
    .C(_01173_),
    .ZN(_02072_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06317_ (.A1(_02070_),
    .A2(_01737_),
    .B1(_02072_),
    .B2(_01361_),
    .ZN(_02073_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06318_ (.A1(\dp.rf.rf[27][18] ),
    .A2(_01569_),
    .Z(_02074_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _06319_ (.A1(_01211_),
    .A2(_01511_),
    .B1(_01571_),
    .B2(\dp.rf.rf[26][18] ),
    .C(_02074_),
    .ZN(_02075_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06320_ (.I0(\dp.rf.rf[30][18] ),
    .I1(\dp.rf.rf[31][18] ),
    .S(_01645_),
    .Z(_02076_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _06321_ (.A1(_01568_),
    .A2(_02076_),
    .B(_01511_),
    .C(_01456_),
    .ZN(_02077_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06322_ (.I0(\dp.rf.rf[24][18] ),
    .I1(\dp.rf.rf[25][18] ),
    .I2(\dp.rf.rf[28][18] ),
    .I3(\dp.rf.rf[29][18] ),
    .S0(_01345_),
    .S1(_01210_),
    .Z(_02078_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06323_ (.A1(_01576_),
    .A2(_02078_),
    .B(_01237_),
    .ZN(_02079_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06324_ (.A1(_02075_),
    .A2(_02077_),
    .B(_02079_),
    .ZN(_02080_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _06325_ (.A1(_02069_),
    .A2(_02073_),
    .B(net205),
    .C(_02080_),
    .ZN(_02081_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _06326_ (.A1(_02064_),
    .A2(_02081_),
    .ZN(_04936_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _06327_ (.I(_04936_),
    .ZN(_04940_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06328_ (.A1(_01530_),
    .A2(_01300_),
    .B1(_01296_),
    .B2(_01211_),
    .ZN(_02082_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06329_ (.A1(_01293_),
    .A2(_02082_),
    .B(_01303_),
    .ZN(_02083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06330_ (.I0(_02029_),
    .I1(_02083_),
    .S(net240),
    .Z(_05146_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06331_ (.I(_05146_),
    .ZN(_02084_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06332_ (.I0(\dp.rf.rf[24][17] ),
    .I1(\dp.rf.rf[25][17] ),
    .I2(\dp.rf.rf[26][17] ),
    .I3(\dp.rf.rf[27][17] ),
    .S0(_01919_),
    .S1(_01819_),
    .Z(_02085_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06333_ (.I0(\dp.rf.rf[16][17] ),
    .I1(\dp.rf.rf[17][17] ),
    .I2(\dp.rf.rf[18][17] ),
    .I3(\dp.rf.rf[19][17] ),
    .S0(_01919_),
    .S1(_01819_),
    .Z(_02086_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06334_ (.I0(\dp.rf.rf[28][17] ),
    .I1(\dp.rf.rf[29][17] ),
    .I2(\dp.rf.rf[30][17] ),
    .I3(\dp.rf.rf[31][17] ),
    .S0(_01919_),
    .S1(_01819_),
    .Z(_02087_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06335_ (.I0(\dp.rf.rf[20][17] ),
    .I1(\dp.rf.rf[21][17] ),
    .I2(\dp.rf.rf[22][17] ),
    .I3(\dp.rf.rf[23][17] ),
    .S0(_01919_),
    .S1(_01819_),
    .Z(_02088_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _06336_ (.I0(_02085_),
    .I1(_02086_),
    .I2(_02087_),
    .I3(_02088_),
    .S0(_01311_),
    .S1(_01312_),
    .Z(_02089_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06337_ (.I0(\dp.rf.rf[8][17] ),
    .I1(\dp.rf.rf[9][17] ),
    .I2(\dp.rf.rf[10][17] ),
    .I3(\dp.rf.rf[11][17] ),
    .S0(_01919_),
    .S1(_01819_),
    .Z(_02090_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06338_ (.I0(\dp.rf.rf[0][17] ),
    .I1(\dp.rf.rf[1][17] ),
    .I2(\dp.rf.rf[2][17] ),
    .I3(\dp.rf.rf[3][17] ),
    .S0(_01919_),
    .S1(_01819_),
    .Z(_02091_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06339_ (.I0(\dp.rf.rf[12][17] ),
    .I1(\dp.rf.rf[13][17] ),
    .I2(\dp.rf.rf[14][17] ),
    .I3(\dp.rf.rf[15][17] ),
    .S0(_01919_),
    .S1(_01306_),
    .Z(_02092_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06340_ (.I0(\dp.rf.rf[4][17] ),
    .I1(\dp.rf.rf[5][17] ),
    .I2(\dp.rf.rf[6][17] ),
    .I3(\dp.rf.rf[7][17] ),
    .S0(_01919_),
    .S1(_01819_),
    .Z(_02093_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06341_ (.I0(_02090_),
    .I1(_02091_),
    .I2(_02092_),
    .I3(_02093_),
    .S0(_01311_),
    .S1(_01312_),
    .Z(_02094_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _06342_ (.A1(_01111_),
    .A2(_02089_),
    .B1(_02094_),
    .B2(_01112_),
    .ZN(_02095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06343_ (.I0(_02084_),
    .I1(_02095_),
    .S(_01546_),
    .Z(_02096_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06344_ (.A1(_01086_),
    .A2(_02096_),
    .Z(_04945_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06345_ (.I(_04945_),
    .ZN(_04949_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06346_ (.I0(\dp.rf.rf[30][17] ),
    .I1(\dp.rf.rf[31][17] ),
    .S(_01532_),
    .Z(_02097_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06347_ (.A1(\dp.rf.rf[26][17] ),
    .A2(_01626_),
    .Z(_02098_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06348_ (.A1(\dp.rf.rf[27][17] ),
    .A2(_01569_),
    .ZN(_02099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06349_ (.A1(_01224_),
    .A2(_02099_),
    .ZN(_02100_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _06350_ (.A1(_01568_),
    .A2(_02097_),
    .B1(_02098_),
    .B2(_02100_),
    .C(_01335_),
    .ZN(_02101_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06351_ (.I0(\dp.rf.rf[24][17] ),
    .I1(\dp.rf.rf[25][17] ),
    .I2(\dp.rf.rf[28][17] ),
    .I3(\dp.rf.rf[29][17] ),
    .S0(_01345_),
    .S1(_01458_),
    .Z(_02102_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06352_ (.A1(_01500_),
    .A2(_02102_),
    .B(_01237_),
    .ZN(_02103_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06353_ (.I0(\dp.rf.rf[18][17] ),
    .I1(\dp.rf.rf[19][17] ),
    .I2(\dp.rf.rf[22][17] ),
    .I3(\dp.rf.rf[23][17] ),
    .S0(_01135_),
    .S1(_01369_),
    .Z(_02104_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06354_ (.I0(\dp.rf.rf[16][17] ),
    .I1(\dp.rf.rf[17][17] ),
    .I2(\dp.rf.rf[20][17] ),
    .I3(\dp.rf.rf[21][17] ),
    .S0(_01135_),
    .S1(_01369_),
    .Z(_02105_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06355_ (.I0(_02104_),
    .I1(_02105_),
    .S(_01193_),
    .Z(_02106_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06356_ (.A1(_01178_),
    .A2(_02106_),
    .ZN(_02107_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _06357_ (.A1(_02103_),
    .A2(_02101_),
    .B(_01455_),
    .C(_02107_),
    .ZN(_02108_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06358_ (.I0(\dp.rf.rf[2][17] ),
    .I1(\dp.rf.rf[3][17] ),
    .I2(\dp.rf.rf[6][17] ),
    .I3(\dp.rf.rf[7][17] ),
    .S0(_01238_),
    .S1(_01209_),
    .Z(_02109_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06359_ (.I(_02109_),
    .ZN(_02110_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06360_ (.I0(\dp.rf.rf[1][17] ),
    .I1(\dp.rf.rf[5][17] ),
    .S(_01200_),
    .Z(_02111_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _06361_ (.A1(\dp.rf.rf[4][17] ),
    .A2(_01496_),
    .B1(_02111_),
    .B2(_01328_),
    .ZN(_02112_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06362_ (.I0(_02110_),
    .I1(_02112_),
    .S(_01430_),
    .Z(_02113_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06363_ (.I0(\dp.rf.rf[14][17] ),
    .I1(\dp.rf.rf[15][17] ),
    .S(_01157_),
    .Z(_02114_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06364_ (.A1(\dp.rf.rf[10][17] ),
    .A2(net202),
    .Z(_02115_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06365_ (.A1(\dp.rf.rf[11][17] ),
    .A2(_01532_),
    .ZN(_02116_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06366_ (.A1(_01344_),
    .A2(_02116_),
    .ZN(_02117_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _06367_ (.A1(_01339_),
    .A2(_02114_),
    .B1(_02115_),
    .B2(_02117_),
    .C(_01334_),
    .ZN(_02118_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06368_ (.I0(\dp.rf.rf[8][17] ),
    .I1(\dp.rf.rf[9][17] ),
    .I2(\dp.rf.rf[12][17] ),
    .I3(\dp.rf.rf[13][17] ),
    .S0(_01340_),
    .S1(_01169_),
    .Z(_02119_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06369_ (.A1(_01889_),
    .A2(_02119_),
    .B(_01176_),
    .ZN(_02120_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _06370_ (.A1(_01361_),
    .A2(_02113_),
    .B1(_02118_),
    .B2(_02120_),
    .C(net189),
    .ZN(_02121_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _06371_ (.A1(_02108_),
    .A2(_02121_),
    .Z(_02122_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _06372_ (.I(_02122_),
    .Z(_04944_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _06373_ (.I(_04944_),
    .ZN(_04948_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06374_ (.A1(_01504_),
    .A2(_01300_),
    .B1(_01296_),
    .B2(_01530_),
    .ZN(_02123_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06375_ (.A1(_01293_),
    .A2(_02123_),
    .B(_01303_),
    .ZN(_02124_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06376_ (.I0(_02083_),
    .I1(_02124_),
    .S(net240),
    .Z(_05142_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06377_ (.I(_05142_),
    .ZN(_02125_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06378_ (.I0(\dp.rf.rf[28][16] ),
    .I1(\dp.rf.rf[29][16] ),
    .I2(\dp.rf.rf[30][16] ),
    .I3(\dp.rf.rf[31][16] ),
    .S0(_02032_),
    .S1(_01317_),
    .Z(_02126_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06379_ (.I0(\dp.rf.rf[20][16] ),
    .I1(\dp.rf.rf[21][16] ),
    .I2(\dp.rf.rf[22][16] ),
    .I3(\dp.rf.rf[23][16] ),
    .S0(_02032_),
    .S1(_01317_),
    .Z(_02127_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06380_ (.I0(\dp.rf.rf[24][16] ),
    .I1(\dp.rf.rf[25][16] ),
    .I2(\dp.rf.rf[26][16] ),
    .I3(\dp.rf.rf[27][16] ),
    .S0(_02032_),
    .S1(_01317_),
    .Z(_02128_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06381_ (.I0(\dp.rf.rf[16][16] ),
    .I1(\dp.rf.rf[17][16] ),
    .I2(\dp.rf.rf[18][16] ),
    .I3(\dp.rf.rf[19][16] ),
    .S0(_02032_),
    .S1(_01317_),
    .Z(_02129_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06382_ (.I0(_02126_),
    .I1(_02127_),
    .I2(_02128_),
    .I3(_02129_),
    .S0(_01311_),
    .S1(_01669_),
    .Z(_02130_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06383_ (.I0(\dp.rf.rf[12][16] ),
    .I1(\dp.rf.rf[13][16] ),
    .I2(\dp.rf.rf[14][16] ),
    .I3(\dp.rf.rf[15][16] ),
    .S0(_01305_),
    .S1(_01306_),
    .Z(_02131_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06384_ (.I0(\dp.rf.rf[8][16] ),
    .I1(\dp.rf.rf[9][16] ),
    .I2(\dp.rf.rf[10][16] ),
    .I3(\dp.rf.rf[11][16] ),
    .S0(_01305_),
    .S1(_01306_),
    .Z(_02132_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06385_ (.I0(_02131_),
    .I1(_02132_),
    .S(_01669_),
    .Z(_02133_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06386_ (.I0(\dp.rf.rf[4][16] ),
    .I1(\dp.rf.rf[5][16] ),
    .I2(\dp.rf.rf[6][16] ),
    .I3(\dp.rf.rf[7][16] ),
    .S0(_01484_),
    .S1(_01485_),
    .Z(_02134_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06387_ (.I0(\dp.rf.rf[0][16] ),
    .I1(\dp.rf.rf[1][16] ),
    .I2(\dp.rf.rf[2][16] ),
    .I3(\dp.rf.rf[3][16] ),
    .S0(_01484_),
    .S1(_01485_),
    .Z(_02135_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06388_ (.I0(_02134_),
    .I1(_02135_),
    .S(_01779_),
    .Z(_02136_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _06389_ (.A1(net223),
    .A2(_02136_),
    .Z(_02137_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06390_ (.A1(_01608_),
    .A2(_02137_),
    .Z(_02138_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _06391_ (.A1(_01656_),
    .A2(_02130_),
    .B1(_02133_),
    .B2(_01672_),
    .C(_02138_),
    .ZN(_02139_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06392_ (.I0(_02125_),
    .I1(_02139_),
    .S(_01546_),
    .Z(_02140_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06393_ (.A1(_01086_),
    .A2(_02140_),
    .Z(_04953_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06394_ (.I(_04953_),
    .ZN(_04957_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06395_ (.I0(\dp.rf.rf[26][16] ),
    .I1(\dp.rf.rf[27][16] ),
    .I2(\dp.rf.rf[30][16] ),
    .I3(\dp.rf.rf[31][16] ),
    .S0(_01157_),
    .S1(_01458_),
    .Z(_02141_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06396_ (.I0(\dp.rf.rf[24][16] ),
    .I1(\dp.rf.rf[25][16] ),
    .I2(\dp.rf.rf[28][16] ),
    .I3(\dp.rf.rf[29][16] ),
    .S0(_01157_),
    .S1(_01139_),
    .Z(_02142_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06397_ (.I0(_02141_),
    .I1(_02142_),
    .S(_01889_),
    .Z(_02143_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06398_ (.A1(_01415_),
    .A2(_02143_),
    .ZN(_02144_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06399_ (.I0(\dp.rf.rf[18][16] ),
    .I1(\dp.rf.rf[19][16] ),
    .I2(\dp.rf.rf[22][16] ),
    .I3(\dp.rf.rf[23][16] ),
    .S0(_01429_),
    .S1(_01146_),
    .Z(_02145_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06400_ (.I0(\dp.rf.rf[17][16] ),
    .I1(\dp.rf.rf[21][16] ),
    .S(_01201_),
    .Z(_02146_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06401_ (.A1(_01693_),
    .A2(_02146_),
    .ZN(_02147_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06402_ (.A1(\dp.rf.rf[20][16] ),
    .A2(_01504_),
    .A3(_01339_),
    .B(_01889_),
    .ZN(_02148_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _06403_ (.A1(_02147_),
    .A2(_02148_),
    .B(_01415_),
    .C(_01511_),
    .ZN(_02149_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06404_ (.I(\dp.rf.rf[16][16] ),
    .ZN(_02150_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06405_ (.A1(_02150_),
    .A2(_01737_),
    .ZN(_02151_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06406_ (.A1(_01335_),
    .A2(_02145_),
    .B1(_02149_),
    .B2(_02151_),
    .ZN(_02152_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06407_ (.I0(\dp.rf.rf[14][16] ),
    .I1(\dp.rf.rf[15][16] ),
    .S(_01136_),
    .Z(_02153_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06408_ (.I(_02153_),
    .ZN(_02154_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06409_ (.A1(_01211_),
    .A2(_02154_),
    .B(_02019_),
    .ZN(_02155_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _06410_ (.A1(_01154_),
    .A2(_01155_),
    .A3(_01090_),
    .A4(\dp.rf.rf[10][16] ),
    .ZN(_02156_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06411_ (.I(\dp.rf.rf[10][16] ),
    .ZN(_02157_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _06412_ (.A1(_01028_),
    .A2(_01185_),
    .A3(_02156_),
    .B1(_02157_),
    .B2(_01645_),
    .ZN(_02158_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06413_ (.A1(\dp.rf.rf[11][16] ),
    .A2(_01600_),
    .Z(_02159_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _06414_ (.A1(_01164_),
    .A2(_01166_),
    .A3(_02158_),
    .A4(_02159_),
    .Z(_02160_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06415_ (.I0(\dp.rf.rf[8][16] ),
    .I1(\dp.rf.rf[9][16] ),
    .I2(\dp.rf.rf[12][16] ),
    .I3(\dp.rf.rf[13][16] ),
    .S0(_01577_),
    .S1(_01578_),
    .Z(_02161_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _06416_ (.A1(_02155_),
    .A2(_02160_),
    .B1(_02161_),
    .B2(_01576_),
    .C(_01580_),
    .ZN(_02162_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06417_ (.I0(\dp.rf.rf[2][16] ),
    .I1(\dp.rf.rf[3][16] ),
    .I2(\dp.rf.rf[6][16] ),
    .I3(\dp.rf.rf[7][16] ),
    .S0(_01157_),
    .S1(_01139_),
    .Z(_02163_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06418_ (.A1(_01456_),
    .A2(_02163_),
    .ZN(_02164_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06419_ (.I0(\dp.rf.rf[1][16] ),
    .I1(\dp.rf.rf[5][16] ),
    .S(_01381_),
    .Z(_02165_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06420_ (.A1(\dp.rf.rf[4][16] ),
    .A2(_01497_),
    .B1(_02165_),
    .B2(_01422_),
    .C(_01889_),
    .ZN(_02166_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _06421_ (.A1(_01361_),
    .A2(_02164_),
    .A3(_02166_),
    .Z(_02167_));
 gf180mcu_fd_sc_mcu9t5v0__oai33_4 _06422_ (.A1(_02152_),
    .A2(_02144_),
    .A3(_01455_),
    .B1(_02162_),
    .B2(_02167_),
    .B3(_01589_),
    .ZN(_02168_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _06423_ (.I(_02168_),
    .Z(_04952_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _06424_ (.I(_04952_),
    .ZN(_04956_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _06425_ (.A1(_01292_),
    .A2(_01291_),
    .B(net20),
    .ZN(_02169_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _06426_ (.I(net6),
    .Z(_02170_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06427_ (.A1(_02170_),
    .A2(_01300_),
    .B1(_01296_),
    .B2(_01504_),
    .ZN(_02171_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06428_ (.A1(_02169_),
    .A2(_02171_),
    .ZN(_02172_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06429_ (.I0(_02124_),
    .I1(_02172_),
    .S(net240),
    .Z(_05138_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06430_ (.I(_05138_),
    .ZN(_02173_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06431_ (.I0(\dp.rf.rf[24][15] ),
    .I1(\dp.rf.rf[25][15] ),
    .I2(\dp.rf.rf[26][15] ),
    .I3(\dp.rf.rf[27][15] ),
    .S0(_01928_),
    .S1(_01929_),
    .Z(_02174_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 _06432_ (.I(_01657_),
    .Z(_02175_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _06433_ (.I(_01549_),
    .Z(_02176_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06434_ (.I0(\dp.rf.rf[16][15] ),
    .I1(\dp.rf.rf[17][15] ),
    .I2(\dp.rf.rf[18][15] ),
    .I3(\dp.rf.rf[19][15] ),
    .S0(_02175_),
    .S1(_02176_),
    .Z(_02177_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06435_ (.I0(\dp.rf.rf[28][15] ),
    .I1(\dp.rf.rf[29][15] ),
    .I2(\dp.rf.rf[30][15] ),
    .I3(\dp.rf.rf[31][15] ),
    .S0(_01928_),
    .S1(_01929_),
    .Z(_02178_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06436_ (.I0(\dp.rf.rf[20][15] ),
    .I1(\dp.rf.rf[21][15] ),
    .I2(\dp.rf.rf[22][15] ),
    .I3(\dp.rf.rf[23][15] ),
    .S0(_01928_),
    .S1(_01929_),
    .Z(_02179_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06437_ (.I0(_02174_),
    .I1(_02177_),
    .I2(_02178_),
    .I3(_02179_),
    .S0(_01666_),
    .S1(_01400_),
    .Z(_02180_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06438_ (.I0(\dp.rf.rf[8][15] ),
    .I1(\dp.rf.rf[9][15] ),
    .I2(\dp.rf.rf[10][15] ),
    .I3(\dp.rf.rf[11][15] ),
    .S0(_01928_),
    .S1(_01929_),
    .Z(_02181_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06439_ (.I0(\dp.rf.rf[0][15] ),
    .I1(\dp.rf.rf[1][15] ),
    .I2(\dp.rf.rf[2][15] ),
    .I3(\dp.rf.rf[3][15] ),
    .S0(_02175_),
    .S1(_02176_),
    .Z(_02182_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06440_ (.I0(\dp.rf.rf[12][15] ),
    .I1(\dp.rf.rf[13][15] ),
    .I2(\dp.rf.rf[14][15] ),
    .I3(\dp.rf.rf[15][15] ),
    .S0(net249),
    .S1(_01929_),
    .Z(_02183_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06441_ (.I0(\dp.rf.rf[4][15] ),
    .I1(\dp.rf.rf[5][15] ),
    .I2(\dp.rf.rf[6][15] ),
    .I3(\dp.rf.rf[7][15] ),
    .S0(_01928_),
    .S1(_01929_),
    .Z(_02184_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06442_ (.I0(_02181_),
    .I1(_02182_),
    .I2(_02183_),
    .I3(_02184_),
    .S0(_01272_),
    .S1(_01400_),
    .Z(_02185_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06443_ (.I0(_02180_),
    .I1(_02185_),
    .S(_01058_),
    .Z(_02186_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _06444_ (.A1(net192),
    .A2(_02186_),
    .ZN(_02187_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06445_ (.I0(_02173_),
    .I1(_02187_),
    .S(_01546_),
    .Z(_02188_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06446_ (.A1(_01086_),
    .A2(_02188_),
    .Z(_04961_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06447_ (.I(_04961_),
    .ZN(_04965_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06448_ (.I0(\dp.rf.rf[22][15] ),
    .I1(\dp.rf.rf[23][15] ),
    .S(_01429_),
    .Z(_02189_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06449_ (.A1(_01568_),
    .A2(_02189_),
    .ZN(_02190_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06450_ (.A1(_02019_),
    .A2(_02190_),
    .ZN(_02191_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06451_ (.A1(\dp.rf.rf[18][15] ),
    .A2(_01571_),
    .Z(_02192_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06452_ (.A1(\dp.rf.rf[19][15] ),
    .A2(_01504_),
    .Z(_02193_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _06453_ (.A1(_01593_),
    .A2(_02192_),
    .A3(_02193_),
    .Z(_02194_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06454_ (.I0(\dp.rf.rf[17][15] ),
    .I1(\dp.rf.rf[21][15] ),
    .S(_01169_),
    .Z(_02195_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06455_ (.A1(\dp.rf.rf[20][15] ),
    .A2(_01497_),
    .B1(_02195_),
    .B2(_01693_),
    .C(_01500_),
    .ZN(_02196_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06456_ (.A1(net206),
    .A2(_01355_),
    .B(\dp.rf.rf[16][15] ),
    .ZN(_02197_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06457_ (.A1(_01361_),
    .A2(_02196_),
    .B(_02197_),
    .ZN(_02198_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06458_ (.A1(_02191_),
    .A2(_02194_),
    .B(_02198_),
    .ZN(_02199_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06459_ (.I0(\dp.rf.rf[30][15] ),
    .I1(\dp.rf.rf[31][15] ),
    .S(_01577_),
    .Z(_02200_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _06460_ (.A1(_01568_),
    .A2(_02200_),
    .B(net206),
    .C(_01530_),
    .ZN(_02201_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06461_ (.A1(\dp.rf.rf[27][15] ),
    .A2(_01569_),
    .Z(_02202_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _06462_ (.A1(_01211_),
    .A2(_01511_),
    .B1(_01571_),
    .B2(\dp.rf.rf[26][15] ),
    .C(_02202_),
    .ZN(_02203_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06463_ (.A1(net206),
    .A2(_01377_),
    .B(\dp.rf.rf[24][15] ),
    .ZN(_02204_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06464_ (.I0(\dp.rf.rf[25][15] ),
    .I1(\dp.rf.rf[29][15] ),
    .S(_01201_),
    .Z(_02205_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06465_ (.A1(\dp.rf.rf[28][15] ),
    .A2(_01497_),
    .B1(_02205_),
    .B2(_01693_),
    .C(_01889_),
    .ZN(_02206_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06466_ (.A1(_02201_),
    .A2(_02203_),
    .B1(_02204_),
    .B2(_02206_),
    .C(_01385_),
    .ZN(_02207_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06467_ (.A1(_01207_),
    .A2(_02207_),
    .ZN(_02208_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06468_ (.I0(\dp.rf.rf[14][15] ),
    .I1(\dp.rf.rf[15][15] ),
    .S(_01577_),
    .Z(_02209_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06469_ (.I(_02209_),
    .ZN(_02210_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06470_ (.A1(\dp.rf.rf[10][15] ),
    .A2(_01571_),
    .ZN(_02211_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06471_ (.A1(\dp.rf.rf[11][15] ),
    .A2(_01504_),
    .B1(_01146_),
    .B2(_01435_),
    .ZN(_02212_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _06472_ (.A1(_01211_),
    .A2(_02210_),
    .B1(_02211_),
    .B2(_02212_),
    .C(_02019_),
    .ZN(_02213_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06473_ (.I0(\dp.rf.rf[8][15] ),
    .I1(\dp.rf.rf[9][15] ),
    .I2(\dp.rf.rf[12][15] ),
    .I3(\dp.rf.rf[13][15] ),
    .S0(_01577_),
    .S1(_01146_),
    .Z(_02214_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06474_ (.A1(_01576_),
    .A2(_02214_),
    .Z(_02215_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _06475_ (.A1(_01580_),
    .A2(_02213_),
    .A3(_02215_),
    .ZN(_02216_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06476_ (.I0(\dp.rf.rf[1][15] ),
    .I1(\dp.rf.rf[5][15] ),
    .S(_01381_),
    .Z(_02217_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06477_ (.A1(_01422_),
    .A2(_02217_),
    .ZN(_02218_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06478_ (.A1(\dp.rf.rf[4][15] ),
    .A2(_01429_),
    .A3(_01505_),
    .B(_01430_),
    .ZN(_02219_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06479_ (.A1(_02218_),
    .A2(_02219_),
    .B(_01435_),
    .ZN(_02220_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06480_ (.I(\dp.rf.rf[0][15] ),
    .ZN(_02221_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06481_ (.A1(_02221_),
    .A2(_02012_),
    .ZN(_02222_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06482_ (.I0(\dp.rf.rf[2][15] ),
    .I1(\dp.rf.rf[3][15] ),
    .I2(\dp.rf.rf[6][15] ),
    .I3(\dp.rf.rf[7][15] ),
    .S0(_01520_),
    .S1(_01364_),
    .Z(_02223_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06483_ (.A1(_01362_),
    .A2(_02223_),
    .ZN(_02224_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06484_ (.A1(_01337_),
    .A2(_02224_),
    .ZN(_02225_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06485_ (.A1(_02220_),
    .A2(_02222_),
    .B1(_02225_),
    .B2(net206),
    .ZN(_02226_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _06486_ (.A1(_01589_),
    .A2(_02226_),
    .Z(_02227_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _06487_ (.A1(_02208_),
    .A2(_02199_),
    .B1(_02216_),
    .B2(_02227_),
    .ZN(_02228_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _06488_ (.I(net243),
    .ZN(_04964_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _06489_ (.I(_01085_),
    .Z(_02229_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06490_ (.A1(net5),
    .A2(_01300_),
    .B1(_01296_),
    .B2(_02170_),
    .ZN(_02230_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06491_ (.A1(_02169_),
    .A2(_02230_),
    .ZN(_02231_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06492_ (.I0(_02172_),
    .I1(_02231_),
    .S(net240),
    .Z(_05134_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _06493_ (.I(_01102_),
    .Z(_02232_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06494_ (.I0(\dp.rf.rf[24][14] ),
    .I1(\dp.rf.rf[25][14] ),
    .I2(\dp.rf.rf[26][14] ),
    .I3(\dp.rf.rf[27][14] ),
    .S0(_01661_),
    .S1(_02232_),
    .Z(_02233_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06495_ (.I0(\dp.rf.rf[16][14] ),
    .I1(\dp.rf.rf[17][14] ),
    .I2(\dp.rf.rf[18][14] ),
    .I3(\dp.rf.rf[19][14] ),
    .S0(_01661_),
    .S1(_02232_),
    .Z(_02234_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06496_ (.I0(\dp.rf.rf[28][14] ),
    .I1(\dp.rf.rf[29][14] ),
    .I2(\dp.rf.rf[30][14] ),
    .I3(\dp.rf.rf[31][14] ),
    .S0(_01661_),
    .S1(_01391_),
    .Z(_02235_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06497_ (.I0(\dp.rf.rf[20][14] ),
    .I1(\dp.rf.rf[21][14] ),
    .I2(\dp.rf.rf[22][14] ),
    .I3(\dp.rf.rf[23][14] ),
    .S0(_01661_),
    .S1(_02232_),
    .Z(_02236_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _06498_ (.I0(_02233_),
    .I1(_02234_),
    .I2(_02235_),
    .I3(_02236_),
    .S0(_01394_),
    .S1(net194),
    .Z(_02237_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06499_ (.I0(\dp.rf.rf[8][14] ),
    .I1(\dp.rf.rf[9][14] ),
    .I2(\dp.rf.rf[10][14] ),
    .I3(\dp.rf.rf[11][14] ),
    .S0(_01390_),
    .S1(_01403_),
    .Z(_02238_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06500_ (.I0(\dp.rf.rf[0][14] ),
    .I1(\dp.rf.rf[1][14] ),
    .I2(\dp.rf.rf[2][14] ),
    .I3(\dp.rf.rf[3][14] ),
    .S0(_01390_),
    .S1(_01391_),
    .Z(_02239_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06501_ (.I0(\dp.rf.rf[12][14] ),
    .I1(\dp.rf.rf[13][14] ),
    .I2(\dp.rf.rf[14][14] ),
    .I3(\dp.rf.rf[15][14] ),
    .S0(_01402_),
    .S1(_01403_),
    .Z(_02240_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06502_ (.I0(\dp.rf.rf[4][14] ),
    .I1(\dp.rf.rf[5][14] ),
    .I2(\dp.rf.rf[6][14] ),
    .I3(\dp.rf.rf[7][14] ),
    .S0(_01390_),
    .S1(_01403_),
    .Z(_02241_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _06503_ (.I0(_02238_),
    .I1(_02239_),
    .I2(_02240_),
    .I3(_02241_),
    .S0(_01394_),
    .S1(net194),
    .Z(_02242_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _06504_ (.A1(_01037_),
    .A2(_02237_),
    .B1(_02242_),
    .B2(_01061_),
    .ZN(_02243_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _06505_ (.I(_02243_),
    .ZN(_02244_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06506_ (.I0(_05134_),
    .I1(_02244_),
    .S(_01289_),
    .Z(_02245_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _06507_ (.A1(_02229_),
    .A2(_02245_),
    .ZN(_04969_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06508_ (.I(_04969_),
    .ZN(_04973_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06509_ (.A1(\dp.rf.rf[11][14] ),
    .A2(_01340_),
    .Z(_02246_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _06510_ (.A1(_01578_),
    .A2(net168),
    .B1(_01626_),
    .B2(\dp.rf.rf[10][14] ),
    .C(_02246_),
    .ZN(_02247_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06511_ (.I0(\dp.rf.rf[14][14] ),
    .I1(\dp.rf.rf[15][14] ),
    .S(_01160_),
    .Z(_02248_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06512_ (.A1(_01505_),
    .A2(_02248_),
    .ZN(_02249_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06513_ (.I0(\dp.rf.rf[8][14] ),
    .I1(\dp.rf.rf[9][14] ),
    .I2(\dp.rf.rf[12][14] ),
    .I3(\dp.rf.rf[13][14] ),
    .S0(_01363_),
    .S1(_01364_),
    .Z(_02250_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06514_ (.A1(_01889_),
    .A2(_02250_),
    .ZN(_02251_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06515_ (.A1(_02019_),
    .A2(_02247_),
    .A3(_02249_),
    .B(_02251_),
    .ZN(_02252_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06516_ (.I0(\dp.rf.rf[2][14] ),
    .I1(\dp.rf.rf[3][14] ),
    .I2(\dp.rf.rf[6][14] ),
    .I3(\dp.rf.rf[7][14] ),
    .S0(_01508_),
    .S1(_01201_),
    .Z(_02253_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06517_ (.A1(_01362_),
    .A2(_02253_),
    .ZN(_02254_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06518_ (.I0(\dp.rf.rf[1][14] ),
    .I1(\dp.rf.rf[5][14] ),
    .S(_01457_),
    .Z(_02255_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06519_ (.A1(\dp.rf.rf[4][14] ),
    .A2(_01368_),
    .B1(_02255_),
    .B2(_01442_),
    .C(_01430_),
    .ZN(_02256_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _06520_ (.A1(_01361_),
    .A2(_02254_),
    .A3(_02256_),
    .ZN(_02257_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _06521_ (.A1(_01580_),
    .A2(_02252_),
    .B(_02257_),
    .C(_01376_),
    .ZN(_02258_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06522_ (.I0(\dp.rf.rf[22][14] ),
    .I1(\dp.rf.rf[23][14] ),
    .S(_01428_),
    .Z(_02259_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06523_ (.I(_02259_),
    .ZN(_02260_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06524_ (.A1(\dp.rf.rf[18][14] ),
    .A2(_01571_),
    .ZN(_02261_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06525_ (.A1(\dp.rf.rf[19][14] ),
    .A2(_01429_),
    .B1(_01210_),
    .B2(_01192_),
    .ZN(_02262_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _06526_ (.A1(_01211_),
    .A2(_02260_),
    .B1(_02261_),
    .B2(_02262_),
    .C(_01151_),
    .ZN(_02263_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06527_ (.I(\dp.rf.rf[16][14] ),
    .ZN(_02264_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06528_ (.I0(\dp.rf.rf[17][14] ),
    .I1(\dp.rf.rf[21][14] ),
    .S(_01369_),
    .Z(_02265_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06529_ (.A1(\dp.rf.rf[20][14] ),
    .A2(_01368_),
    .B1(_02265_),
    .B2(_01442_),
    .C(_01372_),
    .ZN(_02266_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06530_ (.A1(_02264_),
    .A2(_01737_),
    .B1(_02266_),
    .B2(_01854_),
    .ZN(_02267_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06531_ (.I0(\dp.rf.rf[26][14] ),
    .I1(\dp.rf.rf[27][14] ),
    .S(_01531_),
    .Z(_02268_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06532_ (.I0(\dp.rf.rf[30][14] ),
    .I1(\dp.rf.rf[31][14] ),
    .S(_01520_),
    .Z(_02269_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _06533_ (.A1(_01164_),
    .A2(_01166_),
    .A3(_02268_),
    .B1(_02269_),
    .B2(_01505_),
    .ZN(_02270_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06534_ (.I0(\dp.rf.rf[24][14] ),
    .I1(\dp.rf.rf[25][14] ),
    .I2(\dp.rf.rf[28][14] ),
    .I3(\dp.rf.rf[29][14] ),
    .S0(_01121_),
    .S1(_01432_),
    .Z(_02271_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06535_ (.A1(_01506_),
    .A2(_02271_),
    .ZN(_02272_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _06536_ (.A1(_01173_),
    .A2(_02270_),
    .B(_02272_),
    .C(_01385_),
    .ZN(_02273_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _06537_ (.A1(_02263_),
    .A2(_02267_),
    .B(net205),
    .C(_02273_),
    .ZN(_02274_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _06538_ (.A1(_02258_),
    .A2(_02274_),
    .ZN(_04968_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _06539_ (.I(_04968_),
    .ZN(_04972_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06540_ (.A1(net4),
    .A2(_01300_),
    .B1(_01296_),
    .B2(net5),
    .ZN(_02275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06541_ (.A1(_02169_),
    .A2(_02275_),
    .ZN(_02276_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06542_ (.I0(_02231_),
    .I1(_02276_),
    .S(net240),
    .Z(_05130_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06543_ (.I(_05130_),
    .ZN(_02277_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _06544_ (.I(_01408_),
    .Z(_02278_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06545_ (.I0(\dp.rf.rf[24][13] ),
    .I1(\dp.rf.rf[25][13] ),
    .I2(\dp.rf.rf[26][13] ),
    .I3(\dp.rf.rf[27][13] ),
    .S0(_01658_),
    .S1(_02278_),
    .Z(_02279_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06546_ (.I0(\dp.rf.rf[16][13] ),
    .I1(\dp.rf.rf[17][13] ),
    .I2(\dp.rf.rf[18][13] ),
    .I3(\dp.rf.rf[19][13] ),
    .S0(_01658_),
    .S1(_02278_),
    .Z(_02280_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06547_ (.I0(\dp.rf.rf[28][13] ),
    .I1(\dp.rf.rf[29][13] ),
    .I2(\dp.rf.rf[30][13] ),
    .I3(\dp.rf.rf[31][13] ),
    .S0(_01820_),
    .S1(_02278_),
    .Z(_02281_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06548_ (.I0(\dp.rf.rf[20][13] ),
    .I1(\dp.rf.rf[21][13] ),
    .I2(\dp.rf.rf[22][13] ),
    .I3(\dp.rf.rf[23][13] ),
    .S0(_01820_),
    .S1(_02278_),
    .Z(_02282_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _06549_ (.I0(_02279_),
    .I1(_02280_),
    .I2(_02281_),
    .I3(_02282_),
    .S0(_01666_),
    .S1(_01478_),
    .Z(_02283_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06550_ (.I0(\dp.rf.rf[8][13] ),
    .I1(\dp.rf.rf[9][13] ),
    .I2(\dp.rf.rf[10][13] ),
    .I3(\dp.rf.rf[11][13] ),
    .S0(_01820_),
    .S1(_02278_),
    .Z(_02284_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06551_ (.I0(\dp.rf.rf[0][13] ),
    .I1(\dp.rf.rf[1][13] ),
    .I2(\dp.rf.rf[2][13] ),
    .I3(\dp.rf.rf[3][13] ),
    .S0(_01820_),
    .S1(_02278_),
    .Z(_02285_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06552_ (.I0(\dp.rf.rf[12][13] ),
    .I1(\dp.rf.rf[13][13] ),
    .I2(\dp.rf.rf[14][13] ),
    .I3(\dp.rf.rf[15][13] ),
    .S0(_01820_),
    .S1(_02278_),
    .Z(_02286_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06553_ (.I0(\dp.rf.rf[4][13] ),
    .I1(\dp.rf.rf[5][13] ),
    .I2(\dp.rf.rf[6][13] ),
    .I3(\dp.rf.rf[7][13] ),
    .S0(_01820_),
    .S1(_02278_),
    .Z(_02287_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _06554_ (.I0(_02284_),
    .I1(_02285_),
    .I2(_02286_),
    .I3(_02287_),
    .S0(_01666_),
    .S1(_01478_),
    .Z(_02288_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _06555_ (.A1(_01111_),
    .A2(_02283_),
    .B1(_02288_),
    .B2(_01112_),
    .ZN(_02289_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06556_ (.I0(_02277_),
    .I1(_02289_),
    .S(_01546_),
    .Z(_02290_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06557_ (.A1(_01086_),
    .A2(_02290_),
    .Z(_04977_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06558_ (.I(_04977_),
    .ZN(_04981_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06559_ (.I0(\dp.rf.rf[17][13] ),
    .I1(\dp.rf.rf[21][13] ),
    .S(_01144_),
    .Z(_02291_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06560_ (.A1(_01636_),
    .A2(_02291_),
    .ZN(_02292_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06561_ (.A1(\dp.rf.rf[20][13] ),
    .A2(_01600_),
    .A3(_01196_),
    .B(_01193_),
    .ZN(_02293_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _06562_ (.A1(_02292_),
    .A2(_02293_),
    .B(_01228_),
    .C(_01077_),
    .ZN(_02294_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06563_ (.I(\dp.rf.rf[16][13] ),
    .ZN(_02295_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06564_ (.A1(_02295_),
    .A2(_01737_),
    .ZN(_02296_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06565_ (.I0(\dp.rf.rf[18][13] ),
    .I1(\dp.rf.rf[19][13] ),
    .S(_01238_),
    .Z(_02297_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06566_ (.I(_02297_),
    .ZN(_02298_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06567_ (.I0(\dp.rf.rf[22][13] ),
    .I1(\dp.rf.rf[23][13] ),
    .S(_01194_),
    .Z(_02299_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06568_ (.A1(_01182_),
    .A2(_02299_),
    .B(_01118_),
    .ZN(_02300_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06569_ (.A1(_01224_),
    .A2(_02298_),
    .B(_02300_),
    .ZN(_02301_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06570_ (.A1(_02294_),
    .A2(_02296_),
    .B(_02301_),
    .ZN(_02302_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _06571_ (.I0(\dp.rf.rf[26][13] ),
    .I1(\dp.rf.rf[27][13] ),
    .I2(\dp.rf.rf[30][13] ),
    .I3(\dp.rf.rf[31][13] ),
    .S0(_01508_),
    .S1(_01201_),
    .Z(_02303_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06572_ (.I0(\dp.rf.rf[24][13] ),
    .I1(\dp.rf.rf[25][13] ),
    .I2(\dp.rf.rf[28][13] ),
    .I3(\dp.rf.rf[29][13] ),
    .S0(_01582_),
    .S1(_01124_),
    .Z(_02304_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _06573_ (.A1(_01334_),
    .A2(_02303_),
    .B1(_02304_),
    .B2(_01506_),
    .C(_01199_),
    .ZN(_02305_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _06574_ (.A1(\dp.rf.rf[4][13] ),
    .A2(_01532_),
    .A3(_01182_),
    .ZN(_02306_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06575_ (.I0(\dp.rf.rf[1][13] ),
    .I1(\dp.rf.rf[5][13] ),
    .S(_01200_),
    .Z(_02307_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06576_ (.A1(_01636_),
    .A2(_02307_),
    .ZN(_02308_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06577_ (.I0(\dp.rf.rf[2][13] ),
    .I1(\dp.rf.rf[3][13] ),
    .I2(\dp.rf.rf[6][13] ),
    .I3(\dp.rf.rf[7][13] ),
    .S0(_01194_),
    .S1(_01369_),
    .Z(_02309_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06578_ (.A1(_01213_),
    .A2(_02309_),
    .ZN(_02310_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06579_ (.A1(_01119_),
    .A2(_02306_),
    .A3(_02308_),
    .B(_02310_),
    .ZN(_02311_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06580_ (.I0(\dp.rf.rf[10][13] ),
    .I1(\dp.rf.rf[11][13] ),
    .I2(\dp.rf.rf[14][13] ),
    .I3(\dp.rf.rf[15][13] ),
    .S0(_01427_),
    .S1(_01168_),
    .Z(_02312_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06581_ (.I0(\dp.rf.rf[8][13] ),
    .I1(\dp.rf.rf[9][13] ),
    .I2(\dp.rf.rf[12][13] ),
    .I3(\dp.rf.rf[13][13] ),
    .S0(_01427_),
    .S1(_01168_),
    .Z(_02313_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06582_ (.I0(_02312_),
    .I1(_02313_),
    .S(_01218_),
    .Z(_02314_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _06583_ (.A1(_01541_),
    .A2(_02311_),
    .B1(_02314_),
    .B2(_01176_),
    .C(_01375_),
    .ZN(_02315_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _06584_ (.A1(net211),
    .A2(_02302_),
    .A3(_02305_),
    .B(_02315_),
    .ZN(_04976_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _06585_ (.I(_04976_),
    .ZN(_04980_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06586_ (.A1(net4),
    .A2(_01296_),
    .ZN(_02316_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06587_ (.A1(_01293_),
    .A2(_02316_),
    .ZN(_02317_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06588_ (.I0(_02276_),
    .I1(_02317_),
    .S(net240),
    .Z(_05126_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06589_ (.I(_05126_),
    .ZN(_02318_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06590_ (.I0(\dp.rf.rf[28][12] ),
    .I1(\dp.rf.rf[29][12] ),
    .I2(\dp.rf.rf[30][12] ),
    .I3(\dp.rf.rf[31][12] ),
    .S0(_01390_),
    .S1(_01403_),
    .Z(_02319_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06591_ (.I0(\dp.rf.rf[20][12] ),
    .I1(\dp.rf.rf[21][12] ),
    .I2(\dp.rf.rf[22][12] ),
    .I3(\dp.rf.rf[23][12] ),
    .S0(_01402_),
    .S1(_01403_),
    .Z(_02320_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06592_ (.I0(_02319_),
    .I1(_02320_),
    .S(_01398_),
    .Z(_02321_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06593_ (.I0(\dp.rf.rf[24][12] ),
    .I1(\dp.rf.rf[25][12] ),
    .I2(\dp.rf.rf[26][12] ),
    .I3(\dp.rf.rf[27][12] ),
    .S0(_01402_),
    .S1(_01403_),
    .Z(_02322_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06594_ (.I0(\dp.rf.rf[16][12] ),
    .I1(\dp.rf.rf[17][12] ),
    .I2(\dp.rf.rf[18][12] ),
    .I3(\dp.rf.rf[19][12] ),
    .S0(_01402_),
    .S1(_01403_),
    .Z(_02323_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06595_ (.I0(_02322_),
    .I1(_02323_),
    .S(_01398_),
    .Z(_02324_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06596_ (.I0(_02321_),
    .I1(_02324_),
    .S(_01669_),
    .Z(_02325_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _06597_ (.I(instr[21]),
    .Z(_02326_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06598_ (.I0(\dp.rf.rf[12][12] ),
    .I1(\dp.rf.rf[13][12] ),
    .I2(\dp.rf.rf[14][12] ),
    .I3(\dp.rf.rf[15][12] ),
    .S0(_01260_),
    .S1(_02326_),
    .Z(_02327_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06599_ (.I0(\dp.rf.rf[8][12] ),
    .I1(\dp.rf.rf[9][12] ),
    .I2(\dp.rf.rf[10][12] ),
    .I3(\dp.rf.rf[11][12] ),
    .S0(_01260_),
    .S1(_02326_),
    .Z(_02328_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06600_ (.I0(_02327_),
    .I1(_02328_),
    .S(_01668_),
    .Z(_02329_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _06601_ (.A1(_01672_),
    .A2(_02329_),
    .Z(_02330_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06602_ (.I0(\dp.rf.rf[4][12] ),
    .I1(\dp.rf.rf[5][12] ),
    .I2(\dp.rf.rf[6][12] ),
    .I3(\dp.rf.rf[7][12] ),
    .S0(_01260_),
    .S1(_02326_),
    .Z(_02331_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06603_ (.I0(\dp.rf.rf[0][12] ),
    .I1(\dp.rf.rf[1][12] ),
    .I2(\dp.rf.rf[2][12] ),
    .I3(\dp.rf.rf[3][12] ),
    .S0(_01260_),
    .S1(_02326_),
    .Z(_02332_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06604_ (.I0(_02331_),
    .I1(_02332_),
    .S(_01668_),
    .Z(_02333_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _06605_ (.A1(_01677_),
    .A2(_02333_),
    .Z(_02334_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _06606_ (.A1(net192),
    .A2(_02330_),
    .A3(_02334_),
    .Z(_02335_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _06607_ (.A1(_01656_),
    .A2(_02325_),
    .B(_02335_),
    .ZN(_02336_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06608_ (.I0(_02318_),
    .I1(_02336_),
    .S(_01546_),
    .Z(_02337_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06609_ (.A1(_01086_),
    .A2(_02337_),
    .Z(_04985_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06610_ (.I(_04985_),
    .ZN(_04989_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06611_ (.I0(\dp.rf.rf[8][12] ),
    .I1(\dp.rf.rf[9][12] ),
    .I2(\dp.rf.rf[12][12] ),
    .I3(\dp.rf.rf[13][12] ),
    .S0(_01157_),
    .S1(_01139_),
    .Z(_02338_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06612_ (.I0(\dp.rf.rf[10][12] ),
    .I1(\dp.rf.rf[11][12] ),
    .S(_01186_),
    .Z(_02339_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06613_ (.I(_02339_),
    .ZN(_02340_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06614_ (.I0(\dp.rf.rf[14][12] ),
    .I1(\dp.rf.rf[15][12] ),
    .S(_01427_),
    .Z(_02341_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06615_ (.A1(_01196_),
    .A2(_02341_),
    .ZN(_02342_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _06616_ (.A1(_01344_),
    .A2(_02340_),
    .B(_02342_),
    .C(_01172_),
    .ZN(_02343_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _06617_ (.A1(_01500_),
    .A2(_02338_),
    .B(_02343_),
    .C(_01176_),
    .ZN(_02344_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06618_ (.I0(\dp.rf.rf[2][12] ),
    .I1(\dp.rf.rf[3][12] ),
    .I2(\dp.rf.rf[6][12] ),
    .I3(\dp.rf.rf[7][12] ),
    .S0(_01531_),
    .S1(_01443_),
    .Z(_02345_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06619_ (.A1(_01119_),
    .A2(_02345_),
    .ZN(_02346_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06620_ (.I0(\dp.rf.rf[1][12] ),
    .I1(\dp.rf.rf[5][12] ),
    .S(_01144_),
    .Z(_02347_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06621_ (.A1(\dp.rf.rf[4][12] ),
    .A2(_01496_),
    .B1(_02347_),
    .B2(_01636_),
    .C(_01241_),
    .ZN(_02348_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _06622_ (.A1(_01854_),
    .A2(_02346_),
    .A3(_02348_),
    .Z(_02349_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06623_ (.I0(\dp.rf.rf[26][12] ),
    .I1(\dp.rf.rf[27][12] ),
    .I2(\dp.rf.rf[30][12] ),
    .I3(\dp.rf.rf[31][12] ),
    .S0(_01194_),
    .S1(_01138_),
    .Z(_02350_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06624_ (.I0(\dp.rf.rf[24][12] ),
    .I1(\dp.rf.rf[25][12] ),
    .I2(\dp.rf.rf[28][12] ),
    .I3(\dp.rf.rf[29][12] ),
    .S0(_01194_),
    .S1(_01138_),
    .Z(_02351_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06625_ (.I0(_02350_),
    .I1(_02351_),
    .S(_01193_),
    .Z(_02352_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06626_ (.A1(_01337_),
    .A2(_02352_),
    .ZN(_02353_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06627_ (.I0(\dp.rf.rf[18][12] ),
    .I1(\dp.rf.rf[19][12] ),
    .I2(\dp.rf.rf[22][12] ),
    .I3(\dp.rf.rf[23][12] ),
    .S0(_01428_),
    .S1(_01145_),
    .Z(_02354_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06628_ (.I0(\dp.rf.rf[17][12] ),
    .I1(\dp.rf.rf[21][12] ),
    .S(_01123_),
    .Z(_02355_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06629_ (.A1(_01328_),
    .A2(_02355_),
    .ZN(_02356_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06630_ (.A1(\dp.rf.rf[20][12] ),
    .A2(_01157_),
    .A3(_01196_),
    .B(_01218_),
    .ZN(_02357_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _06631_ (.A1(_02356_),
    .A2(_02357_),
    .B(_01228_),
    .C(net257),
    .ZN(_02358_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06632_ (.I(\dp.rf.rf[16][12] ),
    .ZN(_02359_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06633_ (.A1(_02359_),
    .A2(_01736_),
    .ZN(_02360_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06634_ (.A1(_01334_),
    .A2(_02354_),
    .B1(_02358_),
    .B2(_02360_),
    .ZN(_02361_));
 gf180mcu_fd_sc_mcu9t5v0__oai33_4 _06635_ (.A1(_02349_),
    .A2(_02344_),
    .A3(_01589_),
    .B1(_02353_),
    .B2(_02361_),
    .B3(net210),
    .ZN(_04984_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _06636_ (.I(_04984_),
    .ZN(_04988_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06637_ (.A1(_01079_),
    .A2(_01082_),
    .Z(_02362_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06638_ (.A1(net25),
    .A2(_02362_),
    .B1(_01296_),
    .B2(_01919_),
    .ZN(_02363_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06639_ (.A1(net239),
    .A2(_02169_),
    .B(_02363_),
    .ZN(_05122_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06640_ (.I0(\dp.rf.rf[24][11] ),
    .I1(\dp.rf.rf[25][11] ),
    .I2(\dp.rf.rf[26][11] ),
    .I3(\dp.rf.rf[27][11] ),
    .S0(_02032_),
    .S1(_01317_),
    .Z(_02364_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06641_ (.I0(\dp.rf.rf[16][11] ),
    .I1(\dp.rf.rf[17][11] ),
    .I2(\dp.rf.rf[18][11] ),
    .I3(\dp.rf.rf[19][11] ),
    .S0(_02032_),
    .S1(_01317_),
    .Z(_02365_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06642_ (.I0(\dp.rf.rf[28][11] ),
    .I1(\dp.rf.rf[29][11] ),
    .I2(\dp.rf.rf[30][11] ),
    .I3(\dp.rf.rf[31][11] ),
    .S0(_01773_),
    .S1(_01774_),
    .Z(_02366_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06643_ (.I0(\dp.rf.rf[20][11] ),
    .I1(\dp.rf.rf[21][11] ),
    .I2(\dp.rf.rf[22][11] ),
    .I3(\dp.rf.rf[23][11] ),
    .S0(_02032_),
    .S1(_01317_),
    .Z(_02367_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06644_ (.I0(_02364_),
    .I1(_02365_),
    .I2(_02366_),
    .I3(_02367_),
    .S0(_01311_),
    .S1(_01312_),
    .Z(_02368_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06645_ (.I0(\dp.rf.rf[8][11] ),
    .I1(\dp.rf.rf[9][11] ),
    .I2(\dp.rf.rf[10][11] ),
    .I3(\dp.rf.rf[11][11] ),
    .S0(_01548_),
    .S1(_01550_),
    .Z(_02369_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06646_ (.I0(\dp.rf.rf[0][11] ),
    .I1(\dp.rf.rf[1][11] ),
    .I2(\dp.rf.rf[2][11] ),
    .I3(\dp.rf.rf[3][11] ),
    .S0(_01548_),
    .S1(_01550_),
    .Z(_02370_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06647_ (.I0(\dp.rf.rf[12][11] ),
    .I1(\dp.rf.rf[13][11] ),
    .I2(\dp.rf.rf[14][11] ),
    .I3(\dp.rf.rf[15][11] ),
    .S0(_01553_),
    .S1(_01555_),
    .Z(_02371_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06648_ (.I0(\dp.rf.rf[4][11] ),
    .I1(\dp.rf.rf[5][11] ),
    .I2(\dp.rf.rf[6][11] ),
    .I3(\dp.rf.rf[7][11] ),
    .S0(net249),
    .S1(_01550_),
    .Z(_02372_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06649_ (.I0(_02369_),
    .I1(_02370_),
    .I2(_02371_),
    .I3(_02372_),
    .S0(_01272_),
    .S1(_01400_),
    .Z(_02373_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06650_ (.A1(_01608_),
    .A2(_02373_),
    .Z(_02374_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _06651_ (.I0(_02368_),
    .I1(_02374_),
    .S(_01656_),
    .Z(_02375_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06652_ (.I0(_05122_),
    .I1(_02375_),
    .S(_01289_),
    .Z(_02376_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _06653_ (.A1(_02229_),
    .A2(_02376_),
    .ZN(_04993_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06654_ (.I(_04993_),
    .ZN(_04997_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06655_ (.I0(\dp.rf.rf[1][11] ),
    .I1(\dp.rf.rf[5][11] ),
    .S(_01248_),
    .Z(_02377_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06656_ (.A1(_01190_),
    .A2(_02377_),
    .ZN(_02378_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06657_ (.A1(\dp.rf.rf[4][11] ),
    .A2(_01340_),
    .A3(_01162_),
    .B(_01218_),
    .ZN(_02379_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06658_ (.A1(_02378_),
    .A2(_02379_),
    .B(net257),
    .ZN(_02380_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06659_ (.A1(\dp.rf.rf[0][11] ),
    .A2(_01325_),
    .B(_02380_),
    .ZN(_02381_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06660_ (.I0(\dp.rf.rf[2][11] ),
    .I1(\dp.rf.rf[3][11] ),
    .I2(\dp.rf.rf[6][11] ),
    .I3(\dp.rf.rf[7][11] ),
    .S0(_01128_),
    .S1(_01144_),
    .Z(_02382_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06661_ (.A1(_01353_),
    .A2(_02382_),
    .B(net8),
    .ZN(_02383_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _06662_ (.A1(net199),
    .A2(_02383_),
    .Z(_02384_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06663_ (.I0(\dp.rf.rf[14][11] ),
    .I1(\dp.rf.rf[15][11] ),
    .S(_01121_),
    .Z(_02385_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06664_ (.A1(\dp.rf.rf[10][11] ),
    .A2(net203),
    .Z(_02386_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06665_ (.A1(\dp.rf.rf[11][11] ),
    .A2(_01428_),
    .ZN(_02387_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06666_ (.A1(_01223_),
    .A2(_02387_),
    .ZN(_02388_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06667_ (.A1(_01230_),
    .A2(_02385_),
    .B1(_02386_),
    .B2(_02388_),
    .C(_01334_),
    .ZN(_02389_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06668_ (.I0(\dp.rf.rf[8][11] ),
    .I1(\dp.rf.rf[9][11] ),
    .I2(\dp.rf.rf[12][11] ),
    .I3(\dp.rf.rf[13][11] ),
    .S0(_01225_),
    .S1(_01443_),
    .Z(_02390_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06669_ (.A1(_01430_),
    .A2(_02390_),
    .B(_01199_),
    .ZN(_02391_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _06670_ (.A1(_02381_),
    .A2(_02384_),
    .B1(_02391_),
    .B2(_02389_),
    .C(net190),
    .ZN(_02392_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06671_ (.I0(\dp.rf.rf[22][11] ),
    .I1(\dp.rf.rf[23][11] ),
    .S(_01428_),
    .Z(_02393_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06672_ (.A1(\dp.rf.rf[18][11] ),
    .A2(net203),
    .Z(_02394_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06673_ (.A1(\dp.rf.rf[19][11] ),
    .A2(_01212_),
    .ZN(_02395_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06674_ (.A1(_01344_),
    .A2(_02395_),
    .ZN(_02396_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06675_ (.A1(_01339_),
    .A2(_02393_),
    .B1(_02394_),
    .B2(_02396_),
    .C(_01334_),
    .ZN(_02397_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06676_ (.I(\dp.rf.rf[20][11] ),
    .ZN(_02398_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06677_ (.I0(\dp.rf.rf[17][11] ),
    .I1(\dp.rf.rf[21][11] ),
    .S(_01129_),
    .Z(_02399_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06678_ (.A1(_01190_),
    .A2(_02399_),
    .ZN(_02400_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _06679_ (.A1(_02398_),
    .A2(_01249_),
    .B(_02400_),
    .C(_01353_),
    .ZN(_02401_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _06680_ (.A1(\dp.rf.rf[16][11] ),
    .A2(_01356_),
    .B1(_02401_),
    .B2(net229),
    .ZN(_02402_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06681_ (.I0(\dp.rf.rf[26][11] ),
    .I1(\dp.rf.rf[27][11] ),
    .I2(\dp.rf.rf[30][11] ),
    .I3(\dp.rf.rf[31][11] ),
    .S0(_01202_),
    .S1(_01200_),
    .Z(_02403_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06682_ (.I0(\dp.rf.rf[24][11] ),
    .I1(\dp.rf.rf[25][11] ),
    .I2(\dp.rf.rf[28][11] ),
    .I3(\dp.rf.rf[29][11] ),
    .S0(_01202_),
    .S1(_01200_),
    .Z(_02404_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06683_ (.I0(_02403_),
    .I1(_02404_),
    .S(_01171_),
    .Z(_02405_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06684_ (.A1(_01228_),
    .A2(_02405_),
    .B(net177),
    .ZN(_02406_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06685_ (.A1(_02397_),
    .A2(_02402_),
    .B(_02406_),
    .ZN(_02407_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _06686_ (.A1(_02392_),
    .A2(_02407_),
    .Z(_04992_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06687_ (.I(net237),
    .ZN(_02408_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _06688_ (.I(_02408_),
    .Z(_04996_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _06689_ (.I(_01078_),
    .Z(_02409_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06690_ (.A1(net19),
    .A2(_02409_),
    .Z(_05118_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06691_ (.I0(\dp.rf.rf[6][10] ),
    .I1(\dp.rf.rf[7][10] ),
    .I2(\dp.rf.rf[14][10] ),
    .I3(\dp.rf.rf[15][10] ),
    .S0(_01820_),
    .S1(_01761_),
    .Z(_02410_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06692_ (.I0(\dp.rf.rf[2][10] ),
    .I1(\dp.rf.rf[3][10] ),
    .I2(\dp.rf.rf[10][10] ),
    .I3(\dp.rf.rf[11][10] ),
    .S0(_01820_),
    .S1(_01761_),
    .Z(_02411_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06693_ (.I0(\dp.rf.rf[4][10] ),
    .I1(\dp.rf.rf[5][10] ),
    .I2(\dp.rf.rf[12][10] ),
    .I3(\dp.rf.rf[13][10] ),
    .S0(_02175_),
    .S1(_01763_),
    .Z(_02412_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06694_ (.I0(\dp.rf.rf[0][10] ),
    .I1(\dp.rf.rf[1][10] ),
    .I2(\dp.rf.rf[8][10] ),
    .I3(\dp.rf.rf[9][10] ),
    .S0(_01820_),
    .S1(_01761_),
    .Z(_02413_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06695_ (.I0(_02410_),
    .I1(_02411_),
    .I2(_02412_),
    .I3(_02413_),
    .S0(_01779_),
    .S1(_01766_),
    .Z(_02414_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06696_ (.A1(_01112_),
    .A2(_02414_),
    .Z(_02415_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06697_ (.I0(\dp.rf.rf[24][10] ),
    .I1(\dp.rf.rf[25][10] ),
    .I2(\dp.rf.rf[26][10] ),
    .I3(\dp.rf.rf[27][10] ),
    .S0(_01662_),
    .S1(_01659_),
    .Z(_02416_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _06698_ (.A1(_01311_),
    .A2(_02416_),
    .Z(_02417_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06699_ (.I0(\dp.rf.rf[18][10] ),
    .I1(\dp.rf.rf[19][10] ),
    .S(_01658_),
    .Z(_02418_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _06700_ (.A1(_01766_),
    .A2(_01761_),
    .A3(_02418_),
    .Z(_02419_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06701_ (.I0(\dp.rf.rf[16][10] ),
    .I1(\dp.rf.rf[17][10] ),
    .S(_01658_),
    .Z(_02420_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _06702_ (.A1(_01819_),
    .A2(_01761_),
    .A3(_02420_),
    .Z(_02421_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _06703_ (.A1(_01780_),
    .A2(_02417_),
    .A3(_02419_),
    .A4(_02421_),
    .Z(_02422_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06704_ (.I0(\dp.rf.rf[28][10] ),
    .I1(\dp.rf.rf[29][10] ),
    .I2(\dp.rf.rf[30][10] ),
    .I3(\dp.rf.rf[31][10] ),
    .S0(_01658_),
    .S1(_02278_),
    .Z(_02423_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06705_ (.I0(\dp.rf.rf[20][10] ),
    .I1(\dp.rf.rf[21][10] ),
    .I2(\dp.rf.rf[22][10] ),
    .I3(\dp.rf.rf[23][10] ),
    .S0(_01658_),
    .S1(_02278_),
    .Z(_02424_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06706_ (.I0(_02423_),
    .I1(_02424_),
    .S(_01666_),
    .Z(_02425_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06707_ (.A1(net213),
    .A2(_02425_),
    .Z(_02426_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _06708_ (.A1(_02422_),
    .A2(_02415_),
    .A3(_02426_),
    .Z(_02427_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06709_ (.I0(_05118_),
    .I1(_02427_),
    .S(_01289_),
    .Z(_02428_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _06710_ (.A1(_02229_),
    .A2(_02428_),
    .ZN(_05001_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06711_ (.I(_05001_),
    .ZN(_05005_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06712_ (.A1(\dp.rf.rf[2][10] ),
    .A2(_01118_),
    .B(_01355_),
    .ZN(_02429_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06713_ (.A1(net199),
    .A2(_02429_),
    .ZN(_02430_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06714_ (.A1(\dp.rf.rf[0][10] ),
    .A2(_02430_),
    .ZN(_02431_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06715_ (.I0(\dp.rf.rf[10][10] ),
    .I1(\dp.rf.rf[11][10] ),
    .I2(\dp.rf.rf[14][10] ),
    .I3(\dp.rf.rf[15][10] ),
    .S0(_01202_),
    .S1(_01123_),
    .Z(_02432_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06716_ (.I0(\dp.rf.rf[8][10] ),
    .I1(\dp.rf.rf[9][10] ),
    .I2(\dp.rf.rf[12][10] ),
    .I3(\dp.rf.rf[13][10] ),
    .S0(_01202_),
    .S1(_01123_),
    .Z(_02433_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06717_ (.I0(_02432_),
    .I1(_02433_),
    .S(_01171_),
    .Z(_02434_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06718_ (.A1(_01199_),
    .A2(_02434_),
    .ZN(_02435_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06719_ (.I0(\dp.rf.rf[2][10] ),
    .I1(\dp.rf.rf[3][10] ),
    .I2(\dp.rf.rf[6][10] ),
    .I3(\dp.rf.rf[7][10] ),
    .S0(_01128_),
    .S1(_01144_),
    .Z(_02436_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06720_ (.A1(_01353_),
    .A2(_02436_),
    .ZN(_02437_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06721_ (.I0(\dp.rf.rf[1][10] ),
    .I1(\dp.rf.rf[5][10] ),
    .S(_01129_),
    .Z(_02438_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06722_ (.A1(\dp.rf.rf[4][10] ),
    .A2(_01367_),
    .B1(_02438_),
    .B2(_01190_),
    .C(_01218_),
    .ZN(_02439_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _06723_ (.A1(_01360_),
    .A2(_02437_),
    .A3(_02439_),
    .Z(_02440_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _06724_ (.A1(net189),
    .A2(_02431_),
    .A3(_02435_),
    .A4(_02440_),
    .Z(_02441_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06725_ (.A1(\dp.rf.rf[18][10] ),
    .A2(_01571_),
    .ZN(_02442_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06726_ (.A1(\dp.rf.rf[19][10] ),
    .A2(_01429_),
    .B1(_01578_),
    .B2(_01077_),
    .ZN(_02443_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06727_ (.I0(\dp.rf.rf[22][10] ),
    .I1(\dp.rf.rf[23][10] ),
    .S(_01582_),
    .Z(_02444_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06728_ (.A1(_01230_),
    .A2(_02444_),
    .ZN(_02445_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _06729_ (.A1(_02442_),
    .A2(_02443_),
    .B(_01151_),
    .C(_02445_),
    .ZN(_02446_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06730_ (.I(\dp.rf.rf[16][10] ),
    .ZN(_02447_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06731_ (.I0(\dp.rf.rf[17][10] ),
    .I1(\dp.rf.rf[21][10] ),
    .S(_01168_),
    .Z(_02448_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06732_ (.A1(\dp.rf.rf[20][10] ),
    .A2(_01496_),
    .B1(_02448_),
    .B2(_01371_),
    .C(_01172_),
    .ZN(_02449_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06733_ (.A1(_02447_),
    .A2(_01737_),
    .B1(_02449_),
    .B2(_01854_),
    .ZN(_02450_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06734_ (.I0(\dp.rf.rf[30][10] ),
    .I1(\dp.rf.rf[31][10] ),
    .S(_01202_),
    .Z(_02451_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06735_ (.I(_02451_),
    .ZN(_02452_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06736_ (.I0(\dp.rf.rf[26][10] ),
    .I1(\dp.rf.rf[27][10] ),
    .S(_01120_),
    .Z(_02453_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06737_ (.I(_02453_),
    .ZN(_02454_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06738_ (.A1(_01169_),
    .A2(_02452_),
    .B1(_02454_),
    .B2(_01223_),
    .ZN(_02455_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06739_ (.I0(\dp.rf.rf[24][10] ),
    .I1(\dp.rf.rf[25][10] ),
    .I2(\dp.rf.rf[28][10] ),
    .I3(\dp.rf.rf[29][10] ),
    .S0(_01225_),
    .S1(_01443_),
    .Z(_02456_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06740_ (.I0(_02455_),
    .I1(_02456_),
    .S(_01172_),
    .Z(_02457_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _06741_ (.A1(_02446_),
    .A2(_02450_),
    .B1(_02457_),
    .B2(_01237_),
    .C(_01207_),
    .ZN(_02458_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _06742_ (.A1(_02441_),
    .A2(_02458_),
    .ZN(_05000_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06743_ (.I(_05000_),
    .ZN(_02459_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _06744_ (.I(_02459_),
    .Z(_05004_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06745_ (.A1(net18),
    .A2(_02409_),
    .Z(_05114_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06746_ (.I0(\dp.rf.rf[24][9] ),
    .I1(\dp.rf.rf[25][9] ),
    .I2(\dp.rf.rf[26][9] ),
    .I3(\dp.rf.rf[27][9] ),
    .S0(_01484_),
    .S1(_01485_),
    .Z(_02460_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06747_ (.I0(\dp.rf.rf[16][9] ),
    .I1(\dp.rf.rf[17][9] ),
    .I2(\dp.rf.rf[18][9] ),
    .I3(\dp.rf.rf[19][9] ),
    .S0(_01484_),
    .S1(_01485_),
    .Z(_02461_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06748_ (.I0(_02460_),
    .I1(_02461_),
    .S(_01394_),
    .Z(_02462_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06749_ (.I0(\dp.rf.rf[28][9] ),
    .I1(\dp.rf.rf[29][9] ),
    .I2(\dp.rf.rf[30][9] ),
    .I3(\dp.rf.rf[31][9] ),
    .S0(_01484_),
    .S1(_01485_),
    .Z(_02463_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06750_ (.I0(\dp.rf.rf[20][9] ),
    .I1(\dp.rf.rf[21][9] ),
    .I2(\dp.rf.rf[22][9] ),
    .I3(\dp.rf.rf[23][9] ),
    .S0(_01484_),
    .S1(_02232_),
    .Z(_02464_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06751_ (.I0(_02463_),
    .I1(_02464_),
    .S(_01394_),
    .Z(_02465_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06752_ (.I0(_02462_),
    .I1(_02465_),
    .S(_01478_),
    .Z(_02466_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06753_ (.I0(\dp.rf.rf[4][9] ),
    .I1(\dp.rf.rf[5][9] ),
    .I2(\dp.rf.rf[6][9] ),
    .I3(\dp.rf.rf[7][9] ),
    .S0(net261),
    .S1(_01549_),
    .Z(_02467_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06754_ (.I0(\dp.rf.rf[0][9] ),
    .I1(\dp.rf.rf[1][9] ),
    .I2(\dp.rf.rf[2][9] ),
    .I3(\dp.rf.rf[3][9] ),
    .S0(net261),
    .S1(_01549_),
    .Z(_02468_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06755_ (.I0(_02467_),
    .I1(_02468_),
    .S(_01668_),
    .Z(_02469_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _06756_ (.A1(_01677_),
    .A2(_02469_),
    .Z(_02470_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06757_ (.I0(\dp.rf.rf[12][9] ),
    .I1(\dp.rf.rf[13][9] ),
    .I2(\dp.rf.rf[14][9] ),
    .I3(\dp.rf.rf[15][9] ),
    .S0(net261),
    .S1(_01549_),
    .Z(_02471_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06758_ (.I0(\dp.rf.rf[8][9] ),
    .I1(\dp.rf.rf[9][9] ),
    .I2(\dp.rf.rf[10][9] ),
    .I3(\dp.rf.rf[11][9] ),
    .S0(_01098_),
    .S1(_01554_),
    .Z(_02472_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06759_ (.I0(_02471_),
    .I1(_02472_),
    .S(_01668_),
    .Z(_02473_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _06760_ (.A1(_01672_),
    .A2(_02473_),
    .Z(_02474_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _06761_ (.A1(_01608_),
    .A2(_02470_),
    .A3(_02474_),
    .Z(_02475_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _06762_ (.A1(_01656_),
    .A2(_02466_),
    .B(_02475_),
    .ZN(_02476_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _06763_ (.I(_02476_),
    .ZN(_02477_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06764_ (.I0(_05114_),
    .I1(_02477_),
    .S(_01289_),
    .Z(_02478_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _06765_ (.A1(_02478_),
    .A2(_02229_),
    .ZN(_05009_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06766_ (.I(_05009_),
    .ZN(_05013_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06767_ (.I0(\dp.rf.rf[8][9] ),
    .I1(\dp.rf.rf[9][9] ),
    .I2(\dp.rf.rf[12][9] ),
    .I3(\dp.rf.rf[13][9] ),
    .S0(_01136_),
    .S1(_01169_),
    .Z(_02479_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06768_ (.I0(\dp.rf.rf[10][9] ),
    .I1(\dp.rf.rf[11][9] ),
    .S(_01135_),
    .Z(_02480_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06769_ (.I(_02480_),
    .ZN(_02481_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06770_ (.I0(\dp.rf.rf[14][9] ),
    .I1(\dp.rf.rf[15][9] ),
    .S(_01427_),
    .Z(_02482_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06771_ (.A1(_01196_),
    .A2(_02482_),
    .ZN(_02483_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _06772_ (.A1(_01344_),
    .A2(_02481_),
    .B(_02483_),
    .C(_01241_),
    .ZN(_02484_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _06773_ (.A1(_01173_),
    .A2(_02479_),
    .B(_02484_),
    .C(_01176_),
    .ZN(_02485_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06774_ (.I0(\dp.rf.rf[2][9] ),
    .I1(\dp.rf.rf[3][9] ),
    .I2(\dp.rf.rf[6][9] ),
    .I3(\dp.rf.rf[7][9] ),
    .S0(_01179_),
    .S1(_01209_),
    .Z(_02486_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06775_ (.A1(_01119_),
    .A2(_02486_),
    .ZN(_02487_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06776_ (.I0(\dp.rf.rf[1][9] ),
    .I1(\dp.rf.rf[5][9] ),
    .S(_01144_),
    .Z(_02488_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06777_ (.A1(\dp.rf.rf[4][9] ),
    .A2(_01496_),
    .B1(_02488_),
    .B2(_01636_),
    .C(_01241_),
    .ZN(_02489_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _06778_ (.A1(_01854_),
    .A2(_02487_),
    .A3(_02489_),
    .Z(_02490_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06779_ (.I0(\dp.rf.rf[18][9] ),
    .I1(\dp.rf.rf[19][9] ),
    .I2(\dp.rf.rf[22][9] ),
    .I3(\dp.rf.rf[23][9] ),
    .S0(_01121_),
    .S1(_01432_),
    .Z(_02491_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06780_ (.I0(\dp.rf.rf[16][9] ),
    .I1(\dp.rf.rf[17][9] ),
    .I2(\dp.rf.rf[20][9] ),
    .I3(\dp.rf.rf[21][9] ),
    .S0(_01121_),
    .S1(_01432_),
    .Z(_02492_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06781_ (.I0(_02491_),
    .I1(_02492_),
    .S(_01372_),
    .Z(_02493_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06782_ (.A1(_01178_),
    .A2(_02493_),
    .B(_01207_),
    .ZN(_02494_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06783_ (.I0(\dp.rf.rf[24][9] ),
    .I1(\dp.rf.rf[25][9] ),
    .I2(\dp.rf.rf[28][9] ),
    .I3(\dp.rf.rf[29][9] ),
    .S0(_01645_),
    .S1(_01578_),
    .Z(_02495_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06784_ (.I0(\dp.rf.rf[26][9] ),
    .I1(\dp.rf.rf[27][9] ),
    .S(_01582_),
    .Z(_02496_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06785_ (.I(_02496_),
    .ZN(_02497_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06786_ (.I0(\dp.rf.rf[30][9] ),
    .I1(\dp.rf.rf[31][9] ),
    .S(_01179_),
    .Z(_02498_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06787_ (.A1(_01182_),
    .A2(_02498_),
    .ZN(_02499_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _06788_ (.A1(_01224_),
    .A2(_02497_),
    .B(_02499_),
    .C(_01506_),
    .ZN(_02500_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _06789_ (.A1(_01576_),
    .A2(_02495_),
    .B(_02500_),
    .C(_01237_),
    .ZN(_02501_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _06790_ (.A1(_02490_),
    .A2(_02485_),
    .A3(_01589_),
    .B1(_02494_),
    .B2(_02501_),
    .ZN(_05008_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _06791_ (.I(net184),
    .ZN(_05012_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06792_ (.A1(net17),
    .A2(_02409_),
    .Z(_05110_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06793_ (.I0(\dp.rf.rf[28][8] ),
    .I1(\dp.rf.rf[29][8] ),
    .I2(\dp.rf.rf[30][8] ),
    .I3(\dp.rf.rf[31][8] ),
    .S0(_01548_),
    .S1(_01550_),
    .Z(_02502_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06794_ (.I0(\dp.rf.rf[20][8] ),
    .I1(\dp.rf.rf[21][8] ),
    .I2(\dp.rf.rf[22][8] ),
    .I3(\dp.rf.rf[23][8] ),
    .S0(_01548_),
    .S1(_01550_),
    .Z(_02503_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06795_ (.I0(\dp.rf.rf[24][8] ),
    .I1(\dp.rf.rf[25][8] ),
    .I2(\dp.rf.rf[26][8] ),
    .I3(\dp.rf.rf[27][8] ),
    .S0(_01553_),
    .S1(_01555_),
    .Z(_02504_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06796_ (.I0(\dp.rf.rf[16][8] ),
    .I1(\dp.rf.rf[17][8] ),
    .I2(\dp.rf.rf[18][8] ),
    .I3(\dp.rf.rf[19][8] ),
    .S0(_01548_),
    .S1(_01550_),
    .Z(_02505_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _06797_ (.I0(_02502_),
    .I1(_02503_),
    .I2(_02504_),
    .I3(_02505_),
    .S0(_01272_),
    .S1(_01669_),
    .Z(_02506_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06798_ (.I0(\dp.rf.rf[12][8] ),
    .I1(\dp.rf.rf[13][8] ),
    .I2(\dp.rf.rf[14][8] ),
    .I3(\dp.rf.rf[15][8] ),
    .S0(_02175_),
    .S1(_02176_),
    .Z(_02507_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06799_ (.I0(\dp.rf.rf[8][8] ),
    .I1(\dp.rf.rf[9][8] ),
    .I2(\dp.rf.rf[10][8] ),
    .I3(\dp.rf.rf[11][8] ),
    .S0(_02175_),
    .S1(_02176_),
    .Z(_02508_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06800_ (.I0(_02507_),
    .I1(_02508_),
    .S(_01779_),
    .Z(_02509_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06801_ (.I0(\dp.rf.rf[4][8] ),
    .I1(\dp.rf.rf[5][8] ),
    .I2(\dp.rf.rf[6][8] ),
    .I3(\dp.rf.rf[7][8] ),
    .S0(_01266_),
    .S1(_01262_),
    .Z(_02510_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06802_ (.I0(\dp.rf.rf[0][8] ),
    .I1(\dp.rf.rf[1][8] ),
    .I2(\dp.rf.rf[2][8] ),
    .I3(\dp.rf.rf[3][8] ),
    .S0(_01266_),
    .S1(_01262_),
    .Z(_02511_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06803_ (.I0(_02510_),
    .I1(_02511_),
    .S(_01668_),
    .Z(_02512_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _06804_ (.A1(_01677_),
    .A2(_02512_),
    .Z(_02513_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06805_ (.A1(_01607_),
    .A2(_02513_),
    .Z(_02514_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _06806_ (.A1(_01656_),
    .A2(_02506_),
    .B1(_02509_),
    .B2(_01672_),
    .C(_02514_),
    .ZN(_02515_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _06807_ (.I(_02515_),
    .ZN(_02516_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06808_ (.I0(_05110_),
    .I1(_02516_),
    .S(_01289_),
    .Z(_02517_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _06809_ (.A1(_02517_),
    .A2(_02229_),
    .ZN(_05017_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06810_ (.I(_05017_),
    .ZN(_05021_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06811_ (.I0(\dp.rf.rf[14][8] ),
    .I1(\dp.rf.rf[15][8] ),
    .S(_01179_),
    .Z(_02518_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06812_ (.I(_02518_),
    .ZN(_02519_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06813_ (.A1(_01578_),
    .A2(_02519_),
    .B(_01151_),
    .ZN(_02520_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _06814_ (.A1(\dp.rf.rf[10][8] ),
    .A2(_01154_),
    .A3(_01155_),
    .A4(_01034_),
    .ZN(_02521_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06815_ (.I(\dp.rf.rf[10][8] ),
    .ZN(_02522_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _06816_ (.A1(_01028_),
    .A2(_01153_),
    .A3(_02521_),
    .B1(_01520_),
    .B2(_02522_),
    .ZN(_02523_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06817_ (.A1(\dp.rf.rf[11][8] ),
    .A2(_01225_),
    .Z(_02524_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _06818_ (.A1(_01164_),
    .A2(_01166_),
    .A3(_02523_),
    .A4(_02524_),
    .Z(_02525_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06819_ (.I0(\dp.rf.rf[8][8] ),
    .I1(\dp.rf.rf[9][8] ),
    .I2(\dp.rf.rf[12][8] ),
    .I3(\dp.rf.rf[13][8] ),
    .S0(_01508_),
    .S1(_01145_),
    .Z(_02526_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _06820_ (.A1(_02520_),
    .A2(_02525_),
    .B1(_02526_),
    .B2(_01889_),
    .C(_01176_),
    .ZN(_02527_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06821_ (.I0(\dp.rf.rf[2][8] ),
    .I1(\dp.rf.rf[3][8] ),
    .I2(\dp.rf.rf[6][8] ),
    .I3(\dp.rf.rf[7][8] ),
    .S0(_01179_),
    .S1(_01209_),
    .Z(_02528_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06822_ (.A1(_01529_),
    .A2(_02528_),
    .ZN(_02529_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06823_ (.I0(\dp.rf.rf[1][8] ),
    .I1(\dp.rf.rf[5][8] ),
    .S(_01200_),
    .Z(_02530_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06824_ (.A1(\dp.rf.rf[4][8] ),
    .A2(_01496_),
    .B1(_02530_),
    .B2(_01636_),
    .C(_01241_),
    .ZN(_02531_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _06825_ (.A1(_01854_),
    .A2(_02529_),
    .A3(_02531_),
    .Z(_02532_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06826_ (.I0(\dp.rf.rf[26][8] ),
    .I1(\dp.rf.rf[27][8] ),
    .I2(\dp.rf.rf[30][8] ),
    .I3(\dp.rf.rf[31][8] ),
    .S0(_01147_),
    .S1(_01432_),
    .Z(_02533_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06827_ (.I0(\dp.rf.rf[24][8] ),
    .I1(\dp.rf.rf[25][8] ),
    .I2(\dp.rf.rf[28][8] ),
    .I3(\dp.rf.rf[29][8] ),
    .S0(_01147_),
    .S1(_01381_),
    .Z(_02534_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06828_ (.I0(_02533_),
    .I1(_02534_),
    .S(_01372_),
    .Z(_02535_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06829_ (.A1(_01415_),
    .A2(_02535_),
    .B(_01207_),
    .ZN(_02536_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06830_ (.I0(\dp.rf.rf[22][8] ),
    .I1(\dp.rf.rf[23][8] ),
    .S(_01160_),
    .Z(_02537_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06831_ (.I(_02537_),
    .ZN(_02538_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06832_ (.A1(_01146_),
    .A2(_02538_),
    .B(_02019_),
    .ZN(_02539_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _06833_ (.A1(\dp.rf.rf[18][8] ),
    .A2(_01154_),
    .A3(_01155_),
    .A4(_01090_),
    .ZN(_02540_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06834_ (.I(\dp.rf.rf[18][8] ),
    .ZN(_02541_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _06835_ (.A1(_01028_),
    .A2(_01185_),
    .A3(_02540_),
    .B1(_01345_),
    .B2(_02541_),
    .ZN(_02542_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06836_ (.A1(\dp.rf.rf[19][8] ),
    .A2(_01136_),
    .Z(_02543_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _06837_ (.A1(_01164_),
    .A2(_01166_),
    .A3(_02542_),
    .A4(_02543_),
    .Z(_02544_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06838_ (.I0(\dp.rf.rf[17][8] ),
    .I1(\dp.rf.rf[21][8] ),
    .S(_01457_),
    .Z(_02545_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06839_ (.A1(_01442_),
    .A2(_02545_),
    .ZN(_02546_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06840_ (.A1(\dp.rf.rf[20][8] ),
    .A2(_01569_),
    .A3(_01230_),
    .B(_01172_),
    .ZN(_02547_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _06841_ (.A1(_02546_),
    .A2(_02547_),
    .B(_01337_),
    .C(_01435_),
    .ZN(_02548_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06842_ (.I(\dp.rf.rf[16][8] ),
    .ZN(_02549_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06843_ (.A1(_02549_),
    .A2(_01737_),
    .ZN(_02550_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06844_ (.A1(_02539_),
    .A2(_02544_),
    .B1(_02548_),
    .B2(_02550_),
    .ZN(_02551_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _06845_ (.A1(_02532_),
    .A2(_02527_),
    .A3(_01589_),
    .B1(_02536_),
    .B2(_02551_),
    .ZN(_05016_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _06846_ (.I(net170),
    .ZN(_05020_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06847_ (.I0(\dp.rf.rf[24][7] ),
    .I1(\dp.rf.rf[25][7] ),
    .I2(\dp.rf.rf[26][7] ),
    .I3(\dp.rf.rf[27][7] ),
    .S0(_02175_),
    .S1(_02176_),
    .Z(_02552_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06848_ (.I0(\dp.rf.rf[16][7] ),
    .I1(\dp.rf.rf[17][7] ),
    .I2(\dp.rf.rf[18][7] ),
    .I3(\dp.rf.rf[19][7] ),
    .S0(_02175_),
    .S1(_02176_),
    .Z(_02553_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06849_ (.I0(\dp.rf.rf[28][7] ),
    .I1(\dp.rf.rf[29][7] ),
    .I2(\dp.rf.rf[30][7] ),
    .I3(\dp.rf.rf[31][7] ),
    .S0(_01928_),
    .S1(_01929_),
    .Z(_02554_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06850_ (.I0(\dp.rf.rf[20][7] ),
    .I1(\dp.rf.rf[21][7] ),
    .I2(\dp.rf.rf[22][7] ),
    .I3(\dp.rf.rf[23][7] ),
    .S0(_02175_),
    .S1(_02176_),
    .Z(_02555_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06851_ (.I0(_02552_),
    .I1(_02553_),
    .I2(_02554_),
    .I3(_02555_),
    .S0(_01666_),
    .S1(_01478_),
    .Z(_02556_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06852_ (.I0(\dp.rf.rf[8][7] ),
    .I1(\dp.rf.rf[9][7] ),
    .I2(\dp.rf.rf[10][7] ),
    .I3(\dp.rf.rf[11][7] ),
    .S0(_02175_),
    .S1(_02176_),
    .Z(_02557_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06853_ (.I0(\dp.rf.rf[0][7] ),
    .I1(\dp.rf.rf[1][7] ),
    .I2(\dp.rf.rf[2][7] ),
    .I3(\dp.rf.rf[3][7] ),
    .S0(_02175_),
    .S1(_02176_),
    .Z(_02558_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06854_ (.I0(\dp.rf.rf[12][7] ),
    .I1(\dp.rf.rf[13][7] ),
    .I2(\dp.rf.rf[14][7] ),
    .I3(\dp.rf.rf[15][7] ),
    .S0(_01928_),
    .S1(_01929_),
    .Z(_02559_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06855_ (.I0(\dp.rf.rf[4][7] ),
    .I1(\dp.rf.rf[5][7] ),
    .I2(\dp.rf.rf[6][7] ),
    .I3(\dp.rf.rf[7][7] ),
    .S0(_01928_),
    .S1(_02176_),
    .Z(_02560_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06856_ (.I0(_02557_),
    .I1(_02558_),
    .I2(_02559_),
    .I3(_02560_),
    .S0(_01666_),
    .S1(_01400_),
    .Z(_02561_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06857_ (.I0(_02556_),
    .I1(_02561_),
    .S(_01058_),
    .Z(_02562_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _06858_ (.A1(_01608_),
    .A2(_02562_),
    .Z(net157));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06859_ (.A1(net16),
    .A2(_02409_),
    .Z(_05106_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06860_ (.I0(net157),
    .I1(_05106_),
    .S(_01605_),
    .Z(_02563_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _06861_ (.A1(_02229_),
    .A2(_02563_),
    .ZN(_05025_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06862_ (.I(_05025_),
    .ZN(_05029_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06863_ (.I0(\dp.rf.rf[2][7] ),
    .I1(\dp.rf.rf[3][7] ),
    .I2(\dp.rf.rf[6][7] ),
    .I3(\dp.rf.rf[7][7] ),
    .S0(_01363_),
    .S1(_01364_),
    .Z(_02564_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06864_ (.A1(_01362_),
    .A2(_02564_),
    .ZN(_02565_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06865_ (.I0(\dp.rf.rf[1][7] ),
    .I1(\dp.rf.rf[5][7] ),
    .S(_01138_),
    .Z(_02566_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06866_ (.A1(\dp.rf.rf[4][7] ),
    .A2(_01368_),
    .B1(_02566_),
    .B2(_01371_),
    .C(_01372_),
    .ZN(_02567_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _06867_ (.A1(_01854_),
    .A2(_02565_),
    .A3(_02567_),
    .ZN(_02568_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06868_ (.I0(\dp.rf.rf[10][7] ),
    .I1(\dp.rf.rf[11][7] ),
    .I2(\dp.rf.rf[14][7] ),
    .I3(\dp.rf.rf[15][7] ),
    .S0(_01128_),
    .S1(_01200_),
    .Z(_02569_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06869_ (.I0(\dp.rf.rf[8][7] ),
    .I1(\dp.rf.rf[9][7] ),
    .I2(\dp.rf.rf[12][7] ),
    .I3(\dp.rf.rf[13][7] ),
    .S0(_01128_),
    .S1(_01200_),
    .Z(_02570_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06870_ (.I0(_02569_),
    .I1(_02570_),
    .S(_01218_),
    .Z(_02571_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _06871_ (.A1(_01176_),
    .A2(_02571_),
    .Z(_02572_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _06872_ (.A1(_01376_),
    .A2(_02568_),
    .A3(_02572_),
    .Z(_02573_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06873_ (.I0(\dp.rf.rf[22][7] ),
    .I1(\dp.rf.rf[23][7] ),
    .S(_01600_),
    .Z(_02574_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06874_ (.I0(\dp.rf.rf[18][7] ),
    .I1(\dp.rf.rf[19][7] ),
    .S(_01212_),
    .Z(_02575_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06875_ (.A1(_01568_),
    .A2(_02574_),
    .B1(_02575_),
    .B2(_01593_),
    .C(_01456_),
    .ZN(_02576_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06876_ (.I(\dp.rf.rf[20][7] ),
    .ZN(_02577_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06877_ (.I0(\dp.rf.rf[17][7] ),
    .I1(\dp.rf.rf[21][7] ),
    .S(_01123_),
    .Z(_02578_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06878_ (.A1(_01328_),
    .A2(_02578_),
    .ZN(_02579_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _06879_ (.A1(_02577_),
    .A2(_01327_),
    .B(_02579_),
    .C(_01529_),
    .ZN(_02580_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _06880_ (.A1(\dp.rf.rf[16][7] ),
    .A2(_01356_),
    .B1(_02580_),
    .B2(net227),
    .ZN(_02581_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06881_ (.I0(\dp.rf.rf[30][7] ),
    .I1(\dp.rf.rf[31][7] ),
    .S(_01212_),
    .Z(_02582_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06882_ (.A1(\dp.rf.rf[26][7] ),
    .A2(net200),
    .Z(_02583_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06883_ (.A1(\dp.rf.rf[27][7] ),
    .A2(_01532_),
    .ZN(_02584_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06884_ (.A1(_01344_),
    .A2(_02584_),
    .ZN(_02585_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06885_ (.A1(_01339_),
    .A2(_02582_),
    .B1(_02583_),
    .B2(_02585_),
    .C(_01334_),
    .ZN(_02586_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06886_ (.I0(\dp.rf.rf[24][7] ),
    .I1(\dp.rf.rf[25][7] ),
    .I2(\dp.rf.rf[28][7] ),
    .I3(\dp.rf.rf[29][7] ),
    .S0(_01340_),
    .S1(_01169_),
    .Z(_02587_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06887_ (.A1(_01173_),
    .A2(_02587_),
    .B(_01176_),
    .ZN(_02588_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _06888_ (.A1(_02576_),
    .A2(_02581_),
    .B1(_02586_),
    .B2(_02588_),
    .C(net209),
    .ZN(_02589_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _06889_ (.A1(_02589_),
    .A2(_02573_),
    .Z(_05024_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _06890_ (.I(_05024_),
    .ZN(_05028_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06891_ (.I0(\dp.rf.rf[24][6] ),
    .I1(\dp.rf.rf[25][6] ),
    .I2(\dp.rf.rf[26][6] ),
    .I3(\dp.rf.rf[27][6] ),
    .S0(_01267_),
    .S1(_01263_),
    .Z(_02590_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06892_ (.I0(\dp.rf.rf[16][6] ),
    .I1(\dp.rf.rf[17][6] ),
    .I2(\dp.rf.rf[18][6] ),
    .I3(\dp.rf.rf[19][6] ),
    .S0(_01267_),
    .S1(_01268_),
    .Z(_02591_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06893_ (.I0(_02590_),
    .I1(_02591_),
    .S(_01282_),
    .Z(_02592_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06894_ (.I0(\dp.rf.rf[28][6] ),
    .I1(\dp.rf.rf[29][6] ),
    .I2(\dp.rf.rf[30][6] ),
    .I3(\dp.rf.rf[31][6] ),
    .S0(_01267_),
    .S1(_01268_),
    .Z(_02593_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06895_ (.I0(\dp.rf.rf[20][6] ),
    .I1(\dp.rf.rf[21][6] ),
    .I2(\dp.rf.rf[22][6] ),
    .I3(\dp.rf.rf[23][6] ),
    .S0(_01267_),
    .S1(_01268_),
    .Z(_02594_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06896_ (.I0(_02593_),
    .I1(_02594_),
    .S(_01282_),
    .Z(_02595_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06897_ (.I0(_02592_),
    .I1(_02595_),
    .S(_01478_),
    .Z(_02596_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06898_ (.I0(\dp.rf.rf[8][6] ),
    .I1(\dp.rf.rf[9][6] ),
    .I2(\dp.rf.rf[10][6] ),
    .I3(\dp.rf.rf[11][6] ),
    .S0(_01279_),
    .S1(_01276_),
    .Z(_02597_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06899_ (.I0(\dp.rf.rf[0][6] ),
    .I1(\dp.rf.rf[1][6] ),
    .I2(\dp.rf.rf[2][6] ),
    .I3(\dp.rf.rf[3][6] ),
    .S0(_01279_),
    .S1(_01276_),
    .Z(_02598_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06900_ (.I0(_02597_),
    .I1(_02598_),
    .S(_01282_),
    .Z(_02599_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06901_ (.I0(\dp.rf.rf[12][6] ),
    .I1(\dp.rf.rf[13][6] ),
    .I2(\dp.rf.rf[14][6] ),
    .I3(\dp.rf.rf[15][6] ),
    .S0(_01471_),
    .S1(_01316_),
    .Z(_02600_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06902_ (.I0(\dp.rf.rf[4][6] ),
    .I1(\dp.rf.rf[5][6] ),
    .I2(\dp.rf.rf[6][6] ),
    .I3(\dp.rf.rf[7][6] ),
    .S0(_01471_),
    .S1(_01316_),
    .Z(_02601_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06903_ (.I0(_02600_),
    .I1(_02601_),
    .S(_01282_),
    .Z(_02602_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06904_ (.I0(_02599_),
    .I1(_02602_),
    .S(_01478_),
    .Z(_02603_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _06905_ (.A1(_01111_),
    .A2(_02596_),
    .B1(_02603_),
    .B2(_01112_),
    .ZN(_02604_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06906_ (.I(_02604_),
    .ZN(net156));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06907_ (.A1(net15),
    .A2(_02409_),
    .Z(_05102_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06908_ (.I0(net156),
    .I1(_05102_),
    .S(_01605_),
    .Z(_02605_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _06909_ (.A1(_02229_),
    .A2(_02605_),
    .ZN(_05033_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06910_ (.I(_05033_),
    .ZN(_05037_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06911_ (.I0(\dp.rf.rf[17][6] ),
    .I1(\dp.rf.rf[21][6] ),
    .S(_01145_),
    .Z(_02606_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06912_ (.A1(_01693_),
    .A2(_02606_),
    .ZN(_02607_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _06913_ (.A1(\dp.rf.rf[16][6] ),
    .A2(_01600_),
    .A3(_01145_),
    .Z(_02608_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06914_ (.A1(\dp.rf.rf[20][6] ),
    .A2(_01504_),
    .A3(_01339_),
    .B(_02608_),
    .ZN(_02609_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06915_ (.A1(_01530_),
    .A2(_02607_),
    .A3(_02609_),
    .B(_01415_),
    .ZN(_02610_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06916_ (.I0(\dp.rf.rf[18][6] ),
    .I1(\dp.rf.rf[19][6] ),
    .I2(\dp.rf.rf[22][6] ),
    .I3(\dp.rf.rf[23][6] ),
    .S0(_01157_),
    .S1(_01139_),
    .Z(_02611_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _06917_ (.A1(_01456_),
    .A2(_01244_),
    .A3(_01435_),
    .A4(_02611_),
    .Z(_02612_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06918_ (.A1(net205),
    .A2(_02610_),
    .B(_02612_),
    .ZN(_02613_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06919_ (.I0(\dp.rf.rf[30][6] ),
    .I1(\dp.rf.rf[31][6] ),
    .S(_01600_),
    .Z(_02614_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06920_ (.I(_02614_),
    .ZN(_02615_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06921_ (.A1(_01211_),
    .A2(_02615_),
    .B(_02019_),
    .ZN(_02616_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _06922_ (.A1(\dp.rf.rf[26][6] ),
    .A2(_01154_),
    .A3(_01155_),
    .A4(_01090_),
    .ZN(_02617_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06923_ (.I(\dp.rf.rf[26][6] ),
    .ZN(_02618_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _06924_ (.A1(_01028_),
    .A2(_01185_),
    .A3(_02617_),
    .B1(_01569_),
    .B2(_02618_),
    .ZN(_02619_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06925_ (.A1(\dp.rf.rf[27][6] ),
    .A2(_01645_),
    .Z(_02620_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _06926_ (.A1(_01164_),
    .A2(_01166_),
    .A3(_02619_),
    .A4(_02620_),
    .Z(_02621_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06927_ (.I0(\dp.rf.rf[24][6] ),
    .I1(\dp.rf.rf[25][6] ),
    .I2(\dp.rf.rf[28][6] ),
    .I3(\dp.rf.rf[29][6] ),
    .S0(_01569_),
    .S1(_01146_),
    .Z(_02622_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _06928_ (.A1(_02616_),
    .A2(_02621_),
    .B1(_02622_),
    .B2(_01576_),
    .C(_01580_),
    .ZN(_02623_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06929_ (.I0(\dp.rf.rf[10][6] ),
    .I1(\dp.rf.rf[11][6] ),
    .I2(\dp.rf.rf[14][6] ),
    .I3(\dp.rf.rf[15][6] ),
    .S0(_01136_),
    .S1(_01139_),
    .Z(_02624_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06930_ (.I0(\dp.rf.rf[8][6] ),
    .I1(\dp.rf.rf[9][6] ),
    .I2(\dp.rf.rf[12][6] ),
    .I3(\dp.rf.rf[13][6] ),
    .S0(_01136_),
    .S1(_01139_),
    .Z(_02625_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06931_ (.I0(_02624_),
    .I1(_02625_),
    .S(_01889_),
    .Z(_02626_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _06932_ (.A1(\dp.rf.rf[4][6] ),
    .A2(_01504_),
    .A3(_01505_),
    .ZN(_02627_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06933_ (.I0(\dp.rf.rf[1][6] ),
    .I1(\dp.rf.rf[5][6] ),
    .S(_01432_),
    .Z(_02628_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06934_ (.A1(_01422_),
    .A2(_02628_),
    .ZN(_02629_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06935_ (.I0(\dp.rf.rf[2][6] ),
    .I1(\dp.rf.rf[3][6] ),
    .I2(\dp.rf.rf[6][6] ),
    .I3(\dp.rf.rf[7][6] ),
    .S0(_01160_),
    .S1(_01145_),
    .Z(_02630_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06936_ (.A1(_01456_),
    .A2(_02630_),
    .ZN(_02631_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06937_ (.A1(_01530_),
    .A2(_02627_),
    .A3(_02629_),
    .B(_02631_),
    .ZN(_02632_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _06938_ (.A1(_01580_),
    .A2(_02626_),
    .B1(_02632_),
    .B2(_01541_),
    .C(_01376_),
    .ZN(_02633_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _06939_ (.A1(_02613_),
    .A2(_02623_),
    .B(_02633_),
    .ZN(_05032_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _06940_ (.I(_05032_),
    .ZN(_05036_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06941_ (.I0(\dp.rf.rf[24][5] ),
    .I1(\dp.rf.rf[25][5] ),
    .I2(\dp.rf.rf[26][5] ),
    .I3(\dp.rf.rf[27][5] ),
    .S0(_01098_),
    .S1(_01554_),
    .Z(_02634_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06942_ (.I0(\dp.rf.rf[16][5] ),
    .I1(\dp.rf.rf[17][5] ),
    .I2(\dp.rf.rf[18][5] ),
    .I3(\dp.rf.rf[19][5] ),
    .S0(_01098_),
    .S1(_01554_),
    .Z(_02635_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06943_ (.I0(\dp.rf.rf[28][5] ),
    .I1(\dp.rf.rf[29][5] ),
    .I2(\dp.rf.rf[30][5] ),
    .I3(\dp.rf.rf[31][5] ),
    .S0(_01098_),
    .S1(_01554_),
    .Z(_02636_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06944_ (.I0(\dp.rf.rf[20][5] ),
    .I1(\dp.rf.rf[21][5] ),
    .I2(\dp.rf.rf[22][5] ),
    .I3(\dp.rf.rf[23][5] ),
    .S0(_01098_),
    .S1(_01554_),
    .Z(_02637_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06945_ (.I0(_02634_),
    .I1(_02635_),
    .I2(_02636_),
    .I3(_02637_),
    .S0(_01398_),
    .S1(net194),
    .Z(_02638_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06946_ (.I0(\dp.rf.rf[8][5] ),
    .I1(\dp.rf.rf[9][5] ),
    .I2(\dp.rf.rf[10][5] ),
    .I3(\dp.rf.rf[11][5] ),
    .S0(_01098_),
    .S1(_01554_),
    .Z(_02639_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06947_ (.I0(\dp.rf.rf[0][5] ),
    .I1(\dp.rf.rf[1][5] ),
    .I2(\dp.rf.rf[2][5] ),
    .I3(\dp.rf.rf[3][5] ),
    .S0(_01098_),
    .S1(_01554_),
    .Z(_02640_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06948_ (.I0(\dp.rf.rf[12][5] ),
    .I1(\dp.rf.rf[13][5] ),
    .I2(\dp.rf.rf[14][5] ),
    .I3(\dp.rf.rf[15][5] ),
    .S0(_01260_),
    .S1(_02326_),
    .Z(_02641_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06949_ (.I0(\dp.rf.rf[4][5] ),
    .I1(\dp.rf.rf[5][5] ),
    .I2(\dp.rf.rf[6][5] ),
    .I3(\dp.rf.rf[7][5] ),
    .S0(_01098_),
    .S1(_01554_),
    .Z(_02642_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06950_ (.I0(_02639_),
    .I1(_02640_),
    .I2(_02641_),
    .I3(_02642_),
    .S0(_01271_),
    .S1(net194),
    .Z(_02643_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06951_ (.I0(_02638_),
    .I1(_02643_),
    .S(_01058_),
    .Z(_02644_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _06952_ (.A1(net192),
    .A2(_02644_),
    .Z(net155));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06953_ (.A1(net14),
    .A2(_02409_),
    .Z(_05098_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06954_ (.I0(net155),
    .I1(_05098_),
    .S(_01605_),
    .Z(_02645_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _06955_ (.A1(_02229_),
    .A2(_02645_),
    .ZN(_05041_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06956_ (.I(_05041_),
    .ZN(_05045_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06957_ (.I0(\dp.rf.rf[17][5] ),
    .I1(\dp.rf.rf[21][5] ),
    .S(_01200_),
    .Z(_02646_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06958_ (.A1(_01636_),
    .A2(_02646_),
    .ZN(_02647_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06959_ (.A1(\dp.rf.rf[20][5] ),
    .A2(_01600_),
    .A3(_01196_),
    .B(_01193_),
    .ZN(_02648_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _06960_ (.A1(_02647_),
    .A2(_02648_),
    .B(_01228_),
    .C(_01192_),
    .ZN(_02649_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06961_ (.I(\dp.rf.rf[16][5] ),
    .ZN(_02650_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06962_ (.A1(_02650_),
    .A2(_01736_),
    .ZN(_02651_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06963_ (.I0(\dp.rf.rf[18][5] ),
    .I1(\dp.rf.rf[19][5] ),
    .S(_01186_),
    .Z(_02652_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06964_ (.I(_02652_),
    .ZN(_02653_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06965_ (.I0(\dp.rf.rf[22][5] ),
    .I1(\dp.rf.rf[23][5] ),
    .S(_01427_),
    .Z(_02654_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06966_ (.A1(_01182_),
    .A2(_02654_),
    .B(_01118_),
    .ZN(_02655_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06967_ (.A1(_01344_),
    .A2(_02653_),
    .B(_02655_),
    .ZN(_02656_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06968_ (.A1(_02649_),
    .A2(_02651_),
    .B(_02656_),
    .ZN(_02657_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06969_ (.I0(\dp.rf.rf[26][5] ),
    .I1(\dp.rf.rf[27][5] ),
    .I2(\dp.rf.rf[30][5] ),
    .I3(\dp.rf.rf[31][5] ),
    .S0(_01427_),
    .S1(_01168_),
    .Z(_02658_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06970_ (.I0(\dp.rf.rf[24][5] ),
    .I1(\dp.rf.rf[25][5] ),
    .I2(\dp.rf.rf[28][5] ),
    .I3(\dp.rf.rf[29][5] ),
    .S0(_01427_),
    .S1(_01168_),
    .Z(_02659_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06971_ (.I0(_02658_),
    .I1(_02659_),
    .S(_01218_),
    .Z(_02660_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06972_ (.A1(_01337_),
    .A2(_02660_),
    .ZN(_02661_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _06973_ (.A1(\dp.rf.rf[4][5] ),
    .A2(_01645_),
    .A3(_01182_),
    .ZN(_02662_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06974_ (.I0(\dp.rf.rf[1][5] ),
    .I1(\dp.rf.rf[5][5] ),
    .S(_01144_),
    .Z(_02663_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06975_ (.A1(_01371_),
    .A2(_02663_),
    .ZN(_02664_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06976_ (.I0(\dp.rf.rf[2][5] ),
    .I1(\dp.rf.rf[3][5] ),
    .I2(\dp.rf.rf[6][5] ),
    .I3(\dp.rf.rf[7][5] ),
    .S0(_01194_),
    .S1(_01369_),
    .Z(_02665_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06977_ (.A1(_01213_),
    .A2(_02665_),
    .ZN(_02666_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06978_ (.A1(_01416_),
    .A2(_02662_),
    .A3(_02664_),
    .B(_02666_),
    .ZN(_02667_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06979_ (.I0(\dp.rf.rf[10][5] ),
    .I1(\dp.rf.rf[11][5] ),
    .I2(\dp.rf.rf[14][5] ),
    .I3(\dp.rf.rf[15][5] ),
    .S0(_01194_),
    .S1(_01138_),
    .Z(_02668_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06980_ (.I0(\dp.rf.rf[8][5] ),
    .I1(\dp.rf.rf[9][5] ),
    .I2(\dp.rf.rf[12][5] ),
    .I3(\dp.rf.rf[13][5] ),
    .S0(_01194_),
    .S1(_01138_),
    .Z(_02669_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06981_ (.I0(_02668_),
    .I1(_02669_),
    .S(_01218_),
    .Z(_02670_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _06982_ (.A1(_01541_),
    .A2(_02667_),
    .B1(_02670_),
    .B2(_01176_),
    .C(_01376_),
    .ZN(_02671_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _06983_ (.A1(net209),
    .A2(_02657_),
    .A3(_02661_),
    .B(_02671_),
    .ZN(_05040_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _06984_ (.I(_05040_),
    .ZN(_05044_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _06985_ (.I(net3),
    .ZN(_02672_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06986_ (.A1(_02672_),
    .A2(net94),
    .Z(_02673_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _06987_ (.A1(_01111_),
    .A2(_01291_),
    .B(_01109_),
    .C(_01078_),
    .ZN(_02674_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _06988_ (.A1(_01438_),
    .A2(net231),
    .A3(_01081_),
    .Z(_02675_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _06989_ (.A1(_01037_),
    .A2(net21),
    .A3(_01090_),
    .ZN(_02676_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06990_ (.A1(_02672_),
    .A2(_01064_),
    .B(_02676_),
    .ZN(_02677_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06991_ (.A1(_02675_),
    .A2(_02677_),
    .ZN(_02678_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _06992_ (.A1(_02673_),
    .A2(_02674_),
    .B(_02678_),
    .ZN(_05094_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06993_ (.I0(\dp.rf.rf[4][4] ),
    .I1(\dp.rf.rf[5][4] ),
    .I2(\dp.rf.rf[6][4] ),
    .I3(\dp.rf.rf[7][4] ),
    .S0(_01484_),
    .S1(_02232_),
    .Z(_02679_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06994_ (.I0(\dp.rf.rf[0][4] ),
    .I1(\dp.rf.rf[1][4] ),
    .I2(\dp.rf.rf[2][4] ),
    .I3(\dp.rf.rf[3][4] ),
    .S0(_01661_),
    .S1(_02232_),
    .Z(_02680_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06995_ (.I0(_02679_),
    .I1(_02680_),
    .S(_01779_),
    .Z(_02681_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06996_ (.A1(_01677_),
    .A2(_02681_),
    .B(_01607_),
    .ZN(_02682_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06997_ (.I(_01778_),
    .ZN(_02683_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06998_ (.I0(\dp.rf.rf[22][4] ),
    .I1(\dp.rf.rf[23][4] ),
    .I2(\dp.rf.rf[30][4] ),
    .I3(\dp.rf.rf[31][4] ),
    .S0(_01402_),
    .S1(_01671_),
    .Z(_02684_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06999_ (.I0(\dp.rf.rf[20][4] ),
    .I1(\dp.rf.rf[21][4] ),
    .I2(\dp.rf.rf[28][4] ),
    .I3(\dp.rf.rf[29][4] ),
    .S0(_01402_),
    .S1(_01671_),
    .Z(_02685_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07000_ (.I0(_02684_),
    .I1(_02685_),
    .S(_01766_),
    .Z(_02686_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07001_ (.I0(\dp.rf.rf[24][4] ),
    .I1(\dp.rf.rf[25][4] ),
    .I2(\dp.rf.rf[26][4] ),
    .I3(\dp.rf.rf[27][4] ),
    .S0(_01657_),
    .S1(_01408_),
    .Z(_02687_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07002_ (.I0(\dp.rf.rf[16][4] ),
    .I1(\dp.rf.rf[17][4] ),
    .I2(\dp.rf.rf[18][4] ),
    .I3(\dp.rf.rf[19][4] ),
    .S0(_01657_),
    .S1(_01408_),
    .Z(_02688_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07003_ (.I0(_02687_),
    .I1(_02688_),
    .S(_01398_),
    .Z(_02689_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07004_ (.A1(_01037_),
    .A2(_01779_),
    .ZN(_02690_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _07005_ (.A1(_02683_),
    .A2(_02686_),
    .B1(_02689_),
    .B2(_02690_),
    .ZN(_02691_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07006_ (.I0(\dp.rf.rf[12][4] ),
    .I1(\dp.rf.rf[13][4] ),
    .I2(\dp.rf.rf[14][4] ),
    .I3(\dp.rf.rf[15][4] ),
    .S0(_01661_),
    .S1(_02232_),
    .Z(_02692_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07007_ (.I0(\dp.rf.rf[8][4] ),
    .I1(\dp.rf.rf[9][4] ),
    .I2(\dp.rf.rf[10][4] ),
    .I3(\dp.rf.rf[11][4] ),
    .S0(_01661_),
    .S1(_02232_),
    .Z(_02693_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07008_ (.I0(_02692_),
    .I1(_02693_),
    .S(_01779_),
    .Z(_02694_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07009_ (.A1(_01672_),
    .A2(_02694_),
    .ZN(_02695_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _07010_ (.A1(_02682_),
    .A2(_02691_),
    .A3(_02695_),
    .Z(_02696_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07011_ (.I(_02696_),
    .ZN(net154));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _07012_ (.I0(_05094_),
    .I1(net154),
    .S(_01289_),
    .Z(_02697_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer22 (.I(_05008_),
    .Z(net181));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07014_ (.I(_02697_),
    .Z(_02699_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _07015_ (.A1(_02229_),
    .A2(_02699_),
    .ZN(_05049_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07016_ (.I(_05049_),
    .ZN(_05053_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07017_ (.I0(\dp.rf.rf[2][4] ),
    .I1(\dp.rf.rf[3][4] ),
    .I2(\dp.rf.rf[6][4] ),
    .I3(\dp.rf.rf[7][4] ),
    .S0(_01225_),
    .S1(_01381_),
    .Z(_02700_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07018_ (.A1(_01119_),
    .A2(_02700_),
    .Z(_02701_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07019_ (.I(\dp.rf.rf[4][4] ),
    .ZN(_02702_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07020_ (.I0(\dp.rf.rf[1][4] ),
    .I1(\dp.rf.rf[5][4] ),
    .S(_01200_),
    .Z(_02703_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07021_ (.A1(_01636_),
    .A2(_02703_),
    .ZN(_02704_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _07022_ (.A1(_02702_),
    .A2(_01327_),
    .B(_02704_),
    .C(_01529_),
    .ZN(_02705_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07023_ (.I0(\dp.rf.rf[10][4] ),
    .I1(\dp.rf.rf[11][4] ),
    .I2(\dp.rf.rf[14][4] ),
    .I3(\dp.rf.rf[15][4] ),
    .S0(_01120_),
    .S1(_01129_),
    .Z(_02706_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07024_ (.I0(\dp.rf.rf[8][4] ),
    .I1(\dp.rf.rf[9][4] ),
    .I2(\dp.rf.rf[12][4] ),
    .I3(\dp.rf.rf[13][4] ),
    .S0(_01120_),
    .S1(_01129_),
    .Z(_02707_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07025_ (.I0(_02706_),
    .I1(_02707_),
    .S(_01171_),
    .Z(_02708_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07026_ (.A1(_01199_),
    .A2(_02708_),
    .Z(_02709_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07027_ (.A1(_01541_),
    .A2(_02701_),
    .A3(_02705_),
    .B(_02709_),
    .ZN(_02710_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07028_ (.I0(\dp.rf.rf[17][4] ),
    .I1(\dp.rf.rf[21][4] ),
    .S(_01138_),
    .Z(_02711_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07029_ (.A1(_01442_),
    .A2(_02711_),
    .ZN(_02712_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07030_ (.A1(\dp.rf.rf[20][4] ),
    .A2(_01577_),
    .A3(_01182_),
    .B(_01241_),
    .ZN(_02713_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07031_ (.A1(_02712_),
    .A2(_02713_),
    .B(_01228_),
    .C(net168),
    .ZN(_02714_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07032_ (.I(\dp.rf.rf[16][4] ),
    .ZN(_02715_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07033_ (.A1(_02715_),
    .A2(_01737_),
    .ZN(_02716_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07034_ (.I0(\dp.rf.rf[18][4] ),
    .I1(\dp.rf.rf[19][4] ),
    .S(_01225_),
    .Z(_02717_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07035_ (.I(_02717_),
    .ZN(_02718_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07036_ (.I0(\dp.rf.rf[22][4] ),
    .I1(\dp.rf.rf[23][4] ),
    .S(_01135_),
    .Z(_02719_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07037_ (.A1(_01182_),
    .A2(_02719_),
    .ZN(_02720_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _07038_ (.A1(_01224_),
    .A2(_02718_),
    .B(_02720_),
    .C(_01151_),
    .ZN(_02721_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07039_ (.A1(_02714_),
    .A2(_02716_),
    .B(_02721_),
    .ZN(_02722_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07040_ (.I0(\dp.rf.rf[26][4] ),
    .I1(\dp.rf.rf[27][4] ),
    .I2(\dp.rf.rf[30][4] ),
    .I3(\dp.rf.rf[31][4] ),
    .S0(_01186_),
    .S1(_01457_),
    .Z(_02723_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07041_ (.I0(\dp.rf.rf[24][4] ),
    .I1(\dp.rf.rf[25][4] ),
    .I2(\dp.rf.rf[28][4] ),
    .I3(\dp.rf.rf[29][4] ),
    .S0(_01186_),
    .S1(_01457_),
    .Z(_02724_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07042_ (.I0(_02723_),
    .I1(_02724_),
    .S(_01241_),
    .Z(_02725_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07043_ (.A1(_01415_),
    .A2(_02725_),
    .B(_01206_),
    .ZN(_02726_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _07044_ (.A1(_01589_),
    .A2(_02710_),
    .B1(_02722_),
    .B2(_02726_),
    .ZN(_05048_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _07045_ (.I(_05048_),
    .ZN(_05052_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07046_ (.A1(net21),
    .A2(_01034_),
    .Z(_02727_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07047_ (.A1(net2),
    .A2(_01035_),
    .B1(_02727_),
    .B2(_01761_),
    .ZN(_02728_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07048_ (.A1(_01107_),
    .A2(_02728_),
    .ZN(_02729_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07049_ (.A1(_01028_),
    .A2(_01029_),
    .ZN(_02730_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07050_ (.A1(net230),
    .A2(_01035_),
    .B1(_01294_),
    .B2(net24),
    .ZN(_02731_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _07051_ (.A1(_02730_),
    .A2(_02731_),
    .B(_01078_),
    .ZN(_02732_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07052_ (.A1(net2),
    .A2(_01078_),
    .B1(_02675_),
    .B2(_02677_),
    .ZN(_02733_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _07053_ (.A1(_01030_),
    .A2(_01095_),
    .B(_01245_),
    .C(_01761_),
    .ZN(_02734_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _07054_ (.A1(_02732_),
    .A2(_02733_),
    .B(_02734_),
    .C(net236),
    .ZN(_02735_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07055_ (.A1(_02729_),
    .A2(_02735_),
    .Z(_05088_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07056_ (.I0(\dp.rf.rf[24][3] ),
    .I1(\dp.rf.rf[25][3] ),
    .I2(\dp.rf.rf[26][3] ),
    .I3(\dp.rf.rf[27][3] ),
    .S0(_01275_),
    .S1(_01268_),
    .Z(_02736_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07057_ (.I0(\dp.rf.rf[16][3] ),
    .I1(\dp.rf.rf[17][3] ),
    .I2(\dp.rf.rf[18][3] ),
    .I3(\dp.rf.rf[19][3] ),
    .S0(_01267_),
    .S1(_01268_),
    .Z(_02737_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07058_ (.I0(\dp.rf.rf[28][3] ),
    .I1(\dp.rf.rf[29][3] ),
    .I2(\dp.rf.rf[30][3] ),
    .I3(\dp.rf.rf[31][3] ),
    .S0(_01279_),
    .S1(_01276_),
    .Z(_02738_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07059_ (.I0(\dp.rf.rf[20][3] ),
    .I1(\dp.rf.rf[21][3] ),
    .I2(\dp.rf.rf[22][3] ),
    .I3(\dp.rf.rf[23][3] ),
    .S0(_01275_),
    .S1(_01268_),
    .Z(_02739_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07060_ (.I0(_02736_),
    .I1(_02737_),
    .I2(_02738_),
    .I3(_02739_),
    .S0(_01282_),
    .S1(net194),
    .Z(_02740_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07061_ (.I0(\dp.rf.rf[8][3] ),
    .I1(\dp.rf.rf[9][3] ),
    .I2(\dp.rf.rf[10][3] ),
    .I3(\dp.rf.rf[11][3] ),
    .S0(_01275_),
    .S1(_01276_),
    .Z(_02741_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07062_ (.I0(\dp.rf.rf[0][3] ),
    .I1(\dp.rf.rf[1][3] ),
    .I2(\dp.rf.rf[2][3] ),
    .I3(\dp.rf.rf[3][3] ),
    .S0(_01275_),
    .S1(_01268_),
    .Z(_02742_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07063_ (.I0(\dp.rf.rf[12][3] ),
    .I1(\dp.rf.rf[13][3] ),
    .I2(\dp.rf.rf[14][3] ),
    .I3(\dp.rf.rf[15][3] ),
    .S0(_01279_),
    .S1(_01276_),
    .Z(_02743_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07064_ (.I0(\dp.rf.rf[4][3] ),
    .I1(\dp.rf.rf[5][3] ),
    .I2(\dp.rf.rf[6][3] ),
    .I3(\dp.rf.rf[7][3] ),
    .S0(_01279_),
    .S1(_01276_),
    .Z(_02744_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07065_ (.I0(_02741_),
    .I1(_02742_),
    .I2(_02743_),
    .I3(_02744_),
    .S0(_01282_),
    .S1(net194),
    .Z(_02745_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07066_ (.I0(_02740_),
    .I1(_02745_),
    .S(_01058_),
    .Z(_02746_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07067_ (.A1(_01608_),
    .A2(_02746_),
    .Z(net153));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _07068_ (.A1(_02735_),
    .A2(_02729_),
    .B(_01093_),
    .ZN(_02747_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _07069_ (.A1(net153),
    .A2(_01259_),
    .ZN(_02748_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _07070_ (.A1(_02747_),
    .A2(_02748_),
    .ZN(_02749_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _07071_ (.I(_02749_),
    .Z(_02750_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 split9 (.I(_01077_),
    .Z(net168));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 split28 (.I(net253),
    .Z(net187));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _07074_ (.A1(_02229_),
    .A2(_02750_),
    .ZN(_05057_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07075_ (.I(_05057_),
    .ZN(_05061_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07076_ (.I0(\dp.rf.rf[30][3] ),
    .I1(\dp.rf.rf[31][3] ),
    .S(_01212_),
    .Z(_02753_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07077_ (.A1(\dp.rf.rf[26][3] ),
    .A2(_01626_),
    .Z(_02754_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07078_ (.A1(\dp.rf.rf[27][3] ),
    .A2(_01532_),
    .ZN(_02755_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07079_ (.A1(_01344_),
    .A2(_02755_),
    .ZN(_02756_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _07080_ (.A1(_01339_),
    .A2(_02753_),
    .B1(_02754_),
    .B2(_02756_),
    .C(_01334_),
    .ZN(_02757_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07081_ (.I0(\dp.rf.rf[24][3] ),
    .I1(\dp.rf.rf[25][3] ),
    .I2(\dp.rf.rf[28][3] ),
    .I3(\dp.rf.rf[29][3] ),
    .S0(_01340_),
    .S1(_01169_),
    .Z(_02758_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07082_ (.A1(_01173_),
    .A2(_02758_),
    .B(net209),
    .ZN(_02759_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07083_ (.A1(_02757_),
    .A2(_02759_),
    .Z(_02760_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07084_ (.I0(\dp.rf.rf[9][3] ),
    .I1(\dp.rf.rf[13][3] ),
    .S(_01369_),
    .Z(_02761_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _07085_ (.A1(\dp.rf.rf[12][3] ),
    .A2(_01368_),
    .B1(_02761_),
    .B2(_01442_),
    .C(_01430_),
    .ZN(_02762_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07086_ (.A1(_01141_),
    .A2(_01130_),
    .ZN(_02763_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07087_ (.A1(_01077_),
    .A2(_02763_),
    .ZN(_02764_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07088_ (.I(\dp.rf.rf[8][3] ),
    .ZN(_02765_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07089_ (.A1(net267),
    .A2(_02762_),
    .B1(_02764_),
    .B2(_02765_),
    .ZN(_02766_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07090_ (.A1(\dp.rf.rf[11][3] ),
    .A2(_01340_),
    .Z(_02767_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _07091_ (.A1(_01578_),
    .A2(_01077_),
    .B1(_01626_),
    .B2(\dp.rf.rf[10][3] ),
    .C(_02767_),
    .ZN(_02768_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07092_ (.I0(\dp.rf.rf[14][3] ),
    .I1(\dp.rf.rf[15][3] ),
    .S(_01160_),
    .Z(_02769_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07093_ (.A1(_01505_),
    .A2(_02769_),
    .ZN(_02770_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _07094_ (.A1(_01500_),
    .A2(_02768_),
    .A3(_02770_),
    .ZN(_02771_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07095_ (.A1(_02766_),
    .A2(_02771_),
    .B(_01385_),
    .ZN(_02772_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07096_ (.A1(_01530_),
    .A2(_02763_),
    .B(_01361_),
    .ZN(_02773_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07097_ (.I0(\dp.rf.rf[6][3] ),
    .I1(\dp.rf.rf[7][3] ),
    .S(_01508_),
    .Z(_02774_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07098_ (.A1(_01505_),
    .A2(_02774_),
    .ZN(_02775_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07099_ (.A1(\dp.rf.rf[3][3] ),
    .A2(_01428_),
    .Z(_02776_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _07100_ (.A1(_01533_),
    .A2(_01192_),
    .B1(_01626_),
    .B2(\dp.rf.rf[2][3] ),
    .C(_02776_),
    .ZN(_02777_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _07101_ (.A1(_02019_),
    .A2(_02775_),
    .A3(_02777_),
    .ZN(_02778_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07102_ (.I(\dp.rf.rf[0][3] ),
    .ZN(_02779_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07103_ (.I0(\dp.rf.rf[1][3] ),
    .I1(\dp.rf.rf[5][3] ),
    .S(_01168_),
    .Z(_02780_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _07104_ (.A1(\dp.rf.rf[4][3] ),
    .A2(_01496_),
    .B1(_02780_),
    .B2(_01371_),
    .C(_01172_),
    .ZN(_02781_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07105_ (.A1(_02779_),
    .A2(_02764_),
    .B1(_02781_),
    .B2(net267),
    .ZN(_02782_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07106_ (.A1(\dp.rf.rf[19][3] ),
    .A2(_01508_),
    .Z(_02783_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _07107_ (.A1(_01210_),
    .A2(_01192_),
    .B1(_01626_),
    .B2(\dp.rf.rf[18][3] ),
    .C(_02783_),
    .ZN(_02784_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07108_ (.I0(\dp.rf.rf[22][3] ),
    .I1(\dp.rf.rf[23][3] ),
    .S(_01363_),
    .Z(_02785_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07109_ (.A1(_01505_),
    .A2(_02785_),
    .ZN(_02786_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07110_ (.I0(\dp.rf.rf[16][3] ),
    .I1(\dp.rf.rf[17][3] ),
    .I2(\dp.rf.rf[20][3] ),
    .I3(\dp.rf.rf[21][3] ),
    .S0(_01531_),
    .S1(_01443_),
    .Z(_02787_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07111_ (.A1(_01430_),
    .A2(_02787_),
    .B(net207),
    .ZN(_02788_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07112_ (.A1(_02019_),
    .A2(_02784_),
    .A3(_02786_),
    .B(_02788_),
    .ZN(_02789_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07113_ (.A1(_02778_),
    .A2(_02782_),
    .B(_02789_),
    .ZN(_02790_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _07114_ (.A1(_02760_),
    .A2(_02772_),
    .B1(_02790_),
    .B2(_02773_),
    .ZN(_05056_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _07115_ (.I(_05056_),
    .ZN(_05060_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07116_ (.A1(net27),
    .A2(_01035_),
    .B1(_02727_),
    .B2(_01047_),
    .ZN(_02791_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07117_ (.A1(_01107_),
    .A2(_02791_),
    .ZN(_02792_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _07118_ (.I(net27),
    .ZN(_02793_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _07119_ (.A1(_02793_),
    .A2(_01245_),
    .B1(_01107_),
    .B2(_02728_),
    .ZN(_02794_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07120_ (.I0(_01312_),
    .I1(_02794_),
    .S(_02732_),
    .Z(_02795_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07121_ (.A1(_01109_),
    .A2(_02795_),
    .Z(_02796_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07122_ (.A1(_02792_),
    .A2(_02796_),
    .Z(_05084_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07123_ (.I0(\dp.rf.rf[24][2] ),
    .I1(\dp.rf.rf[25][2] ),
    .I2(\dp.rf.rf[26][2] ),
    .I3(\dp.rf.rf[27][2] ),
    .S0(_01260_),
    .S1(_02326_),
    .Z(_02797_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07124_ (.I0(\dp.rf.rf[16][2] ),
    .I1(\dp.rf.rf[17][2] ),
    .I2(\dp.rf.rf[18][2] ),
    .I3(\dp.rf.rf[19][2] ),
    .S0(_01260_),
    .S1(_02326_),
    .Z(_02798_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07125_ (.I0(_02797_),
    .I1(_02798_),
    .S(_01271_),
    .Z(_02799_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07126_ (.I0(\dp.rf.rf[28][2] ),
    .I1(\dp.rf.rf[29][2] ),
    .I2(\dp.rf.rf[30][2] ),
    .I3(\dp.rf.rf[31][2] ),
    .S0(_01260_),
    .S1(_02326_),
    .Z(_02800_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07127_ (.I0(\dp.rf.rf[20][2] ),
    .I1(\dp.rf.rf[21][2] ),
    .I2(\dp.rf.rf[22][2] ),
    .I3(\dp.rf.rf[23][2] ),
    .S0(_01266_),
    .S1(_02326_),
    .Z(_02801_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07128_ (.I0(_02800_),
    .I1(_02801_),
    .S(_01271_),
    .Z(_02802_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07129_ (.I0(_02799_),
    .I1(_02802_),
    .S(net194),
    .Z(_02803_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07130_ (.I0(\dp.rf.rf[8][2] ),
    .I1(\dp.rf.rf[9][2] ),
    .I2(\dp.rf.rf[10][2] ),
    .I3(\dp.rf.rf[11][2] ),
    .S0(_01266_),
    .S1(_02326_),
    .Z(_02804_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07131_ (.I0(\dp.rf.rf[0][2] ),
    .I1(\dp.rf.rf[1][2] ),
    .I2(\dp.rf.rf[2][2] ),
    .I3(\dp.rf.rf[3][2] ),
    .S0(_01266_),
    .S1(_01262_),
    .Z(_02805_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07132_ (.I0(_02804_),
    .I1(_02805_),
    .S(_01271_),
    .Z(_02806_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07133_ (.I0(\dp.rf.rf[12][2] ),
    .I1(\dp.rf.rf[13][2] ),
    .I2(\dp.rf.rf[14][2] ),
    .I3(\dp.rf.rf[15][2] ),
    .S0(_01266_),
    .S1(_01262_),
    .Z(_02807_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07134_ (.I0(\dp.rf.rf[4][2] ),
    .I1(\dp.rf.rf[5][2] ),
    .I2(\dp.rf.rf[6][2] ),
    .I3(\dp.rf.rf[7][2] ),
    .S0(_01266_),
    .S1(_01262_),
    .Z(_02808_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07135_ (.I0(_02807_),
    .I1(_02808_),
    .S(_01271_),
    .Z(_02809_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07136_ (.I0(_02806_),
    .I1(_02809_),
    .S(net194),
    .Z(_02810_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _07137_ (.A1(_01037_),
    .A2(_02803_),
    .B1(_02810_),
    .B2(_01061_),
    .ZN(_02811_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07138_ (.I(_02811_),
    .ZN(net150));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _07139_ (.A1(_02795_),
    .A2(_01109_),
    .B(_02792_),
    .C(_01259_),
    .ZN(_02812_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07140_ (.A1(_01259_),
    .A2(_02811_),
    .Z(_02813_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _07141_ (.A1(_02812_),
    .A2(_02813_),
    .ZN(_02814_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 split16 (.I(_02816_),
    .Z(net175));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 _07143_ (.I(_02814_),
    .Z(_02816_));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer5 (.I(_02891_),
    .Z(net164));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _07145_ (.A1(net245),
    .A2(_02816_),
    .ZN(_05065_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07146_ (.I(_05065_),
    .ZN(_05069_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07147_ (.I0(\dp.rf.rf[6][2] ),
    .I1(\dp.rf.rf[7][2] ),
    .S(_01135_),
    .Z(_02818_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07148_ (.I(_02818_),
    .ZN(_02819_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07149_ (.A1(_01533_),
    .A2(_02819_),
    .B(_01151_),
    .ZN(_02820_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _07150_ (.A1(\dp.rf.rf[2][2] ),
    .A2(net10),
    .A3(net1),
    .A4(_01033_),
    .ZN(_02821_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07151_ (.I(\dp.rf.rf[2][2] ),
    .ZN(_02822_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _07152_ (.A1(_01028_),
    .A2(_01153_),
    .A3(_02821_),
    .B1(_01147_),
    .B2(_02822_),
    .ZN(_02823_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07153_ (.A1(\dp.rf.rf[3][2] ),
    .A2(_01179_),
    .Z(_02824_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _07154_ (.A1(_01163_),
    .A2(_01165_),
    .A3(_02823_),
    .A4(_02824_),
    .Z(_02825_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07155_ (.I0(\dp.rf.rf[1][2] ),
    .I1(\dp.rf.rf[5][2] ),
    .S(_01248_),
    .Z(_02826_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07156_ (.A1(_01328_),
    .A2(_02826_),
    .ZN(_02827_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07157_ (.A1(\dp.rf.rf[4][2] ),
    .A2(_01340_),
    .A3(_01162_),
    .B(_01218_),
    .ZN(_02828_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07158_ (.A1(_02827_),
    .A2(_02828_),
    .B(_01228_),
    .C(_01324_),
    .ZN(_02829_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07159_ (.I(\dp.rf.rf[0][2] ),
    .ZN(_02830_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07160_ (.A1(_02830_),
    .A2(_01736_),
    .ZN(_02831_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07161_ (.A1(_02820_),
    .A2(_02825_),
    .B1(_02829_),
    .B2(_02831_),
    .ZN(_02832_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07162_ (.I0(\dp.rf.rf[10][2] ),
    .I1(\dp.rf.rf[11][2] ),
    .I2(\dp.rf.rf[14][2] ),
    .I3(\dp.rf.rf[15][2] ),
    .S0(_01508_),
    .S1(_01145_),
    .Z(_02833_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07163_ (.I0(\dp.rf.rf[9][2] ),
    .I1(\dp.rf.rf[13][2] ),
    .S(_01122_),
    .Z(_02834_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _07164_ (.A1(_01225_),
    .A2(_01133_),
    .A3(_02834_),
    .Z(_02835_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07165_ (.A1(_01128_),
    .A2(net7),
    .ZN(_02836_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07166_ (.I0(\dp.rf.rf[8][2] ),
    .I1(\dp.rf.rf[12][2] ),
    .S(_01137_),
    .Z(_02837_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07167_ (.A1(_02836_),
    .A2(_02837_),
    .Z(_02838_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07168_ (.A1(_01175_),
    .A2(_02835_),
    .A3(_02838_),
    .Z(_02839_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07169_ (.A1(_01362_),
    .A2(_02833_),
    .B(_02839_),
    .ZN(_02840_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07170_ (.I0(\dp.rf.rf[22][2] ),
    .I1(\dp.rf.rf[23][2] ),
    .S(_01427_),
    .Z(_02841_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07171_ (.I(_02841_),
    .ZN(_02842_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07172_ (.A1(_01458_),
    .A2(_02842_),
    .B(_01150_),
    .ZN(_02843_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _07173_ (.A1(\dp.rf.rf[18][2] ),
    .A2(net10),
    .A3(net1),
    .A4(_01033_),
    .ZN(_02844_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07174_ (.I(\dp.rf.rf[18][2] ),
    .ZN(_02845_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _07175_ (.A1(_01028_),
    .A2(_01153_),
    .A3(_02844_),
    .B1(_01179_),
    .B2(_02845_),
    .ZN(_02846_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07176_ (.A1(\dp.rf.rf[19][2] ),
    .A2(_01135_),
    .Z(_02847_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _07177_ (.A1(_01163_),
    .A2(_01165_),
    .A3(_02846_),
    .A4(_02847_),
    .Z(_02848_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07178_ (.I0(\dp.rf.rf[17][2] ),
    .I1(\dp.rf.rf[21][2] ),
    .S(_01129_),
    .Z(_02849_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07179_ (.A1(_01190_),
    .A2(_02849_),
    .ZN(_02850_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07180_ (.A1(\dp.rf.rf[20][2] ),
    .A2(_01160_),
    .A3(_01162_),
    .B(_01171_),
    .ZN(_02851_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07181_ (.A1(_02850_),
    .A2(_02851_),
    .B(_01228_),
    .C(net257),
    .ZN(_02852_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07182_ (.I(\dp.rf.rf[16][2] ),
    .ZN(_02853_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07183_ (.A1(_02853_),
    .A2(_01736_),
    .ZN(_02854_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07184_ (.A1(_02843_),
    .A2(_02848_),
    .B1(_02852_),
    .B2(_02854_),
    .ZN(_02855_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07185_ (.I0(\dp.rf.rf[26][2] ),
    .I1(\dp.rf.rf[27][2] ),
    .I2(\dp.rf.rf[30][2] ),
    .I3(\dp.rf.rf[31][2] ),
    .S0(_01121_),
    .S1(_01124_),
    .Z(_02856_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07186_ (.I0(\dp.rf.rf[25][2] ),
    .I1(\dp.rf.rf[29][2] ),
    .S(_01122_),
    .Z(_02857_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _07187_ (.A1(_01238_),
    .A2(_01133_),
    .A3(_02857_),
    .Z(_02858_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07188_ (.I0(\dp.rf.rf[24][2] ),
    .I1(\dp.rf.rf[28][2] ),
    .S(_01122_),
    .Z(_02859_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07189_ (.A1(_02836_),
    .A2(_02859_),
    .Z(_02860_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07190_ (.A1(_01175_),
    .A2(_02858_),
    .A3(_02860_),
    .Z(_02861_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07191_ (.A1(_01416_),
    .A2(_02856_),
    .B(_02861_),
    .ZN(_02862_));
 gf180mcu_fd_sc_mcu9t5v0__oai33_4 _07192_ (.A1(net188),
    .A2(_02832_),
    .A3(_02840_),
    .B1(_02862_),
    .B2(_02855_),
    .B3(_01358_),
    .ZN(_05064_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07193_ (.I(net266),
    .ZN(_05068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07194_ (.A1(_01082_),
    .A2(_01104_),
    .ZN(_02863_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _07195_ (.A1(_01101_),
    .A2(_01097_),
    .A3(_02030_),
    .B1(_02791_),
    .B2(_01107_),
    .ZN(_02864_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07196_ (.A1(_02730_),
    .A2(_02731_),
    .B(_01324_),
    .C(_01766_),
    .ZN(_02865_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _07197_ (.A1(_01292_),
    .A2(_02864_),
    .B(_02865_),
    .C(_01109_),
    .ZN(_02866_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _07198_ (.A1(_02863_),
    .A2(_02866_),
    .ZN(_04821_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07199_ (.I0(\dp.rf.rf[26][1] ),
    .I1(\dp.rf.rf[27][1] ),
    .S(_01260_),
    .Z(_02867_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07200_ (.A1(_01823_),
    .A2(_02867_),
    .Z(_02868_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07201_ (.I0(\dp.rf.rf[18][1] ),
    .I1(\dp.rf.rf[19][1] ),
    .S(_01059_),
    .Z(_02869_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07202_ (.A1(_01103_),
    .A2(_01671_),
    .A3(_02869_),
    .Z(_02870_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07203_ (.I0(\dp.rf.rf[16][1] ),
    .I1(\dp.rf.rf[17][1] ),
    .S(_01059_),
    .Z(_02871_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07204_ (.A1(_02232_),
    .A2(_01671_),
    .A3(_02871_),
    .Z(_02872_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07205_ (.I0(\dp.rf.rf[24][1] ),
    .I1(\dp.rf.rf[25][1] ),
    .S(_01059_),
    .Z(_02873_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07206_ (.A1(_02232_),
    .A2(_01271_),
    .A3(_02873_),
    .Z(_02874_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _07207_ (.A1(_02868_),
    .A2(_02870_),
    .A3(_02872_),
    .A4(_02874_),
    .ZN(_02875_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _07208_ (.A1(_01057_),
    .A2(_01103_),
    .A3(_01060_),
    .Z(_02876_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07209_ (.I0(\dp.rf.rf[1][1] ),
    .I1(\dp.rf.rf[5][1] ),
    .I2(\dp.rf.rf[9][1] ),
    .I3(\dp.rf.rf[13][1] ),
    .S0(_01047_),
    .S1(_01671_),
    .Z(_02877_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07210_ (.I0(\dp.rf.rf[0][1] ),
    .I1(\dp.rf.rf[4][1] ),
    .I2(\dp.rf.rf[8][1] ),
    .I3(\dp.rf.rf[12][1] ),
    .S0(net11),
    .S1(_01671_),
    .Z(_02878_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07211_ (.I0(_02877_),
    .I1(_02878_),
    .S(_01099_),
    .Z(_02879_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07212_ (.I0(\dp.rf.rf[6][1] ),
    .I1(\dp.rf.rf[7][1] ),
    .I2(\dp.rf.rf[14][1] ),
    .I3(\dp.rf.rf[15][1] ),
    .S0(_01038_),
    .S1(net12),
    .Z(_02880_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07213_ (.I0(\dp.rf.rf[2][1] ),
    .I1(\dp.rf.rf[3][1] ),
    .I2(\dp.rf.rf[10][1] ),
    .I3(\dp.rf.rf[11][1] ),
    .S0(net264),
    .S1(net12),
    .Z(_02881_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07214_ (.I0(_02880_),
    .I1(_02881_),
    .S(_01667_),
    .Z(_02882_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07215_ (.A1(_01057_),
    .A2(_01485_),
    .Z(_02883_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _07216_ (.A1(_02876_),
    .A2(_02879_),
    .B1(_02882_),
    .B2(_02883_),
    .ZN(_02884_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07217_ (.I0(\dp.rf.rf[28][1] ),
    .I1(\dp.rf.rf[29][1] ),
    .I2(\dp.rf.rf[30][1] ),
    .I3(\dp.rf.rf[31][1] ),
    .S0(_01038_),
    .S1(_01102_),
    .Z(_02885_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07218_ (.I0(\dp.rf.rf[20][1] ),
    .I1(\dp.rf.rf[21][1] ),
    .I2(\dp.rf.rf[22][1] ),
    .I3(\dp.rf.rf[23][1] ),
    .S0(_01038_),
    .S1(_01102_),
    .Z(_02886_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07219_ (.I0(_02885_),
    .I1(_02886_),
    .S(_01271_),
    .Z(_02887_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07220_ (.A1(_01778_),
    .A2(_02887_),
    .ZN(_02888_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _07221_ (.A1(_02690_),
    .A2(_02875_),
    .B(_02884_),
    .C(_02888_),
    .ZN(net139));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _07222_ (.A1(_01093_),
    .A2(_02863_),
    .A3(_02866_),
    .Z(_02889_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _07223_ (.A1(_01093_),
    .A2(net139),
    .ZN(_02890_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _07224_ (.A1(_02890_),
    .A2(_02889_),
    .ZN(_02891_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _07225_ (.I(_02891_),
    .Z(_02892_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer8 (.I(_01073_),
    .Z(net167));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _07227_ (.A1(_01085_),
    .A2(_02892_),
    .ZN(_04816_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07228_ (.I(_04816_),
    .ZN(_05075_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07229_ (.I0(\dp.rf.rf[14][1] ),
    .I1(\dp.rf.rf[15][1] ),
    .S(_01147_),
    .Z(_02894_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07230_ (.A1(_01230_),
    .A2(_02894_),
    .ZN(_02895_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07231_ (.A1(_01151_),
    .A2(_02895_),
    .ZN(_02896_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _07232_ (.A1(\dp.rf.rf[10][1] ),
    .A2(_01154_),
    .A3(_01155_),
    .A4(_01034_),
    .ZN(_02897_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07233_ (.I(\dp.rf.rf[10][1] ),
    .ZN(_02898_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _07234_ (.A1(_01028_),
    .A2(_01153_),
    .A3(_02897_),
    .B1(_01136_),
    .B2(_02898_),
    .ZN(_02899_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07235_ (.A1(\dp.rf.rf[11][1] ),
    .A2(_01160_),
    .Z(_02900_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _07236_ (.A1(_01164_),
    .A2(_01166_),
    .A3(_02899_),
    .A4(_02900_),
    .Z(_02901_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07237_ (.I0(\dp.rf.rf[8][1] ),
    .I1(\dp.rf.rf[9][1] ),
    .I2(\dp.rf.rf[12][1] ),
    .I3(\dp.rf.rf[13][1] ),
    .S0(_01157_),
    .S1(_01139_),
    .Z(_02902_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _07238_ (.A1(_02896_),
    .A2(_02901_),
    .B1(_02902_),
    .B2(_01173_),
    .C(_01237_),
    .ZN(_02903_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07239_ (.I0(\dp.rf.rf[2][1] ),
    .I1(\dp.rf.rf[3][1] ),
    .I2(\dp.rf.rf[6][1] ),
    .I3(\dp.rf.rf[7][1] ),
    .S0(_01582_),
    .S1(_01124_),
    .Z(_02904_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07240_ (.A1(_01119_),
    .A2(_02904_),
    .Z(_02905_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07241_ (.I(\dp.rf.rf[4][1] ),
    .ZN(_02906_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07242_ (.I0(\dp.rf.rf[1][1] ),
    .I1(\dp.rf.rf[5][1] ),
    .S(_01144_),
    .Z(_02907_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07243_ (.A1(_01371_),
    .A2(_02907_),
    .ZN(_02908_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _07244_ (.A1(_02906_),
    .A2(_01327_),
    .B(_02908_),
    .C(_01119_),
    .ZN(_02909_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07245_ (.A1(_01541_),
    .A2(_02905_),
    .A3(_02909_),
    .B(_01376_),
    .ZN(_02910_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07246_ (.A1(_02903_),
    .A2(_02910_),
    .Z(_02911_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07247_ (.I0(\dp.rf.rf[24][1] ),
    .I1(\dp.rf.rf[25][1] ),
    .I2(\dp.rf.rf[28][1] ),
    .I3(\dp.rf.rf[29][1] ),
    .S0(_01363_),
    .S1(_01364_),
    .Z(_02912_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07248_ (.I0(\dp.rf.rf[26][1] ),
    .I1(\dp.rf.rf[27][1] ),
    .S(_01520_),
    .Z(_02913_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07249_ (.I(_02913_),
    .ZN(_02914_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07250_ (.I0(\dp.rf.rf[30][1] ),
    .I1(\dp.rf.rf[31][1] ),
    .S(_01363_),
    .Z(_02915_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07251_ (.I(_02915_),
    .ZN(_02916_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07252_ (.A1(_01224_),
    .A2(_02914_),
    .B1(_02916_),
    .B2(_01146_),
    .ZN(_02917_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07253_ (.I0(_02912_),
    .I1(_02917_),
    .S(_01530_),
    .Z(_02918_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07254_ (.I0(\dp.rf.rf[22][1] ),
    .I1(\dp.rf.rf[23][1] ),
    .S(_01363_),
    .Z(_02919_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07255_ (.A1(_01505_),
    .A2(_02919_),
    .ZN(_02920_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07256_ (.A1(\dp.rf.rf[19][1] ),
    .A2(_01520_),
    .Z(_02921_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _07257_ (.A1(_01210_),
    .A2(net257),
    .B1(_01626_),
    .B2(\dp.rf.rf[18][1] ),
    .C(_02921_),
    .ZN(_02922_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _07258_ (.A1(_01697_),
    .A2(_02920_),
    .A3(_02922_),
    .ZN(_02923_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07259_ (.I(\dp.rf.rf[16][1] ),
    .ZN(_02924_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07260_ (.I0(\dp.rf.rf[17][1] ),
    .I1(\dp.rf.rf[21][1] ),
    .S(_01123_),
    .Z(_02925_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _07261_ (.A1(\dp.rf.rf[20][1] ),
    .A2(_01497_),
    .B1(_02925_),
    .B2(_01693_),
    .C(_01576_),
    .ZN(_02926_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _07262_ (.A1(_02924_),
    .A2(_01737_),
    .B1(_02926_),
    .B2(_01361_),
    .C(_01455_),
    .ZN(_02927_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _07263_ (.A1(_01580_),
    .A2(_02918_),
    .B1(_02923_),
    .B2(_02927_),
    .ZN(_02928_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _07264_ (.A1(_02928_),
    .A2(_02911_),
    .ZN(_04815_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07265_ (.I(_04815_),
    .ZN(_05074_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07266_ (.I(_04835_),
    .ZN(_02929_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _07267_ (.A1(_01438_),
    .A2(_01036_),
    .ZN(_02930_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _07268_ (.A1(net6),
    .A2(net4),
    .ZN(_02931_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07269_ (.A1(_02930_),
    .A2(_02931_),
    .ZN(_02932_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07270_ (.A1(net22),
    .A2(_01066_),
    .B(_01065_),
    .ZN(_02933_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07271_ (.A1(_01438_),
    .A2(_01068_),
    .B(_01067_),
    .ZN(_02934_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07272_ (.A1(_02933_),
    .A2(_02934_),
    .B(net6),
    .ZN(_02935_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _07273_ (.A1(_01068_),
    .A2(_02932_),
    .B(_02935_),
    .C(_01084_),
    .ZN(_02936_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07274_ (.I(_02936_),
    .Z(_02937_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07275_ (.A1(_01029_),
    .A2(_01031_),
    .B(_01438_),
    .ZN(_02938_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07276_ (.A1(net24),
    .A2(_01066_),
    .B(_02938_),
    .ZN(_02939_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _07277_ (.A1(_01079_),
    .A2(_02939_),
    .B(_01245_),
    .ZN(_02940_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _07278_ (.A1(net5),
    .A2(_02931_),
    .A3(_02940_),
    .ZN(_02941_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07279_ (.I(_02941_),
    .Z(_02942_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _07280_ (.A1(_02170_),
    .A2(_01067_),
    .A3(_01068_),
    .A4(_02933_),
    .Z(_02943_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _07281_ (.A1(_01258_),
    .A2(_01287_),
    .Z(_02944_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07282_ (.A1(_02943_),
    .A2(_02944_),
    .Z(_02945_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _07283_ (.A1(net248),
    .A2(_02945_),
    .ZN(_02946_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _07284_ (.A1(_02929_),
    .A2(_02937_),
    .A3(_02942_),
    .A4(_02946_),
    .Z(_02947_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _07285_ (.A1(_04834_),
    .A2(_04842_),
    .A3(_02937_),
    .A4(_02942_),
    .ZN(_02948_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07286_ (.A1(_02946_),
    .A2(_02948_),
    .ZN(_02949_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _07287_ (.I(_04995_),
    .ZN(_02950_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _07288_ (.I(_05011_),
    .ZN(_02951_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _07289_ (.A1(_05026_),
    .A2(_05019_),
    .B(_05018_),
    .ZN(_02952_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07290_ (.I(_05010_),
    .ZN(_02953_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _07291_ (.A1(_02952_),
    .A2(_02951_),
    .B(_02953_),
    .ZN(_02954_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _07292_ (.A1(_05003_),
    .A2(_02954_),
    .B(_05002_),
    .ZN(_02955_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07293_ (.A1(_04986_),
    .A2(_04994_),
    .ZN(_02956_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _07294_ (.A1(_02955_),
    .A2(_02950_),
    .B(_02956_),
    .ZN(_02957_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07295_ (.I(_04979_),
    .ZN(_02958_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07296_ (.A1(_04986_),
    .A2(_04987_),
    .ZN(_02959_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07297_ (.A1(_02958_),
    .A2(_02959_),
    .ZN(_02960_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07298_ (.I(_05059_),
    .ZN(_02961_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _07299_ (.A1(_05067_),
    .A2(_04817_),
    .B(_05066_),
    .ZN(_02962_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07300_ (.I(_05058_),
    .ZN(_02963_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _07301_ (.A1(_02961_),
    .A2(_02962_),
    .B(_02963_),
    .ZN(_02964_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _07302_ (.A1(_05051_),
    .A2(_02964_),
    .B(_05050_),
    .ZN(_02965_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07303_ (.A1(_05035_),
    .A2(_05043_),
    .ZN(_02966_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07304_ (.A1(_05035_),
    .A2(_05042_),
    .B(_05034_),
    .ZN(_02967_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _07305_ (.A1(_02965_),
    .A2(_02966_),
    .B(_02967_),
    .ZN(_02968_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _07306_ (.A1(_05003_),
    .A2(_05011_),
    .A3(_05019_),
    .A4(_05027_),
    .Z(_02969_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _07307_ (.A1(_04979_),
    .A2(_04987_),
    .A3(_04995_),
    .A4(_02969_),
    .Z(_02970_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _07308_ (.A1(_02957_),
    .A2(_02960_),
    .B1(_02968_),
    .B2(_02970_),
    .C(_04978_),
    .ZN(_02971_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07309_ (.I(_04971_),
    .ZN(_02972_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07310_ (.A1(_04955_),
    .A2(_04963_),
    .ZN(_02973_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07311_ (.A1(_02972_),
    .A2(_02973_),
    .Z(_02974_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _07312_ (.A1(_04970_),
    .A2(_04955_),
    .A3(_04963_),
    .Z(_02975_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07313_ (.A1(_04955_),
    .A2(_04962_),
    .B(_02975_),
    .ZN(_02976_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _07314_ (.A1(net268),
    .A2(_02974_),
    .B(_02976_),
    .ZN(_02977_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _07315_ (.A1(_04939_),
    .A2(_04923_),
    .A3(_04931_),
    .A4(_04947_),
    .Z(_02978_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _07316_ (.I(_04939_),
    .ZN(_02979_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07317_ (.I(_04946_),
    .ZN(_02980_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07318_ (.A1(_04923_),
    .A2(_04931_),
    .ZN(_02981_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07319_ (.I(_04954_),
    .ZN(_02982_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07320_ (.A1(_02982_),
    .A2(_02979_),
    .A3(_02981_),
    .Z(_02983_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _07321_ (.I(_04947_),
    .ZN(_02984_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _07322_ (.A1(_02979_),
    .A2(_02980_),
    .A3(_02981_),
    .B1(_02983_),
    .B2(_02984_),
    .ZN(_02985_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07323_ (.I(_04923_),
    .ZN(_02986_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07324_ (.A1(_04938_),
    .A2(_04931_),
    .B(_04930_),
    .ZN(_02987_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07325_ (.I(_04922_),
    .ZN(_02988_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07326_ (.A1(_02986_),
    .A2(_02987_),
    .B(_02988_),
    .ZN(_02989_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07327_ (.A1(_04906_),
    .A2(_04914_),
    .A3(_02989_),
    .Z(_02990_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _07328_ (.A1(_02977_),
    .A2(_02978_),
    .B(_02985_),
    .C(_02990_),
    .ZN(_02991_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07329_ (.A1(_04906_),
    .A2(_04915_),
    .A3(_04914_),
    .Z(_02992_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07330_ (.A1(_04906_),
    .A2(_04907_),
    .B(_02992_),
    .ZN(_02993_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07331_ (.A1(_04891_),
    .A2(_04883_),
    .Z(_02994_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _07332_ (.A1(_04875_),
    .A2(_04899_),
    .A3(_02994_),
    .Z(_02995_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07333_ (.A1(_04867_),
    .A2(_02995_),
    .ZN(_02996_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07334_ (.I(_04874_),
    .ZN(_02997_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07335_ (.A1(_04890_),
    .A2(_04883_),
    .Z(_02998_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07336_ (.A1(_04898_),
    .A2(_02994_),
    .Z(_02999_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07337_ (.A1(_04882_),
    .A2(_02998_),
    .A3(_02999_),
    .B(_04875_),
    .ZN(_03000_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07338_ (.A1(_02997_),
    .A2(_03000_),
    .ZN(_03001_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07339_ (.A1(_04867_),
    .A2(_03001_),
    .B(_04866_),
    .ZN(_03002_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _07340_ (.A1(_02996_),
    .A2(_02993_),
    .A3(_02991_),
    .B(_03002_),
    .ZN(_03003_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _07341_ (.A1(_04851_),
    .A2(_04859_),
    .A3(_03003_),
    .A4(_04843_),
    .Z(_03004_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _07342_ (.A1(_04851_),
    .A2(_04843_),
    .A3(_04858_),
    .Z(_03005_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _07343_ (.A1(_04843_),
    .A2(_04850_),
    .B(_03004_),
    .C(_03005_),
    .ZN(_03006_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07344_ (.I0(_02947_),
    .I1(_02949_),
    .S(_03006_),
    .Z(_03007_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07345_ (.A1(net4),
    .A2(_01068_),
    .Z(_03008_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _07346_ (.I(_02170_),
    .ZN(_03009_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07347_ (.A1(_03009_),
    .A2(net19),
    .ZN(_03010_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _07348_ (.A1(_02409_),
    .A2(_02930_),
    .A3(_03008_),
    .A4(_03010_),
    .ZN(_03011_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _07349_ (.I(_03011_),
    .Z(_03012_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _07350_ (.I(_02937_),
    .Z(_03013_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _07351_ (.I(_02941_),
    .Z(_03014_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07352_ (.A1(_01067_),
    .A2(_01068_),
    .Z(_03015_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _07353_ (.A1(_02170_),
    .A2(_03015_),
    .A3(_02940_),
    .ZN(_03016_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07354_ (.A1(_02941_),
    .A2(_03016_),
    .Z(_03017_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07355_ (.I(_03017_),
    .Z(_03018_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07356_ (.A1(_04826_),
    .A2(_03018_),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07357_ (.A1(_04830_),
    .A2(_03014_),
    .B(_03019_),
    .ZN(_03020_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07358_ (.A1(_03013_),
    .A2(_03020_),
    .ZN(_03021_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _07359_ (.A1(net5),
    .A2(_02931_),
    .A3(_02940_),
    .Z(_03022_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07360_ (.A1(_02937_),
    .A2(_03022_),
    .Z(_03023_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07361_ (.A1(net247),
    .A2(_03023_),
    .Z(_03024_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _07362_ (.A1(_02936_),
    .A2(_03022_),
    .ZN(_03025_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07363_ (.I(_03025_),
    .Z(_03026_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _07364_ (.A1(_02170_),
    .A2(_03015_),
    .A3(_02940_),
    .Z(_03027_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07365_ (.I(_03027_),
    .Z(_03028_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07366_ (.A1(net247),
    .A2(_03026_),
    .B(_03028_),
    .ZN(_03029_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07367_ (.I0(_03024_),
    .I1(_03029_),
    .S(_04827_),
    .Z(_03030_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07368_ (.I(_02937_),
    .Z(_03031_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07369_ (.A1(_04835_),
    .A2(_04842_),
    .B(_04834_),
    .ZN(_03032_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07370_ (.A1(_04835_),
    .A2(_04834_),
    .Z(_03033_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07371_ (.I0(_03032_),
    .I1(_03033_),
    .S(_02946_),
    .Z(_03034_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07372_ (.A1(_03031_),
    .A2(_02942_),
    .A3(_03034_),
    .Z(_03035_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _07373_ (.A1(_03012_),
    .A2(_03021_),
    .A3(_03030_),
    .A4(_03035_),
    .Z(_03036_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07374_ (.A1(_01259_),
    .A2(net154),
    .Z(_03037_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _07375_ (.A1(_01605_),
    .A2(_05094_),
    .B(_03037_),
    .ZN(_03038_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07376_ (.I(_03038_),
    .Z(_03039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07377_ (.I0(_01062_),
    .I1(_01110_),
    .S(_01093_),
    .Z(_03040_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _07378_ (.I(_03040_),
    .Z(_03041_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07379_ (.I(_03041_),
    .Z(_03042_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _07380_ (.A1(_02889_),
    .A2(_02890_),
    .Z(_03043_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07381_ (.I(_03043_),
    .Z(_03044_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _07382_ (.I(_03044_),
    .Z(_03045_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07383_ (.I0(_04896_),
    .I1(_04904_),
    .I2(_04912_),
    .I3(_04920_),
    .S0(_03042_),
    .S1(_03045_),
    .Z(_03046_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07384_ (.I0(_04936_),
    .I1(_04952_),
    .S(_03044_),
    .Z(_03047_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07385_ (.I0(_04928_),
    .I1(_04944_),
    .S(_03044_),
    .Z(_03048_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07386_ (.I0(_03047_),
    .I1(_03048_),
    .S(_01115_),
    .Z(_03049_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _07387_ (.I(_01388_),
    .Z(_04840_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07388_ (.I(_03044_),
    .Z(_03050_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07389_ (.I0(_01258_),
    .I1(_04840_),
    .I2(_04848_),
    .I3(_04856_),
    .S0(_03042_),
    .S1(_03050_),
    .Z(_03051_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07390_ (.I0(_04864_),
    .I1(_04872_),
    .I2(_04880_),
    .I3(_04888_),
    .S0(_03042_),
    .S1(_03050_),
    .Z(_03052_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _07391_ (.A1(_02812_),
    .A2(_02813_),
    .Z(_03053_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _07392_ (.I(_03053_),
    .Z(_03054_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07393_ (.I0(_03046_),
    .I1(_03049_),
    .I2(_03051_),
    .I3(_03052_),
    .S0(_03054_),
    .S1(_02750_),
    .Z(_03055_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07394_ (.I0(_05028_),
    .I1(_05036_),
    .S(net221),
    .Z(_03056_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07395_ (.I(_03041_),
    .Z(_03057_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07396_ (.I0(_05044_),
    .I1(_05052_),
    .S(_03057_),
    .Z(_03058_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07397_ (.I0(_05060_),
    .I1(_05068_),
    .S(_03057_),
    .Z(_03059_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07398_ (.I0(_04824_),
    .I1(net242),
    .S(_01116_),
    .Z(_03060_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07399_ (.I(_03060_),
    .ZN(_03061_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _07400_ (.I(_03043_),
    .Z(_03062_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _07401_ (.I(_03062_),
    .Z(_03063_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07402_ (.I(_03053_),
    .Z(_03064_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07403_ (.I(_03064_),
    .Z(_03065_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07404_ (.I0(_03056_),
    .I1(_03058_),
    .I2(_03059_),
    .I3(_03061_),
    .S0(_03063_),
    .S1(_03065_),
    .Z(_03066_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07405_ (.I(_02750_),
    .Z(_03067_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07406_ (.I0(net243),
    .I1(_04968_),
    .I2(_04976_),
    .I3(_04984_),
    .S0(_03042_),
    .S1(_03050_),
    .Z(_03068_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07407_ (.I0(net238),
    .I1(_05000_),
    .I2(net181),
    .I3(net174),
    .S0(_03042_),
    .S1(_03050_),
    .Z(_03069_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _07408_ (.I(_03053_),
    .Z(_03070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07409_ (.I0(_03068_),
    .I1(_03069_),
    .S(_03070_),
    .Z(_03071_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07410_ (.A1(_03067_),
    .A2(_03071_),
    .ZN(_03072_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07411_ (.A1(net222),
    .A2(_03066_),
    .B(_03072_),
    .C(_03039_),
    .ZN(_03073_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _07412_ (.A1(_02170_),
    .A2(net4),
    .A3(_01068_),
    .A4(_02930_),
    .Z(_03074_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07413_ (.I(_03074_),
    .Z(_03075_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _07414_ (.I(_03075_),
    .Z(_03076_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _07415_ (.A1(_03039_),
    .A2(_03055_),
    .B(_03073_),
    .C(_03076_),
    .ZN(_03077_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07416_ (.I(_03041_),
    .Z(_03078_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07417_ (.I(_03078_),
    .Z(_03079_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _07418_ (.A1(_03079_),
    .A2(_04824_),
    .A3(_03063_),
    .Z(_03080_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _07419_ (.A1(_02170_),
    .A2(net4),
    .A3(_01068_),
    .A4(_02930_),
    .ZN(_03081_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07420_ (.A1(_03038_),
    .A2(_03081_),
    .Z(_03082_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07421_ (.A1(_02747_),
    .A2(_02748_),
    .Z(_03083_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07422_ (.A1(_03083_),
    .A2(_03054_),
    .Z(_03084_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07423_ (.A1(_03082_),
    .A2(_03084_),
    .Z(_03085_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07424_ (.A1(_03080_),
    .A2(_03085_),
    .B(_03012_),
    .ZN(_03086_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _07425_ (.A1(_03007_),
    .A2(_03036_),
    .B1(_03077_),
    .B2(_03086_),
    .ZN(net61));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07426_ (.A1(_01029_),
    .A2(_02930_),
    .Z(_03087_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _07427_ (.I(_03087_),
    .ZN(_03088_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _07428_ (.I(_03088_),
    .Z(_03089_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _07429_ (.I(_03089_),
    .Z(net93));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07430_ (.A1(net250),
    .A2(_03075_),
    .ZN(_03090_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07431_ (.I0(_04896_),
    .I1(_04912_),
    .S(_03062_),
    .Z(_03091_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07432_ (.I0(_04888_),
    .I1(_04904_),
    .S(_03062_),
    .Z(_03092_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07433_ (.I0(_04920_),
    .I1(_04936_),
    .S(_03062_),
    .Z(_03093_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07434_ (.I0(_03091_),
    .I1(_03048_),
    .I2(_03092_),
    .I3(_03093_),
    .S0(_03053_),
    .S1(_01116_),
    .Z(_03094_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07435_ (.I(_03094_),
    .ZN(_03095_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07436_ (.I(_02814_),
    .Z(_03096_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07437_ (.I(_03044_),
    .Z(_03097_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07438_ (.I0(_04856_),
    .I1(_04864_),
    .I2(_04872_),
    .I3(_04880_),
    .S0(_03042_),
    .S1(_03097_),
    .Z(_03098_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07439_ (.A1(_03078_),
    .A2(_04848_),
    .ZN(_03099_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07440_ (.A1(_01359_),
    .A2(_01387_),
    .B(_01115_),
    .ZN(_03100_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07441_ (.I(net164),
    .Z(_03101_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07442_ (.I(_03101_),
    .Z(_03102_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07443_ (.A1(_03099_),
    .A2(_03100_),
    .B(_03102_),
    .ZN(_03103_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07444_ (.A1(_01093_),
    .A2(net139),
    .Z(_03104_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _07445_ (.A1(_01259_),
    .A2(_04821_),
    .B(_03104_),
    .C(_01258_),
    .ZN(_03105_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07446_ (.A1(net163),
    .A2(_03105_),
    .ZN(_03106_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _07447_ (.A1(_03096_),
    .A2(_03098_),
    .B1(_03103_),
    .B2(_03106_),
    .ZN(_03107_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07448_ (.A1(_02889_),
    .A2(_02890_),
    .B(_01469_),
    .ZN(_03108_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07449_ (.A1(_03105_),
    .A2(_03108_),
    .Z(_03109_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07450_ (.I0(_04868_),
    .I1(_04884_),
    .S(_03044_),
    .Z(_03110_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07451_ (.A1(_04840_),
    .A2(_03097_),
    .ZN(_03111_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07452_ (.I0(_04860_),
    .I1(_04876_),
    .S(_03043_),
    .Z(_03112_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07453_ (.I0(_03109_),
    .I1(_03110_),
    .I2(_03111_),
    .I3(_03112_),
    .S0(_03053_),
    .S1(_01115_),
    .Z(_03113_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _07454_ (.I(net19),
    .ZN(_03114_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07455_ (.I0(_03107_),
    .I1(_03113_),
    .S(_03114_),
    .Z(_03115_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _07456_ (.I(_02749_),
    .Z(_03116_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07457_ (.I0(_03095_),
    .I1(_03115_),
    .S(_03116_),
    .Z(_03117_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _07458_ (.A1(_03038_),
    .A2(_03075_),
    .ZN(_03118_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07459_ (.I0(_04964_),
    .I1(_04980_),
    .S(_03062_),
    .Z(_03119_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07460_ (.I0(_04956_),
    .I1(_04972_),
    .S(_03044_),
    .Z(_03120_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07461_ (.I0(_03119_),
    .I1(_03120_),
    .S(_01115_),
    .Z(_03121_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07462_ (.I0(_04988_),
    .I1(_04996_),
    .I2(_05004_),
    .I3(_05012_),
    .S0(net221),
    .S1(_03097_),
    .Z(_03122_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07463_ (.I0(_03121_),
    .I1(_03122_),
    .S(_03054_),
    .Z(_03123_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07464_ (.I0(_05020_),
    .I1(_05028_),
    .I2(_05036_),
    .I3(_05044_),
    .S0(_03042_),
    .S1(_03097_),
    .Z(_03124_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07465_ (.I0(_05052_),
    .I1(_05060_),
    .I2(_05068_),
    .I3(_05074_),
    .S0(_03057_),
    .S1(_03063_),
    .Z(_03125_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07466_ (.I0(_03124_),
    .I1(_03125_),
    .S(_03064_),
    .Z(_03126_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07467_ (.I(_03083_),
    .Z(_03127_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07468_ (.I0(_03123_),
    .I1(_03126_),
    .S(_03127_),
    .Z(_03128_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _07469_ (.A1(_03041_),
    .A2(_04824_),
    .Z(_03129_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _07470_ (.A1(_01115_),
    .A2(net242),
    .B(_03129_),
    .C(_03097_),
    .ZN(_03130_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07471_ (.I(_03130_),
    .ZN(_03131_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07472_ (.A1(_03085_),
    .A2(_03131_),
    .B(_03011_),
    .ZN(_03132_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _07473_ (.A1(_03090_),
    .A2(_03117_),
    .B1(_03118_),
    .B2(_03128_),
    .C(_03132_),
    .ZN(_03133_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07474_ (.A1(_03031_),
    .A2(_03022_),
    .ZN(_03134_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _07475_ (.A1(_02409_),
    .A2(_02930_),
    .A3(_03008_),
    .A4(_03010_),
    .Z(_03135_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07476_ (.I(_03135_),
    .Z(_03136_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07477_ (.A1(_05073_),
    .A2(_03028_),
    .B(_03136_),
    .ZN(_03137_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _07478_ (.I(_03017_),
    .Z(_03138_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07479_ (.I(_03138_),
    .Z(_03139_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07480_ (.I(_04818_),
    .ZN(_03140_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07481_ (.I0(_03140_),
    .I1(_05072_),
    .S(_02937_),
    .Z(_03141_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07482_ (.A1(_03139_),
    .A2(_03141_),
    .ZN(_03142_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07483_ (.A1(_05076_),
    .A2(_03134_),
    .B(_03137_),
    .C(_03142_),
    .ZN(_03143_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07484_ (.A1(_03133_),
    .A2(_03143_),
    .Z(net72));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _07485_ (.I(_03028_),
    .Z(_03144_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07486_ (.A1(_05067_),
    .A2(_03144_),
    .B(_03136_),
    .ZN(_03145_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _07487_ (.A1(_04817_),
    .A2(_05067_),
    .Z(_03146_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07488_ (.I0(_03146_),
    .I1(_05066_),
    .S(_02937_),
    .Z(_03147_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07489_ (.A1(_03139_),
    .A2(_03147_),
    .ZN(_03148_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07490_ (.A1(_05070_),
    .A2(_03134_),
    .B(_03145_),
    .C(_03148_),
    .ZN(_03149_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07491_ (.I(_03070_),
    .Z(_03150_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07492_ (.I0(_04852_),
    .I1(_04860_),
    .I2(_04868_),
    .I3(_04876_),
    .S0(_03078_),
    .S1(_03045_),
    .Z(_03151_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07493_ (.A1(_03150_),
    .A2(_03151_),
    .ZN(_03152_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07494_ (.A1(net178),
    .A2(_03152_),
    .Z(_03153_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07495_ (.A1(_03042_),
    .A2(_01258_),
    .ZN(_03154_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _07496_ (.A1(_01114_),
    .A2(_01359_),
    .A3(_01387_),
    .ZN(_03155_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07497_ (.A1(net271),
    .A2(_03154_),
    .A3(_03155_),
    .Z(_03156_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07498_ (.A1(net175),
    .A2(_03156_),
    .Z(_03157_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07499_ (.A1(_03114_),
    .A2(_03105_),
    .B(_03157_),
    .ZN(_03158_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _07500_ (.I(_03083_),
    .Z(_03159_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _07501_ (.I(_03159_),
    .Z(_03160_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07502_ (.I0(_04912_),
    .I1(_04928_),
    .S(_03062_),
    .Z(_03161_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07503_ (.I0(_04880_),
    .I1(_04896_),
    .S(_03097_),
    .Z(_03162_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07504_ (.I0(_03093_),
    .I1(_03092_),
    .I2(_03161_),
    .I3(_03162_),
    .S0(_03096_),
    .S1(_01116_),
    .Z(_03163_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07505_ (.A1(_03160_),
    .A2(_03163_),
    .Z(_03164_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07506_ (.A1(_03153_),
    .A2(_03158_),
    .B(_03164_),
    .ZN(_03165_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07507_ (.I0(_05012_),
    .I1(_05020_),
    .S(net221),
    .Z(_03166_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07508_ (.I0(_03166_),
    .I1(_03056_),
    .S(_03097_),
    .Z(_03167_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07509_ (.I0(_03058_),
    .I1(_03059_),
    .S(_03063_),
    .Z(_03168_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07510_ (.I0(_04944_),
    .I1(_04952_),
    .I2(net243),
    .I3(_04968_),
    .S0(net221),
    .S1(_03062_),
    .Z(_03169_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07511_ (.I(_03169_),
    .ZN(_03170_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07512_ (.I0(_04980_),
    .I1(_04996_),
    .S(_03043_),
    .Z(_03171_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07513_ (.I0(_04988_),
    .I1(_05004_),
    .S(_03043_),
    .Z(_03172_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07514_ (.I0(_03171_),
    .I1(_03172_),
    .S(_03042_),
    .Z(_03173_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07515_ (.I0(_03167_),
    .I1(_03168_),
    .I2(_03170_),
    .I3(_03173_),
    .S0(_03065_),
    .S1(net178),
    .Z(_03174_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07516_ (.I0(_04824_),
    .I1(net258),
    .S(_03044_),
    .Z(_03175_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07517_ (.A1(_03063_),
    .A2(net242),
    .Z(_03176_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07518_ (.I0(_03175_),
    .I1(_03176_),
    .S(_01116_),
    .Z(_03177_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07519_ (.I(_03011_),
    .Z(_03178_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07520_ (.A1(_03085_),
    .A2(_03177_),
    .B(_03178_),
    .ZN(_03179_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _07521_ (.A1(_03090_),
    .A2(_03165_),
    .B1(_03174_),
    .B2(_03118_),
    .C(_03179_),
    .ZN(_03180_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07522_ (.A1(_03149_),
    .A2(_03180_),
    .Z(net83));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07523_ (.A1(net246),
    .A2(_03041_),
    .ZN(_03181_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07524_ (.A1(_03181_),
    .A2(_03129_),
    .Z(_04814_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _07525_ (.I(_03178_),
    .Z(_03182_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _07526_ (.I(_03031_),
    .Z(_03183_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07527_ (.I(_02942_),
    .Z(_03184_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07528_ (.A1(_05058_),
    .A2(_03139_),
    .ZN(_03185_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07529_ (.A1(_05062_),
    .A2(_03184_),
    .B(_03185_),
    .ZN(_03186_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07530_ (.A1(_03183_),
    .A2(_03186_),
    .ZN(_03187_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07531_ (.A1(_03182_),
    .A2(_03187_),
    .ZN(_03188_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07532_ (.I(_03023_),
    .Z(_03189_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07533_ (.I(_05066_),
    .ZN(_03190_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07534_ (.A1(_05073_),
    .A2(_04814_),
    .Z(_03191_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07535_ (.A1(_05072_),
    .A2(_03191_),
    .B(_05067_),
    .ZN(_03192_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07536_ (.A1(_03190_),
    .A2(_03192_),
    .ZN(_03193_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07537_ (.I(_03016_),
    .Z(_03194_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07538_ (.A1(_03189_),
    .A2(_03193_),
    .B(_03194_),
    .ZN(_03195_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07539_ (.A1(_05059_),
    .A2(_03195_),
    .Z(_03196_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _07540_ (.I(_03026_),
    .Z(_03197_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _07541_ (.A1(_02961_),
    .A2(_03197_),
    .A3(_03193_),
    .Z(_03198_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07542_ (.I(_03079_),
    .Z(_03199_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07543_ (.I0(_05032_),
    .I1(_05040_),
    .I2(_05048_),
    .I3(_05056_),
    .S0(_03199_),
    .S1(_03063_),
    .Z(_03200_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07544_ (.I0(_05004_),
    .I1(_05012_),
    .I2(_05020_),
    .I3(_05028_),
    .S0(_03078_),
    .S1(_03045_),
    .Z(_03201_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07545_ (.A1(_03065_),
    .A2(_03201_),
    .ZN(_03202_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07546_ (.A1(_03065_),
    .A2(_03200_),
    .B(_03202_),
    .ZN(_03203_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07547_ (.I0(_04972_),
    .I1(_04988_),
    .S(_03045_),
    .Z(_03204_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07548_ (.I0(_04940_),
    .I1(_04956_),
    .S(_03045_),
    .Z(_03205_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07549_ (.I0(_04948_),
    .I1(_04964_),
    .S(_03045_),
    .Z(_03206_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07550_ (.I0(_03204_),
    .I1(_03205_),
    .I2(_03171_),
    .I3(_03206_),
    .S0(net179),
    .S1(_03199_),
    .Z(_03207_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07551_ (.I0(_03203_),
    .I1(_03207_),
    .S(_03067_),
    .Z(_03208_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07552_ (.I0(_04908_),
    .I1(_04924_),
    .S(_03050_),
    .Z(_03209_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07553_ (.I0(_04876_),
    .I1(_04892_),
    .S(_03050_),
    .Z(_03210_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07554_ (.I0(_04916_),
    .I1(_04932_),
    .S(_03050_),
    .Z(_03211_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07555_ (.I0(_04884_),
    .I1(_04900_),
    .S(_03097_),
    .Z(_03212_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07556_ (.I(_03078_),
    .Z(_03213_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07557_ (.I0(_03209_),
    .I1(_03210_),
    .I2(_03211_),
    .I3(_03212_),
    .S0(_03096_),
    .S1(_03213_),
    .Z(_03214_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07558_ (.A1(_03160_),
    .A2(_03214_),
    .ZN(_03215_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07559_ (.I0(_04840_),
    .I1(_04848_),
    .I2(_04856_),
    .I3(_04864_),
    .S0(_03057_),
    .S1(_03063_),
    .Z(_03216_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07560_ (.A1(_03150_),
    .A2(_03216_),
    .ZN(_03217_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07561_ (.A1(_03078_),
    .A2(_03045_),
    .Z(_03218_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _07562_ (.I(_01258_),
    .Z(_04833_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07563_ (.A1(net19),
    .A2(_03218_),
    .B(_02816_),
    .C(_04833_),
    .ZN(_03219_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _07564_ (.A1(_03116_),
    .A2(_03217_),
    .A3(_03219_),
    .Z(_03220_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07565_ (.A1(_03090_),
    .A2(_03220_),
    .ZN(_03221_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07566_ (.I0(net219),
    .I1(_04815_),
    .S(_02891_),
    .Z(_03222_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _07567_ (.I0(_03175_),
    .I1(_03222_),
    .S(_03078_),
    .Z(_03223_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _07568_ (.A1(_03215_),
    .A2(_03221_),
    .B1(_03223_),
    .B2(_03085_),
    .C(_03178_),
    .ZN(_03224_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07569_ (.A1(_03118_),
    .A2(_03208_),
    .B(_03224_),
    .ZN(_03225_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _07570_ (.A1(_03188_),
    .A2(_03196_),
    .A3(_03198_),
    .B(_03225_),
    .ZN(_03226_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07571_ (.I(_03226_),
    .ZN(net86));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07572_ (.A1(_02750_),
    .A2(_03052_),
    .B(net179),
    .C(_04833_),
    .ZN(_03227_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07573_ (.I0(_03046_),
    .I1(_03052_),
    .S(_03096_),
    .Z(_03228_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _07574_ (.A1(_02749_),
    .A2(_03064_),
    .A3(_03051_),
    .Z(_03229_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07575_ (.A1(_03127_),
    .A2(_03228_),
    .B(_03229_),
    .ZN(_03230_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07576_ (.A1(_03114_),
    .A2(_03227_),
    .B(_03230_),
    .ZN(_03231_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _07577_ (.A1(_02699_),
    .A2(_03076_),
    .A3(_03231_),
    .ZN(_03232_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07578_ (.I(_03127_),
    .Z(_03233_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07579_ (.I0(_05060_),
    .I1(_05074_),
    .S(_02892_),
    .Z(_03234_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07580_ (.I0(_05052_),
    .I1(_05068_),
    .S(_02892_),
    .Z(_03235_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07581_ (.I0(_03234_),
    .I1(_03235_),
    .S(_03079_),
    .Z(_03236_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07582_ (.A1(_02816_),
    .A2(_03080_),
    .ZN(_03237_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07583_ (.I(_03081_),
    .Z(_03238_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07584_ (.A1(net175),
    .A2(_03236_),
    .B(_03237_),
    .C(_03238_),
    .ZN(_03239_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07585_ (.I0(_03068_),
    .I1(_03049_),
    .S(_02816_),
    .Z(_03240_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07586_ (.A1(_03233_),
    .A2(_03239_),
    .B1(_03240_),
    .B2(_03076_),
    .ZN(_03241_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07587_ (.A1(_02699_),
    .A2(_03241_),
    .Z(_03242_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07588_ (.A1(_03038_),
    .A2(_03075_),
    .Z(_03243_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07589_ (.I0(_03056_),
    .I1(_03058_),
    .S(_03063_),
    .Z(_03244_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07590_ (.A1(_03065_),
    .A2(_03244_),
    .ZN(_03245_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07591_ (.A1(_03065_),
    .A2(_03069_),
    .B(_03245_),
    .ZN(_03246_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _07592_ (.A1(_03233_),
    .A2(_03243_),
    .A3(_03246_),
    .Z(_03247_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07593_ (.A1(_03232_),
    .A2(_03242_),
    .B(_03247_),
    .ZN(_03248_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07594_ (.A1(_05050_),
    .A2(_03138_),
    .ZN(_03249_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07595_ (.A1(_05054_),
    .A2(_02942_),
    .B(_03249_),
    .ZN(_03250_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07596_ (.A1(_03031_),
    .A2(_03250_),
    .Z(_03251_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07597_ (.A1(_02964_),
    .A2(_03026_),
    .Z(_03252_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07598_ (.I(_03023_),
    .Z(_03253_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07599_ (.A1(_02964_),
    .A2(_03253_),
    .B(_03016_),
    .ZN(_03254_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07600_ (.I0(_03252_),
    .I1(_03254_),
    .S(_05051_),
    .Z(_03255_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07601_ (.A1(_03251_),
    .A2(_03255_),
    .Z(_03256_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07602_ (.I0(_03248_),
    .I1(_03256_),
    .S(_03182_),
    .Z(net87));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _07603_ (.A1(_03053_),
    .A2(_03050_),
    .B(_04837_),
    .ZN(_03257_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _07604_ (.A1(_03099_),
    .A2(_03100_),
    .B(net163),
    .C(_03102_),
    .ZN(_03258_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07605_ (.A1(_03257_),
    .A2(_03258_),
    .ZN(_03259_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _07606_ (.A1(_03078_),
    .A2(_03105_),
    .A3(_03108_),
    .Z(_03260_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07607_ (.A1(_04840_),
    .A2(_03045_),
    .B(_03078_),
    .ZN(_03261_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07608_ (.A1(_03096_),
    .A2(_03260_),
    .A3(_03261_),
    .Z(_03262_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07609_ (.I0(_03259_),
    .I1(_03262_),
    .S(_03114_),
    .Z(_03263_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07610_ (.I0(_04900_),
    .I1(_04916_),
    .S(_03044_),
    .Z(_03264_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07611_ (.I0(_04892_),
    .I1(_04908_),
    .S(_03044_),
    .Z(_03265_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07612_ (.I0(_03264_),
    .I1(_03110_),
    .I2(_03265_),
    .I3(_03112_),
    .S0(net244),
    .S1(_01116_),
    .Z(_03266_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07613_ (.A1(_03159_),
    .A2(_03266_),
    .Z(_03267_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _07614_ (.A1(_03116_),
    .A2(_03263_),
    .B(_03267_),
    .C(_03081_),
    .ZN(_03268_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _07615_ (.I(_03038_),
    .Z(_03269_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07616_ (.I(net164),
    .Z(_03270_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07617_ (.I0(_05044_),
    .I1(_05052_),
    .I2(_05060_),
    .I3(_05068_),
    .S0(_01114_),
    .S1(_03270_),
    .Z(_03271_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07618_ (.I0(_03122_),
    .I1(_03124_),
    .I2(_03130_),
    .I3(_03271_),
    .S0(_03070_),
    .S1(_03081_),
    .Z(_03272_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07619_ (.I0(_04932_),
    .I1(_04948_),
    .S(_03062_),
    .Z(_03273_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07620_ (.I0(_04924_),
    .I1(_04940_),
    .S(_03062_),
    .Z(_03274_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07621_ (.I0(_03119_),
    .I1(_03273_),
    .I2(_03120_),
    .I3(_03274_),
    .S0(net244),
    .S1(_01116_),
    .Z(_03275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07622_ (.A1(_02749_),
    .A2(_03075_),
    .ZN(_03276_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _07623_ (.A1(net178),
    .A2(_03272_),
    .B1(_03275_),
    .B2(_03276_),
    .ZN(_03277_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07624_ (.A1(_03269_),
    .A2(_03277_),
    .Z(_03278_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07625_ (.A1(net187),
    .A2(_03268_),
    .B(_03278_),
    .ZN(_03279_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07626_ (.I(_03025_),
    .Z(_03280_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07627_ (.A1(_05073_),
    .A2(_05072_),
    .B(_05067_),
    .ZN(_03281_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07628_ (.A1(_03190_),
    .A2(_03281_),
    .ZN(_03282_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _07629_ (.A1(_05051_),
    .A2(_05059_),
    .A3(_03282_),
    .Z(_03283_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07630_ (.A1(_04814_),
    .A2(_03283_),
    .ZN(_03284_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07631_ (.A1(_05072_),
    .A2(_05067_),
    .B(_05066_),
    .ZN(_03285_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07632_ (.I(_03285_),
    .ZN(_03286_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _07633_ (.A1(_05058_),
    .A2(_05051_),
    .B1(_03283_),
    .B2(_03286_),
    .C(_05050_),
    .ZN(_03287_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07634_ (.A1(_03284_),
    .A2(_03287_),
    .Z(_03288_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _07635_ (.A1(_05043_),
    .A2(_03288_),
    .ZN(_03289_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07636_ (.A1(_05042_),
    .A2(_03017_),
    .ZN(_03290_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07637_ (.A1(_05046_),
    .A2(_02941_),
    .B(_03290_),
    .ZN(_03291_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _07638_ (.A1(_05043_),
    .A2(_03028_),
    .B1(_03280_),
    .B2(_03289_),
    .C1(_03291_),
    .C2(_02937_),
    .ZN(_03292_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07639_ (.I0(_03279_),
    .I1(_03292_),
    .S(_03178_),
    .Z(_03293_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07640_ (.I(_03293_),
    .ZN(net88));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07641_ (.I(_03136_),
    .Z(_03294_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07642_ (.I(_03112_),
    .ZN(_03295_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07643_ (.I0(_04848_),
    .I1(_04864_),
    .S(_03050_),
    .Z(_03296_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07644_ (.I0(_03092_),
    .I1(_03295_),
    .I2(_03162_),
    .I3(_03296_),
    .S0(_03096_),
    .S1(_01116_),
    .Z(_03297_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07645_ (.A1(net19),
    .A2(_03257_),
    .Z(_03298_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _07646_ (.A1(net163),
    .A2(_02892_),
    .A3(_03154_),
    .A4(_03155_),
    .ZN(_03299_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07647_ (.A1(_03083_),
    .A2(_03298_),
    .A3(_03299_),
    .Z(_03300_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07648_ (.A1(_03116_),
    .A2(_03297_),
    .B(_03300_),
    .C(_03075_),
    .ZN(_03301_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07649_ (.A1(_01115_),
    .A2(_04815_),
    .Z(_03302_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07650_ (.A1(_03057_),
    .A2(_03175_),
    .B1(_03302_),
    .B2(_03045_),
    .ZN(_03303_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07651_ (.I0(_05044_),
    .I1(_05060_),
    .S(net165),
    .Z(_03304_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07652_ (.I0(_05036_),
    .I1(_05052_),
    .S(net165),
    .Z(_03305_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07653_ (.I0(_03304_),
    .I1(_03305_),
    .S(_03042_),
    .Z(_03306_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07654_ (.I0(_03303_),
    .I1(_03173_),
    .I2(_03306_),
    .I3(_03167_),
    .S0(_03075_),
    .S1(_03054_),
    .Z(_03307_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07655_ (.I0(_03093_),
    .I1(_03161_),
    .S(_01115_),
    .Z(_03308_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07656_ (.A1(_03096_),
    .A2(_03169_),
    .Z(_03309_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07657_ (.A1(_03064_),
    .A2(_03308_),
    .B(_03309_),
    .C(_03075_),
    .ZN(_03310_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07658_ (.I0(_03307_),
    .I1(_03310_),
    .S(net178),
    .Z(_03311_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07659_ (.I0(_03301_),
    .I1(_03311_),
    .S(_03269_),
    .Z(_03312_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07660_ (.A1(_05034_),
    .A2(_03017_),
    .ZN(_03313_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07661_ (.A1(_05038_),
    .A2(_02941_),
    .B(_03313_),
    .ZN(_03314_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07662_ (.A1(_02937_),
    .A2(_03314_),
    .ZN(_03315_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07663_ (.I(_05043_),
    .ZN(_03316_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07664_ (.A1(_03316_),
    .A2(_02965_),
    .ZN(_03317_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07665_ (.A1(_05042_),
    .A2(_03317_),
    .ZN(_03318_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07666_ (.A1(_03025_),
    .A2(_03318_),
    .Z(_03319_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07667_ (.A1(_03028_),
    .A2(_03319_),
    .B(_05035_),
    .ZN(_03320_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07668_ (.A1(_05035_),
    .A2(_03023_),
    .A3(_03318_),
    .Z(_03321_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _07669_ (.A1(_03178_),
    .A2(_03315_),
    .A3(_03320_),
    .A4(_03321_),
    .Z(_03322_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07670_ (.A1(_03294_),
    .A2(_03312_),
    .B(_03322_),
    .ZN(net89));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07671_ (.I0(_05032_),
    .I1(_05048_),
    .S(_03101_),
    .Z(_03323_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07672_ (.I0(_05024_),
    .I1(_05040_),
    .S(_03101_),
    .Z(_03324_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07673_ (.I0(_03323_),
    .I1(_03324_),
    .S(_03057_),
    .Z(_03325_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _07674_ (.I0(_03223_),
    .I1(_03325_),
    .S(_03054_),
    .Z(_03326_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07675_ (.I0(_04972_),
    .I1(_04980_),
    .I2(_04988_),
    .I3(_04996_),
    .S0(_03057_),
    .S1(_03063_),
    .Z(_03327_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07676_ (.I0(_03201_),
    .I1(_03327_),
    .S(net179),
    .Z(_03328_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07677_ (.A1(_03238_),
    .A2(_03328_),
    .ZN(_03329_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07678_ (.A1(_03238_),
    .A2(_03326_),
    .B(_03329_),
    .ZN(_03330_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07679_ (.I0(_04904_),
    .I1(_04920_),
    .S(_03097_),
    .Z(_03331_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _07680_ (.I(_02228_),
    .Z(_04960_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07681_ (.I0(_04944_),
    .I1(_04960_),
    .S(_03062_),
    .Z(_03332_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07682_ (.I0(_03331_),
    .I1(_03047_),
    .I2(_03161_),
    .I3(_03332_),
    .S0(_03070_),
    .S1(_03213_),
    .Z(_03333_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07683_ (.I(_03333_),
    .ZN(_03334_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07684_ (.A1(_03269_),
    .A2(_03135_),
    .Z(_03335_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _07685_ (.A1(net222),
    .A2(_03330_),
    .B1(_03334_),
    .B2(_03276_),
    .C(_03335_),
    .ZN(_03336_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07686_ (.I0(_04844_),
    .I1(_04860_),
    .S(_03050_),
    .Z(_03337_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07687_ (.I0(_04852_),
    .I1(_04868_),
    .S(_03097_),
    .Z(_03338_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07688_ (.I0(_03337_),
    .I1(_03210_),
    .I2(_03338_),
    .I3(_03212_),
    .S0(_03070_),
    .S1(_03213_),
    .Z(_03339_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _07689_ (.A1(_01258_),
    .A2(_03070_),
    .A3(_03218_),
    .ZN(_03340_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07690_ (.I0(_04837_),
    .I1(_03340_),
    .S(_03114_),
    .Z(_03341_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07691_ (.I0(_03339_),
    .I1(_03341_),
    .S(_03116_),
    .Z(_03342_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07692_ (.A1(net187),
    .A2(_03136_),
    .Z(_03343_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07693_ (.A1(_03238_),
    .A2(_03342_),
    .B(_03343_),
    .ZN(_03344_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07694_ (.A1(_03336_),
    .A2(_03344_),
    .Z(_03345_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07695_ (.I(_05027_),
    .ZN(_03346_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _07696_ (.A1(_05035_),
    .A2(_05043_),
    .A3(_03283_),
    .ZN(_03347_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _07697_ (.A1(net247),
    .A2(net221),
    .B(_03347_),
    .ZN(_03348_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _07698_ (.A1(_03287_),
    .A2(_02966_),
    .B(_02967_),
    .ZN(_03349_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _07699_ (.A1(_03129_),
    .A2(_03348_),
    .B(_03349_),
    .ZN(_03350_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _07700_ (.A1(_03346_),
    .A2(net252),
    .ZN(_03351_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07701_ (.A1(_05026_),
    .A2(_03138_),
    .ZN(_03352_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07702_ (.A1(_05030_),
    .A2(_02942_),
    .B(_03352_),
    .ZN(_03353_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07703_ (.A1(_05027_),
    .A2(_03028_),
    .B1(_03353_),
    .B2(_03031_),
    .ZN(_03354_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07704_ (.A1(_03189_),
    .A2(_03351_),
    .B(_03354_),
    .C(_03178_),
    .ZN(_03355_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07705_ (.A1(_03345_),
    .A2(_03355_),
    .Z(net90));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _07706_ (.I(_03082_),
    .Z(_03356_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07707_ (.I0(_05028_),
    .I1(_05044_),
    .S(_02892_),
    .Z(_03357_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07708_ (.I0(_05020_),
    .I1(_05036_),
    .S(_03101_),
    .Z(_03358_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07709_ (.I0(_03234_),
    .I1(_03235_),
    .I2(_03357_),
    .I3(_03358_),
    .S0(_03079_),
    .S1(_03070_),
    .Z(_03359_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07710_ (.A1(_03150_),
    .A2(_03080_),
    .ZN(_03360_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07711_ (.I0(_03359_),
    .I1(_03360_),
    .S(_02750_),
    .Z(_03361_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07712_ (.I0(_03051_),
    .I1(_03052_),
    .S(_03064_),
    .Z(_03362_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _07713_ (.A1(net19),
    .A2(_03074_),
    .ZN(_03363_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _07714_ (.A1(_02747_),
    .A2(_02748_),
    .B(_01258_),
    .ZN(_03364_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _07715_ (.A1(_03114_),
    .A2(net166),
    .A3(_02748_),
    .A4(_03074_),
    .ZN(_03365_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _07716_ (.A1(_03363_),
    .A2(_03364_),
    .B(_03365_),
    .ZN(_03366_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07717_ (.A1(net222),
    .A2(_03362_),
    .B(_03366_),
    .ZN(_03367_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07718_ (.I0(_03046_),
    .I1(_03049_),
    .S(_03150_),
    .Z(_03368_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07719_ (.A1(_03159_),
    .A2(_03071_),
    .Z(_03369_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _07720_ (.A1(net178),
    .A2(_03368_),
    .B(_03118_),
    .C(_03369_),
    .ZN(_03370_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _07721_ (.A1(_03356_),
    .A2(_03361_),
    .B1(_03367_),
    .B2(net187),
    .C(_03370_),
    .ZN(_03371_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07722_ (.I(_05019_),
    .ZN(_03372_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07723_ (.A1(_05027_),
    .A2(_02968_),
    .B(_05026_),
    .ZN(_03373_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07724_ (.A1(_03197_),
    .A2(_03373_),
    .B(_03028_),
    .ZN(_03374_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07725_ (.A1(_05019_),
    .A2(_03253_),
    .A3(_03373_),
    .Z(_03375_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07726_ (.A1(_05018_),
    .A2(_03138_),
    .ZN(_03376_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07727_ (.A1(_05022_),
    .A2(_02942_),
    .B(_03376_),
    .ZN(_03377_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07728_ (.A1(_03031_),
    .A2(_03377_),
    .ZN(_03378_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07729_ (.A1(_03372_),
    .A2(_03374_),
    .B(_03375_),
    .C(_03378_),
    .ZN(_03379_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07730_ (.I0(_03371_),
    .I1(_03379_),
    .S(_03012_),
    .Z(net91));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _07731_ (.I(_03136_),
    .Z(_03380_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07732_ (.I(_05026_),
    .ZN(_03381_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07733_ (.A1(_03346_),
    .A2(_03350_),
    .B(_03381_),
    .ZN(_03382_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07734_ (.A1(_05019_),
    .A2(_03382_),
    .B(_05018_),
    .ZN(_03383_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _07735_ (.A1(_05011_),
    .A2(_03383_),
    .ZN(_03384_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07736_ (.A1(_05010_),
    .A2(_03018_),
    .ZN(_03385_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07737_ (.A1(_05014_),
    .A2(_03184_),
    .B(_03385_),
    .ZN(_03386_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_4 _07738_ (.A1(_05011_),
    .A2(_03144_),
    .B1(_03197_),
    .B2(_03384_),
    .C1(_03386_),
    .C2(_03183_),
    .ZN(_03387_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07739_ (.A1(_03160_),
    .A2(_03107_),
    .Z(_03388_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07740_ (.A1(_03363_),
    .A2(_03364_),
    .Z(_03389_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _07741_ (.A1(_03113_),
    .A2(_03365_),
    .B1(_03388_),
    .B2(_03389_),
    .C(_02699_),
    .ZN(_03390_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07742_ (.I0(_05012_),
    .I1(_05028_),
    .S(_03101_),
    .Z(_03391_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07743_ (.I0(_03235_),
    .I1(_03304_),
    .I2(_03358_),
    .I3(_03391_),
    .S0(_03199_),
    .S1(_03150_),
    .Z(_03392_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07744_ (.A1(net175),
    .A2(_03130_),
    .ZN(_03393_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07745_ (.A1(_03067_),
    .A2(_03393_),
    .ZN(_03394_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07746_ (.A1(net222),
    .A2(_03392_),
    .B(_03394_),
    .C(_03356_),
    .ZN(_03395_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07747_ (.A1(_03067_),
    .A2(_03094_),
    .ZN(_03396_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07748_ (.A1(net222),
    .A2(_03123_),
    .B(_03396_),
    .C(_03243_),
    .ZN(_03397_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _07749_ (.A1(_03380_),
    .A2(_03390_),
    .A3(_03395_),
    .A4(_03397_),
    .ZN(_03398_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _07750_ (.A1(_03380_),
    .A2(_03387_),
    .B(_03398_),
    .ZN(net92));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07751_ (.A1(_05002_),
    .A2(_03138_),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07752_ (.A1(_05006_),
    .A2(_03014_),
    .B(_03399_),
    .ZN(_03400_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07753_ (.I(_05018_),
    .ZN(_03401_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07754_ (.A1(_03372_),
    .A2(_03373_),
    .B(_03401_),
    .ZN(_03402_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07755_ (.A1(_05011_),
    .A2(_03402_),
    .B(_05010_),
    .ZN(_03403_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07756_ (.A1(_03026_),
    .A2(_03403_),
    .ZN(_03404_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07757_ (.A1(_03194_),
    .A2(_03404_),
    .ZN(_03405_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _07758_ (.A1(_05003_),
    .A2(_03253_),
    .A3(_03403_),
    .ZN(_03406_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _07759_ (.A1(_03013_),
    .A2(_03400_),
    .B1(_03405_),
    .B2(_05003_),
    .C(_03406_),
    .ZN(_03407_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _07760_ (.A1(_03038_),
    .A2(_03081_),
    .ZN(_03408_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07761_ (.A1(_02750_),
    .A2(_03150_),
    .ZN(_03409_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07762_ (.I0(_05004_),
    .I1(_05020_),
    .S(_03270_),
    .Z(_03410_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07763_ (.I0(_03304_),
    .I1(_03305_),
    .I2(_03391_),
    .I3(_03410_),
    .S0(_03079_),
    .S1(_03054_),
    .Z(_03411_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _07764_ (.A1(_03303_),
    .A2(_03409_),
    .B1(_03411_),
    .B2(net178),
    .ZN(_03412_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07765_ (.I0(_04976_),
    .I1(_04984_),
    .I2(net237),
    .I3(_05000_),
    .S0(_03078_),
    .S1(_03045_),
    .Z(_03413_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07766_ (.I0(_03169_),
    .I1(_03413_),
    .S(_03054_),
    .Z(_03414_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07767_ (.I0(_03163_),
    .I1(_03414_),
    .S(_03159_),
    .Z(_03415_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07768_ (.A1(net271),
    .A2(_03154_),
    .A3(_03155_),
    .B(net179),
    .ZN(_03416_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07769_ (.A1(net19),
    .A2(_03074_),
    .Z(_03417_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _07770_ (.A1(_01258_),
    .A2(net271),
    .A3(_03417_),
    .Z(_03418_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07771_ (.A1(_03416_),
    .A2(_03366_),
    .B(_03418_),
    .ZN(_03419_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07772_ (.A1(_03064_),
    .A2(_03151_),
    .Z(_03420_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _07773_ (.A1(_03127_),
    .A2(_03389_),
    .B1(_03419_),
    .B2(_03420_),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _07774_ (.A1(_03408_),
    .A2(_03412_),
    .B1(_03415_),
    .B2(_03118_),
    .C1(_03421_),
    .C2(_03269_),
    .ZN(_03422_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07775_ (.I0(_03407_),
    .I1(_03422_),
    .S(_03294_),
    .Z(_03423_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _07776_ (.I(_03423_),
    .ZN(net62));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07777_ (.I0(_04996_),
    .I1(_05012_),
    .S(_03270_),
    .Z(_03424_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07778_ (.I0(_03305_),
    .I1(_03357_),
    .I2(_03410_),
    .I3(_03424_),
    .S0(_03213_),
    .S1(_03064_),
    .Z(_03425_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07779_ (.A1(_03065_),
    .A2(_03223_),
    .B(_03160_),
    .ZN(_03426_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _07780_ (.A1(_03233_),
    .A2(_03425_),
    .B(_03426_),
    .ZN(_03427_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07781_ (.I0(_03214_),
    .I1(_03207_),
    .S(_03127_),
    .Z(_03428_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07782_ (.A1(_03243_),
    .A2(_03428_),
    .ZN(_03429_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _07783_ (.A1(_04833_),
    .A2(net179),
    .A3(_03218_),
    .ZN(_03430_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07784_ (.A1(_03217_),
    .A2(_03430_),
    .Z(_03431_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07785_ (.I0(_04833_),
    .I1(_03216_),
    .S(_03150_),
    .Z(_03432_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _07786_ (.A1(_03363_),
    .A2(_03364_),
    .ZN(_03433_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07787_ (.A1(net178),
    .A2(_03432_),
    .B(_03433_),
    .ZN(_03434_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07788_ (.A1(_03365_),
    .A2(_03431_),
    .B(_03434_),
    .C(_02699_),
    .ZN(_03435_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _07789_ (.A1(_03408_),
    .A2(_03427_),
    .B(_03429_),
    .C(_03435_),
    .ZN(_03436_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07790_ (.I(_02969_),
    .ZN(_03437_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07791_ (.A1(_03437_),
    .A2(_03350_),
    .B(_02955_),
    .ZN(_03438_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _07792_ (.A1(_02950_),
    .A2(_03438_),
    .ZN(_03439_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07793_ (.A1(_04994_),
    .A2(_03138_),
    .ZN(_03440_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07794_ (.A1(_04998_),
    .A2(_02942_),
    .B(_03440_),
    .ZN(_03441_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _07795_ (.A1(_04995_),
    .A2(_03144_),
    .B1(_03280_),
    .B2(_03439_),
    .C1(_03441_),
    .C2(_03031_),
    .ZN(_03442_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07796_ (.A1(_03012_),
    .A2(_03442_),
    .Z(_03443_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _07797_ (.A1(_03380_),
    .A2(_03436_),
    .B(_03443_),
    .ZN(net63));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07798_ (.A1(_04986_),
    .A2(_03139_),
    .ZN(_03444_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07799_ (.A1(_04990_),
    .A2(_03184_),
    .B(_03444_),
    .ZN(_03445_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07800_ (.A1(_02968_),
    .A2(_02969_),
    .ZN(_03446_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07801_ (.A1(_02955_),
    .A2(_03446_),
    .B(_02950_),
    .ZN(_03447_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07802_ (.A1(_04994_),
    .A2(_03447_),
    .Z(_03448_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07803_ (.A1(_03026_),
    .A2(_03448_),
    .Z(_03449_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07804_ (.A1(_03253_),
    .A2(_03448_),
    .B(_03194_),
    .ZN(_03450_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07805_ (.I0(_03449_),
    .I1(_03450_),
    .S(_04987_),
    .Z(_03451_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07806_ (.A1(_03183_),
    .A2(_03445_),
    .B(_03451_),
    .ZN(_03452_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07807_ (.A1(_03380_),
    .A2(_03452_),
    .ZN(_03453_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07808_ (.I0(_03228_),
    .I1(_03240_),
    .S(_03127_),
    .Z(_03454_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07809_ (.A1(_03118_),
    .A2(_03454_),
    .Z(_03455_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _07810_ (.A1(net175),
    .A2(_03236_),
    .B(_03237_),
    .ZN(_03456_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07811_ (.I0(_04988_),
    .I1(_05004_),
    .S(_03101_),
    .Z(_03457_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07812_ (.I0(_03357_),
    .I1(_03358_),
    .I2(_03424_),
    .I3(_03457_),
    .S0(_03079_),
    .S1(_03054_),
    .Z(_03458_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07813_ (.A1(_03116_),
    .A2(_03458_),
    .ZN(_03459_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _07814_ (.A1(net178),
    .A2(_03456_),
    .B(_03459_),
    .C(_03076_),
    .ZN(_03460_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _07815_ (.A1(_03076_),
    .A2(_03051_),
    .A3(_03084_),
    .ZN(_03461_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _07816_ (.A1(_04833_),
    .A2(_03417_),
    .ZN(_03462_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07817_ (.A1(_03269_),
    .A2(_03084_),
    .A3(_03462_),
    .Z(_03463_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07818_ (.A1(_02699_),
    .A2(_03460_),
    .B(_03461_),
    .C(_03463_),
    .ZN(_03464_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _07819_ (.A1(_03294_),
    .A2(_03455_),
    .A3(_03464_),
    .Z(_03465_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07820_ (.A1(_03453_),
    .A2(_03465_),
    .Z(net64));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _07821_ (.A1(_04995_),
    .A2(_03438_),
    .B(_04994_),
    .C(_04986_),
    .ZN(_03466_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07822_ (.A1(_02959_),
    .A2(_03466_),
    .B(_03197_),
    .ZN(_03467_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07823_ (.A1(_03194_),
    .A2(_03467_),
    .B(_02958_),
    .ZN(_03468_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07824_ (.A1(_04978_),
    .A2(_03018_),
    .ZN(_03469_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07825_ (.A1(_04982_),
    .A2(_03014_),
    .B(_03469_),
    .ZN(_03470_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07826_ (.A1(_03013_),
    .A2(_03470_),
    .ZN(_03471_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _07827_ (.A1(_04979_),
    .A2(_02959_),
    .A3(_03253_),
    .A4(_03466_),
    .Z(_03472_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07828_ (.A1(_03471_),
    .A2(_03472_),
    .ZN(_03473_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07829_ (.I0(_03130_),
    .I1(_03271_),
    .S(_03070_),
    .Z(_03474_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07830_ (.I0(_04980_),
    .I1(_04996_),
    .S(_02892_),
    .Z(_03475_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07831_ (.I0(_03358_),
    .I1(_03391_),
    .I2(_03457_),
    .I3(_03475_),
    .S0(_03057_),
    .S1(_03070_),
    .Z(_03476_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07832_ (.I0(_03474_),
    .I1(_03476_),
    .S(_03083_),
    .Z(_03477_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07833_ (.I0(_03266_),
    .I1(_03275_),
    .S(_03159_),
    .Z(_03478_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07834_ (.A1(_02749_),
    .A2(_03257_),
    .A3(_03258_),
    .B(_03433_),
    .ZN(_03479_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _07835_ (.A1(_02816_),
    .A2(_03260_),
    .A3(_03261_),
    .A4(_03365_),
    .Z(_03480_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _07836_ (.A1(net253),
    .A2(_03479_),
    .A3(_03480_),
    .Z(_03481_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _07837_ (.A1(_03356_),
    .A2(_03477_),
    .B1(_03478_),
    .B2(_03243_),
    .C(_03481_),
    .ZN(_03482_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07838_ (.A1(_03178_),
    .A2(_03482_),
    .Z(_03483_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07839_ (.A1(_03380_),
    .A2(_03468_),
    .A3(_03473_),
    .B(_03483_),
    .ZN(_03484_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07840_ (.I(_03484_),
    .ZN(net65));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _07841_ (.A1(_03199_),
    .A2(_03175_),
    .B1(_03302_),
    .B2(_03063_),
    .C(_03064_),
    .ZN(_03485_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _07842_ (.A1(_03065_),
    .A2(_03306_),
    .B(_03485_),
    .ZN(_03486_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07843_ (.I0(_03308_),
    .I1(_03169_),
    .S(_03150_),
    .Z(_03487_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07844_ (.I0(net176),
    .I1(_05024_),
    .S(_03102_),
    .Z(_03488_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07845_ (.I0(_05000_),
    .I1(net173),
    .S(_03270_),
    .Z(_03489_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07846_ (.I0(_04976_),
    .I1(net237),
    .S(_03102_),
    .Z(_03490_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07847_ (.I0(_04968_),
    .I1(_04984_),
    .S(_03270_),
    .Z(_03491_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07848_ (.I0(_03488_),
    .I1(_03489_),
    .I2(_03490_),
    .I3(_03491_),
    .S0(_03213_),
    .S1(_03064_),
    .Z(_03492_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07849_ (.I0(_03297_),
    .I1(_03486_),
    .I2(_03487_),
    .I3(_03492_),
    .S0(_03238_),
    .S1(_03233_),
    .Z(_03493_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07850_ (.A1(_02699_),
    .A2(_03493_),
    .ZN(_03494_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07851_ (.A1(_03067_),
    .A2(_03257_),
    .Z(_03495_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _07852_ (.A1(_03299_),
    .A2(_03366_),
    .B1(_03495_),
    .B2(_03433_),
    .C(_03039_),
    .ZN(_03496_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07853_ (.A1(_02971_),
    .A2(_03197_),
    .B(_03028_),
    .ZN(_03497_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07854_ (.A1(_04971_),
    .A2(_02971_),
    .A3(_03253_),
    .Z(_03498_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07855_ (.A1(_04970_),
    .A2(_03138_),
    .ZN(_03499_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07856_ (.A1(_04974_),
    .A2(_03014_),
    .B(_03499_),
    .ZN(_03500_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07857_ (.A1(_03013_),
    .A2(_03500_),
    .ZN(_03501_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07858_ (.A1(_02972_),
    .A2(_03497_),
    .B(_03498_),
    .C(_03501_),
    .ZN(_03502_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07859_ (.A1(_03182_),
    .A2(_03502_),
    .ZN(_03503_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _07860_ (.A1(_03182_),
    .A2(_03494_),
    .A3(_03496_),
    .B(_03503_),
    .ZN(net66));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07861_ (.I(_02970_),
    .ZN(_03504_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _07862_ (.A1(_02957_),
    .A2(_02960_),
    .B(_04978_),
    .ZN(_03505_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07863_ (.A1(_03504_),
    .A2(_03350_),
    .B(_03505_),
    .ZN(_03506_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07864_ (.A1(_04971_),
    .A2(_03506_),
    .B(_04970_),
    .ZN(_03507_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _07865_ (.A1(_04963_),
    .A2(_03507_),
    .ZN(_03508_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07866_ (.A1(_04962_),
    .A2(_03018_),
    .ZN(_03509_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07867_ (.A1(_04966_),
    .A2(_03014_),
    .B(_03509_),
    .ZN(_03510_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_4 _07868_ (.A1(_04963_),
    .A2(_03144_),
    .B1(_03197_),
    .B2(_03508_),
    .C1(_03510_),
    .C2(_03013_),
    .ZN(_03511_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07869_ (.A1(_03182_),
    .A2(_03511_),
    .ZN(_03512_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07870_ (.I0(net237),
    .I1(net176),
    .S(_03270_),
    .Z(_03513_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07871_ (.I0(net243),
    .I1(_04976_),
    .S(_03270_),
    .Z(_03514_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07872_ (.I0(_03489_),
    .I1(_03513_),
    .I2(_03491_),
    .I3(_03514_),
    .S0(_03213_),
    .S1(_03054_),
    .Z(_03515_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07873_ (.I0(_03326_),
    .I1(_03515_),
    .S(_03159_),
    .Z(_03516_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07874_ (.A1(_03356_),
    .A2(_03516_),
    .Z(_03517_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07875_ (.I0(_03334_),
    .I1(_03339_),
    .S(_02750_),
    .Z(_03518_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07876_ (.A1(_03118_),
    .A2(_03518_),
    .ZN(_03519_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07877_ (.A1(_03340_),
    .A2(_03365_),
    .Z(_03520_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07878_ (.A1(_03039_),
    .A2(_03518_),
    .B1(_03520_),
    .B2(_03462_),
    .ZN(_03521_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _07879_ (.A1(_03012_),
    .A2(_03517_),
    .A3(_03519_),
    .A4(_03521_),
    .Z(_03522_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07880_ (.A1(_03512_),
    .A2(_03522_),
    .Z(net67));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07881_ (.A1(_03075_),
    .A2(_03055_),
    .Z(_03523_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07882_ (.I0(_04964_),
    .I1(_04980_),
    .I2(_04996_),
    .I3(_05012_),
    .S0(_03270_),
    .S1(_02814_),
    .Z(_03524_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07883_ (.I0(_04956_),
    .I1(_04972_),
    .I2(_04988_),
    .I3(_05004_),
    .S0(_02892_),
    .S1(_02814_),
    .Z(_03525_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07884_ (.I0(_03524_),
    .I1(_03525_),
    .S(_03079_),
    .Z(_03526_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07885_ (.I0(_03359_),
    .I1(_03526_),
    .S(_03159_),
    .Z(_03527_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07886_ (.A1(_03076_),
    .A2(_03527_),
    .ZN(_03528_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07887_ (.A1(_03083_),
    .A2(_03081_),
    .Z(_03529_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07888_ (.I(_03529_),
    .ZN(_03530_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07889_ (.A1(_03360_),
    .A2(_03530_),
    .B(_03462_),
    .C(net187),
    .ZN(_03531_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07890_ (.A1(net250),
    .A2(_03523_),
    .A3(_03528_),
    .B(_03531_),
    .ZN(_03532_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07891_ (.I(_04970_),
    .ZN(_03533_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07892_ (.A1(_02972_),
    .A2(_02971_),
    .B(_03533_),
    .ZN(_03534_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _07893_ (.A1(_04963_),
    .A2(_03534_),
    .B(_04962_),
    .C(_04955_),
    .ZN(_03535_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07894_ (.A1(_02977_),
    .A2(_03535_),
    .ZN(_03536_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07895_ (.A1(_04954_),
    .A2(_03138_),
    .ZN(_03537_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07896_ (.A1(_04958_),
    .A2(_02942_),
    .B(_03537_),
    .ZN(_03538_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _07897_ (.A1(_04955_),
    .A2(_03144_),
    .B1(_03280_),
    .B2(_03536_),
    .C1(_03538_),
    .C2(_03031_),
    .ZN(_03539_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07898_ (.I0(_03532_),
    .I1(_03539_),
    .S(_03178_),
    .Z(_03540_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07899_ (.I(_03540_),
    .ZN(net68));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _07900_ (.A1(_04955_),
    .A2(_04962_),
    .B(_04954_),
    .ZN(_03541_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07901_ (.A1(_02973_),
    .A2(_03507_),
    .B(_03541_),
    .ZN(_03542_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _07902_ (.A1(_02984_),
    .A2(_03542_),
    .ZN(_03543_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07903_ (.A1(_04946_),
    .A2(_03018_),
    .ZN(_03544_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07904_ (.A1(_04950_),
    .A2(_03014_),
    .B(_03544_),
    .ZN(_03545_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_4 _07905_ (.A1(_04947_),
    .A2(_03144_),
    .B1(_03197_),
    .B2(_03543_),
    .C1(_03545_),
    .C2(_03013_),
    .ZN(_03546_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _07906_ (.A1(_04837_),
    .A2(net254),
    .B(_03363_),
    .ZN(_03547_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07907_ (.A1(_03393_),
    .A2(_03529_),
    .B(_03547_),
    .ZN(_03548_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07908_ (.I(_03462_),
    .ZN(_03549_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07909_ (.I0(_04944_),
    .I1(_04960_),
    .I2(_04976_),
    .I3(net237),
    .S0(_03102_),
    .S1(_02814_),
    .Z(_03550_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07910_ (.A1(_03199_),
    .A2(_03550_),
    .ZN(_03551_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07911_ (.A1(_03199_),
    .A2(_03525_),
    .B(_03551_),
    .ZN(_03552_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07912_ (.I0(_03094_),
    .I1(_03552_),
    .S(_03081_),
    .Z(_03553_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07913_ (.A1(_03094_),
    .A2(_03549_),
    .B1(_03553_),
    .B2(_03039_),
    .ZN(_03554_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07914_ (.A1(_04833_),
    .A2(_03038_),
    .B(_03417_),
    .ZN(_03555_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07915_ (.A1(_03114_),
    .A2(_03074_),
    .ZN(_03556_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _07916_ (.A1(net253),
    .A2(_03556_),
    .Z(_03557_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _07917_ (.A1(_03408_),
    .A2(_03392_),
    .B1(_03555_),
    .B2(_03107_),
    .C1(_03557_),
    .C2(_03113_),
    .ZN(_03558_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07918_ (.A1(net222),
    .A2(_03558_),
    .ZN(_03559_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _07919_ (.A1(_03039_),
    .A2(_03548_),
    .B1(_03554_),
    .B2(net222),
    .C(_03559_),
    .ZN(_03560_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07920_ (.A1(_03182_),
    .A2(_03560_),
    .ZN(_03561_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07921_ (.A1(_03182_),
    .A2(_03546_),
    .B(_03561_),
    .ZN(net69));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _07922_ (.A1(_03105_),
    .A2(_03157_),
    .B(_03420_),
    .C(_03233_),
    .ZN(_03562_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _07923_ (.A1(_02699_),
    .A2(_03164_),
    .A3(_03562_),
    .B(_03547_),
    .ZN(_03563_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _07924_ (.I(_03557_),
    .ZN(_03564_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _07925_ (.A1(_02750_),
    .A2(_03152_),
    .A3(_03416_),
    .Z(_03565_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07926_ (.A1(_03164_),
    .A2(_03565_),
    .Z(_03566_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07927_ (.A1(_02750_),
    .A2(_03411_),
    .Z(_03567_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07928_ (.I0(_04936_),
    .I1(_04952_),
    .I2(_04968_),
    .I3(_04984_),
    .S0(net271),
    .S1(_03096_),
    .Z(_03568_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07929_ (.I0(_03550_),
    .I1(_03568_),
    .S(_03199_),
    .Z(_03569_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07930_ (.A1(_03067_),
    .A2(_03569_),
    .ZN(_03570_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07931_ (.A1(_02697_),
    .A2(_03081_),
    .Z(_03571_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07932_ (.A1(_03084_),
    .A2(_03571_),
    .Z(_03572_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07933_ (.A1(_03177_),
    .A2(_03572_),
    .B(_03011_),
    .ZN(_03573_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07934_ (.A1(_03408_),
    .A2(_03567_),
    .A3(_03570_),
    .B(_03573_),
    .ZN(_03574_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _07935_ (.A1(_03564_),
    .A2(_03566_),
    .B(_03574_),
    .ZN(_03575_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07936_ (.A1(_04938_),
    .A2(_03139_),
    .ZN(_03576_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07937_ (.A1(_04942_),
    .A2(_03184_),
    .B(_03576_),
    .ZN(_03577_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07938_ (.A1(_03183_),
    .A2(_03577_),
    .B(_03380_),
    .ZN(_03578_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07939_ (.A1(_02971_),
    .A2(_02974_),
    .B(_02976_),
    .C(_02982_),
    .ZN(_03579_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07940_ (.A1(_03579_),
    .A2(_04947_),
    .B(_04946_),
    .ZN(_03580_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07941_ (.A1(_03580_),
    .A2(_03197_),
    .Z(_03581_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07942_ (.A1(_03580_),
    .A2(_03189_),
    .B(_02979_),
    .ZN(_03582_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07943_ (.A1(_02979_),
    .A2(_03144_),
    .A3(_03581_),
    .B(_03582_),
    .ZN(_03583_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _07944_ (.A1(_03563_),
    .A2(_03575_),
    .B1(_03578_),
    .B2(_03583_),
    .ZN(net70));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07945_ (.A1(_03067_),
    .A2(_03432_),
    .ZN(_03584_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07946_ (.A1(net222),
    .A2(_03214_),
    .B(_03584_),
    .C(_03039_),
    .ZN(_03585_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07947_ (.A1(net222),
    .A2(_03431_),
    .B(_03557_),
    .ZN(_03586_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07948_ (.I0(_04940_),
    .I1(_04956_),
    .I2(_04972_),
    .I3(_04988_),
    .S0(_03102_),
    .S1(_03096_),
    .Z(_03587_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07949_ (.I0(_04932_),
    .I1(_04948_),
    .I2(_04964_),
    .I3(_04980_),
    .S0(_03102_),
    .S1(net163),
    .Z(_03588_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07950_ (.I0(_03587_),
    .I1(_03588_),
    .S(_03213_),
    .Z(_03589_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07951_ (.I0(_03425_),
    .I1(_03589_),
    .S(_03127_),
    .Z(_03590_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07952_ (.A1(_03223_),
    .A2(_03572_),
    .ZN(_03591_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07953_ (.A1(_03408_),
    .A2(_03590_),
    .B(_03591_),
    .C(_03136_),
    .ZN(_03592_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _07954_ (.A1(_03547_),
    .A2(_03585_),
    .B1(_03586_),
    .B2(_03215_),
    .C(_03592_),
    .ZN(_03593_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07955_ (.A1(_04930_),
    .A2(_03018_),
    .ZN(_03594_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07956_ (.A1(_04934_),
    .A2(_03014_),
    .B(_03594_),
    .ZN(_03595_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07957_ (.A1(_03013_),
    .A2(_03595_),
    .ZN(_03596_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07958_ (.A1(_02973_),
    .A2(_03541_),
    .B(_02984_),
    .ZN(_03597_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07959_ (.A1(_04946_),
    .A2(_03597_),
    .Z(_03598_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07960_ (.A1(_04939_),
    .A2(_03598_),
    .B(_04938_),
    .ZN(_03599_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07961_ (.I(_04938_),
    .ZN(_03600_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07962_ (.A1(_02984_),
    .A2(_03541_),
    .B(_02980_),
    .ZN(_03601_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07963_ (.A1(_04939_),
    .A2(_03601_),
    .ZN(_03602_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _07964_ (.A1(_03600_),
    .A2(_03505_),
    .A3(_03533_),
    .A4(_03602_),
    .ZN(_03603_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _07965_ (.A1(_03129_),
    .A2(_03348_),
    .B(_03349_),
    .C(_03603_),
    .ZN(_03604_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07966_ (.A1(_03600_),
    .A2(_03602_),
    .ZN(_03605_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07967_ (.A1(_04970_),
    .A2(_02970_),
    .A3(_03605_),
    .Z(_03606_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07968_ (.I(_03505_),
    .ZN(_03607_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _07969_ (.A1(_04970_),
    .A2(_04971_),
    .A3(_03605_),
    .B1(_03606_),
    .B2(_03607_),
    .ZN(_03608_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07970_ (.A1(_03599_),
    .A2(_03604_),
    .A3(_03608_),
    .Z(_03609_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07971_ (.A1(_03280_),
    .A2(_03609_),
    .Z(_03610_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07972_ (.A1(_03144_),
    .A2(_03610_),
    .B(_04931_),
    .ZN(_03611_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07973_ (.A1(_04931_),
    .A2(_03189_),
    .A3(_03609_),
    .Z(_03612_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _07974_ (.A1(_03012_),
    .A2(_03596_),
    .A3(_03611_),
    .A4(_03612_),
    .Z(_03613_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _07975_ (.A1(_03593_),
    .A2(_03613_),
    .ZN(net71));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07976_ (.A1(_02979_),
    .A2(_03580_),
    .B(_03600_),
    .ZN(_03614_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07977_ (.A1(_04931_),
    .A2(_03614_),
    .B(_04930_),
    .ZN(_03615_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07978_ (.A1(_03197_),
    .A2(_03615_),
    .ZN(_03616_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07979_ (.A1(_03194_),
    .A2(_03616_),
    .B(_02986_),
    .ZN(_03617_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07980_ (.A1(_04922_),
    .A2(_03138_),
    .ZN(_03618_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07981_ (.A1(_04926_),
    .A2(_02942_),
    .B(_03618_),
    .ZN(_03619_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07982_ (.A1(_03031_),
    .A2(_03619_),
    .ZN(_03620_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07983_ (.A1(_04923_),
    .A2(_03189_),
    .A3(_03615_),
    .B(_03620_),
    .ZN(_03621_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07984_ (.I0(_04928_),
    .I1(_04944_),
    .S(_03101_),
    .Z(_03622_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07985_ (.I0(_04920_),
    .I1(_04936_),
    .S(_02892_),
    .Z(_03623_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07986_ (.I0(_03622_),
    .I1(_03623_),
    .S(_03057_),
    .Z(_03624_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07987_ (.I0(net263),
    .I1(_04968_),
    .S(_02892_),
    .Z(_03625_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07988_ (.I0(_03514_),
    .I1(_03625_),
    .S(_03079_),
    .Z(_03626_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07989_ (.I0(_03624_),
    .I1(_03626_),
    .S(net175),
    .Z(_03627_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07990_ (.I0(_03456_),
    .I1(_03627_),
    .S(_03269_),
    .Z(_03628_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07991_ (.A1(_03529_),
    .A2(_03628_),
    .Z(_03629_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07992_ (.A1(_03118_),
    .A2(_03462_),
    .B(_03230_),
    .ZN(_03630_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07993_ (.A1(_03269_),
    .A2(_03227_),
    .B(_03555_),
    .ZN(_03631_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _07994_ (.A1(_03160_),
    .A2(_03408_),
    .A3(_03458_),
    .ZN(_03632_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _07995_ (.A1(_03178_),
    .A2(_03630_),
    .A3(_03631_),
    .A4(_03632_),
    .Z(_03633_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _07996_ (.A1(_03617_),
    .A2(_03621_),
    .A3(_03380_),
    .B1(_03629_),
    .B2(_03633_),
    .ZN(_03634_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07997_ (.I(_03634_),
    .ZN(net73));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07998_ (.I0(_04912_),
    .I1(_04928_),
    .I2(_04944_),
    .I3(_04960_),
    .S0(net271),
    .S1(_03096_),
    .Z(_03635_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07999_ (.I0(_03625_),
    .I1(_03623_),
    .S(_03070_),
    .Z(_03636_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08000_ (.I0(_03635_),
    .I1(_03636_),
    .S(_01116_),
    .Z(_03637_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08001_ (.A1(_03269_),
    .A2(_03075_),
    .A3(_03474_),
    .ZN(_03638_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08002_ (.A1(_03266_),
    .A2(_03557_),
    .ZN(_03639_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08003_ (.A1(_03356_),
    .A2(_03637_),
    .B(_03638_),
    .C(_03639_),
    .ZN(_03640_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _08004_ (.A1(_03408_),
    .A2(_03476_),
    .B1(_03557_),
    .B2(_03262_),
    .ZN(_03641_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08005_ (.I(_03641_),
    .ZN(_03642_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08006_ (.I0(_03640_),
    .I1(_03642_),
    .S(net222),
    .Z(_03643_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08007_ (.I0(_03259_),
    .I1(_03266_),
    .S(_03160_),
    .Z(_03644_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08008_ (.A1(_03039_),
    .A2(_03644_),
    .ZN(_03645_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08009_ (.A1(_03547_),
    .A2(_03645_),
    .B(_03012_),
    .ZN(_03646_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08010_ (.A1(_02981_),
    .A2(_03599_),
    .Z(_03647_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08011_ (.A1(_04923_),
    .A2(_04930_),
    .B(_04922_),
    .ZN(_03648_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _08012_ (.A1(_03647_),
    .A2(_03608_),
    .A3(_03604_),
    .B(_03648_),
    .ZN(_03649_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08013_ (.A1(_03189_),
    .A2(_03649_),
    .B(_03194_),
    .ZN(_03650_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08014_ (.A1(_04914_),
    .A2(_03018_),
    .ZN(_03651_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08015_ (.A1(_04918_),
    .A2(_03184_),
    .B(_03651_),
    .ZN(_03652_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08016_ (.I(_04915_),
    .ZN(_03653_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08017_ (.A1(_03653_),
    .A2(_03280_),
    .A3(net265),
    .Z(_03654_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _08018_ (.A1(_04915_),
    .A2(_03650_),
    .B1(_03652_),
    .B2(_03183_),
    .C(_03654_),
    .ZN(_03655_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _08019_ (.A1(_03643_),
    .A2(_03646_),
    .B1(_03655_),
    .B2(_03182_),
    .ZN(net74));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08020_ (.A1(_04906_),
    .A2(_03139_),
    .ZN(_03656_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08021_ (.A1(_04910_),
    .A2(_03184_),
    .B(_03656_),
    .ZN(_03657_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08022_ (.A1(_02977_),
    .A2(_02978_),
    .B(_02985_),
    .C(_02989_),
    .ZN(_03658_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08023_ (.I(_04914_),
    .ZN(_03659_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08024_ (.A1(_03653_),
    .A2(_03658_),
    .B(_03659_),
    .ZN(_03660_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08025_ (.A1(_03660_),
    .A2(_03026_),
    .Z(_03661_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08026_ (.A1(_03660_),
    .A2(_03253_),
    .B(_03194_),
    .ZN(_03662_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08027_ (.I0(_03661_),
    .I1(_03662_),
    .S(_04907_),
    .Z(_03663_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08028_ (.A1(_03183_),
    .A2(_03657_),
    .B(_03663_),
    .ZN(_03664_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _08029_ (.A1(net253),
    .A2(_03083_),
    .A3(_03257_),
    .A4(_03299_),
    .Z(_03665_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08030_ (.A1(_03038_),
    .A2(_03083_),
    .ZN(_03666_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08031_ (.A1(_03547_),
    .A2(_03665_),
    .A3(_03666_),
    .Z(_03667_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08032_ (.A1(_03127_),
    .A2(_03564_),
    .Z(_03668_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08033_ (.A1(_03547_),
    .A2(_03665_),
    .Z(_03669_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _08034_ (.A1(_03297_),
    .A2(_03667_),
    .B1(_03668_),
    .B2(_03669_),
    .ZN(_03670_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08035_ (.I0(_04904_),
    .I1(_04920_),
    .I2(_04936_),
    .I3(net263),
    .S0(_03270_),
    .S1(net163),
    .Z(_03671_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08036_ (.I0(_03635_),
    .I1(_03671_),
    .S(_03199_),
    .Z(_03672_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08037_ (.A1(_03160_),
    .A2(_03672_),
    .Z(_03673_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08038_ (.A1(_03116_),
    .A2(_03492_),
    .Z(_03674_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08039_ (.A1(_03673_),
    .A2(_03674_),
    .B(_03356_),
    .ZN(_03675_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08040_ (.A1(_03159_),
    .A2(_03571_),
    .Z(_03676_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08041_ (.A1(_03116_),
    .A2(_03299_),
    .A3(_03564_),
    .Z(_03677_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08042_ (.A1(_03486_),
    .A2(_03676_),
    .B(_03677_),
    .ZN(_03678_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08043_ (.A1(_03294_),
    .A2(_03670_),
    .A3(_03675_),
    .A4(_03678_),
    .Z(_03679_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08044_ (.A1(_03182_),
    .A2(_03664_),
    .B(_03679_),
    .ZN(net75));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08045_ (.A1(_03159_),
    .A2(_03564_),
    .ZN(_03680_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08046_ (.A1(_03038_),
    .A2(_03083_),
    .Z(_03681_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08047_ (.A1(_04833_),
    .A2(_03681_),
    .B(_03417_),
    .ZN(_03682_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08048_ (.A1(_03680_),
    .A2(_03682_),
    .B(_03339_),
    .ZN(_03683_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08049_ (.A1(_03340_),
    .A2(_03557_),
    .B(_03682_),
    .ZN(_03684_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08050_ (.A1(_03666_),
    .A2(_03684_),
    .Z(_03685_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08051_ (.A1(_03326_),
    .A2(_03676_),
    .Z(_03686_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _08052_ (.A1(_03178_),
    .A2(_03683_),
    .A3(_03685_),
    .A4(_03686_),
    .Z(_03687_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08053_ (.I0(_04896_),
    .I1(_04912_),
    .S(_03101_),
    .Z(_03688_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08054_ (.I0(_03622_),
    .I1(_03688_),
    .S(_03053_),
    .Z(_03689_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08055_ (.I0(_03671_),
    .I1(_03689_),
    .S(_03213_),
    .Z(_03690_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08056_ (.A1(_03233_),
    .A2(_03690_),
    .ZN(_03691_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08057_ (.A1(_03067_),
    .A2(_03515_),
    .ZN(_03692_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08058_ (.A1(_03691_),
    .A2(_03692_),
    .B(_03408_),
    .ZN(_03693_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08059_ (.A1(_03687_),
    .A2(_03693_),
    .Z(_03694_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08060_ (.I(_04899_),
    .ZN(_03695_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08061_ (.A1(_04907_),
    .A2(_04915_),
    .Z(_03696_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _08062_ (.A1(_04907_),
    .A2(_04914_),
    .B1(_03649_),
    .B2(_03696_),
    .C(_04906_),
    .ZN(_03697_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08063_ (.A1(_03197_),
    .A2(_03697_),
    .B(_03144_),
    .ZN(_03698_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08064_ (.A1(_04899_),
    .A2(_03189_),
    .A3(_03697_),
    .Z(_03699_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08065_ (.A1(_04898_),
    .A2(_03018_),
    .ZN(_03700_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08066_ (.A1(_04902_),
    .A2(_03014_),
    .B(_03700_),
    .ZN(_03701_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08067_ (.A1(_03013_),
    .A2(_03701_),
    .B(_03294_),
    .ZN(_03702_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08068_ (.A1(_03695_),
    .A2(_03698_),
    .B(_03699_),
    .C(_03702_),
    .ZN(_03703_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08069_ (.A1(_03694_),
    .A2(_03703_),
    .Z(net76));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08070_ (.I(_03526_),
    .ZN(_03704_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08071_ (.I0(_04888_),
    .I1(_04904_),
    .S(_03270_),
    .Z(_03705_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08072_ (.I0(_03688_),
    .I1(_03705_),
    .S(_03079_),
    .Z(_03706_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08073_ (.I0(_03624_),
    .I1(_03706_),
    .S(_03150_),
    .Z(_03707_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08074_ (.I0(_03704_),
    .I1(_03707_),
    .S(_03160_),
    .Z(_03708_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08075_ (.I(_03367_),
    .ZN(_03709_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08076_ (.A1(_03238_),
    .A2(_03708_),
    .B(_03709_),
    .ZN(_03710_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08077_ (.A1(_03076_),
    .A2(_03361_),
    .Z(_03711_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08078_ (.A1(_03462_),
    .A2(_03711_),
    .Z(_03712_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08079_ (.I0(_03710_),
    .I1(_03712_),
    .S(_02699_),
    .Z(_03713_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08080_ (.A1(_04890_),
    .A2(_03139_),
    .ZN(_03714_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08081_ (.A1(_04894_),
    .A2(_03184_),
    .B(_03714_),
    .ZN(_03715_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08082_ (.I(_04898_),
    .ZN(_03716_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _08083_ (.A1(_03695_),
    .A2(_02991_),
    .A3(_02993_),
    .B(_03716_),
    .ZN(_03717_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08084_ (.A1(_03717_),
    .A2(_03026_),
    .Z(_03718_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08085_ (.A1(_03253_),
    .A2(_03717_),
    .B(_03016_),
    .ZN(_03719_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08086_ (.I0(_03718_),
    .I1(_03719_),
    .S(_04891_),
    .Z(_03720_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08087_ (.A1(_03183_),
    .A2(_03715_),
    .B(_03294_),
    .C(_03720_),
    .ZN(_03721_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08088_ (.A1(_03380_),
    .A2(_03713_),
    .B(_03721_),
    .ZN(net77));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08089_ (.A1(_03113_),
    .A2(_03680_),
    .Z(_03722_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08090_ (.I0(_04912_),
    .I1(_04928_),
    .S(net271),
    .Z(_03723_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08091_ (.I0(_04880_),
    .I1(_04896_),
    .S(_03102_),
    .Z(_03724_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08092_ (.I0(_03623_),
    .I1(_03723_),
    .I2(_03705_),
    .I3(_03724_),
    .S0(_03199_),
    .S1(_03150_),
    .Z(_03725_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08093_ (.A1(_03233_),
    .A2(_03356_),
    .A3(_03725_),
    .ZN(_03726_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08094_ (.A1(_03116_),
    .A2(_03238_),
    .A3(_03393_),
    .Z(_03727_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08095_ (.A1(_03547_),
    .A2(_03727_),
    .B(net187),
    .ZN(_03728_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08096_ (.A1(_03294_),
    .A2(_03722_),
    .A3(_03726_),
    .A4(_03728_),
    .Z(_03729_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08097_ (.A1(_03116_),
    .A2(_03082_),
    .Z(_03730_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08098_ (.A1(_04837_),
    .A2(_03666_),
    .B(_03363_),
    .ZN(_03731_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08099_ (.A1(_03233_),
    .A2(_03107_),
    .ZN(_03732_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _08100_ (.A1(_03039_),
    .A2(_03067_),
    .A3(_03076_),
    .A4(_03392_),
    .ZN(_03733_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _08101_ (.A1(_03552_),
    .A2(_03730_),
    .B1(_03731_),
    .B2(_03732_),
    .C(_03733_),
    .ZN(_03734_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08102_ (.A1(_04882_),
    .A2(_03139_),
    .ZN(_03735_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08103_ (.A1(_04886_),
    .A2(_03184_),
    .B(_03735_),
    .ZN(_03736_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08104_ (.A1(_03183_),
    .A2(_03736_),
    .B(_03380_),
    .ZN(_03737_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08105_ (.I(_04890_),
    .ZN(_03738_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08106_ (.A1(_04907_),
    .A2(_04914_),
    .B(_04906_),
    .ZN(_03739_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08107_ (.A1(_03695_),
    .A2(_03739_),
    .B(_03716_),
    .ZN(_03740_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08108_ (.A1(_04891_),
    .A2(_03740_),
    .ZN(_03741_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08109_ (.A1(_03738_),
    .A2(_03741_),
    .ZN(_03742_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08110_ (.A1(_04891_),
    .A2(_04899_),
    .A3(_03649_),
    .A4(_03696_),
    .Z(_03743_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08111_ (.A1(_03189_),
    .A2(_03742_),
    .A3(_03743_),
    .B(_03194_),
    .ZN(_03744_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08112_ (.I(_03742_),
    .ZN(_03745_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _08113_ (.A1(_04891_),
    .A2(_04899_),
    .A3(_03649_),
    .A4(_03696_),
    .ZN(_03746_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08114_ (.A1(_03745_),
    .A2(_03746_),
    .B(_04883_),
    .C(_03189_),
    .ZN(_03747_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08115_ (.A1(_04883_),
    .A2(_03744_),
    .B(_03747_),
    .ZN(_03748_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08116_ (.A1(_03729_),
    .A2(_03734_),
    .B1(_03737_),
    .B2(_03748_),
    .ZN(net78));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08117_ (.A1(_04874_),
    .A2(_03139_),
    .ZN(_03749_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08118_ (.A1(_04878_),
    .A2(_03184_),
    .B(_03749_),
    .ZN(_03750_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08119_ (.A1(_03183_),
    .A2(_03750_),
    .B(_03294_),
    .ZN(_03751_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08120_ (.A1(_02994_),
    .A2(_03717_),
    .B(_04882_),
    .C(_02998_),
    .ZN(_03752_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08121_ (.A1(_03253_),
    .A2(_03752_),
    .Z(_03753_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08122_ (.A1(_03280_),
    .A2(_03752_),
    .B(_03028_),
    .ZN(_03754_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08123_ (.I0(_03753_),
    .I1(_03754_),
    .S(_04875_),
    .Z(_03755_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08124_ (.I0(_04872_),
    .I1(_04880_),
    .I2(_04888_),
    .I3(_04896_),
    .S0(_01115_),
    .S1(net271),
    .Z(_03756_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08125_ (.I0(_04904_),
    .I1(_04920_),
    .S(_02892_),
    .Z(_03757_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08126_ (.I0(_03723_),
    .I1(_03757_),
    .S(_03079_),
    .Z(_03758_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08127_ (.I0(_03756_),
    .I1(_03758_),
    .S(net175),
    .Z(_03759_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08128_ (.I0(_03569_),
    .I1(_03759_),
    .S(_03127_),
    .Z(_03760_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08129_ (.A1(_03269_),
    .A2(_03136_),
    .ZN(_03761_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08130_ (.A1(_03238_),
    .A2(_03760_),
    .B(_03421_),
    .C(_03761_),
    .ZN(_03762_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08131_ (.A1(_03238_),
    .A2(_03412_),
    .ZN(_03763_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08132_ (.A1(_03259_),
    .A2(_03681_),
    .ZN(_03764_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08133_ (.A1(_03731_),
    .A2(_03764_),
    .B(_03011_),
    .ZN(_03765_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08134_ (.A1(net187),
    .A2(_03763_),
    .A3(_03765_),
    .Z(_03766_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08135_ (.A1(_03751_),
    .A2(_03755_),
    .B(_03762_),
    .C(_03766_),
    .ZN(net79));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08136_ (.I0(_04864_),
    .I1(_04872_),
    .I2(_04880_),
    .I3(_04888_),
    .S0(_01115_),
    .S1(net271),
    .Z(_03767_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08137_ (.I0(_03757_),
    .I1(_03688_),
    .S(_03213_),
    .Z(_03768_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08138_ (.I0(_03767_),
    .I1(_03768_),
    .S(net175),
    .Z(_03769_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08139_ (.A1(_03233_),
    .A2(_03356_),
    .A3(_03769_),
    .Z(_03770_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _08140_ (.A1(_03233_),
    .A2(_03408_),
    .A3(_03589_),
    .B1(_03680_),
    .B2(_03431_),
    .ZN(_03771_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08141_ (.A1(_03012_),
    .A2(_03770_),
    .A3(_03771_),
    .ZN(_03772_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08142_ (.A1(_03427_),
    .A2(_03571_),
    .ZN(_03773_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08143_ (.A1(_03432_),
    .A2(_03666_),
    .B(_03731_),
    .ZN(_03774_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08144_ (.A1(_03772_),
    .A2(_03773_),
    .A3(_03774_),
    .ZN(_03775_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08145_ (.I(_02995_),
    .ZN(_03776_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _08146_ (.A1(_03776_),
    .A2(_03697_),
    .B(_02997_),
    .C(_03000_),
    .ZN(_03777_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08147_ (.A1(_03777_),
    .A2(_04867_),
    .ZN(_03778_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08148_ (.A1(_04866_),
    .A2(_03018_),
    .ZN(_03779_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08149_ (.A1(_04870_),
    .A2(_03014_),
    .B(_03779_),
    .ZN(_03780_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _08150_ (.A1(_04867_),
    .A2(_03144_),
    .B1(_03780_),
    .B2(_03013_),
    .C(_03294_),
    .ZN(_03781_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08151_ (.A1(_03778_),
    .A2(_03189_),
    .B(_03781_),
    .ZN(_03782_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08152_ (.A1(_03782_),
    .A2(_03775_),
    .Z(net80));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08153_ (.A1(_03065_),
    .A2(_03681_),
    .ZN(_03783_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08154_ (.I0(_03051_),
    .I1(_04833_),
    .S(_03783_),
    .Z(_03784_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08155_ (.A1(_03065_),
    .A2(_03051_),
    .A3(_03668_),
    .Z(_03785_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08156_ (.A1(_03417_),
    .A2(_03784_),
    .B(_03785_),
    .C(_03012_),
    .ZN(_03786_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08157_ (.A1(_03067_),
    .A2(_03456_),
    .B(_03459_),
    .C(_03269_),
    .ZN(_03787_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08158_ (.I0(_04856_),
    .I1(_04864_),
    .I2(_04872_),
    .I3(_04880_),
    .S0(_01116_),
    .S1(net271),
    .Z(_03788_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08159_ (.I0(_03624_),
    .I1(_03626_),
    .I2(_03788_),
    .I3(_03706_),
    .S0(net175),
    .S1(_03127_),
    .Z(_03789_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08160_ (.A1(net187),
    .A2(_03789_),
    .ZN(_03790_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08161_ (.A1(_03076_),
    .A2(_03787_),
    .A3(_03790_),
    .Z(_03791_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08162_ (.A1(_04858_),
    .A2(_03139_),
    .ZN(_03792_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08163_ (.A1(_04862_),
    .A2(_03184_),
    .B(_03792_),
    .ZN(_03793_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08164_ (.A1(_03025_),
    .A2(_03003_),
    .Z(_03794_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08165_ (.A1(_03003_),
    .A2(_03253_),
    .B(_03016_),
    .ZN(_03795_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08166_ (.I0(_03794_),
    .I1(_03795_),
    .S(_04859_),
    .Z(_03796_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08167_ (.A1(_03183_),
    .A2(_03793_),
    .B(_03294_),
    .C(_03796_),
    .ZN(_03797_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08168_ (.A1(_03786_),
    .A2(_03791_),
    .B(_03797_),
    .ZN(net81));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08169_ (.A1(_03076_),
    .A2(_03477_),
    .Z(_03798_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08170_ (.A1(_02699_),
    .A2(_03765_),
    .A3(_03798_),
    .Z(_03799_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08171_ (.I0(_04856_),
    .I1(_04872_),
    .S(_03102_),
    .Z(_03800_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08172_ (.I0(_04848_),
    .I1(_04864_),
    .S(_03102_),
    .Z(_03801_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08173_ (.I0(_03705_),
    .I1(_03724_),
    .I2(_03800_),
    .I3(_03801_),
    .S0(_03213_),
    .S1(_03064_),
    .Z(_03802_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08174_ (.A1(_03529_),
    .A2(_03802_),
    .ZN(_03803_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08175_ (.A1(_03480_),
    .A2(_03803_),
    .Z(_03804_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08176_ (.A1(net178),
    .A2(_03238_),
    .A3(_03637_),
    .ZN(_03805_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08177_ (.A1(_03039_),
    .A2(_03765_),
    .A3(_03804_),
    .A4(_03805_),
    .Z(_03806_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08178_ (.A1(_04851_),
    .A2(_03026_),
    .ZN(_03807_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08179_ (.I(_04851_),
    .ZN(_03808_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08180_ (.A1(_03808_),
    .A2(_03026_),
    .ZN(_03809_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08181_ (.I(_04858_),
    .ZN(_03810_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08182_ (.A1(_04883_),
    .A2(_03742_),
    .Z(_03811_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08183_ (.A1(_04882_),
    .A2(_03811_),
    .B(_04875_),
    .ZN(_03812_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08184_ (.A1(_02995_),
    .A2(_03696_),
    .ZN(_03813_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08185_ (.A1(_03648_),
    .A2(_03813_),
    .Z(_03814_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08186_ (.A1(_04866_),
    .A2(_04874_),
    .ZN(_03815_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08187_ (.A1(_03810_),
    .A2(_03812_),
    .A3(_03814_),
    .A4(_03815_),
    .Z(_03816_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08188_ (.A1(_02981_),
    .A2(_03813_),
    .Z(_03817_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _08189_ (.A1(_03599_),
    .A2(_03604_),
    .A3(_03608_),
    .A4(_03817_),
    .Z(_03818_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08190_ (.A1(_04867_),
    .A2(_04866_),
    .B(_04859_),
    .ZN(_03819_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08191_ (.A1(_03816_),
    .A2(_03818_),
    .B1(_03819_),
    .B2(_03810_),
    .ZN(_03820_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08192_ (.I0(_03807_),
    .I1(_03809_),
    .S(_03820_),
    .Z(_03821_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08193_ (.A1(_04850_),
    .A2(_03138_),
    .ZN(_03822_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08194_ (.A1(_04854_),
    .A2(_02941_),
    .B(_03822_),
    .ZN(_03823_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _08195_ (.A1(_04851_),
    .A2(_03028_),
    .B1(_03823_),
    .B2(_02937_),
    .C(_03136_),
    .ZN(_03824_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08196_ (.A1(_03821_),
    .A2(_03824_),
    .Z(_03825_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08197_ (.A1(_03799_),
    .A2(_03806_),
    .A3(_03825_),
    .ZN(net82));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08198_ (.I0(_03486_),
    .I1(_03492_),
    .S(_03160_),
    .Z(_03826_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08199_ (.A1(_03571_),
    .A2(_03826_),
    .ZN(_03827_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08200_ (.A1(_03668_),
    .A2(_03731_),
    .B(_03299_),
    .ZN(_03828_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _08201_ (.A1(_03160_),
    .A2(net175),
    .A3(_03356_),
    .A4(_03756_),
    .ZN(_03829_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08202_ (.A1(_03257_),
    .A2(_03666_),
    .Z(_03830_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08203_ (.I0(_04840_),
    .I1(_04856_),
    .S(_03101_),
    .Z(_03831_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08204_ (.I0(_03801_),
    .I1(_03831_),
    .S(_03199_),
    .Z(_03832_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _08205_ (.A1(_03731_),
    .A2(_03830_),
    .B1(_03832_),
    .B2(_03085_),
    .C(_03011_),
    .ZN(_03833_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08206_ (.A1(_03730_),
    .A2(_03672_),
    .ZN(_03834_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08207_ (.A1(_03828_),
    .A2(_03829_),
    .A3(_03833_),
    .A4(_03834_),
    .Z(_03835_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08208_ (.A1(_04842_),
    .A2(_03017_),
    .ZN(_03836_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08209_ (.A1(_04846_),
    .A2(_02941_),
    .B(_03836_),
    .ZN(_03837_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08210_ (.A1(_03031_),
    .A2(_03837_),
    .B(_03136_),
    .ZN(_03838_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08211_ (.A1(_04851_),
    .A2(_04859_),
    .A3(_03794_),
    .ZN(_03839_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08212_ (.A1(_04851_),
    .A2(_04858_),
    .A3(_03026_),
    .Z(_03840_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08213_ (.A1(_04850_),
    .A2(_03280_),
    .B(_03840_),
    .C(_04843_),
    .ZN(_03841_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08214_ (.A1(_03838_),
    .A2(_03839_),
    .A3(_03841_),
    .Z(_03842_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08215_ (.A1(_04859_),
    .A2(_03003_),
    .B(_04858_),
    .ZN(_03843_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08216_ (.I(_04850_),
    .ZN(_03844_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08217_ (.A1(_03808_),
    .A2(_03843_),
    .B(_03280_),
    .C(_03844_),
    .ZN(_03845_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08218_ (.A1(_04843_),
    .A2(_03194_),
    .A3(_03845_),
    .A4(_03838_),
    .Z(_03846_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08219_ (.A1(_03827_),
    .A2(_03835_),
    .B(_03846_),
    .C(_03842_),
    .ZN(net84));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08220_ (.A1(_04859_),
    .A2(_04866_),
    .B(_04858_),
    .ZN(_03847_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08221_ (.A1(_03808_),
    .A2(_03847_),
    .B(_03844_),
    .ZN(_03848_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08222_ (.A1(_04843_),
    .A2(_03848_),
    .B(_04842_),
    .ZN(_03849_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08223_ (.A1(_04835_),
    .A2(_03280_),
    .A3(_03849_),
    .ZN(_03850_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _08224_ (.A1(_04851_),
    .A2(_04859_),
    .A3(_04867_),
    .A4(_04843_),
    .ZN(_03851_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08225_ (.A1(_04835_),
    .A2(_03023_),
    .A3(_03851_),
    .Z(_03852_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08226_ (.I0(_03850_),
    .I1(_03852_),
    .S(_03777_),
    .Z(_03853_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08227_ (.A1(_04834_),
    .A2(_03018_),
    .ZN(_03854_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08228_ (.A1(_04838_),
    .A2(_03014_),
    .B(_03854_),
    .ZN(_03855_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08229_ (.A1(_04835_),
    .A2(_03851_),
    .Z(_03856_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08230_ (.I0(_02929_),
    .I1(_03856_),
    .S(_03849_),
    .Z(_03857_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08231_ (.A1(_02929_),
    .A2(_03194_),
    .B(_03011_),
    .ZN(_03858_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _08232_ (.A1(_03013_),
    .A2(_03855_),
    .B1(_03857_),
    .B2(_03280_),
    .C(_03858_),
    .ZN(_03859_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08233_ (.I0(_01258_),
    .I1(_04848_),
    .S(_03101_),
    .Z(_03860_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08234_ (.I0(_03831_),
    .I1(_03860_),
    .S(_03057_),
    .Z(_03861_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08235_ (.I0(_03767_),
    .I1(_03861_),
    .S(_03054_),
    .Z(_03862_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08236_ (.I0(_03690_),
    .I1(_03862_),
    .S(_03159_),
    .Z(_03863_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08237_ (.A1(_03340_),
    .A2(_03680_),
    .B(_03462_),
    .C(_03136_),
    .ZN(_03864_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _08238_ (.A1(_03516_),
    .A2(_03571_),
    .B1(_03863_),
    .B2(_03356_),
    .C(_03864_),
    .ZN(_03865_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08239_ (.A1(_03853_),
    .A2(_03859_),
    .B(_03865_),
    .ZN(net85));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_20 _08240_ (.I(net60),
    .ZN(_00000_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08241_ (.A1(_01029_),
    .A2(_02409_),
    .Z(_03866_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08242_ (.A1(_01109_),
    .A2(_03866_),
    .Z(_03867_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08243_ (.I(_03867_),
    .Z(_03868_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08244_ (.I0(net95),
    .I1(_04824_),
    .S(_03868_),
    .Z(_05078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08245_ (.I0(net106),
    .I1(net242),
    .S(_03868_),
    .Z(_04820_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08246_ (.I0(net117),
    .I1(net259),
    .S(_03868_),
    .Z(_05083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08247_ (.I0(net120),
    .I1(_05056_),
    .S(_03868_),
    .Z(_05087_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08248_ (.I0(net121),
    .I1(_05048_),
    .S(_03868_),
    .Z(_05093_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08249_ (.I0(net122),
    .I1(_05040_),
    .S(_03868_),
    .Z(_05097_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08250_ (.I0(net123),
    .I1(_05032_),
    .S(_03868_),
    .Z(_05101_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08251_ (.I0(net124),
    .I1(_05024_),
    .S(_03868_),
    .Z(_05105_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08252_ (.I0(net125),
    .I1(net172),
    .S(_03868_),
    .Z(_05109_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08253_ (.I0(net126),
    .I1(net185),
    .S(_03868_),
    .Z(_05113_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _08254_ (.I(_03867_),
    .Z(_03869_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08255_ (.I0(net96),
    .I1(_05000_),
    .S(_03869_),
    .Z(_05117_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08256_ (.I0(net97),
    .I1(_04992_),
    .S(_03869_),
    .Z(_05121_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08257_ (.I0(net98),
    .I1(_04984_),
    .S(_03869_),
    .Z(_05125_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08258_ (.I0(net99),
    .I1(_04976_),
    .S(_03869_),
    .Z(_05129_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08259_ (.I0(net100),
    .I1(_04968_),
    .S(_03869_),
    .Z(_05133_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08260_ (.I0(net101),
    .I1(_04960_),
    .S(_03869_),
    .Z(_05137_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08261_ (.I0(net102),
    .I1(net263),
    .S(_03869_),
    .Z(_05141_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08262_ (.I0(net103),
    .I1(_04944_),
    .S(_03869_),
    .Z(_05145_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08263_ (.I0(net104),
    .I1(_04936_),
    .S(_03869_),
    .Z(_05149_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08264_ (.I0(net105),
    .I1(_04928_),
    .S(_03869_),
    .Z(_05153_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _08265_ (.I(_03867_),
    .Z(_03870_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08266_ (.I0(net107),
    .I1(_04920_),
    .S(_03870_),
    .Z(_05157_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08267_ (.I0(net108),
    .I1(_04912_),
    .S(_03870_),
    .Z(_05161_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08268_ (.I0(net109),
    .I1(_04904_),
    .S(_03870_),
    .Z(_05165_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08269_ (.I0(net110),
    .I1(_04896_),
    .S(_03870_),
    .Z(_05169_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08270_ (.I0(net111),
    .I1(_04888_),
    .S(_03870_),
    .Z(_05173_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08271_ (.I0(net112),
    .I1(_04880_),
    .S(_03870_),
    .Z(_05177_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08272_ (.I0(net113),
    .I1(_04872_),
    .S(_03870_),
    .Z(_05181_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08273_ (.I0(net114),
    .I1(_04864_),
    .S(_03870_),
    .Z(_05185_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08274_ (.I0(net115),
    .I1(_04856_),
    .S(_03870_),
    .Z(_05189_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08275_ (.I0(net116),
    .I1(_04848_),
    .S(_03870_),
    .Z(_05193_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08276_ (.I0(net118),
    .I1(_04840_),
    .S(_03867_),
    .Z(_05197_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08277_ (.I(_01110_),
    .ZN(_05079_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08278_ (.I(_01922_),
    .ZN(_05158_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08279_ (.A1(_01090_),
    .A2(_02675_),
    .Z(_03871_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _08280_ (.I(_03871_),
    .Z(_03872_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08281_ (.A1(_02243_),
    .A2(_04968_),
    .Z(_03873_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08282_ (.A1(_02336_),
    .A2(_04984_),
    .ZN(_03874_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08283_ (.A1(_02244_),
    .A2(_02258_),
    .A3(_02274_),
    .Z(_03875_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _08284_ (.I(_02289_),
    .ZN(_03876_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08285_ (.A1(_04980_),
    .A2(_03874_),
    .B(_03875_),
    .C(_03876_),
    .ZN(_03877_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08286_ (.A1(_04980_),
    .A2(_03875_),
    .A3(_03874_),
    .ZN(_03878_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08287_ (.A1(_03873_),
    .A2(_03877_),
    .A3(_03878_),
    .Z(_03879_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _08288_ (.A1(_02289_),
    .A2(_04976_),
    .B1(_02336_),
    .B2(_04984_),
    .ZN(_03880_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _08289_ (.A1(_02244_),
    .A2(_04972_),
    .B1(_03876_),
    .B2(_04980_),
    .C(_03880_),
    .ZN(_03881_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08290_ (.A1(_02476_),
    .A2(net183),
    .ZN(_03882_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08291_ (.A1(_02515_),
    .A2(net171),
    .B(_02476_),
    .ZN(_03883_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08292_ (.A1(_02515_),
    .A2(net170),
    .B(net182),
    .ZN(_03884_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _08293_ (.A1(_03882_),
    .A2(_03883_),
    .A3(_03884_),
    .B1(_05004_),
    .B2(_02427_),
    .ZN(_03885_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08294_ (.A1(_02427_),
    .A2(_05004_),
    .ZN(_03886_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08295_ (.A1(_02375_),
    .A2(_04996_),
    .B(_03875_),
    .ZN(_03887_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08296_ (.A1(_03881_),
    .A2(_03885_),
    .A3(_03886_),
    .A4(_03887_),
    .Z(_03888_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08297_ (.A1(_02244_),
    .A2(_04972_),
    .ZN(_03889_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08298_ (.A1(_02375_),
    .A2(_02408_),
    .ZN(_03890_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08299_ (.A1(_03889_),
    .A2(_03881_),
    .A3(_03890_),
    .Z(_03891_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _08300_ (.A1(_04960_),
    .A2(_03879_),
    .A3(_03888_),
    .A4(_03891_),
    .Z(_03892_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08301_ (.A1(_02604_),
    .A2(_05032_),
    .ZN(_03893_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08302_ (.A1(_05028_),
    .A2(_03893_),
    .ZN(_03894_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08303_ (.A1(_05028_),
    .A2(_03893_),
    .B(net157),
    .ZN(_03895_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08304_ (.A1(_02903_),
    .A2(_02910_),
    .ZN(_03896_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08305_ (.A1(_01416_),
    .A2(_02912_),
    .Z(_03897_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08306_ (.A1(_01576_),
    .A2(_02917_),
    .B(_03897_),
    .ZN(_03898_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08307_ (.A1(_01697_),
    .A2(_02920_),
    .A3(_02922_),
    .Z(_03899_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08308_ (.I(\dp.rf.rf[20][1] ),
    .ZN(_03900_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08309_ (.A1(_01328_),
    .A2(_02925_),
    .ZN(_03901_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08310_ (.A1(_03900_),
    .A2(_01327_),
    .B(_03901_),
    .C(_01529_),
    .ZN(_03902_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _08311_ (.A1(\dp.rf.rf[16][1] ),
    .A2(_01356_),
    .B1(_03902_),
    .B2(_01541_),
    .C(_01206_),
    .ZN(_03903_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _08312_ (.A1(_01385_),
    .A2(_03898_),
    .B1(_03899_),
    .B2(_03903_),
    .ZN(_03904_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08313_ (.A1(_02868_),
    .A2(_02870_),
    .A3(_02872_),
    .A4(_02874_),
    .Z(_03905_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08314_ (.A1(_01778_),
    .A2(_02887_),
    .B1(_03905_),
    .B2(_01780_),
    .ZN(_03906_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _08315_ (.A1(_03896_),
    .A2(_03904_),
    .B(_02884_),
    .C(_03906_),
    .ZN(_03907_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08316_ (.A1(_02811_),
    .A2(net260),
    .B(_01062_),
    .C(net169),
    .ZN(_03908_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08317_ (.A1(_02903_),
    .A2(_02910_),
    .B(net139),
    .ZN(_03909_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08318_ (.A1(_02811_),
    .A2(net260),
    .B(_03904_),
    .C(_03909_),
    .ZN(_03910_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08319_ (.A1(_02811_),
    .A2(_05064_),
    .ZN(_03911_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08320_ (.A1(_03907_),
    .A2(_03908_),
    .B(_03910_),
    .C(_03911_),
    .ZN(_03912_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08321_ (.A1(_02696_),
    .A2(_05048_),
    .B(_05040_),
    .ZN(_03913_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08322_ (.A1(_05040_),
    .A2(_02696_),
    .A3(_05048_),
    .ZN(_03914_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08323_ (.A1(net155),
    .A2(_03913_),
    .B(_03914_),
    .C(_05060_),
    .ZN(_03915_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08324_ (.I(net155),
    .ZN(_03916_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08325_ (.A1(_03916_),
    .A2(_05040_),
    .B(_02696_),
    .C(_05048_),
    .ZN(_03917_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08326_ (.A1(net155),
    .A2(_05044_),
    .B(_03917_),
    .ZN(_03918_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _08327_ (.A1(_03894_),
    .A2(_03895_),
    .B1(_03912_),
    .B2(_03915_),
    .C(_03918_),
    .ZN(_03919_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08328_ (.A1(_05040_),
    .A2(_02696_),
    .A3(_05048_),
    .Z(_03920_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08329_ (.A1(net155),
    .A2(_03913_),
    .ZN(_03921_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08330_ (.A1(net153),
    .A2(_05060_),
    .ZN(_03922_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08331_ (.A1(net155),
    .A2(_03913_),
    .B(_03914_),
    .C(net153),
    .ZN(_03923_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _08332_ (.A1(_03920_),
    .A2(_03921_),
    .A3(_03922_),
    .B1(_03923_),
    .B2(_03912_),
    .ZN(_03924_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08333_ (.A1(_02604_),
    .A2(_05032_),
    .ZN(_03925_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08334_ (.A1(_05028_),
    .A2(_03925_),
    .ZN(_03926_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08335_ (.A1(_05028_),
    .A2(_03925_),
    .B(net157),
    .ZN(_03927_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08336_ (.A1(_03926_),
    .A2(_03927_),
    .ZN(_03928_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08337_ (.A1(_03919_),
    .A2(_03924_),
    .B(_03928_),
    .ZN(_03929_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08338_ (.A1(_04960_),
    .A2(_03890_),
    .ZN(_03930_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08339_ (.A1(_02187_),
    .A2(_03890_),
    .ZN(_03931_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08340_ (.A1(_03873_),
    .A2(_03877_),
    .A3(_03878_),
    .ZN(_03932_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08341_ (.A1(_02476_),
    .A2(net181),
    .B(_02515_),
    .C(net170),
    .ZN(_03933_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08342_ (.A1(_05004_),
    .A2(_03882_),
    .A3(_03933_),
    .ZN(_03934_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08343_ (.A1(_02375_),
    .A2(_04996_),
    .ZN(_03935_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08344_ (.A1(_02375_),
    .A2(_04996_),
    .B(_02427_),
    .ZN(_03936_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08345_ (.A1(_03882_),
    .A2(_03933_),
    .B(_02459_),
    .ZN(_03937_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08346_ (.A1(_03934_),
    .A2(_03935_),
    .B1(_03936_),
    .B2(_03937_),
    .ZN(_03938_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08347_ (.A1(_03930_),
    .A2(_03931_),
    .B(_03932_),
    .C(_03938_),
    .ZN(_03939_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08348_ (.I(_02187_),
    .ZN(_03940_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08349_ (.A1(_03940_),
    .A2(_04964_),
    .Z(_03941_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08350_ (.A1(_02187_),
    .A2(_04960_),
    .B1(_03889_),
    .B2(_03881_),
    .ZN(_03942_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08351_ (.A1(_03941_),
    .A2(_03942_),
    .ZN(_03943_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08352_ (.A1(_03892_),
    .A2(_03929_),
    .B(_03939_),
    .C(_03943_),
    .ZN(_03944_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08353_ (.A1(_03919_),
    .A2(_03924_),
    .Z(_03945_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08354_ (.A1(_03879_),
    .A2(_03888_),
    .A3(_03891_),
    .B(_04960_),
    .ZN(_03946_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08355_ (.A1(_03940_),
    .A2(_03928_),
    .Z(_03947_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08356_ (.A1(_03945_),
    .A2(_03946_),
    .A3(_03947_),
    .Z(_03948_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08357_ (.I(_02095_),
    .ZN(_03949_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08358_ (.A1(_02139_),
    .A2(net263),
    .ZN(_03950_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08359_ (.A1(_03949_),
    .A2(_04948_),
    .B(_03950_),
    .ZN(_03951_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _08360_ (.I(_02050_),
    .ZN(_03952_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08361_ (.A1(_03952_),
    .A2(_04940_),
    .B1(_03949_),
    .B2(_04948_),
    .ZN(_03953_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _08362_ (.A1(_01989_),
    .A2(_04928_),
    .B1(_02050_),
    .B2(_04936_),
    .C1(_03951_),
    .C2(_03953_),
    .ZN(_03954_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08363_ (.A1(_01785_),
    .A2(_01817_),
    .Z(_03955_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08364_ (.A1(_01841_),
    .A2(_01871_),
    .ZN(_03956_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08365_ (.A1(_01886_),
    .A2(_01918_),
    .ZN(_03957_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08366_ (.A1(_01886_),
    .A2(_01918_),
    .B(_01938_),
    .C(_01974_),
    .ZN(_03958_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08367_ (.A1(_01841_),
    .A2(_01871_),
    .ZN(_03959_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08368_ (.A1(_03956_),
    .A2(_03957_),
    .A3(_03958_),
    .B(_03959_),
    .ZN(_03960_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08369_ (.A1(_01990_),
    .A2(_04932_),
    .ZN(_03961_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08370_ (.A1(_03955_),
    .A2(_03960_),
    .A3(_03961_),
    .ZN(_03962_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_4 _08371_ (.A1(_01841_),
    .A2(_01871_),
    .B1(_01886_),
    .B2(_01918_),
    .C1(_01938_),
    .C2(_04920_),
    .ZN(_03963_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08372_ (.A1(_01841_),
    .A2(_04904_),
    .B(_01886_),
    .C(_04912_),
    .ZN(_03964_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _08373_ (.A1(_03956_),
    .A2(_03963_),
    .A3(_03964_),
    .ZN(_03965_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08374_ (.A1(_01785_),
    .A2(_04896_),
    .Z(_03966_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08375_ (.A1(_03955_),
    .A2(_03965_),
    .B(_03966_),
    .ZN(_03967_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08376_ (.A1(_03954_),
    .A2(_03962_),
    .B(_03967_),
    .ZN(_03968_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _08377_ (.A1(_01565_),
    .A2(_01590_),
    .A3(_01604_),
    .ZN(_03969_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08378_ (.A1(_01590_),
    .A2(_01604_),
    .B(_01565_),
    .ZN(_03970_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08379_ (.A1(_01622_),
    .A2(_04876_),
    .A3(_03969_),
    .B(_03970_),
    .ZN(_03971_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _08380_ (.A1(_01739_),
    .A2(_01743_),
    .B1(_01753_),
    .B2(_01760_),
    .C(_01726_),
    .ZN(_03972_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08381_ (.A1(_01696_),
    .A2(_01710_),
    .B(_03972_),
    .ZN(_03973_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08382_ (.A1(_01696_),
    .A2(_01710_),
    .A3(_03972_),
    .B(_01683_),
    .ZN(_03974_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _08383_ (.A1(_01622_),
    .A2(_04876_),
    .B1(_03973_),
    .B2(_03974_),
    .C(_03969_),
    .ZN(_03975_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08384_ (.A1(_03971_),
    .A2(_03975_),
    .ZN(_03976_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08385_ (.A1(_01257_),
    .A2(_01284_),
    .ZN(_03977_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08386_ (.A1(_01257_),
    .A2(_01284_),
    .Z(_03978_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _08387_ (.A1(_03977_),
    .A2(_03978_),
    .ZN(_03979_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08388_ (.A1(_01321_),
    .A2(_04840_),
    .Z(_03980_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08389_ (.A1(_01412_),
    .A2(_01469_),
    .ZN(_03981_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _08390_ (.A1(_01412_),
    .A2(_01469_),
    .B(_01489_),
    .C(_01544_),
    .ZN(_03982_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08391_ (.A1(_03981_),
    .A2(_03982_),
    .ZN(_03983_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08392_ (.A1(net5),
    .A2(_02362_),
    .Z(_03984_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08393_ (.I0(_03977_),
    .I1(_03978_),
    .S(_03984_),
    .Z(_03985_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08394_ (.A1(_03979_),
    .A2(_03980_),
    .B(_03983_),
    .C(_03985_),
    .ZN(_03986_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08395_ (.A1(_03976_),
    .A2(_03986_),
    .ZN(_03987_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _08396_ (.I(_03979_),
    .ZN(_03988_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08397_ (.A1(_04844_),
    .A2(_03981_),
    .A3(_03982_),
    .ZN(_03989_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08398_ (.A1(_03981_),
    .A2(_03982_),
    .B(_04844_),
    .ZN(_03990_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08399_ (.A1(_01321_),
    .A2(_03989_),
    .B(_03990_),
    .ZN(_03991_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08400_ (.A1(_04876_),
    .A2(_03969_),
    .ZN(_03992_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08401_ (.A1(_01683_),
    .A2(_01696_),
    .A3(_01710_),
    .ZN(_03993_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08402_ (.A1(_01714_),
    .A2(_01718_),
    .Z(_03994_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08403_ (.A1(_03994_),
    .A2(_01725_),
    .Z(_03995_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08404_ (.A1(_03995_),
    .A2(_04888_),
    .B(_01696_),
    .C(_01710_),
    .ZN(_03996_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08405_ (.A1(_03995_),
    .A2(_04888_),
    .B(_01683_),
    .ZN(_03997_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08406_ (.A1(_03993_),
    .A2(_03996_),
    .A3(_03997_),
    .ZN(_03998_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08407_ (.A1(_01565_),
    .A2(_01590_),
    .A3(_01604_),
    .B(_01621_),
    .ZN(_03999_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _08408_ (.A1(_03993_),
    .A2(_03999_),
    .A3(_03996_),
    .A4(_03997_),
    .ZN(_04000_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08409_ (.A1(_03992_),
    .A2(_03998_),
    .B(_04000_),
    .C(_03971_),
    .ZN(_04001_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08410_ (.I(_03985_),
    .ZN(_04002_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _08411_ (.A1(_03988_),
    .A2(_03991_),
    .B(_04001_),
    .C(_04002_),
    .ZN(_04003_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08412_ (.A1(_03968_),
    .A2(_03987_),
    .B(_04003_),
    .ZN(_04004_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08413_ (.A1(_02170_),
    .A2(_01067_),
    .Z(_04005_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08414_ (.A1(_03944_),
    .A2(_03948_),
    .B(_04004_),
    .C(_04005_),
    .ZN(_04006_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08415_ (.A1(_02139_),
    .A2(net263),
    .ZN(_04007_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08416_ (.A1(_03952_),
    .A2(_04940_),
    .B(_04948_),
    .C(_04007_),
    .ZN(_04008_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _08417_ (.A1(_02108_),
    .A2(_02121_),
    .B1(_02139_),
    .B2(_02168_),
    .ZN(_04009_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08418_ (.A1(_04940_),
    .A2(_03949_),
    .A3(_04009_),
    .ZN(_04010_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08419_ (.A1(_03952_),
    .A2(_03949_),
    .A3(_04009_),
    .ZN(_04011_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08420_ (.A1(_01990_),
    .A2(_04932_),
    .B1(_03952_),
    .B2(_04940_),
    .ZN(_04012_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _08421_ (.A1(_04008_),
    .A2(_04010_),
    .A3(_04011_),
    .A4(_04012_),
    .ZN(_04013_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08422_ (.A1(_01989_),
    .A2(_04928_),
    .B(_03966_),
    .C(_03965_),
    .ZN(_04014_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08423_ (.A1(_03955_),
    .A2(_03960_),
    .B(_03966_),
    .ZN(_04015_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08424_ (.A1(_04013_),
    .A2(_04014_),
    .B(_04015_),
    .ZN(_04016_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08425_ (.A1(_03988_),
    .A2(_03991_),
    .B(_03976_),
    .C(_04002_),
    .ZN(_04017_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08426_ (.A1(_03979_),
    .A2(_03980_),
    .B(_03985_),
    .ZN(_04018_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08427_ (.A1(_01412_),
    .A2(_01469_),
    .B(_01489_),
    .C(_04856_),
    .ZN(_04019_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08428_ (.A1(_01412_),
    .A2(_04848_),
    .ZN(_04020_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08429_ (.A1(_04019_),
    .A2(_04020_),
    .ZN(_04021_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08430_ (.A1(_01321_),
    .A2(_04840_),
    .B(_03979_),
    .C(_04021_),
    .ZN(_04022_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08431_ (.A1(_04018_),
    .A2(_04022_),
    .ZN(_04023_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _08432_ (.A1(_04003_),
    .A2(_04016_),
    .B(_04017_),
    .C(_04023_),
    .ZN(_04024_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _08433_ (.A1(_02931_),
    .A2(_04024_),
    .A3(_03944_),
    .A4(_03948_),
    .Z(_04025_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08434_ (.A1(_02931_),
    .A2(_04024_),
    .A3(_04004_),
    .Z(_04026_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08435_ (.A1(_04024_),
    .A2(_04005_),
    .ZN(_04027_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08436_ (.A1(_04006_),
    .A2(_04025_),
    .A3(_04026_),
    .A4(_04027_),
    .Z(_04028_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08437_ (.A1(_03009_),
    .A2(_03015_),
    .Z(_04029_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08438_ (.I(_04029_),
    .ZN(_04030_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08439_ (.A1(_03009_),
    .A2(_03008_),
    .ZN(_04031_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _08440_ (.A1(_04960_),
    .A2(_03879_),
    .A3(_03888_),
    .A4(_03891_),
    .ZN(_04032_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08441_ (.A1(_03928_),
    .A2(_04032_),
    .B1(_03946_),
    .B2(_03947_),
    .ZN(_04033_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08442_ (.A1(_01321_),
    .A2(_04840_),
    .B(_03988_),
    .C(_03983_),
    .ZN(_04034_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08443_ (.I0(_03978_),
    .I1(_03977_),
    .S(_03984_),
    .Z(_04035_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08444_ (.I(_01321_),
    .ZN(_04036_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08445_ (.A1(_04036_),
    .A2(_04844_),
    .A3(_03979_),
    .Z(_04037_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08446_ (.A1(_04035_),
    .A2(_04037_),
    .Z(_04038_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08447_ (.A1(_02095_),
    .A2(_04944_),
    .B1(_02139_),
    .B2(_02168_),
    .ZN(_04039_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _08448_ (.A1(_02050_),
    .A2(_04936_),
    .B1(_02095_),
    .B2(_02122_),
    .ZN(_04040_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_4 _08449_ (.A1(_01990_),
    .A2(_04932_),
    .B1(_03952_),
    .B2(_04940_),
    .C1(_04039_),
    .C2(_04040_),
    .ZN(_04041_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08450_ (.A1(_03955_),
    .A2(_03960_),
    .A3(_03961_),
    .Z(_04042_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _08451_ (.A1(_03955_),
    .A2(_03965_),
    .B1(_04041_),
    .B2(_04042_),
    .C(_03966_),
    .ZN(_04043_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08452_ (.A1(_03976_),
    .A2(_03986_),
    .Z(_04044_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _08453_ (.A1(_04034_),
    .A2(_04038_),
    .B1(_04043_),
    .B2(_04044_),
    .C(_04001_),
    .ZN(_04045_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08454_ (.A1(_03889_),
    .A2(_03881_),
    .ZN(_04046_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08455_ (.I(_03890_),
    .ZN(_04047_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08456_ (.A1(_03932_),
    .A2(_03938_),
    .A3(_04047_),
    .Z(_04048_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08457_ (.I(net153),
    .ZN(_04049_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08458_ (.A1(_03904_),
    .A2(_03909_),
    .B(_01062_),
    .C(net169),
    .ZN(_04050_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08459_ (.A1(_03907_),
    .A2(_04050_),
    .B(_03911_),
    .ZN(_04051_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _08460_ (.A1(_04049_),
    .A2(net220),
    .B1(net193),
    .B2(_05064_),
    .C(_04051_),
    .ZN(_04052_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08461_ (.A1(_03918_),
    .A2(_03922_),
    .ZN(_04053_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08462_ (.A1(_03941_),
    .A2(_03921_),
    .ZN(_04054_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08463_ (.A1(_04052_),
    .A2(_04053_),
    .B(_04054_),
    .C(_03914_),
    .ZN(_04055_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _08464_ (.A1(_04046_),
    .A2(_04048_),
    .A3(_03945_),
    .A4(_04055_),
    .Z(_04056_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _08465_ (.A1(_04024_),
    .A2(_04033_),
    .A3(_04045_),
    .A4(_04056_),
    .Z(_04057_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08466_ (.I0(_04030_),
    .I1(_04031_),
    .S(_04057_),
    .Z(_04058_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08467_ (.A1(_04028_),
    .A2(_04058_),
    .B(_01083_),
    .ZN(_04059_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08468_ (.A1(_03872_),
    .A2(_04059_),
    .Z(_04060_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _08469_ (.I(_04060_),
    .Z(_04061_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08470_ (.I0(net95),
    .I1(_05080_),
    .S(_04061_),
    .Z(_00001_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08471_ (.I(_04823_),
    .ZN(_04062_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08472_ (.I0(net106),
    .I1(_04062_),
    .S(_04061_),
    .Z(_00002_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08473_ (.I(\dp.rf.rf[0][0] ),
    .Z(_00003_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08474_ (.I(\dp.rf.rf[0][10] ),
    .Z(_00004_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08475_ (.I(\dp.rf.rf[0][11] ),
    .Z(_00005_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08476_ (.I(\dp.rf.rf[0][12] ),
    .Z(_00006_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08477_ (.I(\dp.rf.rf[0][13] ),
    .Z(_00007_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08478_ (.I(\dp.rf.rf[0][14] ),
    .Z(_00008_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08479_ (.I(\dp.rf.rf[0][15] ),
    .Z(_00009_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08480_ (.I(\dp.rf.rf[0][16] ),
    .Z(_00010_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08481_ (.I(\dp.rf.rf[0][17] ),
    .Z(_00011_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08482_ (.I(\dp.rf.rf[0][18] ),
    .Z(_00012_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08483_ (.I(\dp.rf.rf[0][19] ),
    .Z(_00013_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08484_ (.I(\dp.rf.rf[0][1] ),
    .Z(_00014_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08485_ (.I(\dp.rf.rf[0][20] ),
    .Z(_00015_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08486_ (.I(\dp.rf.rf[0][21] ),
    .Z(_00016_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08487_ (.I(\dp.rf.rf[0][22] ),
    .Z(_00017_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08488_ (.I(\dp.rf.rf[0][23] ),
    .Z(_00018_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08489_ (.I(\dp.rf.rf[0][24] ),
    .Z(_00019_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08490_ (.I(\dp.rf.rf[0][25] ),
    .Z(_00020_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08491_ (.I(\dp.rf.rf[0][26] ),
    .Z(_00021_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08492_ (.I(\dp.rf.rf[0][27] ),
    .Z(_00022_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08493_ (.I(\dp.rf.rf[0][28] ),
    .Z(_00023_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08494_ (.I(\dp.rf.rf[0][29] ),
    .Z(_00024_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08495_ (.I(\dp.rf.rf[0][2] ),
    .Z(_00025_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08496_ (.I(\dp.rf.rf[0][30] ),
    .Z(_00026_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08497_ (.I(\dp.rf.rf[0][31] ),
    .Z(_00027_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08498_ (.I(\dp.rf.rf[0][3] ),
    .Z(_00028_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08499_ (.I(\dp.rf.rf[0][4] ),
    .Z(_00029_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08500_ (.I(\dp.rf.rf[0][5] ),
    .Z(_00030_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08501_ (.I(\dp.rf.rf[0][6] ),
    .Z(_00031_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08502_ (.I(\dp.rf.rf[0][7] ),
    .Z(_00032_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08503_ (.I(\dp.rf.rf[0][8] ),
    .Z(_00033_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _08504_ (.I(\dp.rf.rf[0][9] ),
    .Z(_00034_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _08505_ (.I(_03866_),
    .Z(_04063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08506_ (.A1(_01090_),
    .A2(_02675_),
    .ZN(_04064_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _08507_ (.A1(_05080_),
    .A2(_04063_),
    .B1(_04064_),
    .B2(net95),
    .ZN(_04065_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08508_ (.A1(_03866_),
    .A2(_04064_),
    .Z(_04066_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _08509_ (.I(_04066_),
    .Z(_04067_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _08510_ (.I(_03089_),
    .Z(_04068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08511_ (.A1(net28),
    .A2(_04068_),
    .ZN(_04069_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08512_ (.A1(_03089_),
    .A2(_04065_),
    .ZN(_04070_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08513_ (.A1(net61),
    .A2(_04070_),
    .ZN(_04071_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _08514_ (.A1(_04065_),
    .A2(_04067_),
    .B(_04069_),
    .C(_04071_),
    .ZN(_04072_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _08515_ (.I(_04072_),
    .Z(_04073_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08516_ (.A1(_02672_),
    .A2(_02793_),
    .Z(_04074_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08517_ (.A1(net2),
    .A2(_04074_),
    .Z(_04075_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08518_ (.I(net25),
    .ZN(_04076_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08519_ (.A1(_01090_),
    .A2(_01029_),
    .B(_01438_),
    .ZN(_04077_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08520_ (.A1(_01090_),
    .A2(_01082_),
    .B1(_04077_),
    .B2(_01096_),
    .ZN(_04078_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _08521_ (.A1(_01063_),
    .A2(_04078_),
    .ZN(_04079_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08522_ (.A1(_04076_),
    .A2(_04079_),
    .Z(_04080_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08523_ (.A1(net26),
    .A2(_04080_),
    .Z(_04081_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08524_ (.A1(_04075_),
    .A2(_04081_),
    .Z(_04082_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _08525_ (.I(_04082_),
    .Z(_04083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08526_ (.I0(\dp.rf.rf[10][0] ),
    .I1(_04073_),
    .S(_04083_),
    .Z(_00035_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08527_ (.I(net29),
    .ZN(_04084_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08528_ (.A1(_03015_),
    .A2(_03088_),
    .Z(_04085_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _08529_ (.I(_04085_),
    .Z(_04086_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08530_ (.I(_04086_),
    .Z(_04087_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08531_ (.A1(net57),
    .A2(_04029_),
    .ZN(_04088_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08532_ (.A1(_03088_),
    .A2(_04088_),
    .Z(_04089_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08533_ (.I(_04089_),
    .Z(_04090_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08534_ (.I(_04090_),
    .Z(_04091_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08535_ (.A1(_04084_),
    .A2(_04087_),
    .B(_04091_),
    .ZN(_04092_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08536_ (.A1(net93),
    .A2(net62),
    .B(_04067_),
    .C(_04092_),
    .ZN(_04093_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _08537_ (.A1(_01029_),
    .A2(_02409_),
    .ZN(_04094_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _08538_ (.I(_04094_),
    .Z(_04095_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08539_ (.A1(_05108_),
    .A2(_05103_),
    .Z(_04096_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08540_ (.A1(_05107_),
    .A2(_04096_),
    .Z(_04097_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08541_ (.I(_05100_),
    .ZN(_04098_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08542_ (.I(_05090_),
    .ZN(_04099_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08543_ (.A1(_04822_),
    .A2(_05086_),
    .B(_05085_),
    .ZN(_04100_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08544_ (.I(_05089_),
    .ZN(_04101_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08545_ (.A1(_04099_),
    .A2(_04100_),
    .B(_04101_),
    .ZN(_04102_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08546_ (.A1(_05096_),
    .A2(_04102_),
    .B(_05095_),
    .ZN(_04103_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08547_ (.I(_05099_),
    .ZN(_04104_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08548_ (.A1(_04098_),
    .A2(_04103_),
    .B(_04104_),
    .ZN(_04105_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08549_ (.A1(_05108_),
    .A2(_05112_),
    .Z(_04106_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08550_ (.A1(_05104_),
    .A2(_04106_),
    .Z(_04107_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _08551_ (.A1(_05112_),
    .A2(_04097_),
    .B1(_04105_),
    .B2(_04107_),
    .C(_05111_),
    .ZN(_04108_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08552_ (.I(_04108_),
    .ZN(_04109_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08553_ (.A1(_05116_),
    .A2(_04109_),
    .Z(_04110_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08554_ (.A1(_05115_),
    .A2(_04110_),
    .Z(_04111_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08555_ (.A1(_05120_),
    .A2(_04111_),
    .Z(_04112_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08556_ (.A1(net121),
    .A2(_05091_),
    .A3(net122),
    .Z(_04113_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08557_ (.A1(net123),
    .A2(net124),
    .A3(net125),
    .A4(net126),
    .Z(_04114_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08558_ (.A1(_04113_),
    .A2(_04114_),
    .Z(_04115_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08559_ (.I(_04115_),
    .Z(_04116_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08560_ (.A1(net96),
    .A2(_04116_),
    .Z(_04117_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08561_ (.A1(_04095_),
    .A2(_04112_),
    .B1(_04117_),
    .B2(_03872_),
    .ZN(_04118_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08562_ (.A1(_04093_),
    .A2(_04118_),
    .ZN(_04119_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _08563_ (.I(_04119_),
    .Z(_04120_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08564_ (.I0(\dp.rf.rf[10][10] ),
    .I1(_04120_),
    .S(_04083_),
    .Z(_00036_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08565_ (.A1(_03088_),
    .A2(_04088_),
    .ZN(_04121_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08566_ (.A1(net30),
    .A2(_01069_),
    .Z(_04122_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _08567_ (.I(_04066_),
    .Z(_04123_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _08568_ (.A1(_04068_),
    .A2(net63),
    .B1(_04121_),
    .B2(_04122_),
    .C(_04123_),
    .ZN(_04124_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08569_ (.I(_05096_),
    .ZN(_04125_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08570_ (.I(_05086_),
    .ZN(_04126_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08571_ (.A1(_04819_),
    .A2(_05082_),
    .B(_05081_),
    .ZN(_04127_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08572_ (.I(_05085_),
    .ZN(_04128_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08573_ (.A1(_04126_),
    .A2(_04127_),
    .B(_04128_),
    .ZN(_04129_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08574_ (.A1(_05090_),
    .A2(_04129_),
    .B(_05089_),
    .ZN(_04130_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08575_ (.I(_05095_),
    .ZN(_04131_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08576_ (.A1(_04125_),
    .A2(_04130_),
    .B(_04131_),
    .ZN(_04132_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08577_ (.A1(_05100_),
    .A2(_04132_),
    .B(_05099_),
    .ZN(_04133_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08578_ (.A1(_05104_),
    .A2(_05116_),
    .A3(_04106_),
    .ZN(_04134_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08579_ (.A1(_05112_),
    .A2(_05107_),
    .Z(_04135_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08580_ (.A1(_05111_),
    .A2(_04135_),
    .Z(_04136_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08581_ (.A1(_05116_),
    .A2(_05103_),
    .Z(_04137_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08582_ (.A1(_05116_),
    .A2(_04136_),
    .B1(_04137_),
    .B2(_04106_),
    .ZN(_04138_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08583_ (.A1(_04133_),
    .A2(_04134_),
    .B(_04138_),
    .ZN(_04139_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08584_ (.A1(_05115_),
    .A2(_04139_),
    .Z(_04140_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08585_ (.A1(_05120_),
    .A2(_04140_),
    .B(_05119_),
    .ZN(_04141_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08586_ (.A1(_05124_),
    .A2(_04141_),
    .ZN(_04142_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08587_ (.A1(net117),
    .A2(net120),
    .A3(net121),
    .A4(net122),
    .Z(_04143_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08588_ (.A1(_04114_),
    .A2(_04143_),
    .Z(_04144_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08589_ (.I(_04144_),
    .Z(_04145_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08590_ (.A1(net96),
    .A2(_04145_),
    .ZN(_04146_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08591_ (.A1(net97),
    .A2(_04146_),
    .ZN(_04147_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08592_ (.A1(_04095_),
    .A2(_04142_),
    .B1(_04147_),
    .B2(_03872_),
    .ZN(_04148_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08593_ (.A1(_04124_),
    .A2(_04148_),
    .ZN(_04149_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _08594_ (.I(_04149_),
    .Z(_04150_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08595_ (.I0(\dp.rf.rf[10][11] ),
    .I1(_04150_),
    .S(_04083_),
    .Z(_00037_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08596_ (.A1(_04063_),
    .A2(_04064_),
    .ZN(_04151_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08597_ (.A1(_03089_),
    .A2(_03453_),
    .A3(_03465_),
    .ZN(_04152_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08598_ (.A1(net31),
    .A2(_01069_),
    .B(_04121_),
    .ZN(_04153_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _08599_ (.I(_04094_),
    .Z(_04154_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08600_ (.A1(_05120_),
    .A2(_04111_),
    .Z(_04155_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08601_ (.A1(_05119_),
    .A2(_04155_),
    .Z(_04156_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08602_ (.A1(_05124_),
    .A2(_04156_),
    .B(_05123_),
    .ZN(_04157_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08603_ (.A1(_05128_),
    .A2(_04157_),
    .ZN(_04158_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08604_ (.A1(net96),
    .A2(net97),
    .A3(_04115_),
    .Z(_04159_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08605_ (.A1(net98),
    .A2(_04159_),
    .Z(_04160_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _08606_ (.I(_03871_),
    .Z(_04161_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08607_ (.A1(_04154_),
    .A2(_04158_),
    .B1(_04160_),
    .B2(_04161_),
    .ZN(_04162_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _08608_ (.A1(_04151_),
    .A2(_04152_),
    .A3(_04153_),
    .B(_04162_),
    .ZN(_04163_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _08609_ (.I(_04163_),
    .Z(_04164_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08610_ (.I0(\dp.rf.rf[10][12] ),
    .I1(_04164_),
    .S(_04083_),
    .Z(_00038_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08611_ (.I(_03087_),
    .Z(_04165_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08612_ (.A1(net32),
    .A2(_01069_),
    .B(_04121_),
    .ZN(_04166_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08613_ (.A1(_04165_),
    .A2(_03484_),
    .B(_04151_),
    .C(_04166_),
    .ZN(_04167_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08614_ (.I(_05127_),
    .ZN(_04168_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08615_ (.I(_05124_),
    .ZN(_04169_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08616_ (.A1(_04169_),
    .A2(_04141_),
    .ZN(_04170_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08617_ (.A1(_05123_),
    .A2(_04170_),
    .B(_05128_),
    .ZN(_04171_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08618_ (.A1(_04168_),
    .A2(_04171_),
    .ZN(_04172_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08619_ (.A1(_05132_),
    .A2(_04172_),
    .ZN(_04173_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08620_ (.A1(net96),
    .A2(net97),
    .A3(net98),
    .A4(_04145_),
    .Z(_04174_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08621_ (.A1(net99),
    .A2(_04174_),
    .ZN(_04175_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _08622_ (.A1(_04063_),
    .A2(_04173_),
    .B1(_04175_),
    .B2(_04064_),
    .ZN(_04176_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08623_ (.A1(_04167_),
    .A2(_04176_),
    .Z(_04177_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _08624_ (.I(_04177_),
    .Z(_04178_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08625_ (.I0(\dp.rf.rf[10][13] ),
    .I1(_04178_),
    .S(_04083_),
    .Z(_00039_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08626_ (.I(net33),
    .ZN(_04179_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08627_ (.A1(_04179_),
    .A2(_04087_),
    .B(_04091_),
    .ZN(_04180_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _08628_ (.A1(net93),
    .A2(net66),
    .B(_04067_),
    .C(_04180_),
    .ZN(_04181_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _08629_ (.I(_03871_),
    .Z(_04182_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08630_ (.A1(net96),
    .A2(net97),
    .A3(net98),
    .A4(net99),
    .Z(_04183_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08631_ (.A1(_04116_),
    .A2(_04183_),
    .ZN(_04184_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08632_ (.A1(net100),
    .A2(_04184_),
    .ZN(_04185_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08633_ (.A1(_05120_),
    .A2(_05124_),
    .A3(_05128_),
    .A4(_05132_),
    .Z(_04186_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08634_ (.A1(_05116_),
    .A2(_04186_),
    .ZN(_04187_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08635_ (.A1(_05124_),
    .A2(_05119_),
    .Z(_04188_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08636_ (.A1(_05123_),
    .A2(_04188_),
    .B(_05128_),
    .ZN(_04189_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08637_ (.A1(_04168_),
    .A2(_04189_),
    .ZN(_04190_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _08638_ (.A1(_05132_),
    .A2(_04190_),
    .B1(_04186_),
    .B2(_05115_),
    .C(_05131_),
    .ZN(_04191_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08639_ (.A1(_04108_),
    .A2(_04187_),
    .B(_04191_),
    .ZN(_04192_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08640_ (.A1(_05136_),
    .A2(_04192_),
    .Z(_04193_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08641_ (.A1(_04182_),
    .A2(_04185_),
    .B1(_04193_),
    .B2(_04154_),
    .ZN(_04194_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08642_ (.A1(_04181_),
    .A2(_04194_),
    .ZN(_04195_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _08643_ (.I(_04195_),
    .Z(_04196_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08644_ (.I0(\dp.rf.rf[10][14] ),
    .I1(_04196_),
    .S(_04083_),
    .Z(_00040_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08645_ (.A1(_04139_),
    .A2(_04186_),
    .ZN(_04197_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08646_ (.A1(_04191_),
    .A2(_04197_),
    .ZN(_04198_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08647_ (.A1(_05136_),
    .A2(_04198_),
    .B(_05135_),
    .ZN(_04199_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08648_ (.A1(_05140_),
    .A2(_04199_),
    .ZN(_04200_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08649_ (.A1(_04095_),
    .A2(_04200_),
    .ZN(_04201_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08650_ (.A1(net100),
    .A2(_04145_),
    .A3(_04183_),
    .Z(_04202_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08651_ (.A1(net101),
    .A2(_04202_),
    .Z(_04203_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08652_ (.A1(_03012_),
    .A2(_04165_),
    .Z(_04204_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08653_ (.A1(net34),
    .A2(_01069_),
    .B(_04121_),
    .ZN(_04205_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08654_ (.A1(_03511_),
    .A2(_04204_),
    .B(_04205_),
    .C(_04151_),
    .ZN(_04206_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08655_ (.A1(_04182_),
    .A2(_04203_),
    .B1(_04206_),
    .B2(_03522_),
    .ZN(_04207_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08656_ (.A1(_04201_),
    .A2(_04207_),
    .ZN(_04208_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _08657_ (.I(_04208_),
    .Z(_04209_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08658_ (.I0(\dp.rf.rf[10][15] ),
    .I1(_04209_),
    .S(_04083_),
    .Z(_00041_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08659_ (.A1(_04165_),
    .A2(_03540_),
    .Z(_04210_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08660_ (.A1(_03008_),
    .A2(_03088_),
    .ZN(_04211_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08661_ (.I(_04211_),
    .Z(_04212_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08662_ (.I(_04211_),
    .ZN(_04213_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08663_ (.A1(_03009_),
    .A2(net34),
    .A3(_04213_),
    .Z(_04214_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08664_ (.I(_04214_),
    .Z(_04215_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08665_ (.A1(net35),
    .A2(_04212_),
    .B(_04215_),
    .ZN(_04216_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08666_ (.A1(_04087_),
    .A2(_04216_),
    .B(_04091_),
    .ZN(_04217_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08667_ (.A1(_04067_),
    .A2(_04217_),
    .ZN(_04218_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08668_ (.A1(net100),
    .A2(net101),
    .A3(_04116_),
    .A4(_04183_),
    .Z(_04219_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08669_ (.A1(net102),
    .A2(_04219_),
    .Z(_04220_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08670_ (.A1(_05136_),
    .A2(_04192_),
    .Z(_04221_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08671_ (.A1(_05135_),
    .A2(_04221_),
    .Z(_04222_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08672_ (.A1(_05140_),
    .A2(_04222_),
    .B(_05139_),
    .ZN(_04223_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08673_ (.A1(_05144_),
    .A2(_04223_),
    .ZN(_04224_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08674_ (.A1(_04161_),
    .A2(_04220_),
    .B1(_04224_),
    .B2(_04154_),
    .ZN(_04225_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08675_ (.A1(_04210_),
    .A2(_04218_),
    .B(_04225_),
    .ZN(_04226_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08676_ (.I(_04226_),
    .Z(_04227_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08677_ (.I0(\dp.rf.rf[10][16] ),
    .I1(_04227_),
    .S(_04083_),
    .Z(_00042_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08678_ (.A1(net36),
    .A2(_04212_),
    .B(_04215_),
    .ZN(_04228_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08679_ (.A1(_04086_),
    .A2(_04228_),
    .B(_04090_),
    .ZN(_04229_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08680_ (.A1(_04123_),
    .A2(_04229_),
    .ZN(_04230_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08681_ (.A1(_03546_),
    .A2(_04204_),
    .Z(_04231_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08682_ (.A1(net100),
    .A2(net101),
    .A3(net102),
    .A4(_04183_),
    .Z(_04232_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08683_ (.A1(_04145_),
    .A2(_04232_),
    .ZN(_04233_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08684_ (.A1(net103),
    .A2(_04233_),
    .ZN(_04234_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08685_ (.A1(_05136_),
    .A2(_05140_),
    .A3(_05144_),
    .Z(_04235_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08686_ (.I(_05143_),
    .ZN(_04236_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08687_ (.A1(_05140_),
    .A2(_05135_),
    .Z(_04237_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08688_ (.A1(_05139_),
    .A2(_04237_),
    .B(_05144_),
    .ZN(_04238_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08689_ (.A1(_04236_),
    .A2(_04238_),
    .ZN(_04239_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08690_ (.A1(_04198_),
    .A2(_04235_),
    .B(_04239_),
    .ZN(_04240_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08691_ (.A1(_05148_),
    .A2(_04240_),
    .ZN(_04241_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08692_ (.A1(_04161_),
    .A2(_04234_),
    .B1(_04241_),
    .B2(_04154_),
    .ZN(_04242_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _08693_ (.A1(_03561_),
    .A2(_04230_),
    .A3(_04231_),
    .B(_04242_),
    .ZN(_04243_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _08694_ (.I(_04243_),
    .Z(_04244_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _08695_ (.I(_04082_),
    .Z(_04245_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08696_ (.I0(\dp.rf.rf[10][17] ),
    .I1(_04244_),
    .S(_04245_),
    .Z(_00043_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08697_ (.A1(net57),
    .A2(_04086_),
    .B1(_04213_),
    .B2(net34),
    .ZN(_04246_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08698_ (.A1(net5),
    .A2(net37),
    .ZN(_04247_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _08699_ (.A1(_02170_),
    .A2(_04246_),
    .B(_04247_),
    .C(_03089_),
    .ZN(_04248_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _08700_ (.A1(net93),
    .A2(net70),
    .B(_04067_),
    .C(_04248_),
    .ZN(_04249_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08701_ (.A1(net103),
    .A2(_04116_),
    .A3(_04232_),
    .Z(_04250_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08702_ (.A1(net104),
    .A2(_04250_),
    .Z(_04251_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08703_ (.I(_05148_),
    .ZN(_04252_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08704_ (.A1(_04192_),
    .A2(_04235_),
    .B(_04239_),
    .ZN(_04253_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08705_ (.I(_05147_),
    .ZN(_04254_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08706_ (.A1(_04252_),
    .A2(_04253_),
    .B(_04254_),
    .ZN(_04255_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08707_ (.A1(_05152_),
    .A2(_04255_),
    .Z(_04256_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08708_ (.A1(_04182_),
    .A2(_04251_),
    .B1(_04256_),
    .B2(_04154_),
    .ZN(_04257_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08709_ (.A1(_04249_),
    .A2(_04257_),
    .ZN(_04258_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _08710_ (.I(_04258_),
    .Z(_04259_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08711_ (.I0(\dp.rf.rf[10][18] ),
    .I1(_04259_),
    .S(_04245_),
    .Z(_00044_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08712_ (.A1(net38),
    .A2(_04212_),
    .B(_04215_),
    .ZN(_04260_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08713_ (.A1(_04087_),
    .A2(_04260_),
    .B(_04091_),
    .ZN(_04261_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _08714_ (.A1(net93),
    .A2(net71),
    .B(_04123_),
    .C(_04261_),
    .ZN(_04262_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08715_ (.A1(net103),
    .A2(net104),
    .A3(_04145_),
    .A4(_04232_),
    .Z(_04263_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08716_ (.A1(net105),
    .A2(_04263_),
    .Z(_04264_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08717_ (.A1(_04252_),
    .A2(_04240_),
    .B(_04254_),
    .ZN(_04265_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08718_ (.A1(_05152_),
    .A2(_04265_),
    .B(_05151_),
    .ZN(_04266_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08719_ (.A1(_05156_),
    .A2(_04266_),
    .ZN(_04267_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08720_ (.A1(_04182_),
    .A2(_04264_),
    .B1(_04267_),
    .B2(_04154_),
    .ZN(_04268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08721_ (.A1(_04262_),
    .A2(_04268_),
    .ZN(_04269_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _08722_ (.I(_04269_),
    .Z(_04270_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08723_ (.I0(\dp.rf.rf[10][19] ),
    .I1(_04270_),
    .S(_04245_),
    .Z(_00045_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08724_ (.A1(net106),
    .A2(_04064_),
    .ZN(_04271_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08725_ (.A1(net39),
    .A2(_03089_),
    .Z(_04272_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08726_ (.A1(_04165_),
    .A2(net72),
    .B(_04151_),
    .C(_04272_),
    .ZN(_04273_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08727_ (.A1(_04823_),
    .A2(_04095_),
    .B(_04271_),
    .C(_04273_),
    .ZN(_04274_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08728_ (.I(_04274_),
    .Z(_04275_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08729_ (.I0(\dp.rf.rf[10][1] ),
    .I1(_04275_),
    .S(_04245_),
    .Z(_00046_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08730_ (.A1(_04165_),
    .A2(_03634_),
    .Z(_04276_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08731_ (.A1(net40),
    .A2(_04212_),
    .B(_04215_),
    .ZN(_04277_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08732_ (.A1(_04087_),
    .A2(_04277_),
    .B(_04091_),
    .ZN(_04278_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08733_ (.A1(_04067_),
    .A2(_04278_),
    .ZN(_04279_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08734_ (.A1(_05148_),
    .A2(_05152_),
    .A3(_04192_),
    .A4(_04235_),
    .Z(_04280_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08735_ (.A1(_05148_),
    .A2(_05152_),
    .A3(_04239_),
    .Z(_04281_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08736_ (.A1(_05152_),
    .A2(_05147_),
    .Z(_04282_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08737_ (.A1(_04281_),
    .A2(_04282_),
    .Z(_04283_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08738_ (.A1(_05151_),
    .A2(_04280_),
    .A3(_04283_),
    .Z(_04284_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08739_ (.A1(_05156_),
    .A2(_04284_),
    .B(_05155_),
    .ZN(_04285_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08740_ (.A1(_05160_),
    .A2(_04285_),
    .ZN(_04286_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08741_ (.A1(net103),
    .A2(net104),
    .A3(net105),
    .A4(_04232_),
    .Z(_04287_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08742_ (.A1(_04116_),
    .A2(_04287_),
    .ZN(_04288_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08743_ (.A1(net107),
    .A2(_04288_),
    .ZN(_04289_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08744_ (.A1(_04154_),
    .A2(_04286_),
    .B1(_04289_),
    .B2(_04161_),
    .ZN(_04290_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08745_ (.A1(_04276_),
    .A2(_04279_),
    .B(_04290_),
    .ZN(_04291_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _08746_ (.I(_04291_),
    .Z(_04292_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08747_ (.I0(\dp.rf.rf[10][20] ),
    .I1(_04292_),
    .S(_04245_),
    .Z(_00047_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08748_ (.A1(net41),
    .A2(_04212_),
    .B(_04215_),
    .ZN(_04293_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08749_ (.A1(_04087_),
    .A2(_04293_),
    .B(_04091_),
    .ZN(_04294_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08750_ (.A1(net93),
    .A2(net74),
    .B(_04123_),
    .C(_04294_),
    .ZN(_04295_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08751_ (.I(_05160_),
    .ZN(_04296_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08752_ (.A1(_05148_),
    .A2(_04186_),
    .A3(_04235_),
    .Z(_04297_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08753_ (.A1(_05148_),
    .A2(_04235_),
    .ZN(_04298_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08754_ (.A1(_05148_),
    .A2(_04239_),
    .ZN(_04299_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08755_ (.A1(_04191_),
    .A2(_04298_),
    .B(_04299_),
    .ZN(_04300_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08756_ (.A1(_05147_),
    .A2(_05151_),
    .A3(_05155_),
    .Z(_04301_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08757_ (.A1(_04139_),
    .A2(_04297_),
    .B(_04300_),
    .C(_04301_),
    .ZN(_04302_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08758_ (.A1(_05152_),
    .A2(_05151_),
    .Z(_04303_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08759_ (.A1(_05156_),
    .A2(_04303_),
    .B(_05155_),
    .ZN(_04304_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08760_ (.I(_05159_),
    .ZN(_04305_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08761_ (.A1(_04296_),
    .A2(_04302_),
    .A3(_04304_),
    .B(_04305_),
    .ZN(_04306_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08762_ (.A1(_05164_),
    .A2(_04306_),
    .Z(_04307_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08763_ (.A1(net107),
    .A2(_04287_),
    .Z(_04308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08764_ (.A1(_04145_),
    .A2(_04308_),
    .ZN(_04309_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08765_ (.A1(net108),
    .A2(_04309_),
    .ZN(_04310_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08766_ (.A1(_04095_),
    .A2(_04307_),
    .B1(_04310_),
    .B2(_03872_),
    .ZN(_04311_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08767_ (.A1(_04295_),
    .A2(_04311_),
    .ZN(_04312_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _08768_ (.I(_04312_),
    .Z(_04313_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08769_ (.I0(\dp.rf.rf[10][21] ),
    .I1(_04313_),
    .S(_04245_),
    .Z(_00048_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08770_ (.A1(net42),
    .A2(_04212_),
    .B(_04215_),
    .ZN(_04314_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08771_ (.A1(_04087_),
    .A2(_04314_),
    .B(_04091_),
    .ZN(_04315_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08772_ (.A1(net93),
    .A2(net75),
    .B(_04123_),
    .C(_04315_),
    .ZN(_04316_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08773_ (.A1(_05151_),
    .A2(_05155_),
    .Z(_04317_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08774_ (.A1(_05156_),
    .A2(_05155_),
    .Z(_04318_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08775_ (.A1(_05160_),
    .A2(_04318_),
    .Z(_04319_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _08776_ (.A1(_04280_),
    .A2(_04283_),
    .A3(_04317_),
    .B(_04319_),
    .ZN(_04320_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08777_ (.A1(_04305_),
    .A2(_04320_),
    .ZN(_04321_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08778_ (.A1(_05164_),
    .A2(_04321_),
    .B(_05163_),
    .ZN(_04322_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08779_ (.A1(_05168_),
    .A2(_04322_),
    .ZN(_04323_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08780_ (.A1(net108),
    .A2(_04116_),
    .A3(_04308_),
    .Z(_04324_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08781_ (.A1(net109),
    .A2(_04324_),
    .Z(_04325_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08782_ (.A1(_04095_),
    .A2(_04323_),
    .B1(_04325_),
    .B2(_03872_),
    .ZN(_04326_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08783_ (.A1(_04316_),
    .A2(_04326_),
    .ZN(_04327_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _08784_ (.I(_04327_),
    .Z(_04328_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08785_ (.I0(\dp.rf.rf[10][22] ),
    .I1(_04328_),
    .S(_04245_),
    .Z(_00049_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08786_ (.I(_05167_),
    .ZN(_04329_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08787_ (.A1(_05164_),
    .A2(_04306_),
    .Z(_04330_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08788_ (.A1(_05163_),
    .A2(_04330_),
    .B(_05168_),
    .ZN(_04331_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08789_ (.A1(_04329_),
    .A2(_04331_),
    .ZN(_04332_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08790_ (.A1(_05172_),
    .A2(_04332_),
    .ZN(_04333_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08791_ (.A1(net43),
    .A2(_04211_),
    .B(_04214_),
    .ZN(_04334_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08792_ (.A1(_04086_),
    .A2(_04334_),
    .B(_04090_),
    .ZN(_04335_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08793_ (.A1(_04123_),
    .A2(_04335_),
    .ZN(_04336_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08794_ (.A1(_03694_),
    .A2(_03703_),
    .B(_03089_),
    .ZN(_04337_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08795_ (.A1(net108),
    .A2(net109),
    .Z(_04338_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08796_ (.A1(_04145_),
    .A2(_04308_),
    .A3(_04338_),
    .Z(_04339_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08797_ (.A1(net110),
    .A2(_04339_),
    .ZN(_04340_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_4 _08798_ (.A1(_04063_),
    .A2(_04333_),
    .B1(_04336_),
    .B2(_04337_),
    .C1(_04340_),
    .C2(_04064_),
    .ZN(_04341_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _08799_ (.I(_04341_),
    .Z(_04342_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08800_ (.I0(\dp.rf.rf[10][23] ),
    .I1(_04342_),
    .S(_04245_),
    .Z(_00050_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08801_ (.A1(_03335_),
    .A2(_03710_),
    .B(_03721_),
    .ZN(_04343_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08802_ (.A1(_04068_),
    .A2(_04343_),
    .ZN(_04344_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08803_ (.A1(net44),
    .A2(_04212_),
    .B(_04215_),
    .ZN(_04345_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08804_ (.A1(_04087_),
    .A2(_04345_),
    .B(_04091_),
    .ZN(_04346_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08805_ (.A1(_03343_),
    .A2(_03712_),
    .ZN(_04347_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08806_ (.A1(_04067_),
    .A2(_04346_),
    .A3(_04347_),
    .ZN(_04348_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _08807_ (.A1(net110),
    .A2(_04116_),
    .A3(_04308_),
    .A4(_04338_),
    .ZN(_04349_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08808_ (.A1(net111),
    .A2(_04349_),
    .ZN(_04350_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08809_ (.A1(_05159_),
    .A2(_05163_),
    .A3(_05167_),
    .ZN(_04351_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08810_ (.A1(_05164_),
    .A2(_05163_),
    .Z(_04352_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08811_ (.A1(_05168_),
    .A2(_04352_),
    .B(_05167_),
    .ZN(_04353_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08812_ (.A1(_04320_),
    .A2(_04351_),
    .B(_04353_),
    .ZN(_04354_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08813_ (.A1(_05172_),
    .A2(_04354_),
    .B(_05171_),
    .ZN(_04355_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08814_ (.A1(_05176_),
    .A2(_04355_),
    .ZN(_04356_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _08815_ (.A1(_04161_),
    .A2(_04350_),
    .B1(_04356_),
    .B2(_04154_),
    .ZN(_04357_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08816_ (.A1(_04344_),
    .A2(_04348_),
    .B(_04357_),
    .ZN(_04358_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _08817_ (.I(_04358_),
    .Z(_04359_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08818_ (.I0(\dp.rf.rf[10][24] ),
    .I1(_04359_),
    .S(_04245_),
    .Z(_00051_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08819_ (.A1(net45),
    .A2(_04212_),
    .B(_04215_),
    .ZN(_04360_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08820_ (.A1(_04087_),
    .A2(_04360_),
    .B(_04091_),
    .ZN(_04361_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08821_ (.A1(net93),
    .A2(net78),
    .B(_04123_),
    .C(_04361_),
    .ZN(_04362_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08822_ (.A1(net110),
    .A2(net111),
    .A3(_04308_),
    .A4(_04338_),
    .Z(_04363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08823_ (.A1(_04145_),
    .A2(_04363_),
    .ZN(_04364_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08824_ (.A1(net112),
    .A2(_04364_),
    .ZN(_04365_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08825_ (.A1(_05168_),
    .A2(_05172_),
    .A3(_05176_),
    .Z(_04366_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08826_ (.A1(_05160_),
    .A2(_05164_),
    .A3(_04366_),
    .ZN(_04367_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08827_ (.A1(_04302_),
    .A2(_04304_),
    .A3(_04367_),
    .Z(_04368_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08828_ (.I(_05171_),
    .ZN(_04369_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08829_ (.A1(_05168_),
    .A2(_05163_),
    .Z(_04370_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08830_ (.A1(_05167_),
    .A2(_04370_),
    .B(_05172_),
    .ZN(_04371_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08831_ (.A1(_04369_),
    .A2(_04371_),
    .ZN(_04372_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08832_ (.A1(_05164_),
    .A2(_05159_),
    .A3(_04366_),
    .Z(_04373_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08833_ (.A1(_05176_),
    .A2(_04372_),
    .B(_04373_),
    .C(_05175_),
    .ZN(_04374_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08834_ (.I(_05180_),
    .ZN(_04375_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08835_ (.A1(_04368_),
    .A2(_04374_),
    .B(_04375_),
    .ZN(_04376_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08836_ (.A1(_04375_),
    .A2(_04368_),
    .A3(_04374_),
    .Z(_04377_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08837_ (.A1(_04376_),
    .A2(_04377_),
    .ZN(_04378_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08838_ (.A1(_03872_),
    .A2(_04365_),
    .B1(_04378_),
    .B2(_04154_),
    .ZN(_04379_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08839_ (.A1(_04362_),
    .A2(_04379_),
    .ZN(_04380_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _08840_ (.I(_04380_),
    .Z(_04381_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08841_ (.I0(\dp.rf.rf[10][25] ),
    .I1(_04381_),
    .S(_04245_),
    .Z(_00052_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08842_ (.I(_05184_),
    .ZN(_04382_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08843_ (.A1(_05171_),
    .A2(_05175_),
    .A3(_05179_),
    .Z(_04383_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08844_ (.A1(_05172_),
    .A2(_05171_),
    .B(_05176_),
    .ZN(_04384_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08845_ (.A1(_05175_),
    .A2(_05179_),
    .ZN(_04385_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08846_ (.A1(_04384_),
    .A2(_04385_),
    .ZN(_04386_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _08847_ (.A1(_05180_),
    .A2(_05179_),
    .B1(_04354_),
    .B2(_04383_),
    .C(_04386_),
    .ZN(_04387_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08848_ (.A1(_04382_),
    .A2(_04387_),
    .ZN(_04388_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08849_ (.A1(net112),
    .A2(_04116_),
    .A3(_04363_),
    .Z(_04389_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08850_ (.A1(net113),
    .A2(_04389_),
    .ZN(_04390_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08851_ (.A1(net46),
    .A2(_04211_),
    .B(_04214_),
    .ZN(_04391_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08852_ (.A1(_04086_),
    .A2(_04391_),
    .B(_04090_),
    .ZN(_04392_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08853_ (.A1(_04068_),
    .A2(net79),
    .B(_04066_),
    .C(_04392_),
    .ZN(_04393_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _08854_ (.A1(_04063_),
    .A2(_04388_),
    .B1(_04390_),
    .B2(_04064_),
    .C(_04393_),
    .ZN(_04394_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _08855_ (.I(_04394_),
    .Z(_04395_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _08856_ (.I(_04082_),
    .Z(_04396_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08857_ (.I0(\dp.rf.rf[10][26] ),
    .I1(_04395_),
    .S(_04396_),
    .Z(_00053_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08858_ (.A1(_03775_),
    .A2(_03782_),
    .B(_04068_),
    .ZN(_04397_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08859_ (.A1(net47),
    .A2(_04212_),
    .B(_04215_),
    .ZN(_04398_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08860_ (.A1(_04087_),
    .A2(_04398_),
    .B(_04091_),
    .ZN(_04399_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08861_ (.A1(_04067_),
    .A2(_04399_),
    .ZN(_04400_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08862_ (.I(_05183_),
    .ZN(_04401_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08863_ (.A1(_05179_),
    .A2(_04376_),
    .B(_05184_),
    .ZN(_04402_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08864_ (.A1(_04401_),
    .A2(_04402_),
    .Z(_04403_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08865_ (.A1(_05188_),
    .A2(_04403_),
    .ZN(_04404_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08866_ (.A1(net112),
    .A2(net113),
    .A3(_04145_),
    .A4(_04363_),
    .Z(_04405_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08867_ (.A1(net114),
    .A2(_04405_),
    .Z(_04406_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08868_ (.A1(_04154_),
    .A2(_04404_),
    .B1(_04406_),
    .B2(_04161_),
    .ZN(_04407_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08869_ (.A1(_04397_),
    .A2(_04400_),
    .B(_04407_),
    .ZN(_04408_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _08870_ (.I(_04408_),
    .Z(_04409_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08871_ (.I0(\dp.rf.rf[10][27] ),
    .I1(_04409_),
    .S(_04396_),
    .Z(_00054_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08872_ (.A1(_04382_),
    .A2(_04387_),
    .B(_04401_),
    .ZN(_04410_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08873_ (.A1(_05188_),
    .A2(_04410_),
    .B(_05187_),
    .ZN(_04411_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08874_ (.A1(_05192_),
    .A2(_04411_),
    .Z(_04412_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08875_ (.A1(net112),
    .A2(net113),
    .A3(net114),
    .A4(_04363_),
    .Z(_04413_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08876_ (.A1(_04116_),
    .A2(_04413_),
    .ZN(_04414_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08877_ (.A1(net115),
    .A2(_04414_),
    .ZN(_04415_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08878_ (.A1(_03872_),
    .A2(_04415_),
    .ZN(_04416_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08879_ (.A1(net48),
    .A2(_04211_),
    .B(_04214_),
    .ZN(_04417_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08880_ (.A1(_04086_),
    .A2(_04417_),
    .B(_04090_),
    .ZN(_04418_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08881_ (.A1(_04068_),
    .A2(net81),
    .B(_04066_),
    .C(_04418_),
    .ZN(_04419_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _08882_ (.A1(_04063_),
    .A2(_04412_),
    .B(_04416_),
    .C(_04419_),
    .ZN(_04420_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _08883_ (.I(_04420_),
    .Z(_04421_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08884_ (.I0(\dp.rf.rf[10][28] ),
    .I1(_04421_),
    .S(_04396_),
    .Z(_00055_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08885_ (.A1(_05180_),
    .A2(_05184_),
    .A3(_05188_),
    .ZN(_04422_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08886_ (.A1(_04368_),
    .A2(_04374_),
    .B(_04422_),
    .ZN(_04423_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08887_ (.A1(_05188_),
    .A2(_05183_),
    .Z(_04424_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08888_ (.A1(_05184_),
    .A2(_05188_),
    .A3(_05179_),
    .Z(_04425_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _08889_ (.A1(_05187_),
    .A2(_04423_),
    .A3(_04424_),
    .A4(_04425_),
    .Z(_04426_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08890_ (.A1(_05192_),
    .A2(_04426_),
    .Z(_04427_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08891_ (.A1(_05191_),
    .A2(_04427_),
    .Z(_04428_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08892_ (.A1(_05196_),
    .A2(_04428_),
    .ZN(_04429_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08893_ (.A1(net115),
    .A2(_04413_),
    .Z(_04430_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08894_ (.A1(_04145_),
    .A2(_04430_),
    .ZN(_04431_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08895_ (.A1(net116),
    .A2(_04431_),
    .ZN(_04432_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08896_ (.A1(net49),
    .A2(_04211_),
    .B(_04214_),
    .ZN(_04433_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08897_ (.A1(_04086_),
    .A2(_04433_),
    .B(_04090_),
    .ZN(_04434_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08898_ (.A1(_04066_),
    .A2(_04434_),
    .Z(_04435_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08899_ (.A1(_03799_),
    .A2(_03806_),
    .A3(_03825_),
    .B(_04165_),
    .ZN(_04436_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08900_ (.A1(_04161_),
    .A2(_04432_),
    .B1(_04435_),
    .B2(_04436_),
    .ZN(_04437_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _08901_ (.A1(_04063_),
    .A2(_04182_),
    .A3(_04429_),
    .B(_04437_),
    .ZN(_04438_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _08902_ (.I(_04438_),
    .Z(_04439_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08903_ (.I0(\dp.rf.rf[10][29] ),
    .I1(_04439_),
    .S(_04396_),
    .Z(_00056_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08904_ (.A1(net50),
    .A2(_03089_),
    .Z(_04440_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08905_ (.A1(_04165_),
    .A2(net83),
    .B(_04440_),
    .ZN(_04441_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08906_ (.I(net117),
    .ZN(_04442_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08907_ (.A1(_04822_),
    .A2(_05086_),
    .Z(_04443_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _08908_ (.A1(_04442_),
    .A2(_04064_),
    .B1(_04443_),
    .B2(_04063_),
    .ZN(_04444_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08909_ (.A1(_04067_),
    .A2(_04441_),
    .B(_04444_),
    .ZN(_04445_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _08910_ (.I(_04445_),
    .Z(_04446_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08911_ (.I0(\dp.rf.rf[10][2] ),
    .I1(_04446_),
    .S(_04396_),
    .Z(_00057_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08912_ (.A1(_05184_),
    .A2(_05188_),
    .A3(_05192_),
    .ZN(_04447_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08913_ (.A1(_05188_),
    .A2(_05192_),
    .A3(_05183_),
    .Z(_04448_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08914_ (.A1(_05192_),
    .A2(_05187_),
    .B(_04448_),
    .ZN(_04449_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08915_ (.I(_05191_),
    .ZN(_04450_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08916_ (.A1(_04387_),
    .A2(_04447_),
    .B(_04449_),
    .C(_04450_),
    .ZN(_04451_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08917_ (.A1(_05196_),
    .A2(_04451_),
    .B(_05195_),
    .ZN(_04452_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08918_ (.A1(_05200_),
    .A2(_04452_),
    .Z(_04453_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08919_ (.A1(net51),
    .A2(_04212_),
    .B(_04215_),
    .ZN(_04454_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08920_ (.A1(_04086_),
    .A2(_04454_),
    .B(_04090_),
    .ZN(_04455_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08921_ (.A1(_04068_),
    .A2(net84),
    .B(_04123_),
    .C(_04455_),
    .ZN(_04456_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08922_ (.A1(net116),
    .A2(_04430_),
    .Z(_04457_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08923_ (.A1(_04116_),
    .A2(_04457_),
    .ZN(_04458_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08924_ (.A1(net118),
    .A2(_04458_),
    .ZN(_04459_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08925_ (.A1(_03872_),
    .A2(_04459_),
    .ZN(_04460_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _08926_ (.A1(_04063_),
    .A2(_04453_),
    .B(_04456_),
    .C(_04460_),
    .ZN(_04461_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _08927_ (.I(_04461_),
    .Z(_04462_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08928_ (.I0(\dp.rf.rf[10][30] ),
    .I1(_04462_),
    .S(_04396_),
    .Z(_00058_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08929_ (.I0(net119),
    .I1(_04833_),
    .S(_03867_),
    .Z(_04463_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08930_ (.A1(_05187_),
    .A2(_05191_),
    .Z(_04464_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _08931_ (.A1(_04423_),
    .A2(_04424_),
    .A3(_04425_),
    .A4(_04464_),
    .ZN(_04465_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08932_ (.A1(_05192_),
    .A2(_05191_),
    .B(_05196_),
    .ZN(_04466_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08933_ (.I(_05195_),
    .ZN(_04467_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08934_ (.A1(_04465_),
    .A2(_04466_),
    .B(_04467_),
    .ZN(_04468_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08935_ (.A1(_05200_),
    .A2(_04468_),
    .B(_05199_),
    .ZN(_04469_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _08936_ (.A1(net20),
    .A2(_04463_),
    .A3(_04469_),
    .ZN(_04470_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08937_ (.A1(_04059_),
    .A2(_04470_),
    .B(_04095_),
    .ZN(_04471_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08938_ (.I(_04471_),
    .Z(_04472_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08939_ (.A1(net118),
    .A2(_04144_),
    .A3(_04457_),
    .Z(_04473_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08940_ (.A1(net119),
    .A2(_04473_),
    .Z(_04474_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08941_ (.A1(_03871_),
    .A2(_04474_),
    .ZN(_04475_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08942_ (.A1(_04165_),
    .A2(_03853_),
    .A3(_03859_),
    .A4(_04475_),
    .Z(_04476_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08943_ (.A1(net52),
    .A2(_04211_),
    .B(_04214_),
    .ZN(_04477_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08944_ (.A1(_04086_),
    .A2(_04477_),
    .B(_04090_),
    .ZN(_04478_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08945_ (.A1(_03871_),
    .A2(_04474_),
    .B1(_04478_),
    .B2(_04066_),
    .ZN(_04479_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08946_ (.A1(_04165_),
    .A2(_03865_),
    .A3(_04475_),
    .Z(_04480_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _08947_ (.A1(_04476_),
    .A2(_04479_),
    .A3(_04480_),
    .Z(_04481_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _08948_ (.I(_04481_),
    .Z(_04482_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08949_ (.A1(_04083_),
    .A2(_04482_),
    .Z(_04483_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08950_ (.A1(\dp.rf.rf[10][31] ),
    .A2(_04083_),
    .ZN(_04484_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08951_ (.A1(_04472_),
    .A2(_04483_),
    .B(_04484_),
    .ZN(_00059_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08952_ (.A1(_04099_),
    .A2(_04129_),
    .ZN(_04485_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_4 _08953_ (.A1(net53),
    .A2(_03089_),
    .B1(_04094_),
    .B2(_04485_),
    .C1(_03871_),
    .C2(_05092_),
    .ZN(_04486_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _08954_ (.A1(net93),
    .A2(_03226_),
    .A3(_04151_),
    .B(_04486_),
    .ZN(_04487_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _08955_ (.I(_04487_),
    .Z(_04488_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08956_ (.I0(\dp.rf.rf[10][3] ),
    .I1(_04488_),
    .S(_04396_),
    .Z(_00060_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08957_ (.A1(_03380_),
    .A2(_03256_),
    .Z(_04489_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08958_ (.A1(_03087_),
    .A2(_04066_),
    .Z(_04490_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08959_ (.A1(_03182_),
    .A2(_03248_),
    .B(_04489_),
    .C(_04490_),
    .ZN(_04491_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08960_ (.A1(net121),
    .A2(_05091_),
    .Z(_04492_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08961_ (.A1(_04125_),
    .A2(_04102_),
    .ZN(_04493_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_4 _08962_ (.A1(net54),
    .A2(_04068_),
    .B1(_04161_),
    .B2(_04492_),
    .C1(_04493_),
    .C2(_04094_),
    .ZN(_04494_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08963_ (.A1(_04491_),
    .A2(_04494_),
    .ZN(_04495_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _08964_ (.I(_04495_),
    .Z(_04496_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08965_ (.I0(\dp.rf.rf[10][4] ),
    .I1(_04496_),
    .S(_04396_),
    .Z(_00061_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08966_ (.I(net55),
    .ZN(_04497_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08967_ (.I0(_04497_),
    .I1(_03293_),
    .S(_04165_),
    .Z(_04498_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08968_ (.A1(_04098_),
    .A2(_04132_),
    .ZN(_04499_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08969_ (.A1(net117),
    .A2(net120),
    .A3(net121),
    .Z(_04500_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08970_ (.A1(net122),
    .A2(_04500_),
    .Z(_04501_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _08971_ (.A1(_04063_),
    .A2(_04499_),
    .B1(_04501_),
    .B2(_04064_),
    .ZN(_04502_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08972_ (.A1(_04067_),
    .A2(_04498_),
    .B(_04502_),
    .ZN(_04503_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _08973_ (.I(_04503_),
    .Z(_04504_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08974_ (.I0(\dp.rf.rf[10][5] ),
    .I1(_04504_),
    .S(_04396_),
    .Z(_00062_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08975_ (.A1(_05104_),
    .A2(_04105_),
    .Z(_04505_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08976_ (.A1(_04094_),
    .A2(_04505_),
    .Z(_04506_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08977_ (.A1(net123),
    .A2(_04113_),
    .Z(_04507_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08978_ (.A1(_03871_),
    .A2(_04507_),
    .Z(_04508_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08979_ (.A1(net89),
    .A2(_04490_),
    .Z(_04509_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08980_ (.A1(net56),
    .A2(_03089_),
    .Z(_04510_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _08981_ (.A1(_04506_),
    .A2(_04508_),
    .A3(_04509_),
    .A4(_04510_),
    .Z(_04511_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _08982_ (.I(_04511_),
    .Z(_04512_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08983_ (.I0(\dp.rf.rf[10][6] ),
    .I1(_04512_),
    .S(_04396_),
    .Z(_00063_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08984_ (.I(_04133_),
    .ZN(_04513_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08985_ (.A1(_05104_),
    .A2(_04513_),
    .Z(_04514_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08986_ (.A1(_05103_),
    .A2(_04514_),
    .Z(_04515_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08987_ (.A1(_05108_),
    .A2(_04515_),
    .Z(_04516_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08988_ (.A1(_04095_),
    .A2(_04516_),
    .ZN(_04517_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08989_ (.A1(net123),
    .A2(_04143_),
    .ZN(_04518_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08990_ (.A1(net124),
    .A2(_04518_),
    .ZN(_04519_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08991_ (.A1(_03355_),
    .A2(_04490_),
    .Z(_04520_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_4 _08992_ (.A1(net57),
    .A2(_04068_),
    .B1(_04161_),
    .B2(_04519_),
    .C1(_04520_),
    .C2(_03345_),
    .ZN(_04521_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08993_ (.A1(_04517_),
    .A2(_04521_),
    .ZN(_04522_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _08994_ (.I(_04522_),
    .Z(_04523_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08995_ (.I0(\dp.rf.rf[10][7] ),
    .I1(_04523_),
    .S(_04082_),
    .Z(_00064_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08996_ (.A1(net58),
    .A2(_01069_),
    .Z(_04524_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _08997_ (.A1(_04068_),
    .A2(net91),
    .B1(_04121_),
    .B2(_04524_),
    .C(_04123_),
    .ZN(_04525_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08998_ (.A1(_05104_),
    .A2(_04105_),
    .Z(_04526_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08999_ (.A1(_05103_),
    .A2(_04526_),
    .Z(_04527_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09000_ (.A1(_05108_),
    .A2(_04527_),
    .B(_05107_),
    .ZN(_04528_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09001_ (.A1(_05112_),
    .A2(_04528_),
    .ZN(_04529_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09002_ (.A1(net123),
    .A2(net124),
    .A3(_04113_),
    .Z(_04530_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09003_ (.A1(net125),
    .A2(_04530_),
    .Z(_04531_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _09004_ (.A1(_04095_),
    .A2(_04529_),
    .B1(_04531_),
    .B2(_03872_),
    .ZN(_04532_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09005_ (.A1(_04525_),
    .A2(_04532_),
    .ZN(_04533_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09006_ (.I(_04533_),
    .Z(_04534_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09007_ (.I0(\dp.rf.rf[10][8] ),
    .I1(_04534_),
    .S(_04082_),
    .Z(_00065_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09008_ (.I(net59),
    .ZN(_04535_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09009_ (.A1(_04535_),
    .A2(_04086_),
    .B(_04090_),
    .ZN(_04536_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _09010_ (.A1(net93),
    .A2(net92),
    .B(_04123_),
    .C(_04536_),
    .ZN(_04537_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _09011_ (.A1(_04106_),
    .A2(_04515_),
    .B(_04136_),
    .C(_05116_),
    .ZN(_04538_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09012_ (.A1(_04139_),
    .A2(_04538_),
    .ZN(_04539_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09013_ (.A1(net123),
    .A2(net124),
    .A3(net125),
    .A4(_04143_),
    .Z(_04540_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09014_ (.A1(net126),
    .A2(_04540_),
    .Z(_04541_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09015_ (.A1(_04095_),
    .A2(_04539_),
    .B1(_04541_),
    .B2(_03872_),
    .ZN(_04542_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09016_ (.A1(_04537_),
    .A2(_04542_),
    .ZN(_04543_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09017_ (.I(_04543_),
    .Z(_04544_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09018_ (.I0(\dp.rf.rf[10][9] ),
    .I1(_04544_),
    .S(_04082_),
    .Z(_00066_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _09019_ (.A1(net26),
    .A2(net25),
    .A3(_04079_),
    .Z(_04545_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09020_ (.A1(_04075_),
    .A2(_04545_),
    .Z(_04546_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09021_ (.I(_04546_),
    .Z(_04547_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09022_ (.I0(\dp.rf.rf[11][0] ),
    .I1(_04073_),
    .S(_04547_),
    .Z(_00067_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09023_ (.I0(\dp.rf.rf[11][10] ),
    .I1(_04120_),
    .S(_04547_),
    .Z(_00068_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09024_ (.I0(\dp.rf.rf[11][11] ),
    .I1(_04150_),
    .S(_04547_),
    .Z(_00069_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09025_ (.I0(\dp.rf.rf[11][12] ),
    .I1(_04164_),
    .S(_04547_),
    .Z(_00070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09026_ (.I0(\dp.rf.rf[11][13] ),
    .I1(_04178_),
    .S(_04547_),
    .Z(_00071_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09027_ (.I0(\dp.rf.rf[11][14] ),
    .I1(_04196_),
    .S(_04547_),
    .Z(_00072_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09028_ (.I0(\dp.rf.rf[11][15] ),
    .I1(_04209_),
    .S(_04547_),
    .Z(_00073_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09029_ (.I0(\dp.rf.rf[11][16] ),
    .I1(_04227_),
    .S(_04547_),
    .Z(_00074_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09030_ (.I(_04546_),
    .Z(_04548_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09031_ (.I0(\dp.rf.rf[11][17] ),
    .I1(_04244_),
    .S(_04548_),
    .Z(_00075_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09032_ (.I0(\dp.rf.rf[11][18] ),
    .I1(_04259_),
    .S(_04548_),
    .Z(_00076_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09033_ (.I0(\dp.rf.rf[11][19] ),
    .I1(_04270_),
    .S(_04548_),
    .Z(_00077_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09034_ (.I0(\dp.rf.rf[11][1] ),
    .I1(_04275_),
    .S(_04548_),
    .Z(_00078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09035_ (.I0(\dp.rf.rf[11][20] ),
    .I1(_04292_),
    .S(_04548_),
    .Z(_00079_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09036_ (.I0(\dp.rf.rf[11][21] ),
    .I1(_04313_),
    .S(_04548_),
    .Z(_00080_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09037_ (.I0(\dp.rf.rf[11][22] ),
    .I1(_04328_),
    .S(_04548_),
    .Z(_00081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09038_ (.I0(\dp.rf.rf[11][23] ),
    .I1(_04342_),
    .S(_04548_),
    .Z(_00082_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09039_ (.I0(\dp.rf.rf[11][24] ),
    .I1(_04359_),
    .S(_04548_),
    .Z(_00083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09040_ (.I0(\dp.rf.rf[11][25] ),
    .I1(_04381_),
    .S(_04548_),
    .Z(_00084_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _09041_ (.I(_04546_),
    .Z(_04549_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09042_ (.I0(\dp.rf.rf[11][26] ),
    .I1(_04395_),
    .S(_04549_),
    .Z(_00085_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09043_ (.I0(\dp.rf.rf[11][27] ),
    .I1(_04409_),
    .S(_04549_),
    .Z(_00086_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09044_ (.I0(\dp.rf.rf[11][28] ),
    .I1(_04421_),
    .S(_04549_),
    .Z(_00087_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09045_ (.I0(\dp.rf.rf[11][29] ),
    .I1(_04439_),
    .S(_04549_),
    .Z(_00088_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09046_ (.I0(\dp.rf.rf[11][2] ),
    .I1(_04446_),
    .S(_04549_),
    .Z(_00089_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09047_ (.I0(\dp.rf.rf[11][30] ),
    .I1(_04462_),
    .S(_04549_),
    .Z(_00090_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09048_ (.I(_04481_),
    .Z(_04550_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09049_ (.A1(_04550_),
    .A2(_04547_),
    .Z(_04551_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09050_ (.A1(\dp.rf.rf[11][31] ),
    .A2(_04547_),
    .ZN(_04552_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09051_ (.A1(_04472_),
    .A2(_04551_),
    .B(_04552_),
    .ZN(_00091_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09052_ (.I0(\dp.rf.rf[11][3] ),
    .I1(_04488_),
    .S(_04549_),
    .Z(_00092_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09053_ (.I0(\dp.rf.rf[11][4] ),
    .I1(_04496_),
    .S(_04549_),
    .Z(_00093_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09054_ (.I0(\dp.rf.rf[11][5] ),
    .I1(_04504_),
    .S(_04549_),
    .Z(_00094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09055_ (.I0(\dp.rf.rf[11][6] ),
    .I1(_04512_),
    .S(_04549_),
    .Z(_00095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09056_ (.I0(\dp.rf.rf[11][7] ),
    .I1(_04523_),
    .S(_04546_),
    .Z(_00096_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09057_ (.I0(\dp.rf.rf[11][8] ),
    .I1(_04534_),
    .S(_04546_),
    .Z(_00097_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09058_ (.I0(\dp.rf.rf[11][9] ),
    .I1(_04544_),
    .S(_04546_),
    .Z(_00098_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09059_ (.I(_04072_),
    .Z(_04553_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09060_ (.A1(_02672_),
    .A2(net2),
    .A3(net27),
    .Z(_04554_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09061_ (.I(net2),
    .ZN(_04555_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09062_ (.A1(_04555_),
    .A2(_04074_),
    .Z(_04556_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09063_ (.A1(net26),
    .A2(_04556_),
    .ZN(_04557_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09064_ (.A1(_04080_),
    .A2(_04557_),
    .Z(_04558_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09065_ (.A1(_04554_),
    .A2(_04558_),
    .Z(_04559_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09066_ (.I(_04559_),
    .Z(_04560_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09067_ (.I0(\dp.rf.rf[12][0] ),
    .I1(_04553_),
    .S(_04560_),
    .Z(_00099_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09068_ (.I(_04119_),
    .Z(_04561_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09069_ (.I0(\dp.rf.rf[12][10] ),
    .I1(_04561_),
    .S(_04560_),
    .Z(_00100_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _09070_ (.I(_04149_),
    .Z(_04562_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09071_ (.I0(\dp.rf.rf[12][11] ),
    .I1(_04562_),
    .S(_04560_),
    .Z(_00101_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _09072_ (.I(_04163_),
    .Z(_04563_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09073_ (.I0(\dp.rf.rf[12][12] ),
    .I1(_04563_),
    .S(_04560_),
    .Z(_00102_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09074_ (.I(_04177_),
    .Z(_04564_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09075_ (.I0(\dp.rf.rf[12][13] ),
    .I1(_04564_),
    .S(_04560_),
    .Z(_00103_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _09076_ (.I(_04195_),
    .Z(_04565_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09077_ (.I0(\dp.rf.rf[12][14] ),
    .I1(_04565_),
    .S(_04560_),
    .Z(_00104_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _09078_ (.I(_04208_),
    .Z(_04566_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09079_ (.I0(\dp.rf.rf[12][15] ),
    .I1(_04566_),
    .S(_04560_),
    .Z(_00105_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _09080_ (.I(_04226_),
    .Z(_04567_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09081_ (.I0(\dp.rf.rf[12][16] ),
    .I1(_04567_),
    .S(_04560_),
    .Z(_00106_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09082_ (.I(_04243_),
    .Z(_04568_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _09083_ (.I(_04559_),
    .Z(_04569_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09084_ (.I0(\dp.rf.rf[12][17] ),
    .I1(_04568_),
    .S(_04569_),
    .Z(_00107_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _09085_ (.I(_04258_),
    .Z(_04570_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09086_ (.I0(\dp.rf.rf[12][18] ),
    .I1(_04570_),
    .S(_04569_),
    .Z(_00108_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09087_ (.I(_04269_),
    .Z(_04571_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09088_ (.I0(\dp.rf.rf[12][19] ),
    .I1(_04571_),
    .S(_04569_),
    .Z(_00109_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _09089_ (.I(_04274_),
    .Z(_04572_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09090_ (.I0(\dp.rf.rf[12][1] ),
    .I1(_04572_),
    .S(_04569_),
    .Z(_00110_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _09091_ (.I(_04291_),
    .Z(_04573_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09092_ (.I0(\dp.rf.rf[12][20] ),
    .I1(_04573_),
    .S(_04569_),
    .Z(_00111_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09093_ (.I(_04312_),
    .Z(_04574_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09094_ (.I0(\dp.rf.rf[12][21] ),
    .I1(_04574_),
    .S(_04569_),
    .Z(_00112_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09095_ (.I(_04327_),
    .Z(_04575_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09096_ (.I0(\dp.rf.rf[12][22] ),
    .I1(_04575_),
    .S(_04569_),
    .Z(_00113_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _09097_ (.I(_04341_),
    .Z(_04576_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09098_ (.I0(\dp.rf.rf[12][23] ),
    .I1(_04576_),
    .S(_04569_),
    .Z(_00114_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09099_ (.I(_04358_),
    .Z(_04577_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09100_ (.I0(\dp.rf.rf[12][24] ),
    .I1(_04577_),
    .S(_04569_),
    .Z(_00115_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09101_ (.I(_04380_),
    .Z(_04578_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09102_ (.I0(\dp.rf.rf[12][25] ),
    .I1(_04578_),
    .S(_04569_),
    .Z(_00116_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09103_ (.I(_04394_),
    .Z(_04579_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09104_ (.I(_04559_),
    .Z(_04580_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09105_ (.I0(\dp.rf.rf[12][26] ),
    .I1(_04579_),
    .S(_04580_),
    .Z(_00117_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09106_ (.I(_04408_),
    .Z(_04581_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09107_ (.I0(\dp.rf.rf[12][27] ),
    .I1(_04581_),
    .S(_04580_),
    .Z(_00118_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09108_ (.I(_04420_),
    .Z(_04582_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09109_ (.I0(\dp.rf.rf[12][28] ),
    .I1(_04582_),
    .S(_04580_),
    .Z(_00119_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09110_ (.I(_04438_),
    .Z(_04583_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09111_ (.I0(\dp.rf.rf[12][29] ),
    .I1(_04583_),
    .S(_04580_),
    .Z(_00120_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09112_ (.I(_04445_),
    .Z(_04584_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09113_ (.I0(\dp.rf.rf[12][2] ),
    .I1(_04584_),
    .S(_04580_),
    .Z(_00121_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09114_ (.I(_04461_),
    .Z(_04585_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09115_ (.I0(\dp.rf.rf[12][30] ),
    .I1(_04585_),
    .S(_04580_),
    .Z(_00122_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09116_ (.A1(_04550_),
    .A2(_04560_),
    .Z(_04586_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09117_ (.A1(\dp.rf.rf[12][31] ),
    .A2(_04560_),
    .ZN(_04587_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09118_ (.A1(_04472_),
    .A2(_04586_),
    .B(_04587_),
    .ZN(_00123_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09119_ (.I(_04487_),
    .Z(_04588_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09120_ (.I0(\dp.rf.rf[12][3] ),
    .I1(_04588_),
    .S(_04580_),
    .Z(_00124_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09121_ (.I(_04495_),
    .Z(_04589_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09122_ (.I0(\dp.rf.rf[12][4] ),
    .I1(_04589_),
    .S(_04580_),
    .Z(_00125_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09123_ (.I(_04503_),
    .Z(_04590_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09124_ (.I0(\dp.rf.rf[12][5] ),
    .I1(_04590_),
    .S(_04580_),
    .Z(_00126_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _09125_ (.I(_04511_),
    .Z(_04591_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09126_ (.I0(\dp.rf.rf[12][6] ),
    .I1(_04591_),
    .S(_04580_),
    .Z(_00127_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _09127_ (.I(_04522_),
    .Z(_04592_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09128_ (.I0(\dp.rf.rf[12][7] ),
    .I1(_04592_),
    .S(_04559_),
    .Z(_00128_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _09129_ (.I(_04533_),
    .Z(_04593_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09130_ (.I0(\dp.rf.rf[12][8] ),
    .I1(_04593_),
    .S(_04559_),
    .Z(_00129_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09131_ (.I(_04543_),
    .Z(_04594_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09132_ (.I0(\dp.rf.rf[12][9] ),
    .I1(_04594_),
    .S(_04559_),
    .Z(_00130_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _09133_ (.A1(_01101_),
    .A2(net25),
    .A3(_04079_),
    .Z(_04595_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09134_ (.A1(_04554_),
    .A2(_04595_),
    .ZN(_04596_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09135_ (.I(_04596_),
    .Z(_04597_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09136_ (.I0(_04073_),
    .I1(\dp.rf.rf[13][0] ),
    .S(_04597_),
    .Z(_00131_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09137_ (.I0(_04120_),
    .I1(\dp.rf.rf[13][10] ),
    .S(_04597_),
    .Z(_00132_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09138_ (.I0(_04150_),
    .I1(\dp.rf.rf[13][11] ),
    .S(_04597_),
    .Z(_00133_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09139_ (.I0(_04164_),
    .I1(\dp.rf.rf[13][12] ),
    .S(_04597_),
    .Z(_00134_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09140_ (.I0(_04178_),
    .I1(\dp.rf.rf[13][13] ),
    .S(_04597_),
    .Z(_00135_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09141_ (.I0(_04196_),
    .I1(\dp.rf.rf[13][14] ),
    .S(_04597_),
    .Z(_00136_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09142_ (.I0(_04209_),
    .I1(\dp.rf.rf[13][15] ),
    .S(_04597_),
    .Z(_00137_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09143_ (.I0(_04227_),
    .I1(\dp.rf.rf[13][16] ),
    .S(_04597_),
    .Z(_00138_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09144_ (.I0(_04244_),
    .I1(\dp.rf.rf[13][17] ),
    .S(_04597_),
    .Z(_00139_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _09145_ (.I(_04596_),
    .Z(_04598_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09146_ (.I0(_04259_),
    .I1(\dp.rf.rf[13][18] ),
    .S(_04598_),
    .Z(_00140_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09147_ (.I0(_04270_),
    .I1(\dp.rf.rf[13][19] ),
    .S(_04598_),
    .Z(_00141_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09148_ (.I0(_04275_),
    .I1(\dp.rf.rf[13][1] ),
    .S(_04598_),
    .Z(_00142_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09149_ (.I0(_04292_),
    .I1(\dp.rf.rf[13][20] ),
    .S(_04598_),
    .Z(_00143_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09150_ (.I0(_04313_),
    .I1(\dp.rf.rf[13][21] ),
    .S(_04598_),
    .Z(_00144_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09151_ (.I0(_04328_),
    .I1(\dp.rf.rf[13][22] ),
    .S(_04598_),
    .Z(_00145_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09152_ (.I0(_04342_),
    .I1(\dp.rf.rf[13][23] ),
    .S(_04598_),
    .Z(_00146_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09153_ (.I0(_04359_),
    .I1(\dp.rf.rf[13][24] ),
    .S(_04598_),
    .Z(_00147_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09154_ (.I0(_04381_),
    .I1(\dp.rf.rf[13][25] ),
    .S(_04598_),
    .Z(_00148_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09155_ (.I0(_04395_),
    .I1(\dp.rf.rf[13][26] ),
    .S(_04598_),
    .Z(_00149_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _09156_ (.I(_04596_),
    .Z(_04599_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09157_ (.I0(_04409_),
    .I1(\dp.rf.rf[13][27] ),
    .S(_04599_),
    .Z(_00150_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09158_ (.I0(_04421_),
    .I1(\dp.rf.rf[13][28] ),
    .S(_04599_),
    .Z(_00151_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09159_ (.I0(_04439_),
    .I1(\dp.rf.rf[13][29] ),
    .S(_04599_),
    .Z(_00152_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09160_ (.I0(_04446_),
    .I1(\dp.rf.rf[13][2] ),
    .S(_04599_),
    .Z(_00153_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09161_ (.I0(_04462_),
    .I1(\dp.rf.rf[13][30] ),
    .S(_04599_),
    .Z(_00154_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09162_ (.I(\dp.rf.rf[13][31] ),
    .ZN(_04600_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _09163_ (.I(_04595_),
    .Z(_04601_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09164_ (.A1(_04482_),
    .A2(_04554_),
    .A3(_04601_),
    .Z(_04602_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _09165_ (.I(_04471_),
    .Z(_04603_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09166_ (.A1(_04600_),
    .A2(_04597_),
    .B1(_04602_),
    .B2(_04603_),
    .ZN(_00155_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09167_ (.I0(_04488_),
    .I1(\dp.rf.rf[13][3] ),
    .S(_04599_),
    .Z(_00156_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09168_ (.I0(_04496_),
    .I1(\dp.rf.rf[13][4] ),
    .S(_04599_),
    .Z(_00157_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09169_ (.I0(_04504_),
    .I1(\dp.rf.rf[13][5] ),
    .S(_04599_),
    .Z(_00158_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09170_ (.I0(_04512_),
    .I1(\dp.rf.rf[13][6] ),
    .S(_04599_),
    .Z(_00159_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09171_ (.I0(_04523_),
    .I1(\dp.rf.rf[13][7] ),
    .S(_04599_),
    .Z(_00160_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09172_ (.I0(_04534_),
    .I1(\dp.rf.rf[13][8] ),
    .S(_04596_),
    .Z(_00161_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09173_ (.I0(_04544_),
    .I1(\dp.rf.rf[13][9] ),
    .S(_04596_),
    .Z(_00162_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09174_ (.A1(_04081_),
    .A2(_04554_),
    .Z(_04604_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09175_ (.I(_04604_),
    .Z(_04605_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09176_ (.I0(\dp.rf.rf[14][0] ),
    .I1(_04553_),
    .S(_04605_),
    .Z(_00163_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09177_ (.I0(\dp.rf.rf[14][10] ),
    .I1(_04561_),
    .S(_04605_),
    .Z(_00164_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09178_ (.I0(\dp.rf.rf[14][11] ),
    .I1(_04562_),
    .S(_04605_),
    .Z(_00165_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09179_ (.I0(\dp.rf.rf[14][12] ),
    .I1(_04563_),
    .S(_04605_),
    .Z(_00166_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09180_ (.I0(\dp.rf.rf[14][13] ),
    .I1(_04564_),
    .S(_04605_),
    .Z(_00167_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09181_ (.I0(\dp.rf.rf[14][14] ),
    .I1(_04565_),
    .S(_04605_),
    .Z(_00168_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09182_ (.I0(\dp.rf.rf[14][15] ),
    .I1(_04566_),
    .S(_04605_),
    .Z(_00169_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09183_ (.I0(\dp.rf.rf[14][16] ),
    .I1(_04567_),
    .S(_04605_),
    .Z(_00170_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _09184_ (.I(_04604_),
    .Z(_04606_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09185_ (.I0(\dp.rf.rf[14][17] ),
    .I1(_04568_),
    .S(_04606_),
    .Z(_00171_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09186_ (.I0(\dp.rf.rf[14][18] ),
    .I1(_04570_),
    .S(_04606_),
    .Z(_00172_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09187_ (.I0(\dp.rf.rf[14][19] ),
    .I1(_04571_),
    .S(_04606_),
    .Z(_00173_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09188_ (.I0(\dp.rf.rf[14][1] ),
    .I1(_04572_),
    .S(_04606_),
    .Z(_00174_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09189_ (.I0(\dp.rf.rf[14][20] ),
    .I1(_04573_),
    .S(_04606_),
    .Z(_00175_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09190_ (.I0(\dp.rf.rf[14][21] ),
    .I1(_04574_),
    .S(_04606_),
    .Z(_00176_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09191_ (.I0(\dp.rf.rf[14][22] ),
    .I1(_04575_),
    .S(_04606_),
    .Z(_00177_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09192_ (.I0(\dp.rf.rf[14][23] ),
    .I1(_04576_),
    .S(_04606_),
    .Z(_00178_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09193_ (.I0(\dp.rf.rf[14][24] ),
    .I1(_04577_),
    .S(_04606_),
    .Z(_00179_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09194_ (.I0(\dp.rf.rf[14][25] ),
    .I1(_04578_),
    .S(_04606_),
    .Z(_00180_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09195_ (.I(_04604_),
    .Z(_04607_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09196_ (.I0(\dp.rf.rf[14][26] ),
    .I1(_04579_),
    .S(_04607_),
    .Z(_00181_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09197_ (.I0(\dp.rf.rf[14][27] ),
    .I1(_04581_),
    .S(_04607_),
    .Z(_00182_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09198_ (.I0(\dp.rf.rf[14][28] ),
    .I1(_04582_),
    .S(_04607_),
    .Z(_00183_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09199_ (.I0(\dp.rf.rf[14][29] ),
    .I1(_04583_),
    .S(_04607_),
    .Z(_00184_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09200_ (.I0(\dp.rf.rf[14][2] ),
    .I1(_04584_),
    .S(_04607_),
    .Z(_00185_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09201_ (.I0(\dp.rf.rf[14][30] ),
    .I1(_04585_),
    .S(_04607_),
    .Z(_00186_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09202_ (.A1(_04550_),
    .A2(_04605_),
    .Z(_04608_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09203_ (.A1(\dp.rf.rf[14][31] ),
    .A2(_04605_),
    .ZN(_04609_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09204_ (.A1(_04472_),
    .A2(_04608_),
    .B(_04609_),
    .ZN(_00187_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09205_ (.I0(\dp.rf.rf[14][3] ),
    .I1(_04588_),
    .S(_04607_),
    .Z(_00188_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09206_ (.I0(\dp.rf.rf[14][4] ),
    .I1(_04589_),
    .S(_04607_),
    .Z(_00189_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09207_ (.I0(\dp.rf.rf[14][5] ),
    .I1(_04590_),
    .S(_04607_),
    .Z(_00190_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09208_ (.I0(\dp.rf.rf[14][6] ),
    .I1(_04591_),
    .S(_04607_),
    .Z(_00191_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09209_ (.I0(\dp.rf.rf[14][7] ),
    .I1(_04592_),
    .S(_04604_),
    .Z(_00192_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09210_ (.I0(\dp.rf.rf[14][8] ),
    .I1(_04593_),
    .S(_04604_),
    .Z(_00193_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09211_ (.I0(\dp.rf.rf[14][9] ),
    .I1(_04594_),
    .S(_04604_),
    .Z(_00194_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09212_ (.A1(_04545_),
    .A2(_04554_),
    .Z(_04610_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09213_ (.I(_04610_),
    .Z(_04611_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09214_ (.I0(\dp.rf.rf[15][0] ),
    .I1(_04553_),
    .S(_04611_),
    .Z(_00195_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09215_ (.I0(\dp.rf.rf[15][10] ),
    .I1(_04561_),
    .S(_04611_),
    .Z(_00196_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09216_ (.I0(\dp.rf.rf[15][11] ),
    .I1(_04562_),
    .S(_04611_),
    .Z(_00197_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09217_ (.I0(\dp.rf.rf[15][12] ),
    .I1(_04563_),
    .S(_04611_),
    .Z(_00198_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09218_ (.I0(\dp.rf.rf[15][13] ),
    .I1(_04564_),
    .S(_04611_),
    .Z(_00199_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09219_ (.I0(\dp.rf.rf[15][14] ),
    .I1(_04565_),
    .S(_04611_),
    .Z(_00200_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09220_ (.I0(\dp.rf.rf[15][15] ),
    .I1(_04566_),
    .S(_04611_),
    .Z(_00201_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09221_ (.I0(\dp.rf.rf[15][16] ),
    .I1(_04567_),
    .S(_04611_),
    .Z(_00202_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _09222_ (.I(_04610_),
    .Z(_04612_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09223_ (.I0(\dp.rf.rf[15][17] ),
    .I1(_04568_),
    .S(_04612_),
    .Z(_00203_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09224_ (.I0(\dp.rf.rf[15][18] ),
    .I1(_04570_),
    .S(_04612_),
    .Z(_00204_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09225_ (.I0(\dp.rf.rf[15][19] ),
    .I1(_04571_),
    .S(_04612_),
    .Z(_00205_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09226_ (.I0(\dp.rf.rf[15][1] ),
    .I1(_04572_),
    .S(_04612_),
    .Z(_00206_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09227_ (.I0(\dp.rf.rf[15][20] ),
    .I1(_04573_),
    .S(_04612_),
    .Z(_00207_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09228_ (.I0(\dp.rf.rf[15][21] ),
    .I1(_04574_),
    .S(_04612_),
    .Z(_00208_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09229_ (.I0(\dp.rf.rf[15][22] ),
    .I1(_04575_),
    .S(_04612_),
    .Z(_00209_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09230_ (.I0(\dp.rf.rf[15][23] ),
    .I1(_04576_),
    .S(_04612_),
    .Z(_00210_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09231_ (.I0(\dp.rf.rf[15][24] ),
    .I1(_04577_),
    .S(_04612_),
    .Z(_00211_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09232_ (.I0(\dp.rf.rf[15][25] ),
    .I1(_04578_),
    .S(_04612_),
    .Z(_00212_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09233_ (.I(_04610_),
    .Z(_04613_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09234_ (.I0(\dp.rf.rf[15][26] ),
    .I1(_04579_),
    .S(_04613_),
    .Z(_00213_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09235_ (.I0(\dp.rf.rf[15][27] ),
    .I1(_04581_),
    .S(_04613_),
    .Z(_00214_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09236_ (.I0(\dp.rf.rf[15][28] ),
    .I1(_04582_),
    .S(_04613_),
    .Z(_00215_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09237_ (.I0(\dp.rf.rf[15][29] ),
    .I1(_04583_),
    .S(_04613_),
    .Z(_00216_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09238_ (.I0(\dp.rf.rf[15][2] ),
    .I1(_04584_),
    .S(_04613_),
    .Z(_00217_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09239_ (.I0(\dp.rf.rf[15][30] ),
    .I1(_04585_),
    .S(_04613_),
    .Z(_00218_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09240_ (.A1(_04550_),
    .A2(_04611_),
    .Z(_04614_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09241_ (.A1(\dp.rf.rf[15][31] ),
    .A2(_04611_),
    .ZN(_04615_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09242_ (.A1(_04472_),
    .A2(_04614_),
    .B(_04615_),
    .ZN(_00219_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09243_ (.I0(\dp.rf.rf[15][3] ),
    .I1(_04588_),
    .S(_04613_),
    .Z(_00220_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09244_ (.I0(\dp.rf.rf[15][4] ),
    .I1(_04589_),
    .S(_04613_),
    .Z(_00221_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09245_ (.I0(\dp.rf.rf[15][5] ),
    .I1(_04590_),
    .S(_04613_),
    .Z(_00222_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09246_ (.I0(\dp.rf.rf[15][6] ),
    .I1(_04591_),
    .S(_04613_),
    .Z(_00223_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09247_ (.I0(\dp.rf.rf[15][7] ),
    .I1(_04592_),
    .S(_04610_),
    .Z(_00224_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09248_ (.I0(\dp.rf.rf[15][8] ),
    .I1(_04593_),
    .S(_04610_),
    .Z(_00225_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09249_ (.I0(\dp.rf.rf[15][9] ),
    .I1(_04594_),
    .S(_04610_),
    .Z(_00226_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09250_ (.A1(net3),
    .A2(_04555_),
    .A3(_02793_),
    .Z(_04616_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09251_ (.A1(_04558_),
    .A2(_04616_),
    .Z(_04617_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09252_ (.I(_04617_),
    .Z(_04618_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09253_ (.I0(\dp.rf.rf[16][0] ),
    .I1(_04553_),
    .S(_04618_),
    .Z(_00227_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09254_ (.I0(\dp.rf.rf[16][10] ),
    .I1(_04561_),
    .S(_04618_),
    .Z(_00228_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09255_ (.I0(\dp.rf.rf[16][11] ),
    .I1(_04562_),
    .S(_04618_),
    .Z(_00229_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09256_ (.I0(\dp.rf.rf[16][12] ),
    .I1(_04563_),
    .S(_04618_),
    .Z(_00230_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09257_ (.I0(\dp.rf.rf[16][13] ),
    .I1(_04564_),
    .S(_04618_),
    .Z(_00231_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09258_ (.I0(\dp.rf.rf[16][14] ),
    .I1(_04565_),
    .S(_04618_),
    .Z(_00232_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09259_ (.I0(\dp.rf.rf[16][15] ),
    .I1(_04566_),
    .S(_04618_),
    .Z(_00233_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09260_ (.I0(\dp.rf.rf[16][16] ),
    .I1(_04567_),
    .S(_04618_),
    .Z(_00234_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09261_ (.I(_04617_),
    .Z(_04619_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09262_ (.I0(\dp.rf.rf[16][17] ),
    .I1(_04568_),
    .S(_04619_),
    .Z(_00235_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09263_ (.I0(\dp.rf.rf[16][18] ),
    .I1(_04570_),
    .S(_04619_),
    .Z(_00236_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09264_ (.I0(\dp.rf.rf[16][19] ),
    .I1(_04571_),
    .S(_04619_),
    .Z(_00237_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09265_ (.I0(\dp.rf.rf[16][1] ),
    .I1(_04572_),
    .S(_04619_),
    .Z(_00238_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09266_ (.I0(\dp.rf.rf[16][20] ),
    .I1(_04573_),
    .S(_04619_),
    .Z(_00239_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09267_ (.I0(\dp.rf.rf[16][21] ),
    .I1(_04574_),
    .S(_04619_),
    .Z(_00240_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09268_ (.I0(\dp.rf.rf[16][22] ),
    .I1(_04575_),
    .S(_04619_),
    .Z(_00241_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09269_ (.I0(\dp.rf.rf[16][23] ),
    .I1(_04576_),
    .S(_04619_),
    .Z(_00242_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09270_ (.I0(\dp.rf.rf[16][24] ),
    .I1(_04577_),
    .S(_04619_),
    .Z(_00243_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09271_ (.I0(\dp.rf.rf[16][25] ),
    .I1(_04578_),
    .S(_04619_),
    .Z(_00244_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09272_ (.I(_04617_),
    .Z(_04620_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09273_ (.I0(\dp.rf.rf[16][26] ),
    .I1(_04579_),
    .S(_04620_),
    .Z(_00245_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09274_ (.I0(\dp.rf.rf[16][27] ),
    .I1(_04581_),
    .S(_04620_),
    .Z(_00246_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09275_ (.I0(\dp.rf.rf[16][28] ),
    .I1(_04582_),
    .S(_04620_),
    .Z(_00247_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09276_ (.I0(\dp.rf.rf[16][29] ),
    .I1(_04583_),
    .S(_04620_),
    .Z(_00248_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09277_ (.I0(\dp.rf.rf[16][2] ),
    .I1(_04584_),
    .S(_04620_),
    .Z(_00249_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09278_ (.I0(\dp.rf.rf[16][30] ),
    .I1(_04585_),
    .S(_04620_),
    .Z(_00250_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09279_ (.A1(_04550_),
    .A2(_04618_),
    .Z(_04621_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09280_ (.A1(\dp.rf.rf[16][31] ),
    .A2(_04618_),
    .ZN(_04622_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09281_ (.A1(_04472_),
    .A2(_04621_),
    .B(_04622_),
    .ZN(_00251_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09282_ (.I0(\dp.rf.rf[16][3] ),
    .I1(_04588_),
    .S(_04620_),
    .Z(_00252_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09283_ (.I0(\dp.rf.rf[16][4] ),
    .I1(_04589_),
    .S(_04620_),
    .Z(_00253_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09284_ (.I0(\dp.rf.rf[16][5] ),
    .I1(_04590_),
    .S(_04620_),
    .Z(_00254_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09285_ (.I0(\dp.rf.rf[16][6] ),
    .I1(_04591_),
    .S(_04620_),
    .Z(_00255_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09286_ (.I0(\dp.rf.rf[16][7] ),
    .I1(_04592_),
    .S(_04617_),
    .Z(_00256_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09287_ (.I0(\dp.rf.rf[16][8] ),
    .I1(_04593_),
    .S(_04617_),
    .Z(_00257_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09288_ (.I0(\dp.rf.rf[16][9] ),
    .I1(_04594_),
    .S(_04617_),
    .Z(_00258_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09289_ (.A1(_04601_),
    .A2(_04616_),
    .ZN(_04623_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09290_ (.I(_04623_),
    .Z(_04624_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09291_ (.I0(_04073_),
    .I1(\dp.rf.rf[17][0] ),
    .S(_04624_),
    .Z(_00259_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09292_ (.I0(_04120_),
    .I1(\dp.rf.rf[17][10] ),
    .S(_04624_),
    .Z(_00260_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09293_ (.I0(_04150_),
    .I1(\dp.rf.rf[17][11] ),
    .S(_04624_),
    .Z(_00261_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09294_ (.I0(_04164_),
    .I1(\dp.rf.rf[17][12] ),
    .S(_04624_),
    .Z(_00262_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09295_ (.I0(_04178_),
    .I1(\dp.rf.rf[17][13] ),
    .S(_04624_),
    .Z(_00263_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09296_ (.I0(_04196_),
    .I1(\dp.rf.rf[17][14] ),
    .S(_04624_),
    .Z(_00264_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09297_ (.I0(_04209_),
    .I1(\dp.rf.rf[17][15] ),
    .S(_04624_),
    .Z(_00265_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09298_ (.I0(_04227_),
    .I1(\dp.rf.rf[17][16] ),
    .S(_04624_),
    .Z(_00266_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09299_ (.I0(_04244_),
    .I1(\dp.rf.rf[17][17] ),
    .S(_04624_),
    .Z(_00267_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _09300_ (.I(_04623_),
    .Z(_04625_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09301_ (.I0(_04259_),
    .I1(\dp.rf.rf[17][18] ),
    .S(_04625_),
    .Z(_00268_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09302_ (.I0(_04270_),
    .I1(\dp.rf.rf[17][19] ),
    .S(_04625_),
    .Z(_00269_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09303_ (.I0(_04275_),
    .I1(\dp.rf.rf[17][1] ),
    .S(_04625_),
    .Z(_00270_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09304_ (.I0(_04292_),
    .I1(\dp.rf.rf[17][20] ),
    .S(_04625_),
    .Z(_00271_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09305_ (.I0(_04313_),
    .I1(\dp.rf.rf[17][21] ),
    .S(_04625_),
    .Z(_00272_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09306_ (.I0(_04328_),
    .I1(\dp.rf.rf[17][22] ),
    .S(_04625_),
    .Z(_00273_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09307_ (.I0(_04342_),
    .I1(\dp.rf.rf[17][23] ),
    .S(_04625_),
    .Z(_00274_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09308_ (.I0(_04359_),
    .I1(\dp.rf.rf[17][24] ),
    .S(_04625_),
    .Z(_00275_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09309_ (.I0(_04381_),
    .I1(\dp.rf.rf[17][25] ),
    .S(_04625_),
    .Z(_00276_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09310_ (.I0(_04395_),
    .I1(\dp.rf.rf[17][26] ),
    .S(_04625_),
    .Z(_00277_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09311_ (.I(_04623_),
    .Z(_04626_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09312_ (.I0(_04409_),
    .I1(\dp.rf.rf[17][27] ),
    .S(_04626_),
    .Z(_00278_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09313_ (.I0(_04421_),
    .I1(\dp.rf.rf[17][28] ),
    .S(_04626_),
    .Z(_00279_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09314_ (.I0(_04439_),
    .I1(\dp.rf.rf[17][29] ),
    .S(_04626_),
    .Z(_00280_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09315_ (.I0(_04446_),
    .I1(\dp.rf.rf[17][2] ),
    .S(_04626_),
    .Z(_00281_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09316_ (.I0(_04462_),
    .I1(\dp.rf.rf[17][30] ),
    .S(_04626_),
    .Z(_00282_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09317_ (.I(\dp.rf.rf[17][31] ),
    .ZN(_04627_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09318_ (.A1(_04482_),
    .A2(_04601_),
    .A3(_04616_),
    .Z(_04628_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09319_ (.A1(_04627_),
    .A2(_04624_),
    .B1(_04628_),
    .B2(_04603_),
    .ZN(_00283_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09320_ (.I0(_04488_),
    .I1(\dp.rf.rf[17][3] ),
    .S(_04626_),
    .Z(_00284_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09321_ (.I0(_04496_),
    .I1(\dp.rf.rf[17][4] ),
    .S(_04626_),
    .Z(_00285_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09322_ (.I0(_04504_),
    .I1(\dp.rf.rf[17][5] ),
    .S(_04626_),
    .Z(_00286_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09323_ (.I0(_04512_),
    .I1(\dp.rf.rf[17][6] ),
    .S(_04626_),
    .Z(_00287_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09324_ (.I0(_04523_),
    .I1(\dp.rf.rf[17][7] ),
    .S(_04626_),
    .Z(_00288_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09325_ (.I0(_04534_),
    .I1(\dp.rf.rf[17][8] ),
    .S(_04623_),
    .Z(_00289_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09326_ (.I0(_04544_),
    .I1(\dp.rf.rf[17][9] ),
    .S(_04623_),
    .Z(_00290_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09327_ (.A1(_04081_),
    .A2(_04616_),
    .Z(_04629_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09328_ (.I(_04629_),
    .Z(_04630_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09329_ (.I0(\dp.rf.rf[18][0] ),
    .I1(_04553_),
    .S(_04630_),
    .Z(_00291_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09330_ (.I0(\dp.rf.rf[18][10] ),
    .I1(_04561_),
    .S(_04630_),
    .Z(_00292_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09331_ (.I0(\dp.rf.rf[18][11] ),
    .I1(_04562_),
    .S(_04630_),
    .Z(_00293_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09332_ (.I0(\dp.rf.rf[18][12] ),
    .I1(_04563_),
    .S(_04630_),
    .Z(_00294_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09333_ (.I0(\dp.rf.rf[18][13] ),
    .I1(_04564_),
    .S(_04630_),
    .Z(_00295_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09334_ (.I0(\dp.rf.rf[18][14] ),
    .I1(_04565_),
    .S(_04630_),
    .Z(_00296_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09335_ (.I0(\dp.rf.rf[18][15] ),
    .I1(_04566_),
    .S(_04630_),
    .Z(_00297_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09336_ (.I0(\dp.rf.rf[18][16] ),
    .I1(_04567_),
    .S(_04630_),
    .Z(_00298_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09337_ (.I(_04629_),
    .Z(_04631_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09338_ (.I0(\dp.rf.rf[18][17] ),
    .I1(_04568_),
    .S(_04631_),
    .Z(_00299_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09339_ (.I0(\dp.rf.rf[18][18] ),
    .I1(_04570_),
    .S(_04631_),
    .Z(_00300_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09340_ (.I0(\dp.rf.rf[18][19] ),
    .I1(_04571_),
    .S(_04631_),
    .Z(_00301_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09341_ (.I0(\dp.rf.rf[18][1] ),
    .I1(_04572_),
    .S(_04631_),
    .Z(_00302_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09342_ (.I0(\dp.rf.rf[18][20] ),
    .I1(_04573_),
    .S(_04631_),
    .Z(_00303_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09343_ (.I0(\dp.rf.rf[18][21] ),
    .I1(_04574_),
    .S(_04631_),
    .Z(_00304_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09344_ (.I0(\dp.rf.rf[18][22] ),
    .I1(_04575_),
    .S(_04631_),
    .Z(_00305_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09345_ (.I0(\dp.rf.rf[18][23] ),
    .I1(_04576_),
    .S(_04631_),
    .Z(_00306_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09346_ (.I0(\dp.rf.rf[18][24] ),
    .I1(_04577_),
    .S(_04631_),
    .Z(_00307_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09347_ (.I0(\dp.rf.rf[18][25] ),
    .I1(_04578_),
    .S(_04631_),
    .Z(_00308_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09348_ (.I(_04629_),
    .Z(_04632_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09349_ (.I0(\dp.rf.rf[18][26] ),
    .I1(_04579_),
    .S(_04632_),
    .Z(_00309_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09350_ (.I0(\dp.rf.rf[18][27] ),
    .I1(_04581_),
    .S(_04632_),
    .Z(_00310_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09351_ (.I0(\dp.rf.rf[18][28] ),
    .I1(_04582_),
    .S(_04632_),
    .Z(_00311_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09352_ (.I0(\dp.rf.rf[18][29] ),
    .I1(_04583_),
    .S(_04632_),
    .Z(_00312_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09353_ (.I0(\dp.rf.rf[18][2] ),
    .I1(_04584_),
    .S(_04632_),
    .Z(_00313_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09354_ (.I0(\dp.rf.rf[18][30] ),
    .I1(_04585_),
    .S(_04632_),
    .Z(_00314_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09355_ (.A1(_04550_),
    .A2(_04630_),
    .Z(_04633_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09356_ (.A1(\dp.rf.rf[18][31] ),
    .A2(_04630_),
    .ZN(_04634_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09357_ (.A1(_04472_),
    .A2(_04633_),
    .B(_04634_),
    .ZN(_00315_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09358_ (.I0(\dp.rf.rf[18][3] ),
    .I1(_04588_),
    .S(_04632_),
    .Z(_00316_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09359_ (.I0(\dp.rf.rf[18][4] ),
    .I1(_04589_),
    .S(_04632_),
    .Z(_00317_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09360_ (.I0(\dp.rf.rf[18][5] ),
    .I1(_04590_),
    .S(_04632_),
    .Z(_00318_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09361_ (.I0(\dp.rf.rf[18][6] ),
    .I1(_04591_),
    .S(_04632_),
    .Z(_00319_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09362_ (.I0(\dp.rf.rf[18][7] ),
    .I1(_04592_),
    .S(_04629_),
    .Z(_00320_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09363_ (.I0(\dp.rf.rf[18][8] ),
    .I1(_04593_),
    .S(_04629_),
    .Z(_00321_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09364_ (.I0(\dp.rf.rf[18][9] ),
    .I1(_04594_),
    .S(_04629_),
    .Z(_00322_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09365_ (.A1(_04545_),
    .A2(_04616_),
    .Z(_04635_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09366_ (.I(_04635_),
    .Z(_04636_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09367_ (.I0(\dp.rf.rf[19][0] ),
    .I1(_04553_),
    .S(_04636_),
    .Z(_00323_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09368_ (.I0(\dp.rf.rf[19][10] ),
    .I1(_04561_),
    .S(_04636_),
    .Z(_00324_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09369_ (.I0(\dp.rf.rf[19][11] ),
    .I1(_04562_),
    .S(_04636_),
    .Z(_00325_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09370_ (.I0(\dp.rf.rf[19][12] ),
    .I1(_04563_),
    .S(_04636_),
    .Z(_00326_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09371_ (.I0(\dp.rf.rf[19][13] ),
    .I1(_04564_),
    .S(_04636_),
    .Z(_00327_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09372_ (.I0(\dp.rf.rf[19][14] ),
    .I1(_04565_),
    .S(_04636_),
    .Z(_00328_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09373_ (.I0(\dp.rf.rf[19][15] ),
    .I1(_04566_),
    .S(_04636_),
    .Z(_00329_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09374_ (.I0(\dp.rf.rf[19][16] ),
    .I1(_04567_),
    .S(_04636_),
    .Z(_00330_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09375_ (.I(_04635_),
    .Z(_04637_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09376_ (.I0(\dp.rf.rf[19][17] ),
    .I1(_04568_),
    .S(_04637_),
    .Z(_00331_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09377_ (.I0(\dp.rf.rf[19][18] ),
    .I1(_04570_),
    .S(_04637_),
    .Z(_00332_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09378_ (.I0(\dp.rf.rf[19][19] ),
    .I1(_04571_),
    .S(_04637_),
    .Z(_00333_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09379_ (.I0(\dp.rf.rf[19][1] ),
    .I1(_04572_),
    .S(_04637_),
    .Z(_00334_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09380_ (.I0(\dp.rf.rf[19][20] ),
    .I1(_04573_),
    .S(_04637_),
    .Z(_00335_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09381_ (.I0(\dp.rf.rf[19][21] ),
    .I1(_04574_),
    .S(_04637_),
    .Z(_00336_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09382_ (.I0(\dp.rf.rf[19][22] ),
    .I1(_04575_),
    .S(_04637_),
    .Z(_00337_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09383_ (.I0(\dp.rf.rf[19][23] ),
    .I1(_04576_),
    .S(_04637_),
    .Z(_00338_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09384_ (.I0(\dp.rf.rf[19][24] ),
    .I1(_04577_),
    .S(_04637_),
    .Z(_00339_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09385_ (.I0(\dp.rf.rf[19][25] ),
    .I1(_04578_),
    .S(_04637_),
    .Z(_00340_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09386_ (.I(_04635_),
    .Z(_04638_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09387_ (.I0(\dp.rf.rf[19][26] ),
    .I1(_04579_),
    .S(_04638_),
    .Z(_00341_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09388_ (.I0(\dp.rf.rf[19][27] ),
    .I1(_04581_),
    .S(_04638_),
    .Z(_00342_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09389_ (.I0(\dp.rf.rf[19][28] ),
    .I1(_04582_),
    .S(_04638_),
    .Z(_00343_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09390_ (.I0(\dp.rf.rf[19][29] ),
    .I1(_04583_),
    .S(_04638_),
    .Z(_00344_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09391_ (.I0(\dp.rf.rf[19][2] ),
    .I1(_04584_),
    .S(_04638_),
    .Z(_00345_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09392_ (.I0(\dp.rf.rf[19][30] ),
    .I1(_04585_),
    .S(_04638_),
    .Z(_00346_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09393_ (.A1(_04550_),
    .A2(_04636_),
    .Z(_04639_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09394_ (.A1(\dp.rf.rf[19][31] ),
    .A2(_04636_),
    .ZN(_04640_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09395_ (.A1(_04472_),
    .A2(_04639_),
    .B(_04640_),
    .ZN(_00347_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09396_ (.I0(\dp.rf.rf[19][3] ),
    .I1(_04588_),
    .S(_04638_),
    .Z(_00348_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09397_ (.I0(\dp.rf.rf[19][4] ),
    .I1(_04589_),
    .S(_04638_),
    .Z(_00349_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09398_ (.I0(\dp.rf.rf[19][5] ),
    .I1(_04590_),
    .S(_04638_),
    .Z(_00350_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09399_ (.I0(\dp.rf.rf[19][6] ),
    .I1(_04591_),
    .S(_04638_),
    .Z(_00351_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09400_ (.I0(\dp.rf.rf[19][7] ),
    .I1(_04592_),
    .S(_04635_),
    .Z(_00352_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09401_ (.I0(\dp.rf.rf[19][8] ),
    .I1(_04593_),
    .S(_04635_),
    .Z(_00353_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09402_ (.I0(\dp.rf.rf[19][9] ),
    .I1(_04594_),
    .S(_04635_),
    .Z(_00354_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09403_ (.A1(_04556_),
    .A2(_04595_),
    .ZN(_04641_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09404_ (.I(_04641_),
    .Z(_04642_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09405_ (.I0(_04073_),
    .I1(\dp.rf.rf[1][0] ),
    .S(_04642_),
    .Z(_00355_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09406_ (.I0(_04120_),
    .I1(\dp.rf.rf[1][10] ),
    .S(_04642_),
    .Z(_00356_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09407_ (.I0(_04150_),
    .I1(\dp.rf.rf[1][11] ),
    .S(_04642_),
    .Z(_00357_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09408_ (.I0(_04164_),
    .I1(\dp.rf.rf[1][12] ),
    .S(_04642_),
    .Z(_00358_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09409_ (.I0(_04178_),
    .I1(\dp.rf.rf[1][13] ),
    .S(_04642_),
    .Z(_00359_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09410_ (.I0(_04196_),
    .I1(\dp.rf.rf[1][14] ),
    .S(_04642_),
    .Z(_00360_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09411_ (.I0(_04209_),
    .I1(\dp.rf.rf[1][15] ),
    .S(_04642_),
    .Z(_00361_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09412_ (.I0(_04227_),
    .I1(\dp.rf.rf[1][16] ),
    .S(_04642_),
    .Z(_00362_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09413_ (.I0(_04244_),
    .I1(\dp.rf.rf[1][17] ),
    .S(_04642_),
    .Z(_00363_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09414_ (.I(_04641_),
    .Z(_04643_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09415_ (.I0(_04259_),
    .I1(\dp.rf.rf[1][18] ),
    .S(_04643_),
    .Z(_00364_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09416_ (.I0(_04270_),
    .I1(\dp.rf.rf[1][19] ),
    .S(_04643_),
    .Z(_00365_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09417_ (.I0(_04275_),
    .I1(\dp.rf.rf[1][1] ),
    .S(_04643_),
    .Z(_00366_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09418_ (.I0(_04292_),
    .I1(\dp.rf.rf[1][20] ),
    .S(_04643_),
    .Z(_00367_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09419_ (.I0(_04313_),
    .I1(\dp.rf.rf[1][21] ),
    .S(_04643_),
    .Z(_00368_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09420_ (.I0(_04328_),
    .I1(\dp.rf.rf[1][22] ),
    .S(_04643_),
    .Z(_00369_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09421_ (.I0(_04342_),
    .I1(\dp.rf.rf[1][23] ),
    .S(_04643_),
    .Z(_00370_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09422_ (.I0(_04359_),
    .I1(\dp.rf.rf[1][24] ),
    .S(_04643_),
    .Z(_00371_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09423_ (.I0(_04381_),
    .I1(\dp.rf.rf[1][25] ),
    .S(_04643_),
    .Z(_00372_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09424_ (.I0(_04395_),
    .I1(\dp.rf.rf[1][26] ),
    .S(_04643_),
    .Z(_00373_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09425_ (.I(_04641_),
    .Z(_04644_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09426_ (.I0(_04409_),
    .I1(\dp.rf.rf[1][27] ),
    .S(_04644_),
    .Z(_00374_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09427_ (.I0(_04421_),
    .I1(\dp.rf.rf[1][28] ),
    .S(_04644_),
    .Z(_00375_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09428_ (.I0(_04439_),
    .I1(\dp.rf.rf[1][29] ),
    .S(_04644_),
    .Z(_00376_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09429_ (.I0(_04446_),
    .I1(\dp.rf.rf[1][2] ),
    .S(_04644_),
    .Z(_00377_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09430_ (.I0(_04462_),
    .I1(\dp.rf.rf[1][30] ),
    .S(_04644_),
    .Z(_00378_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09431_ (.I(\dp.rf.rf[1][31] ),
    .ZN(_04645_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09432_ (.A1(_04482_),
    .A2(_04556_),
    .A3(_04601_),
    .Z(_04646_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09433_ (.A1(_04645_),
    .A2(_04642_),
    .B1(_04646_),
    .B2(_04603_),
    .ZN(_00379_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09434_ (.I0(_04488_),
    .I1(\dp.rf.rf[1][3] ),
    .S(_04644_),
    .Z(_00380_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09435_ (.I0(_04496_),
    .I1(\dp.rf.rf[1][4] ),
    .S(_04644_),
    .Z(_00381_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09436_ (.I0(_04504_),
    .I1(\dp.rf.rf[1][5] ),
    .S(_04644_),
    .Z(_00382_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09437_ (.I0(_04512_),
    .I1(\dp.rf.rf[1][6] ),
    .S(_04644_),
    .Z(_00383_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09438_ (.I0(_04523_),
    .I1(\dp.rf.rf[1][7] ),
    .S(_04644_),
    .Z(_00384_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09439_ (.I0(_04534_),
    .I1(\dp.rf.rf[1][8] ),
    .S(_04641_),
    .Z(_00385_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09440_ (.I0(_04544_),
    .I1(\dp.rf.rf[1][9] ),
    .S(_04641_),
    .Z(_00386_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09441_ (.A1(net3),
    .A2(_04555_),
    .A3(net27),
    .Z(_04647_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09442_ (.A1(_04558_),
    .A2(_04647_),
    .Z(_04648_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09443_ (.I(_04648_),
    .Z(_04649_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09444_ (.I0(\dp.rf.rf[20][0] ),
    .I1(_04553_),
    .S(_04649_),
    .Z(_00387_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09445_ (.I0(\dp.rf.rf[20][10] ),
    .I1(_04561_),
    .S(_04649_),
    .Z(_00388_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09446_ (.I0(\dp.rf.rf[20][11] ),
    .I1(_04562_),
    .S(_04649_),
    .Z(_00389_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09447_ (.I0(\dp.rf.rf[20][12] ),
    .I1(_04563_),
    .S(_04649_),
    .Z(_00390_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09448_ (.I0(\dp.rf.rf[20][13] ),
    .I1(_04564_),
    .S(_04649_),
    .Z(_00391_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09449_ (.I0(\dp.rf.rf[20][14] ),
    .I1(_04565_),
    .S(_04649_),
    .Z(_00392_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09450_ (.I0(\dp.rf.rf[20][15] ),
    .I1(_04566_),
    .S(_04649_),
    .Z(_00393_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09451_ (.I0(\dp.rf.rf[20][16] ),
    .I1(_04567_),
    .S(_04649_),
    .Z(_00394_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09452_ (.I(_04648_),
    .Z(_04650_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09453_ (.I0(\dp.rf.rf[20][17] ),
    .I1(_04568_),
    .S(_04650_),
    .Z(_00395_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09454_ (.I0(\dp.rf.rf[20][18] ),
    .I1(_04570_),
    .S(_04650_),
    .Z(_00396_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09455_ (.I0(\dp.rf.rf[20][19] ),
    .I1(_04571_),
    .S(_04650_),
    .Z(_00397_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09456_ (.I0(\dp.rf.rf[20][1] ),
    .I1(_04572_),
    .S(_04650_),
    .Z(_00398_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09457_ (.I0(\dp.rf.rf[20][20] ),
    .I1(_04573_),
    .S(_04650_),
    .Z(_00399_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09458_ (.I0(\dp.rf.rf[20][21] ),
    .I1(_04574_),
    .S(_04650_),
    .Z(_00400_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09459_ (.I0(\dp.rf.rf[20][22] ),
    .I1(_04575_),
    .S(_04650_),
    .Z(_00401_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09460_ (.I0(\dp.rf.rf[20][23] ),
    .I1(_04576_),
    .S(_04650_),
    .Z(_00402_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09461_ (.I0(\dp.rf.rf[20][24] ),
    .I1(_04577_),
    .S(_04650_),
    .Z(_00403_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09462_ (.I0(\dp.rf.rf[20][25] ),
    .I1(_04578_),
    .S(_04650_),
    .Z(_00404_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09463_ (.I(_04648_),
    .Z(_04651_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09464_ (.I0(\dp.rf.rf[20][26] ),
    .I1(_04579_),
    .S(_04651_),
    .Z(_00405_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09465_ (.I0(\dp.rf.rf[20][27] ),
    .I1(_04581_),
    .S(_04651_),
    .Z(_00406_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09466_ (.I0(\dp.rf.rf[20][28] ),
    .I1(_04582_),
    .S(_04651_),
    .Z(_00407_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09467_ (.I0(\dp.rf.rf[20][29] ),
    .I1(_04583_),
    .S(_04651_),
    .Z(_00408_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09468_ (.I0(\dp.rf.rf[20][2] ),
    .I1(_04584_),
    .S(_04651_),
    .Z(_00409_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09469_ (.I0(\dp.rf.rf[20][30] ),
    .I1(_04585_),
    .S(_04651_),
    .Z(_00410_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09470_ (.A1(_04550_),
    .A2(_04649_),
    .Z(_04652_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09471_ (.A1(\dp.rf.rf[20][31] ),
    .A2(_04649_),
    .ZN(_04653_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09472_ (.A1(_04472_),
    .A2(_04652_),
    .B(_04653_),
    .ZN(_00411_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09473_ (.I0(\dp.rf.rf[20][3] ),
    .I1(_04588_),
    .S(_04651_),
    .Z(_00412_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09474_ (.I0(\dp.rf.rf[20][4] ),
    .I1(_04589_),
    .S(_04651_),
    .Z(_00413_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09475_ (.I0(\dp.rf.rf[20][5] ),
    .I1(_04590_),
    .S(_04651_),
    .Z(_00414_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09476_ (.I0(\dp.rf.rf[20][6] ),
    .I1(_04591_),
    .S(_04651_),
    .Z(_00415_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09477_ (.I0(\dp.rf.rf[20][7] ),
    .I1(_04592_),
    .S(_04648_),
    .Z(_00416_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09478_ (.I0(\dp.rf.rf[20][8] ),
    .I1(_04593_),
    .S(_04648_),
    .Z(_00417_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09479_ (.I0(\dp.rf.rf[20][9] ),
    .I1(_04594_),
    .S(_04648_),
    .Z(_00418_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09480_ (.A1(_04601_),
    .A2(_04647_),
    .ZN(_04654_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09481_ (.I(_04654_),
    .Z(_04655_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09482_ (.I0(_04073_),
    .I1(\dp.rf.rf[21][0] ),
    .S(_04655_),
    .Z(_00419_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09483_ (.I0(_04120_),
    .I1(\dp.rf.rf[21][10] ),
    .S(_04655_),
    .Z(_00420_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09484_ (.I0(_04150_),
    .I1(\dp.rf.rf[21][11] ),
    .S(_04655_),
    .Z(_00421_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09485_ (.I0(_04164_),
    .I1(\dp.rf.rf[21][12] ),
    .S(_04655_),
    .Z(_00422_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09486_ (.I0(_04178_),
    .I1(\dp.rf.rf[21][13] ),
    .S(_04655_),
    .Z(_00423_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09487_ (.I0(_04196_),
    .I1(\dp.rf.rf[21][14] ),
    .S(_04655_),
    .Z(_00424_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09488_ (.I0(_04209_),
    .I1(\dp.rf.rf[21][15] ),
    .S(_04655_),
    .Z(_00425_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09489_ (.I0(_04227_),
    .I1(\dp.rf.rf[21][16] ),
    .S(_04655_),
    .Z(_00426_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09490_ (.I0(_04244_),
    .I1(\dp.rf.rf[21][17] ),
    .S(_04655_),
    .Z(_00427_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09491_ (.I(_04654_),
    .Z(_04656_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09492_ (.I0(_04259_),
    .I1(\dp.rf.rf[21][18] ),
    .S(_04656_),
    .Z(_00428_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09493_ (.I0(_04270_),
    .I1(\dp.rf.rf[21][19] ),
    .S(_04656_),
    .Z(_00429_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09494_ (.I0(_04275_),
    .I1(\dp.rf.rf[21][1] ),
    .S(_04656_),
    .Z(_00430_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09495_ (.I0(_04292_),
    .I1(\dp.rf.rf[21][20] ),
    .S(_04656_),
    .Z(_00431_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09496_ (.I0(_04313_),
    .I1(\dp.rf.rf[21][21] ),
    .S(_04656_),
    .Z(_00432_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09497_ (.I0(_04328_),
    .I1(\dp.rf.rf[21][22] ),
    .S(_04656_),
    .Z(_00433_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09498_ (.I0(_04342_),
    .I1(\dp.rf.rf[21][23] ),
    .S(_04656_),
    .Z(_00434_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09499_ (.I0(_04359_),
    .I1(\dp.rf.rf[21][24] ),
    .S(_04656_),
    .Z(_00435_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09500_ (.I0(_04381_),
    .I1(\dp.rf.rf[21][25] ),
    .S(_04656_),
    .Z(_00436_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09501_ (.I0(_04395_),
    .I1(\dp.rf.rf[21][26] ),
    .S(_04656_),
    .Z(_00437_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09502_ (.I(_04654_),
    .Z(_04657_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09503_ (.I0(_04409_),
    .I1(\dp.rf.rf[21][27] ),
    .S(_04657_),
    .Z(_00438_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09504_ (.I0(_04421_),
    .I1(\dp.rf.rf[21][28] ),
    .S(_04657_),
    .Z(_00439_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09505_ (.I0(_04439_),
    .I1(\dp.rf.rf[21][29] ),
    .S(_04657_),
    .Z(_00440_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09506_ (.I0(_04446_),
    .I1(\dp.rf.rf[21][2] ),
    .S(_04657_),
    .Z(_00441_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09507_ (.I0(_04462_),
    .I1(\dp.rf.rf[21][30] ),
    .S(_04657_),
    .Z(_00442_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09508_ (.I(\dp.rf.rf[21][31] ),
    .ZN(_04658_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09509_ (.A1(_04482_),
    .A2(_04601_),
    .A3(_04647_),
    .Z(_04659_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09510_ (.A1(_04658_),
    .A2(_04655_),
    .B1(_04659_),
    .B2(_04603_),
    .ZN(_00443_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09511_ (.I0(_04488_),
    .I1(\dp.rf.rf[21][3] ),
    .S(_04657_),
    .Z(_00444_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09512_ (.I0(_04496_),
    .I1(\dp.rf.rf[21][4] ),
    .S(_04657_),
    .Z(_00445_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09513_ (.I0(_04504_),
    .I1(\dp.rf.rf[21][5] ),
    .S(_04657_),
    .Z(_00446_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09514_ (.I0(_04512_),
    .I1(\dp.rf.rf[21][6] ),
    .S(_04657_),
    .Z(_00447_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09515_ (.I0(_04523_),
    .I1(\dp.rf.rf[21][7] ),
    .S(_04657_),
    .Z(_00448_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09516_ (.I0(_04534_),
    .I1(\dp.rf.rf[21][8] ),
    .S(_04654_),
    .Z(_00449_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09517_ (.I0(_04544_),
    .I1(\dp.rf.rf[21][9] ),
    .S(_04654_),
    .Z(_00450_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09518_ (.A1(_04081_),
    .A2(_04647_),
    .Z(_04660_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09519_ (.I(_04660_),
    .Z(_04661_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09520_ (.I0(\dp.rf.rf[22][0] ),
    .I1(_04553_),
    .S(_04661_),
    .Z(_00451_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09521_ (.I0(\dp.rf.rf[22][10] ),
    .I1(_04561_),
    .S(_04661_),
    .Z(_00452_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09522_ (.I0(\dp.rf.rf[22][11] ),
    .I1(_04562_),
    .S(_04661_),
    .Z(_00453_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09523_ (.I0(\dp.rf.rf[22][12] ),
    .I1(_04563_),
    .S(_04661_),
    .Z(_00454_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09524_ (.I0(\dp.rf.rf[22][13] ),
    .I1(_04564_),
    .S(_04661_),
    .Z(_00455_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09525_ (.I0(\dp.rf.rf[22][14] ),
    .I1(_04565_),
    .S(_04661_),
    .Z(_00456_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09526_ (.I0(\dp.rf.rf[22][15] ),
    .I1(_04566_),
    .S(_04661_),
    .Z(_00457_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09527_ (.I0(\dp.rf.rf[22][16] ),
    .I1(_04567_),
    .S(_04661_),
    .Z(_00458_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09528_ (.I(_04660_),
    .Z(_04662_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09529_ (.I0(\dp.rf.rf[22][17] ),
    .I1(_04568_),
    .S(_04662_),
    .Z(_00459_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09530_ (.I0(\dp.rf.rf[22][18] ),
    .I1(_04570_),
    .S(_04662_),
    .Z(_00460_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09531_ (.I0(\dp.rf.rf[22][19] ),
    .I1(_04571_),
    .S(_04662_),
    .Z(_00461_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09532_ (.I0(\dp.rf.rf[22][1] ),
    .I1(_04572_),
    .S(_04662_),
    .Z(_00462_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09533_ (.I0(\dp.rf.rf[22][20] ),
    .I1(_04573_),
    .S(_04662_),
    .Z(_00463_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09534_ (.I0(\dp.rf.rf[22][21] ),
    .I1(_04574_),
    .S(_04662_),
    .Z(_00464_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09535_ (.I0(\dp.rf.rf[22][22] ),
    .I1(_04575_),
    .S(_04662_),
    .Z(_00465_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09536_ (.I0(\dp.rf.rf[22][23] ),
    .I1(_04576_),
    .S(_04662_),
    .Z(_00466_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09537_ (.I0(\dp.rf.rf[22][24] ),
    .I1(_04577_),
    .S(_04662_),
    .Z(_00467_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09538_ (.I0(\dp.rf.rf[22][25] ),
    .I1(_04578_),
    .S(_04662_),
    .Z(_00468_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09539_ (.I(_04660_),
    .Z(_04663_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09540_ (.I0(\dp.rf.rf[22][26] ),
    .I1(_04579_),
    .S(_04663_),
    .Z(_00469_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09541_ (.I0(\dp.rf.rf[22][27] ),
    .I1(_04581_),
    .S(_04663_),
    .Z(_00470_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09542_ (.I0(\dp.rf.rf[22][28] ),
    .I1(_04582_),
    .S(_04663_),
    .Z(_00471_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09543_ (.I0(\dp.rf.rf[22][29] ),
    .I1(_04583_),
    .S(_04663_),
    .Z(_00472_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09544_ (.I0(\dp.rf.rf[22][2] ),
    .I1(_04584_),
    .S(_04663_),
    .Z(_00473_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09545_ (.I0(\dp.rf.rf[22][30] ),
    .I1(_04585_),
    .S(_04663_),
    .Z(_00474_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09546_ (.A1(_04550_),
    .A2(_04661_),
    .Z(_04664_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09547_ (.A1(\dp.rf.rf[22][31] ),
    .A2(_04661_),
    .ZN(_04665_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09548_ (.A1(_04472_),
    .A2(_04664_),
    .B(_04665_),
    .ZN(_00475_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09549_ (.I0(\dp.rf.rf[22][3] ),
    .I1(_04588_),
    .S(_04663_),
    .Z(_00476_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09550_ (.I0(\dp.rf.rf[22][4] ),
    .I1(_04589_),
    .S(_04663_),
    .Z(_00477_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09551_ (.I0(\dp.rf.rf[22][5] ),
    .I1(_04590_),
    .S(_04663_),
    .Z(_00478_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09552_ (.I0(\dp.rf.rf[22][6] ),
    .I1(_04591_),
    .S(_04663_),
    .Z(_00479_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09553_ (.I0(\dp.rf.rf[22][7] ),
    .I1(_04592_),
    .S(_04660_),
    .Z(_00480_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09554_ (.I0(\dp.rf.rf[22][8] ),
    .I1(_04593_),
    .S(_04660_),
    .Z(_00481_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09555_ (.I0(\dp.rf.rf[22][9] ),
    .I1(_04594_),
    .S(_04660_),
    .Z(_00482_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09556_ (.A1(_04545_),
    .A2(_04647_),
    .Z(_04666_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09557_ (.I(_04666_),
    .Z(_04667_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09558_ (.I0(\dp.rf.rf[23][0] ),
    .I1(_04553_),
    .S(_04667_),
    .Z(_00483_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09559_ (.I0(\dp.rf.rf[23][10] ),
    .I1(_04561_),
    .S(_04667_),
    .Z(_00484_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09560_ (.I0(\dp.rf.rf[23][11] ),
    .I1(_04562_),
    .S(_04667_),
    .Z(_00485_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09561_ (.I0(\dp.rf.rf[23][12] ),
    .I1(_04563_),
    .S(_04667_),
    .Z(_00486_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09562_ (.I0(\dp.rf.rf[23][13] ),
    .I1(_04564_),
    .S(_04667_),
    .Z(_00487_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09563_ (.I0(\dp.rf.rf[23][14] ),
    .I1(_04565_),
    .S(_04667_),
    .Z(_00488_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09564_ (.I0(\dp.rf.rf[23][15] ),
    .I1(_04566_),
    .S(_04667_),
    .Z(_00489_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09565_ (.I0(\dp.rf.rf[23][16] ),
    .I1(_04567_),
    .S(_04667_),
    .Z(_00490_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09566_ (.I(_04666_),
    .Z(_04668_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09567_ (.I0(\dp.rf.rf[23][17] ),
    .I1(_04568_),
    .S(_04668_),
    .Z(_00491_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09568_ (.I0(\dp.rf.rf[23][18] ),
    .I1(_04570_),
    .S(_04668_),
    .Z(_00492_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09569_ (.I0(\dp.rf.rf[23][19] ),
    .I1(_04571_),
    .S(_04668_),
    .Z(_00493_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09570_ (.I0(\dp.rf.rf[23][1] ),
    .I1(_04572_),
    .S(_04668_),
    .Z(_00494_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09571_ (.I0(\dp.rf.rf[23][20] ),
    .I1(_04573_),
    .S(_04668_),
    .Z(_00495_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09572_ (.I0(\dp.rf.rf[23][21] ),
    .I1(_04574_),
    .S(_04668_),
    .Z(_00496_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09573_ (.I0(\dp.rf.rf[23][22] ),
    .I1(_04575_),
    .S(_04668_),
    .Z(_00497_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09574_ (.I0(\dp.rf.rf[23][23] ),
    .I1(_04576_),
    .S(_04668_),
    .Z(_00498_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09575_ (.I0(\dp.rf.rf[23][24] ),
    .I1(_04577_),
    .S(_04668_),
    .Z(_00499_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09576_ (.I0(\dp.rf.rf[23][25] ),
    .I1(_04578_),
    .S(_04668_),
    .Z(_00500_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09577_ (.I(_04666_),
    .Z(_04669_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09578_ (.I0(\dp.rf.rf[23][26] ),
    .I1(_04579_),
    .S(_04669_),
    .Z(_00501_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09579_ (.I0(\dp.rf.rf[23][27] ),
    .I1(_04581_),
    .S(_04669_),
    .Z(_00502_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09580_ (.I0(\dp.rf.rf[23][28] ),
    .I1(_04582_),
    .S(_04669_),
    .Z(_00503_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09581_ (.I0(\dp.rf.rf[23][29] ),
    .I1(_04583_),
    .S(_04669_),
    .Z(_00504_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09582_ (.I0(\dp.rf.rf[23][2] ),
    .I1(_04584_),
    .S(_04669_),
    .Z(_00505_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09583_ (.I0(\dp.rf.rf[23][30] ),
    .I1(_04585_),
    .S(_04669_),
    .Z(_00506_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _09584_ (.I(_04471_),
    .Z(_04670_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09585_ (.A1(_04550_),
    .A2(_04667_),
    .Z(_04671_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09586_ (.A1(\dp.rf.rf[23][31] ),
    .A2(_04667_),
    .ZN(_04672_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09587_ (.A1(_04670_),
    .A2(_04671_),
    .B(_04672_),
    .ZN(_00507_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09588_ (.I0(\dp.rf.rf[23][3] ),
    .I1(_04588_),
    .S(_04669_),
    .Z(_00508_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09589_ (.I0(\dp.rf.rf[23][4] ),
    .I1(_04589_),
    .S(_04669_),
    .Z(_00509_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09590_ (.I0(\dp.rf.rf[23][5] ),
    .I1(_04590_),
    .S(_04669_),
    .Z(_00510_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09591_ (.I0(\dp.rf.rf[23][6] ),
    .I1(_04591_),
    .S(_04669_),
    .Z(_00511_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09592_ (.I0(\dp.rf.rf[23][7] ),
    .I1(_04592_),
    .S(_04666_),
    .Z(_00512_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09593_ (.I0(\dp.rf.rf[23][8] ),
    .I1(_04593_),
    .S(_04666_),
    .Z(_00513_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09594_ (.I0(\dp.rf.rf[23][9] ),
    .I1(_04594_),
    .S(_04666_),
    .Z(_00514_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09595_ (.A1(net3),
    .A2(net2),
    .A3(_02793_),
    .Z(_04673_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09596_ (.A1(_04558_),
    .A2(_04673_),
    .Z(_04674_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09597_ (.I(_04674_),
    .Z(_04675_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09598_ (.I0(\dp.rf.rf[24][0] ),
    .I1(_04553_),
    .S(_04675_),
    .Z(_00515_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09599_ (.I0(\dp.rf.rf[24][10] ),
    .I1(_04561_),
    .S(_04675_),
    .Z(_00516_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09600_ (.I0(\dp.rf.rf[24][11] ),
    .I1(_04562_),
    .S(_04675_),
    .Z(_00517_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09601_ (.I0(\dp.rf.rf[24][12] ),
    .I1(_04563_),
    .S(_04675_),
    .Z(_00518_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09602_ (.I0(\dp.rf.rf[24][13] ),
    .I1(_04564_),
    .S(_04675_),
    .Z(_00519_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09603_ (.I0(\dp.rf.rf[24][14] ),
    .I1(_04565_),
    .S(_04675_),
    .Z(_00520_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09604_ (.I0(\dp.rf.rf[24][15] ),
    .I1(_04566_),
    .S(_04675_),
    .Z(_00521_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09605_ (.I0(\dp.rf.rf[24][16] ),
    .I1(_04567_),
    .S(_04675_),
    .Z(_00522_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09606_ (.I(_04674_),
    .Z(_04676_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09607_ (.I0(\dp.rf.rf[24][17] ),
    .I1(_04568_),
    .S(_04676_),
    .Z(_00523_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09608_ (.I0(\dp.rf.rf[24][18] ),
    .I1(_04570_),
    .S(_04676_),
    .Z(_00524_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09609_ (.I0(\dp.rf.rf[24][19] ),
    .I1(_04571_),
    .S(_04676_),
    .Z(_00525_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09610_ (.I0(\dp.rf.rf[24][1] ),
    .I1(_04572_),
    .S(_04676_),
    .Z(_00526_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09611_ (.I0(\dp.rf.rf[24][20] ),
    .I1(_04573_),
    .S(_04676_),
    .Z(_00527_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09612_ (.I0(\dp.rf.rf[24][21] ),
    .I1(_04574_),
    .S(_04676_),
    .Z(_00528_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09613_ (.I0(\dp.rf.rf[24][22] ),
    .I1(_04575_),
    .S(_04676_),
    .Z(_00529_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09614_ (.I0(\dp.rf.rf[24][23] ),
    .I1(_04576_),
    .S(_04676_),
    .Z(_00530_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09615_ (.I0(\dp.rf.rf[24][24] ),
    .I1(_04577_),
    .S(_04676_),
    .Z(_00531_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09616_ (.I0(\dp.rf.rf[24][25] ),
    .I1(_04578_),
    .S(_04676_),
    .Z(_00532_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09617_ (.I(_04674_),
    .Z(_04677_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09618_ (.I0(\dp.rf.rf[24][26] ),
    .I1(_04579_),
    .S(_04677_),
    .Z(_00533_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09619_ (.I0(\dp.rf.rf[24][27] ),
    .I1(_04581_),
    .S(_04677_),
    .Z(_00534_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09620_ (.I0(\dp.rf.rf[24][28] ),
    .I1(_04582_),
    .S(_04677_),
    .Z(_00535_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09621_ (.I0(\dp.rf.rf[24][29] ),
    .I1(_04583_),
    .S(_04677_),
    .Z(_00536_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09622_ (.I0(\dp.rf.rf[24][2] ),
    .I1(_04584_),
    .S(_04677_),
    .Z(_00537_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09623_ (.I0(\dp.rf.rf[24][30] ),
    .I1(_04585_),
    .S(_04677_),
    .Z(_00538_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _09624_ (.I(_04481_),
    .Z(_04678_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09625_ (.A1(_04678_),
    .A2(_04675_),
    .Z(_04679_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09626_ (.A1(\dp.rf.rf[24][31] ),
    .A2(_04675_),
    .ZN(_04680_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09627_ (.A1(_04670_),
    .A2(_04679_),
    .B(_04680_),
    .ZN(_00539_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09628_ (.I0(\dp.rf.rf[24][3] ),
    .I1(_04588_),
    .S(_04677_),
    .Z(_00540_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09629_ (.I0(\dp.rf.rf[24][4] ),
    .I1(_04589_),
    .S(_04677_),
    .Z(_00541_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09630_ (.I0(\dp.rf.rf[24][5] ),
    .I1(_04590_),
    .S(_04677_),
    .Z(_00542_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09631_ (.I0(\dp.rf.rf[24][6] ),
    .I1(_04591_),
    .S(_04677_),
    .Z(_00543_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09632_ (.I0(\dp.rf.rf[24][7] ),
    .I1(_04592_),
    .S(_04674_),
    .Z(_00544_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09633_ (.I0(\dp.rf.rf[24][8] ),
    .I1(_04593_),
    .S(_04674_),
    .Z(_00545_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09634_ (.I0(\dp.rf.rf[24][9] ),
    .I1(_04594_),
    .S(_04674_),
    .Z(_00546_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09635_ (.A1(_04595_),
    .A2(_04673_),
    .ZN(_04681_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09636_ (.I(_04681_),
    .Z(_04682_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09637_ (.I0(_04073_),
    .I1(\dp.rf.rf[25][0] ),
    .S(_04682_),
    .Z(_00547_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09638_ (.I0(_04120_),
    .I1(\dp.rf.rf[25][10] ),
    .S(_04682_),
    .Z(_00548_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09639_ (.I0(_04150_),
    .I1(\dp.rf.rf[25][11] ),
    .S(_04682_),
    .Z(_00549_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09640_ (.I0(_04164_),
    .I1(\dp.rf.rf[25][12] ),
    .S(_04682_),
    .Z(_00550_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09641_ (.I0(_04178_),
    .I1(\dp.rf.rf[25][13] ),
    .S(_04682_),
    .Z(_00551_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09642_ (.I0(_04196_),
    .I1(\dp.rf.rf[25][14] ),
    .S(_04682_),
    .Z(_00552_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09643_ (.I0(_04209_),
    .I1(\dp.rf.rf[25][15] ),
    .S(_04682_),
    .Z(_00553_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09644_ (.I0(_04227_),
    .I1(\dp.rf.rf[25][16] ),
    .S(_04682_),
    .Z(_00554_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09645_ (.I0(_04244_),
    .I1(\dp.rf.rf[25][17] ),
    .S(_04682_),
    .Z(_00555_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _09646_ (.I(_04681_),
    .Z(_04683_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09647_ (.I0(_04259_),
    .I1(\dp.rf.rf[25][18] ),
    .S(_04683_),
    .Z(_00556_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09648_ (.I0(_04270_),
    .I1(\dp.rf.rf[25][19] ),
    .S(_04683_),
    .Z(_00557_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09649_ (.I0(_04275_),
    .I1(\dp.rf.rf[25][1] ),
    .S(_04683_),
    .Z(_00558_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09650_ (.I0(_04292_),
    .I1(\dp.rf.rf[25][20] ),
    .S(_04683_),
    .Z(_00559_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09651_ (.I0(_04313_),
    .I1(\dp.rf.rf[25][21] ),
    .S(_04683_),
    .Z(_00560_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09652_ (.I0(_04328_),
    .I1(\dp.rf.rf[25][22] ),
    .S(_04683_),
    .Z(_00561_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09653_ (.I0(_04342_),
    .I1(\dp.rf.rf[25][23] ),
    .S(_04683_),
    .Z(_00562_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09654_ (.I0(_04359_),
    .I1(\dp.rf.rf[25][24] ),
    .S(_04683_),
    .Z(_00563_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09655_ (.I0(_04381_),
    .I1(\dp.rf.rf[25][25] ),
    .S(_04683_),
    .Z(_00564_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09656_ (.I0(_04395_),
    .I1(\dp.rf.rf[25][26] ),
    .S(_04683_),
    .Z(_00565_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09657_ (.I(_04681_),
    .Z(_04684_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09658_ (.I0(_04409_),
    .I1(\dp.rf.rf[25][27] ),
    .S(_04684_),
    .Z(_00566_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09659_ (.I0(_04421_),
    .I1(\dp.rf.rf[25][28] ),
    .S(_04684_),
    .Z(_00567_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09660_ (.I0(_04439_),
    .I1(\dp.rf.rf[25][29] ),
    .S(_04684_),
    .Z(_00568_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09661_ (.I0(_04446_),
    .I1(\dp.rf.rf[25][2] ),
    .S(_04684_),
    .Z(_00569_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09662_ (.I0(_04462_),
    .I1(\dp.rf.rf[25][30] ),
    .S(_04684_),
    .Z(_00570_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09663_ (.A1(_04482_),
    .A2(_04601_),
    .A3(_04673_),
    .Z(_04685_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09664_ (.A1(_01216_),
    .A2(_04682_),
    .B1(_04685_),
    .B2(_04603_),
    .ZN(_00571_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09665_ (.I0(_04488_),
    .I1(\dp.rf.rf[25][3] ),
    .S(_04684_),
    .Z(_00572_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09666_ (.I0(_04496_),
    .I1(\dp.rf.rf[25][4] ),
    .S(_04684_),
    .Z(_00573_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09667_ (.I0(_04504_),
    .I1(\dp.rf.rf[25][5] ),
    .S(_04684_),
    .Z(_00574_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09668_ (.I0(_04512_),
    .I1(\dp.rf.rf[25][6] ),
    .S(_04684_),
    .Z(_00575_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09669_ (.I0(_04523_),
    .I1(\dp.rf.rf[25][7] ),
    .S(_04684_),
    .Z(_00576_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09670_ (.I0(_04534_),
    .I1(\dp.rf.rf[25][8] ),
    .S(_04681_),
    .Z(_00577_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09671_ (.I0(_04544_),
    .I1(\dp.rf.rf[25][9] ),
    .S(_04681_),
    .Z(_00578_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09672_ (.I(_04072_),
    .Z(_04686_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09673_ (.A1(_04081_),
    .A2(_04673_),
    .Z(_04687_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09674_ (.I(_04687_),
    .Z(_04688_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09675_ (.I0(\dp.rf.rf[26][0] ),
    .I1(_04686_),
    .S(_04688_),
    .Z(_00579_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09676_ (.I(_04119_),
    .Z(_04689_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09677_ (.I0(\dp.rf.rf[26][10] ),
    .I1(_04689_),
    .S(_04688_),
    .Z(_00580_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _09678_ (.I(_04149_),
    .Z(_04690_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09679_ (.I0(\dp.rf.rf[26][11] ),
    .I1(_04690_),
    .S(_04688_),
    .Z(_00581_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09680_ (.I(_04163_),
    .Z(_04691_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09681_ (.I0(\dp.rf.rf[26][12] ),
    .I1(_04691_),
    .S(_04688_),
    .Z(_00582_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09682_ (.I(_04177_),
    .Z(_04692_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09683_ (.I0(\dp.rf.rf[26][13] ),
    .I1(_04692_),
    .S(_04688_),
    .Z(_00583_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _09684_ (.I(_04195_),
    .Z(_04693_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09685_ (.I0(\dp.rf.rf[26][14] ),
    .I1(_04693_),
    .S(_04688_),
    .Z(_00584_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _09686_ (.I(_04208_),
    .Z(_04694_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09687_ (.I0(\dp.rf.rf[26][15] ),
    .I1(_04694_),
    .S(_04688_),
    .Z(_00585_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _09688_ (.I(_04226_),
    .Z(_04695_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09689_ (.I0(\dp.rf.rf[26][16] ),
    .I1(_04695_),
    .S(_04688_),
    .Z(_00586_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09690_ (.I(_04243_),
    .Z(_04696_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09691_ (.I(_04687_),
    .Z(_04697_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09692_ (.I0(\dp.rf.rf[26][17] ),
    .I1(_04696_),
    .S(_04697_),
    .Z(_00587_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09693_ (.I(_04258_),
    .Z(_04698_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09694_ (.I0(\dp.rf.rf[26][18] ),
    .I1(_04698_),
    .S(_04697_),
    .Z(_00588_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09695_ (.I(_04269_),
    .Z(_04699_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09696_ (.I0(\dp.rf.rf[26][19] ),
    .I1(_04699_),
    .S(_04697_),
    .Z(_00589_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _09697_ (.I(_04274_),
    .Z(_04700_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09698_ (.I0(\dp.rf.rf[26][1] ),
    .I1(_04700_),
    .S(_04697_),
    .Z(_00590_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09699_ (.I(_04291_),
    .Z(_04701_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09700_ (.I0(\dp.rf.rf[26][20] ),
    .I1(_04701_),
    .S(_04697_),
    .Z(_00591_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09701_ (.I(_04312_),
    .Z(_04702_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09702_ (.I0(\dp.rf.rf[26][21] ),
    .I1(_04702_),
    .S(_04697_),
    .Z(_00592_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _09703_ (.I(_04327_),
    .Z(_04703_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09704_ (.I0(\dp.rf.rf[26][22] ),
    .I1(_04703_),
    .S(_04697_),
    .Z(_00593_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _09705_ (.I(_04341_),
    .Z(_04704_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09706_ (.I0(\dp.rf.rf[26][23] ),
    .I1(_04704_),
    .S(_04697_),
    .Z(_00594_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _09707_ (.I(_04358_),
    .Z(_04705_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09708_ (.I0(\dp.rf.rf[26][24] ),
    .I1(_04705_),
    .S(_04697_),
    .Z(_00595_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09709_ (.I(_04380_),
    .Z(_04706_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09710_ (.I0(\dp.rf.rf[26][25] ),
    .I1(_04706_),
    .S(_04697_),
    .Z(_00596_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09711_ (.I(_04394_),
    .Z(_04707_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09712_ (.I(_04687_),
    .Z(_04708_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09713_ (.I0(\dp.rf.rf[26][26] ),
    .I1(_04707_),
    .S(_04708_),
    .Z(_00597_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09714_ (.I(_04408_),
    .Z(_04709_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09715_ (.I0(\dp.rf.rf[26][27] ),
    .I1(_04709_),
    .S(_04708_),
    .Z(_00598_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _09716_ (.I(_04420_),
    .Z(_04710_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09717_ (.I0(\dp.rf.rf[26][28] ),
    .I1(_04710_),
    .S(_04708_),
    .Z(_00599_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _09718_ (.I(_04438_),
    .Z(_04711_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09719_ (.I0(\dp.rf.rf[26][29] ),
    .I1(_04711_),
    .S(_04708_),
    .Z(_00600_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09720_ (.I(_04445_),
    .Z(_04712_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09721_ (.I0(\dp.rf.rf[26][2] ),
    .I1(_04712_),
    .S(_04708_),
    .Z(_00601_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _09722_ (.I(_04461_),
    .Z(_04713_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09723_ (.I0(\dp.rf.rf[26][30] ),
    .I1(_04713_),
    .S(_04708_),
    .Z(_00602_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09724_ (.A1(_04678_),
    .A2(_04688_),
    .Z(_04714_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09725_ (.A1(\dp.rf.rf[26][31] ),
    .A2(_04688_),
    .ZN(_04715_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09726_ (.A1(_04670_),
    .A2(_04714_),
    .B(_04715_),
    .ZN(_00603_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09727_ (.I(_04487_),
    .Z(_04716_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09728_ (.I0(\dp.rf.rf[26][3] ),
    .I1(_04716_),
    .S(_04708_),
    .Z(_00604_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09729_ (.I(_04495_),
    .Z(_04717_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09730_ (.I0(\dp.rf.rf[26][4] ),
    .I1(_04717_),
    .S(_04708_),
    .Z(_00605_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _09731_ (.I(_04503_),
    .Z(_04718_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09732_ (.I0(\dp.rf.rf[26][5] ),
    .I1(_04718_),
    .S(_04708_),
    .Z(_00606_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _09733_ (.I(_04511_),
    .Z(_04719_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09734_ (.I0(\dp.rf.rf[26][6] ),
    .I1(_04719_),
    .S(_04708_),
    .Z(_00607_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _09735_ (.I(_04522_),
    .Z(_04720_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09736_ (.I0(\dp.rf.rf[26][7] ),
    .I1(_04720_),
    .S(_04687_),
    .Z(_00608_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _09737_ (.I(_04533_),
    .Z(_04721_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09738_ (.I0(\dp.rf.rf[26][8] ),
    .I1(_04721_),
    .S(_04687_),
    .Z(_00609_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _09739_ (.I(_04543_),
    .Z(_04722_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09740_ (.I0(\dp.rf.rf[26][9] ),
    .I1(_04722_),
    .S(_04687_),
    .Z(_00610_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09741_ (.A1(_04545_),
    .A2(_04673_),
    .Z(_04723_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09742_ (.I(_04723_),
    .Z(_04724_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09743_ (.I0(\dp.rf.rf[27][0] ),
    .I1(_04686_),
    .S(_04724_),
    .Z(_00611_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09744_ (.I0(\dp.rf.rf[27][10] ),
    .I1(_04689_),
    .S(_04724_),
    .Z(_00612_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09745_ (.I0(\dp.rf.rf[27][11] ),
    .I1(_04690_),
    .S(_04724_),
    .Z(_00613_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09746_ (.I0(\dp.rf.rf[27][12] ),
    .I1(_04691_),
    .S(_04724_),
    .Z(_00614_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09747_ (.I0(\dp.rf.rf[27][13] ),
    .I1(_04692_),
    .S(_04724_),
    .Z(_00615_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09748_ (.I0(\dp.rf.rf[27][14] ),
    .I1(_04693_),
    .S(_04724_),
    .Z(_00616_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09749_ (.I0(\dp.rf.rf[27][15] ),
    .I1(_04694_),
    .S(_04724_),
    .Z(_00617_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09750_ (.I0(\dp.rf.rf[27][16] ),
    .I1(_04695_),
    .S(_04724_),
    .Z(_00618_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09751_ (.I(_04723_),
    .Z(_04725_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09752_ (.I0(\dp.rf.rf[27][17] ),
    .I1(_04696_),
    .S(_04725_),
    .Z(_00619_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09753_ (.I0(\dp.rf.rf[27][18] ),
    .I1(_04698_),
    .S(_04725_),
    .Z(_00620_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09754_ (.I0(\dp.rf.rf[27][19] ),
    .I1(_04699_),
    .S(_04725_),
    .Z(_00621_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09755_ (.I0(\dp.rf.rf[27][1] ),
    .I1(_04700_),
    .S(_04725_),
    .Z(_00622_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09756_ (.I0(\dp.rf.rf[27][20] ),
    .I1(_04701_),
    .S(_04725_),
    .Z(_00623_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09757_ (.I0(\dp.rf.rf[27][21] ),
    .I1(_04702_),
    .S(_04725_),
    .Z(_00624_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09758_ (.I0(\dp.rf.rf[27][22] ),
    .I1(_04703_),
    .S(_04725_),
    .Z(_00625_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09759_ (.I0(\dp.rf.rf[27][23] ),
    .I1(_04704_),
    .S(_04725_),
    .Z(_00626_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09760_ (.I0(\dp.rf.rf[27][24] ),
    .I1(_04705_),
    .S(_04725_),
    .Z(_00627_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09761_ (.I0(\dp.rf.rf[27][25] ),
    .I1(_04706_),
    .S(_04725_),
    .Z(_00628_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09762_ (.I(_04723_),
    .Z(_04726_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09763_ (.I0(\dp.rf.rf[27][26] ),
    .I1(_04707_),
    .S(_04726_),
    .Z(_00629_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09764_ (.I0(\dp.rf.rf[27][27] ),
    .I1(_04709_),
    .S(_04726_),
    .Z(_00630_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09765_ (.I0(\dp.rf.rf[27][28] ),
    .I1(_04710_),
    .S(_04726_),
    .Z(_00631_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09766_ (.I0(\dp.rf.rf[27][29] ),
    .I1(_04711_),
    .S(_04726_),
    .Z(_00632_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09767_ (.I0(\dp.rf.rf[27][2] ),
    .I1(_04712_),
    .S(_04726_),
    .Z(_00633_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09768_ (.I0(\dp.rf.rf[27][30] ),
    .I1(_04713_),
    .S(_04726_),
    .Z(_00634_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09769_ (.A1(_04678_),
    .A2(_04724_),
    .Z(_04727_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09770_ (.A1(\dp.rf.rf[27][31] ),
    .A2(_04724_),
    .ZN(_04728_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09771_ (.A1(_04670_),
    .A2(_04727_),
    .B(_04728_),
    .ZN(_00635_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09772_ (.I0(\dp.rf.rf[27][3] ),
    .I1(_04716_),
    .S(_04726_),
    .Z(_00636_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09773_ (.I0(\dp.rf.rf[27][4] ),
    .I1(_04717_),
    .S(_04726_),
    .Z(_00637_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09774_ (.I0(\dp.rf.rf[27][5] ),
    .I1(_04718_),
    .S(_04726_),
    .Z(_00638_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09775_ (.I0(\dp.rf.rf[27][6] ),
    .I1(_04719_),
    .S(_04726_),
    .Z(_00639_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09776_ (.I0(\dp.rf.rf[27][7] ),
    .I1(_04720_),
    .S(_04723_),
    .Z(_00640_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09777_ (.I0(\dp.rf.rf[27][8] ),
    .I1(_04721_),
    .S(_04723_),
    .Z(_00641_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09778_ (.I0(\dp.rf.rf[27][9] ),
    .I1(_04722_),
    .S(_04723_),
    .Z(_00642_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09779_ (.A1(net3),
    .A2(net2),
    .A3(net27),
    .Z(_04729_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09780_ (.A1(_04558_),
    .A2(_04729_),
    .Z(_04730_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09781_ (.I(_04730_),
    .Z(_04731_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09782_ (.I0(\dp.rf.rf[28][0] ),
    .I1(_04686_),
    .S(_04731_),
    .Z(_00643_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09783_ (.I0(\dp.rf.rf[28][10] ),
    .I1(_04689_),
    .S(_04731_),
    .Z(_00644_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09784_ (.I0(\dp.rf.rf[28][11] ),
    .I1(_04690_),
    .S(_04731_),
    .Z(_00645_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09785_ (.I0(\dp.rf.rf[28][12] ),
    .I1(_04691_),
    .S(_04731_),
    .Z(_00646_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09786_ (.I0(\dp.rf.rf[28][13] ),
    .I1(_04692_),
    .S(_04731_),
    .Z(_00647_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09787_ (.I0(\dp.rf.rf[28][14] ),
    .I1(_04693_),
    .S(_04731_),
    .Z(_00648_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09788_ (.I0(\dp.rf.rf[28][15] ),
    .I1(_04694_),
    .S(_04731_),
    .Z(_00649_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09789_ (.I0(\dp.rf.rf[28][16] ),
    .I1(_04695_),
    .S(_04731_),
    .Z(_00650_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09790_ (.I(_04730_),
    .Z(_04732_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09791_ (.I0(\dp.rf.rf[28][17] ),
    .I1(_04696_),
    .S(_04732_),
    .Z(_00651_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09792_ (.I0(\dp.rf.rf[28][18] ),
    .I1(_04698_),
    .S(_04732_),
    .Z(_00652_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09793_ (.I0(\dp.rf.rf[28][19] ),
    .I1(_04699_),
    .S(_04732_),
    .Z(_00653_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09794_ (.I0(\dp.rf.rf[28][1] ),
    .I1(_04700_),
    .S(_04732_),
    .Z(_00654_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09795_ (.I0(\dp.rf.rf[28][20] ),
    .I1(_04701_),
    .S(_04732_),
    .Z(_00655_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09796_ (.I0(\dp.rf.rf[28][21] ),
    .I1(_04702_),
    .S(_04732_),
    .Z(_00656_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09797_ (.I0(\dp.rf.rf[28][22] ),
    .I1(_04703_),
    .S(_04732_),
    .Z(_00657_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09798_ (.I0(\dp.rf.rf[28][23] ),
    .I1(_04704_),
    .S(_04732_),
    .Z(_00658_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09799_ (.I0(\dp.rf.rf[28][24] ),
    .I1(_04705_),
    .S(_04732_),
    .Z(_00659_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09800_ (.I0(\dp.rf.rf[28][25] ),
    .I1(_04706_),
    .S(_04732_),
    .Z(_00660_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09801_ (.I(_04730_),
    .Z(_04733_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09802_ (.I0(\dp.rf.rf[28][26] ),
    .I1(_04707_),
    .S(_04733_),
    .Z(_00661_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09803_ (.I0(\dp.rf.rf[28][27] ),
    .I1(_04709_),
    .S(_04733_),
    .Z(_00662_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09804_ (.I0(\dp.rf.rf[28][28] ),
    .I1(_04710_),
    .S(_04733_),
    .Z(_00663_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09805_ (.I0(\dp.rf.rf[28][29] ),
    .I1(_04711_),
    .S(_04733_),
    .Z(_00664_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09806_ (.I0(\dp.rf.rf[28][2] ),
    .I1(_04712_),
    .S(_04733_),
    .Z(_00665_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09807_ (.I0(\dp.rf.rf[28][30] ),
    .I1(_04713_),
    .S(_04733_),
    .Z(_00666_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09808_ (.A1(_04678_),
    .A2(_04731_),
    .Z(_04734_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09809_ (.A1(\dp.rf.rf[28][31] ),
    .A2(_04731_),
    .ZN(_04735_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09810_ (.A1(_04670_),
    .A2(_04734_),
    .B(_04735_),
    .ZN(_00667_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09811_ (.I0(\dp.rf.rf[28][3] ),
    .I1(_04716_),
    .S(_04733_),
    .Z(_00668_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09812_ (.I0(\dp.rf.rf[28][4] ),
    .I1(_04717_),
    .S(_04733_),
    .Z(_00669_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09813_ (.I0(\dp.rf.rf[28][5] ),
    .I1(_04718_),
    .S(_04733_),
    .Z(_00670_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09814_ (.I0(\dp.rf.rf[28][6] ),
    .I1(_04719_),
    .S(_04733_),
    .Z(_00671_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09815_ (.I0(\dp.rf.rf[28][7] ),
    .I1(_04720_),
    .S(_04730_),
    .Z(_00672_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09816_ (.I0(\dp.rf.rf[28][8] ),
    .I1(_04721_),
    .S(_04730_),
    .Z(_00673_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09817_ (.I0(\dp.rf.rf[28][9] ),
    .I1(_04722_),
    .S(_04730_),
    .Z(_00674_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09818_ (.A1(_04595_),
    .A2(_04729_),
    .ZN(_04736_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09819_ (.I(_04736_),
    .Z(_04737_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09820_ (.I0(_04073_),
    .I1(\dp.rf.rf[29][0] ),
    .S(_04737_),
    .Z(_00675_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09821_ (.I0(_04120_),
    .I1(\dp.rf.rf[29][10] ),
    .S(_04737_),
    .Z(_00676_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09822_ (.I0(_04150_),
    .I1(\dp.rf.rf[29][11] ),
    .S(_04737_),
    .Z(_00677_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09823_ (.I0(_04164_),
    .I1(\dp.rf.rf[29][12] ),
    .S(_04737_),
    .Z(_00678_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09824_ (.I0(_04178_),
    .I1(\dp.rf.rf[29][13] ),
    .S(_04737_),
    .Z(_00679_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09825_ (.I0(_04196_),
    .I1(\dp.rf.rf[29][14] ),
    .S(_04737_),
    .Z(_00680_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09826_ (.I0(_04209_),
    .I1(\dp.rf.rf[29][15] ),
    .S(_04737_),
    .Z(_00681_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09827_ (.I0(_04227_),
    .I1(\dp.rf.rf[29][16] ),
    .S(_04737_),
    .Z(_00682_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09828_ (.I0(_04244_),
    .I1(\dp.rf.rf[29][17] ),
    .S(_04737_),
    .Z(_00683_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _09829_ (.I(_04736_),
    .Z(_04738_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09830_ (.I0(_04259_),
    .I1(\dp.rf.rf[29][18] ),
    .S(_04738_),
    .Z(_00684_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09831_ (.I0(_04270_),
    .I1(\dp.rf.rf[29][19] ),
    .S(_04738_),
    .Z(_00685_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09832_ (.I0(_04275_),
    .I1(\dp.rf.rf[29][1] ),
    .S(_04738_),
    .Z(_00686_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09833_ (.I0(_04292_),
    .I1(\dp.rf.rf[29][20] ),
    .S(_04738_),
    .Z(_00687_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09834_ (.I0(_04313_),
    .I1(\dp.rf.rf[29][21] ),
    .S(_04738_),
    .Z(_00688_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09835_ (.I0(_04328_),
    .I1(\dp.rf.rf[29][22] ),
    .S(_04738_),
    .Z(_00689_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09836_ (.I0(_04342_),
    .I1(\dp.rf.rf[29][23] ),
    .S(_04738_),
    .Z(_00690_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09837_ (.I0(_04359_),
    .I1(\dp.rf.rf[29][24] ),
    .S(_04738_),
    .Z(_00691_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09838_ (.I0(_04381_),
    .I1(\dp.rf.rf[29][25] ),
    .S(_04738_),
    .Z(_00692_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09839_ (.I0(_04395_),
    .I1(\dp.rf.rf[29][26] ),
    .S(_04738_),
    .Z(_00693_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09840_ (.I(_04736_),
    .Z(_04739_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09841_ (.I0(_04409_),
    .I1(\dp.rf.rf[29][27] ),
    .S(_04739_),
    .Z(_00694_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09842_ (.I0(_04421_),
    .I1(\dp.rf.rf[29][28] ),
    .S(_04739_),
    .Z(_00695_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09843_ (.I0(_04439_),
    .I1(\dp.rf.rf[29][29] ),
    .S(_04739_),
    .Z(_00696_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09844_ (.I0(_04446_),
    .I1(\dp.rf.rf[29][2] ),
    .S(_04739_),
    .Z(_00697_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09845_ (.I0(_04462_),
    .I1(\dp.rf.rf[29][30] ),
    .S(_04739_),
    .Z(_00698_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09846_ (.I(\dp.rf.rf[29][31] ),
    .ZN(_04740_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09847_ (.A1(_04482_),
    .A2(_04601_),
    .A3(_04729_),
    .Z(_04741_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09848_ (.A1(_04740_),
    .A2(_04737_),
    .B1(_04741_),
    .B2(_04603_),
    .ZN(_00699_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09849_ (.I0(_04488_),
    .I1(\dp.rf.rf[29][3] ),
    .S(_04739_),
    .Z(_00700_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09850_ (.I0(_04496_),
    .I1(\dp.rf.rf[29][4] ),
    .S(_04739_),
    .Z(_00701_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09851_ (.I0(_04504_),
    .I1(\dp.rf.rf[29][5] ),
    .S(_04739_),
    .Z(_00702_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09852_ (.I0(_04512_),
    .I1(\dp.rf.rf[29][6] ),
    .S(_04739_),
    .Z(_00703_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09853_ (.I0(_04523_),
    .I1(\dp.rf.rf[29][7] ),
    .S(_04739_),
    .Z(_00704_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09854_ (.I0(_04534_),
    .I1(\dp.rf.rf[29][8] ),
    .S(_04736_),
    .Z(_00705_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09855_ (.I0(_04544_),
    .I1(\dp.rf.rf[29][9] ),
    .S(_04736_),
    .Z(_00706_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09856_ (.A1(_04081_),
    .A2(_04556_),
    .Z(_04742_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _09857_ (.I(_04742_),
    .Z(_04743_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09858_ (.I0(\dp.rf.rf[2][0] ),
    .I1(_04686_),
    .S(_04743_),
    .Z(_00707_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09859_ (.I0(\dp.rf.rf[2][10] ),
    .I1(_04689_),
    .S(_04743_),
    .Z(_00708_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09860_ (.I0(\dp.rf.rf[2][11] ),
    .I1(_04690_),
    .S(_04743_),
    .Z(_00709_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09861_ (.I0(\dp.rf.rf[2][12] ),
    .I1(_04691_),
    .S(_04743_),
    .Z(_00710_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09862_ (.I0(\dp.rf.rf[2][13] ),
    .I1(_04692_),
    .S(_04743_),
    .Z(_00711_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09863_ (.I0(\dp.rf.rf[2][14] ),
    .I1(_04693_),
    .S(_04743_),
    .Z(_00712_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09864_ (.I0(\dp.rf.rf[2][15] ),
    .I1(_04694_),
    .S(_04743_),
    .Z(_00713_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09865_ (.I0(\dp.rf.rf[2][16] ),
    .I1(_04695_),
    .S(_04743_),
    .Z(_00714_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09866_ (.I(_04742_),
    .Z(_04744_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09867_ (.I0(\dp.rf.rf[2][17] ),
    .I1(_04696_),
    .S(_04744_),
    .Z(_00715_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09868_ (.I0(\dp.rf.rf[2][18] ),
    .I1(_04698_),
    .S(_04744_),
    .Z(_00716_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09869_ (.I0(\dp.rf.rf[2][19] ),
    .I1(_04699_),
    .S(_04744_),
    .Z(_00717_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09870_ (.I0(\dp.rf.rf[2][1] ),
    .I1(_04700_),
    .S(_04744_),
    .Z(_00718_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09871_ (.I0(\dp.rf.rf[2][20] ),
    .I1(_04701_),
    .S(_04744_),
    .Z(_00719_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09872_ (.I0(\dp.rf.rf[2][21] ),
    .I1(_04702_),
    .S(_04744_),
    .Z(_00720_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09873_ (.I0(\dp.rf.rf[2][22] ),
    .I1(_04703_),
    .S(_04744_),
    .Z(_00721_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09874_ (.I0(\dp.rf.rf[2][23] ),
    .I1(_04704_),
    .S(_04744_),
    .Z(_00722_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09875_ (.I0(\dp.rf.rf[2][24] ),
    .I1(_04705_),
    .S(_04744_),
    .Z(_00723_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09876_ (.I0(\dp.rf.rf[2][25] ),
    .I1(_04706_),
    .S(_04744_),
    .Z(_00724_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _09877_ (.I(_04742_),
    .Z(_04745_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09878_ (.I0(\dp.rf.rf[2][26] ),
    .I1(_04707_),
    .S(_04745_),
    .Z(_00725_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09879_ (.I0(\dp.rf.rf[2][27] ),
    .I1(_04709_),
    .S(_04745_),
    .Z(_00726_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09880_ (.I0(\dp.rf.rf[2][28] ),
    .I1(_04710_),
    .S(_04745_),
    .Z(_00727_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09881_ (.I0(\dp.rf.rf[2][29] ),
    .I1(_04711_),
    .S(_04745_),
    .Z(_00728_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09882_ (.I0(\dp.rf.rf[2][2] ),
    .I1(_04712_),
    .S(_04745_),
    .Z(_00729_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09883_ (.I0(\dp.rf.rf[2][30] ),
    .I1(_04713_),
    .S(_04745_),
    .Z(_00730_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09884_ (.A1(_04678_),
    .A2(_04743_),
    .Z(_04746_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09885_ (.A1(\dp.rf.rf[2][31] ),
    .A2(_04743_),
    .ZN(_04747_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09886_ (.A1(_04670_),
    .A2(_04746_),
    .B(_04747_),
    .ZN(_00731_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09887_ (.I0(\dp.rf.rf[2][3] ),
    .I1(_04716_),
    .S(_04745_),
    .Z(_00732_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09888_ (.I0(\dp.rf.rf[2][4] ),
    .I1(_04717_),
    .S(_04745_),
    .Z(_00733_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09889_ (.I0(\dp.rf.rf[2][5] ),
    .I1(_04718_),
    .S(_04745_),
    .Z(_00734_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09890_ (.I0(\dp.rf.rf[2][6] ),
    .I1(_04719_),
    .S(_04745_),
    .Z(_00735_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09891_ (.I0(\dp.rf.rf[2][7] ),
    .I1(_04720_),
    .S(_04742_),
    .Z(_00736_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09892_ (.I0(\dp.rf.rf[2][8] ),
    .I1(_04721_),
    .S(_04742_),
    .Z(_00737_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09893_ (.I0(\dp.rf.rf[2][9] ),
    .I1(_04722_),
    .S(_04742_),
    .Z(_00738_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09894_ (.A1(_04081_),
    .A2(_04729_),
    .Z(_04748_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09895_ (.I(_04748_),
    .Z(_04749_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09896_ (.I0(\dp.rf.rf[30][0] ),
    .I1(_04686_),
    .S(_04749_),
    .Z(_00739_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09897_ (.I0(\dp.rf.rf[30][10] ),
    .I1(_04689_),
    .S(_04749_),
    .Z(_00740_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09898_ (.I0(\dp.rf.rf[30][11] ),
    .I1(_04690_),
    .S(_04749_),
    .Z(_00741_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09899_ (.I0(\dp.rf.rf[30][12] ),
    .I1(_04691_),
    .S(_04749_),
    .Z(_00742_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09900_ (.I0(\dp.rf.rf[30][13] ),
    .I1(_04692_),
    .S(_04749_),
    .Z(_00743_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09901_ (.I0(\dp.rf.rf[30][14] ),
    .I1(_04693_),
    .S(_04749_),
    .Z(_00744_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09902_ (.I0(\dp.rf.rf[30][15] ),
    .I1(_04694_),
    .S(_04749_),
    .Z(_00745_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09903_ (.I0(\dp.rf.rf[30][16] ),
    .I1(_04695_),
    .S(_04749_),
    .Z(_00746_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09904_ (.I(_04748_),
    .Z(_04750_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09905_ (.I0(\dp.rf.rf[30][17] ),
    .I1(_04696_),
    .S(_04750_),
    .Z(_00747_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09906_ (.I0(\dp.rf.rf[30][18] ),
    .I1(_04698_),
    .S(_04750_),
    .Z(_00748_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09907_ (.I0(\dp.rf.rf[30][19] ),
    .I1(_04699_),
    .S(_04750_),
    .Z(_00749_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09908_ (.I0(\dp.rf.rf[30][1] ),
    .I1(_04700_),
    .S(_04750_),
    .Z(_00750_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09909_ (.I0(\dp.rf.rf[30][20] ),
    .I1(_04701_),
    .S(_04750_),
    .Z(_00751_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09910_ (.I0(\dp.rf.rf[30][21] ),
    .I1(_04702_),
    .S(_04750_),
    .Z(_00752_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09911_ (.I0(\dp.rf.rf[30][22] ),
    .I1(_04703_),
    .S(_04750_),
    .Z(_00753_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09912_ (.I0(\dp.rf.rf[30][23] ),
    .I1(_04704_),
    .S(_04750_),
    .Z(_00754_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09913_ (.I0(\dp.rf.rf[30][24] ),
    .I1(_04705_),
    .S(_04750_),
    .Z(_00755_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09914_ (.I0(\dp.rf.rf[30][25] ),
    .I1(_04706_),
    .S(_04750_),
    .Z(_00756_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09915_ (.I(_04748_),
    .Z(_04751_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09916_ (.I0(\dp.rf.rf[30][26] ),
    .I1(_04707_),
    .S(_04751_),
    .Z(_00757_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09917_ (.I0(\dp.rf.rf[30][27] ),
    .I1(_04709_),
    .S(_04751_),
    .Z(_00758_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09918_ (.I0(\dp.rf.rf[30][28] ),
    .I1(_04710_),
    .S(_04751_),
    .Z(_00759_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09919_ (.I0(\dp.rf.rf[30][29] ),
    .I1(_04711_),
    .S(_04751_),
    .Z(_00760_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09920_ (.I0(\dp.rf.rf[30][2] ),
    .I1(_04712_),
    .S(_04751_),
    .Z(_00761_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09921_ (.I0(\dp.rf.rf[30][30] ),
    .I1(_04713_),
    .S(_04751_),
    .Z(_00762_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09922_ (.A1(_04678_),
    .A2(_04749_),
    .Z(_04752_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09923_ (.A1(\dp.rf.rf[30][31] ),
    .A2(_04749_),
    .ZN(_04753_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09924_ (.A1(_04670_),
    .A2(_04752_),
    .B(_04753_),
    .ZN(_00763_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09925_ (.I0(\dp.rf.rf[30][3] ),
    .I1(_04716_),
    .S(_04751_),
    .Z(_00764_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09926_ (.I0(\dp.rf.rf[30][4] ),
    .I1(_04717_),
    .S(_04751_),
    .Z(_00765_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09927_ (.I0(\dp.rf.rf[30][5] ),
    .I1(_04718_),
    .S(_04751_),
    .Z(_00766_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09928_ (.I0(\dp.rf.rf[30][6] ),
    .I1(_04719_),
    .S(_04751_),
    .Z(_00767_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09929_ (.I0(\dp.rf.rf[30][7] ),
    .I1(_04720_),
    .S(_04748_),
    .Z(_00768_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09930_ (.I0(\dp.rf.rf[30][8] ),
    .I1(_04721_),
    .S(_04748_),
    .Z(_00769_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09931_ (.I0(\dp.rf.rf[30][9] ),
    .I1(_04722_),
    .S(_04748_),
    .Z(_00770_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09932_ (.A1(_04545_),
    .A2(_04729_),
    .Z(_04754_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09933_ (.I(_04754_),
    .Z(_04755_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09934_ (.I0(\dp.rf.rf[31][0] ),
    .I1(_04686_),
    .S(_04755_),
    .Z(_00771_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09935_ (.I0(\dp.rf.rf[31][10] ),
    .I1(_04689_),
    .S(_04755_),
    .Z(_00772_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09936_ (.I0(\dp.rf.rf[31][11] ),
    .I1(_04690_),
    .S(_04755_),
    .Z(_00773_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09937_ (.I0(\dp.rf.rf[31][12] ),
    .I1(_04691_),
    .S(_04755_),
    .Z(_00774_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09938_ (.I0(\dp.rf.rf[31][13] ),
    .I1(_04692_),
    .S(_04755_),
    .Z(_00775_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09939_ (.I0(\dp.rf.rf[31][14] ),
    .I1(_04693_),
    .S(_04755_),
    .Z(_00776_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09940_ (.I0(\dp.rf.rf[31][15] ),
    .I1(_04694_),
    .S(_04755_),
    .Z(_00777_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09941_ (.I0(\dp.rf.rf[31][16] ),
    .I1(_04695_),
    .S(_04755_),
    .Z(_00778_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09942_ (.I(_04754_),
    .Z(_04756_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09943_ (.I0(\dp.rf.rf[31][17] ),
    .I1(_04696_),
    .S(_04756_),
    .Z(_00779_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09944_ (.I0(\dp.rf.rf[31][18] ),
    .I1(_04698_),
    .S(_04756_),
    .Z(_00780_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09945_ (.I0(\dp.rf.rf[31][19] ),
    .I1(_04699_),
    .S(_04756_),
    .Z(_00781_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09946_ (.I0(\dp.rf.rf[31][1] ),
    .I1(_04700_),
    .S(_04756_),
    .Z(_00782_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09947_ (.I0(\dp.rf.rf[31][20] ),
    .I1(_04701_),
    .S(_04756_),
    .Z(_00783_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09948_ (.I0(\dp.rf.rf[31][21] ),
    .I1(_04702_),
    .S(_04756_),
    .Z(_00784_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09949_ (.I0(\dp.rf.rf[31][22] ),
    .I1(_04703_),
    .S(_04756_),
    .Z(_00785_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09950_ (.I0(\dp.rf.rf[31][23] ),
    .I1(_04704_),
    .S(_04756_),
    .Z(_00786_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09951_ (.I0(\dp.rf.rf[31][24] ),
    .I1(_04705_),
    .S(_04756_),
    .Z(_00787_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09952_ (.I0(\dp.rf.rf[31][25] ),
    .I1(_04706_),
    .S(_04756_),
    .Z(_00788_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09953_ (.I(_04754_),
    .Z(_04757_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09954_ (.I0(\dp.rf.rf[31][26] ),
    .I1(_04707_),
    .S(_04757_),
    .Z(_00789_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09955_ (.I0(\dp.rf.rf[31][27] ),
    .I1(_04709_),
    .S(_04757_),
    .Z(_00790_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09956_ (.I0(\dp.rf.rf[31][28] ),
    .I1(_04710_),
    .S(_04757_),
    .Z(_00791_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09957_ (.I0(\dp.rf.rf[31][29] ),
    .I1(_04711_),
    .S(_04757_),
    .Z(_00792_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09958_ (.I0(\dp.rf.rf[31][2] ),
    .I1(_04712_),
    .S(_04757_),
    .Z(_00793_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09959_ (.I0(\dp.rf.rf[31][30] ),
    .I1(_04713_),
    .S(_04757_),
    .Z(_00794_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09960_ (.A1(_04678_),
    .A2(_04755_),
    .Z(_04758_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09961_ (.A1(\dp.rf.rf[31][31] ),
    .A2(_04755_),
    .ZN(_04759_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09962_ (.A1(_04670_),
    .A2(_04758_),
    .B(_04759_),
    .ZN(_00795_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09963_ (.I0(\dp.rf.rf[31][3] ),
    .I1(_04716_),
    .S(_04757_),
    .Z(_00796_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09964_ (.I0(\dp.rf.rf[31][4] ),
    .I1(_04717_),
    .S(_04757_),
    .Z(_00797_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09965_ (.I0(\dp.rf.rf[31][5] ),
    .I1(_04718_),
    .S(_04757_),
    .Z(_00798_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09966_ (.I0(\dp.rf.rf[31][6] ),
    .I1(_04719_),
    .S(_04757_),
    .Z(_00799_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09967_ (.I0(\dp.rf.rf[31][7] ),
    .I1(_04720_),
    .S(_04754_),
    .Z(_00800_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09968_ (.I0(\dp.rf.rf[31][8] ),
    .I1(_04721_),
    .S(_04754_),
    .Z(_00801_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09969_ (.I0(\dp.rf.rf[31][9] ),
    .I1(_04722_),
    .S(_04754_),
    .Z(_00802_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09970_ (.A1(_04545_),
    .A2(_04556_),
    .Z(_04760_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09971_ (.I(_04760_),
    .Z(_04761_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09972_ (.I0(\dp.rf.rf[3][0] ),
    .I1(_04686_),
    .S(_04761_),
    .Z(_00803_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09973_ (.I0(\dp.rf.rf[3][10] ),
    .I1(_04689_),
    .S(_04761_),
    .Z(_00804_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09974_ (.I0(\dp.rf.rf[3][11] ),
    .I1(_04690_),
    .S(_04761_),
    .Z(_00805_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09975_ (.I0(\dp.rf.rf[3][12] ),
    .I1(_04691_),
    .S(_04761_),
    .Z(_00806_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09976_ (.I0(\dp.rf.rf[3][13] ),
    .I1(_04692_),
    .S(_04761_),
    .Z(_00807_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09977_ (.I0(\dp.rf.rf[3][14] ),
    .I1(_04693_),
    .S(_04761_),
    .Z(_00808_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09978_ (.I0(\dp.rf.rf[3][15] ),
    .I1(_04694_),
    .S(_04761_),
    .Z(_00809_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09979_ (.I0(\dp.rf.rf[3][16] ),
    .I1(_04695_),
    .S(_04761_),
    .Z(_00810_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09980_ (.I(_04760_),
    .Z(_04762_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09981_ (.I0(\dp.rf.rf[3][17] ),
    .I1(_04696_),
    .S(_04762_),
    .Z(_00811_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09982_ (.I0(\dp.rf.rf[3][18] ),
    .I1(_04698_),
    .S(_04762_),
    .Z(_00812_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09983_ (.I0(\dp.rf.rf[3][19] ),
    .I1(_04699_),
    .S(_04762_),
    .Z(_00813_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09984_ (.I0(\dp.rf.rf[3][1] ),
    .I1(_04700_),
    .S(_04762_),
    .Z(_00814_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09985_ (.I0(\dp.rf.rf[3][20] ),
    .I1(_04701_),
    .S(_04762_),
    .Z(_00815_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09986_ (.I0(\dp.rf.rf[3][21] ),
    .I1(_04702_),
    .S(_04762_),
    .Z(_00816_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09987_ (.I0(\dp.rf.rf[3][22] ),
    .I1(_04703_),
    .S(_04762_),
    .Z(_00817_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09988_ (.I0(\dp.rf.rf[3][23] ),
    .I1(_04704_),
    .S(_04762_),
    .Z(_00818_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09989_ (.I0(\dp.rf.rf[3][24] ),
    .I1(_04705_),
    .S(_04762_),
    .Z(_00819_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09990_ (.I0(\dp.rf.rf[3][25] ),
    .I1(_04706_),
    .S(_04762_),
    .Z(_00820_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09991_ (.I(_04760_),
    .Z(_04763_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09992_ (.I0(\dp.rf.rf[3][26] ),
    .I1(_04707_),
    .S(_04763_),
    .Z(_00821_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09993_ (.I0(\dp.rf.rf[3][27] ),
    .I1(_04709_),
    .S(_04763_),
    .Z(_00822_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09994_ (.I0(\dp.rf.rf[3][28] ),
    .I1(_04710_),
    .S(_04763_),
    .Z(_00823_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09995_ (.I0(\dp.rf.rf[3][29] ),
    .I1(_04711_),
    .S(_04763_),
    .Z(_00824_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09996_ (.I0(\dp.rf.rf[3][2] ),
    .I1(_04712_),
    .S(_04763_),
    .Z(_00825_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09997_ (.I0(\dp.rf.rf[3][30] ),
    .I1(_04713_),
    .S(_04763_),
    .Z(_00826_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09998_ (.A1(_04678_),
    .A2(_04761_),
    .Z(_04764_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09999_ (.A1(\dp.rf.rf[3][31] ),
    .A2(_04761_),
    .ZN(_04765_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10000_ (.A1(_04670_),
    .A2(_04764_),
    .B(_04765_),
    .ZN(_00827_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10001_ (.I0(\dp.rf.rf[3][3] ),
    .I1(_04716_),
    .S(_04763_),
    .Z(_00828_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10002_ (.I0(\dp.rf.rf[3][4] ),
    .I1(_04717_),
    .S(_04763_),
    .Z(_00829_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10003_ (.I0(\dp.rf.rf[3][5] ),
    .I1(_04718_),
    .S(_04763_),
    .Z(_00830_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10004_ (.I0(\dp.rf.rf[3][6] ),
    .I1(_04719_),
    .S(_04763_),
    .Z(_00831_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10005_ (.I0(\dp.rf.rf[3][7] ),
    .I1(_04720_),
    .S(_04760_),
    .Z(_00832_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10006_ (.I0(\dp.rf.rf[3][8] ),
    .I1(_04721_),
    .S(_04760_),
    .Z(_00833_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10007_ (.I0(\dp.rf.rf[3][9] ),
    .I1(_04722_),
    .S(_04760_),
    .Z(_00834_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10008_ (.A1(_02672_),
    .A2(_04555_),
    .A3(net27),
    .Z(_04766_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10009_ (.A1(_04558_),
    .A2(_04766_),
    .Z(_04767_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _10010_ (.I(_04767_),
    .Z(_04768_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10011_ (.I0(\dp.rf.rf[4][0] ),
    .I1(_04686_),
    .S(_04768_),
    .Z(_00835_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10012_ (.I0(\dp.rf.rf[4][10] ),
    .I1(_04689_),
    .S(_04768_),
    .Z(_00836_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10013_ (.I0(\dp.rf.rf[4][11] ),
    .I1(_04690_),
    .S(_04768_),
    .Z(_00837_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10014_ (.I0(\dp.rf.rf[4][12] ),
    .I1(_04691_),
    .S(_04768_),
    .Z(_00838_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10015_ (.I0(\dp.rf.rf[4][13] ),
    .I1(_04692_),
    .S(_04768_),
    .Z(_00839_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10016_ (.I0(\dp.rf.rf[4][14] ),
    .I1(_04693_),
    .S(_04768_),
    .Z(_00840_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10017_ (.I0(\dp.rf.rf[4][15] ),
    .I1(_04694_),
    .S(_04768_),
    .Z(_00841_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10018_ (.I0(\dp.rf.rf[4][16] ),
    .I1(_04695_),
    .S(_04768_),
    .Z(_00842_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _10019_ (.I(_04767_),
    .Z(_04769_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10020_ (.I0(\dp.rf.rf[4][17] ),
    .I1(_04696_),
    .S(_04769_),
    .Z(_00843_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10021_ (.I0(\dp.rf.rf[4][18] ),
    .I1(_04698_),
    .S(_04769_),
    .Z(_00844_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10022_ (.I0(\dp.rf.rf[4][19] ),
    .I1(_04699_),
    .S(_04769_),
    .Z(_00845_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10023_ (.I0(\dp.rf.rf[4][1] ),
    .I1(_04700_),
    .S(_04769_),
    .Z(_00846_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10024_ (.I0(\dp.rf.rf[4][20] ),
    .I1(_04701_),
    .S(_04769_),
    .Z(_00847_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10025_ (.I0(\dp.rf.rf[4][21] ),
    .I1(_04702_),
    .S(_04769_),
    .Z(_00848_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10026_ (.I0(\dp.rf.rf[4][22] ),
    .I1(_04703_),
    .S(_04769_),
    .Z(_00849_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10027_ (.I0(\dp.rf.rf[4][23] ),
    .I1(_04704_),
    .S(_04769_),
    .Z(_00850_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10028_ (.I0(\dp.rf.rf[4][24] ),
    .I1(_04705_),
    .S(_04769_),
    .Z(_00851_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10029_ (.I0(\dp.rf.rf[4][25] ),
    .I1(_04706_),
    .S(_04769_),
    .Z(_00852_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _10030_ (.I(_04767_),
    .Z(_04770_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10031_ (.I0(\dp.rf.rf[4][26] ),
    .I1(_04707_),
    .S(_04770_),
    .Z(_00853_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10032_ (.I0(\dp.rf.rf[4][27] ),
    .I1(_04709_),
    .S(_04770_),
    .Z(_00854_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10033_ (.I0(\dp.rf.rf[4][28] ),
    .I1(_04710_),
    .S(_04770_),
    .Z(_00855_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10034_ (.I0(\dp.rf.rf[4][29] ),
    .I1(_04711_),
    .S(_04770_),
    .Z(_00856_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10035_ (.I0(\dp.rf.rf[4][2] ),
    .I1(_04712_),
    .S(_04770_),
    .Z(_00857_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10036_ (.I0(\dp.rf.rf[4][30] ),
    .I1(_04713_),
    .S(_04770_),
    .Z(_00858_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10037_ (.A1(_04678_),
    .A2(_04768_),
    .Z(_04771_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10038_ (.A1(\dp.rf.rf[4][31] ),
    .A2(_04768_),
    .ZN(_04772_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10039_ (.A1(_04670_),
    .A2(_04771_),
    .B(_04772_),
    .ZN(_00859_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10040_ (.I0(\dp.rf.rf[4][3] ),
    .I1(_04716_),
    .S(_04770_),
    .Z(_00860_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10041_ (.I0(\dp.rf.rf[4][4] ),
    .I1(_04717_),
    .S(_04770_),
    .Z(_00861_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10042_ (.I0(\dp.rf.rf[4][5] ),
    .I1(_04718_),
    .S(_04770_),
    .Z(_00862_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10043_ (.I0(\dp.rf.rf[4][6] ),
    .I1(_04719_),
    .S(_04770_),
    .Z(_00863_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10044_ (.I0(\dp.rf.rf[4][7] ),
    .I1(_04720_),
    .S(_04767_),
    .Z(_00864_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10045_ (.I0(\dp.rf.rf[4][8] ),
    .I1(_04721_),
    .S(_04767_),
    .Z(_00865_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10046_ (.I0(\dp.rf.rf[4][9] ),
    .I1(_04722_),
    .S(_04767_),
    .Z(_00866_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10047_ (.A1(_04595_),
    .A2(_04766_),
    .ZN(_04773_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _10048_ (.I(_04773_),
    .Z(_04774_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10049_ (.I0(_04073_),
    .I1(\dp.rf.rf[5][0] ),
    .S(_04774_),
    .Z(_00867_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10050_ (.I0(_04120_),
    .I1(\dp.rf.rf[5][10] ),
    .S(_04774_),
    .Z(_00868_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10051_ (.I0(_04150_),
    .I1(\dp.rf.rf[5][11] ),
    .S(_04774_),
    .Z(_00869_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10052_ (.I0(_04164_),
    .I1(\dp.rf.rf[5][12] ),
    .S(_04774_),
    .Z(_00870_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10053_ (.I0(_04178_),
    .I1(\dp.rf.rf[5][13] ),
    .S(_04774_),
    .Z(_00871_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10054_ (.I0(_04196_),
    .I1(\dp.rf.rf[5][14] ),
    .S(_04774_),
    .Z(_00872_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10055_ (.I0(_04209_),
    .I1(\dp.rf.rf[5][15] ),
    .S(_04774_),
    .Z(_00873_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10056_ (.I0(_04227_),
    .I1(\dp.rf.rf[5][16] ),
    .S(_04774_),
    .Z(_00874_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10057_ (.I0(_04244_),
    .I1(\dp.rf.rf[5][17] ),
    .S(_04774_),
    .Z(_00875_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _10058_ (.I(_04773_),
    .Z(_04775_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10059_ (.I0(_04259_),
    .I1(\dp.rf.rf[5][18] ),
    .S(_04775_),
    .Z(_00876_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10060_ (.I0(_04270_),
    .I1(\dp.rf.rf[5][19] ),
    .S(_04775_),
    .Z(_00877_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10061_ (.I0(_04275_),
    .I1(\dp.rf.rf[5][1] ),
    .S(_04775_),
    .Z(_00878_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10062_ (.I0(_04292_),
    .I1(\dp.rf.rf[5][20] ),
    .S(_04775_),
    .Z(_00879_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10063_ (.I0(_04313_),
    .I1(\dp.rf.rf[5][21] ),
    .S(_04775_),
    .Z(_00880_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10064_ (.I0(_04328_),
    .I1(\dp.rf.rf[5][22] ),
    .S(_04775_),
    .Z(_00881_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10065_ (.I0(_04342_),
    .I1(\dp.rf.rf[5][23] ),
    .S(_04775_),
    .Z(_00882_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10066_ (.I0(_04359_),
    .I1(\dp.rf.rf[5][24] ),
    .S(_04775_),
    .Z(_00883_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10067_ (.I0(_04381_),
    .I1(\dp.rf.rf[5][25] ),
    .S(_04775_),
    .Z(_00884_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10068_ (.I0(_04395_),
    .I1(\dp.rf.rf[5][26] ),
    .S(_04775_),
    .Z(_00885_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _10069_ (.I(_04773_),
    .Z(_04776_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10070_ (.I0(_04409_),
    .I1(\dp.rf.rf[5][27] ),
    .S(_04776_),
    .Z(_00886_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10071_ (.I0(_04421_),
    .I1(\dp.rf.rf[5][28] ),
    .S(_04776_),
    .Z(_00887_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10072_ (.I0(_04439_),
    .I1(\dp.rf.rf[5][29] ),
    .S(_04776_),
    .Z(_00888_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10073_ (.I0(_04446_),
    .I1(\dp.rf.rf[5][2] ),
    .S(_04776_),
    .Z(_00889_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10074_ (.I0(_04462_),
    .I1(\dp.rf.rf[5][30] ),
    .S(_04776_),
    .Z(_00890_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10075_ (.I(\dp.rf.rf[5][31] ),
    .ZN(_04777_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10076_ (.A1(_04482_),
    .A2(_04601_),
    .A3(_04766_),
    .Z(_04778_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10077_ (.A1(_04777_),
    .A2(_04774_),
    .B1(_04778_),
    .B2(_04603_),
    .ZN(_00891_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10078_ (.I0(_04488_),
    .I1(\dp.rf.rf[5][3] ),
    .S(_04776_),
    .Z(_00892_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10079_ (.I0(_04496_),
    .I1(\dp.rf.rf[5][4] ),
    .S(_04776_),
    .Z(_00893_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10080_ (.I0(_04504_),
    .I1(\dp.rf.rf[5][5] ),
    .S(_04776_),
    .Z(_00894_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10081_ (.I0(_04512_),
    .I1(\dp.rf.rf[5][6] ),
    .S(_04776_),
    .Z(_00895_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10082_ (.I0(_04523_),
    .I1(\dp.rf.rf[5][7] ),
    .S(_04776_),
    .Z(_00896_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10083_ (.I0(_04534_),
    .I1(\dp.rf.rf[5][8] ),
    .S(_04773_),
    .Z(_00897_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10084_ (.I0(_04544_),
    .I1(\dp.rf.rf[5][9] ),
    .S(_04773_),
    .Z(_00898_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10085_ (.A1(_04081_),
    .A2(_04766_),
    .Z(_04779_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _10086_ (.I(_04779_),
    .Z(_04780_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10087_ (.I0(\dp.rf.rf[6][0] ),
    .I1(_04686_),
    .S(_04780_),
    .Z(_00899_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10088_ (.I0(\dp.rf.rf[6][10] ),
    .I1(_04689_),
    .S(_04780_),
    .Z(_00900_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10089_ (.I0(\dp.rf.rf[6][11] ),
    .I1(_04690_),
    .S(_04780_),
    .Z(_00901_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10090_ (.I0(\dp.rf.rf[6][12] ),
    .I1(_04691_),
    .S(_04780_),
    .Z(_00902_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10091_ (.I0(\dp.rf.rf[6][13] ),
    .I1(_04692_),
    .S(_04780_),
    .Z(_00903_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10092_ (.I0(\dp.rf.rf[6][14] ),
    .I1(_04693_),
    .S(_04780_),
    .Z(_00904_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10093_ (.I0(\dp.rf.rf[6][15] ),
    .I1(_04694_),
    .S(_04780_),
    .Z(_00905_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10094_ (.I0(\dp.rf.rf[6][16] ),
    .I1(_04695_),
    .S(_04780_),
    .Z(_00906_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _10095_ (.I(_04779_),
    .Z(_04781_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10096_ (.I0(\dp.rf.rf[6][17] ),
    .I1(_04696_),
    .S(_04781_),
    .Z(_00907_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10097_ (.I0(\dp.rf.rf[6][18] ),
    .I1(_04698_),
    .S(_04781_),
    .Z(_00908_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10098_ (.I0(\dp.rf.rf[6][19] ),
    .I1(_04699_),
    .S(_04781_),
    .Z(_00909_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10099_ (.I0(\dp.rf.rf[6][1] ),
    .I1(_04700_),
    .S(_04781_),
    .Z(_00910_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10100_ (.I0(\dp.rf.rf[6][20] ),
    .I1(_04701_),
    .S(_04781_),
    .Z(_00911_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10101_ (.I0(\dp.rf.rf[6][21] ),
    .I1(_04702_),
    .S(_04781_),
    .Z(_00912_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10102_ (.I0(\dp.rf.rf[6][22] ),
    .I1(_04703_),
    .S(_04781_),
    .Z(_00913_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10103_ (.I0(\dp.rf.rf[6][23] ),
    .I1(_04704_),
    .S(_04781_),
    .Z(_00914_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10104_ (.I0(\dp.rf.rf[6][24] ),
    .I1(_04705_),
    .S(_04781_),
    .Z(_00915_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10105_ (.I0(\dp.rf.rf[6][25] ),
    .I1(_04706_),
    .S(_04781_),
    .Z(_00916_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _10106_ (.I(_04779_),
    .Z(_04782_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10107_ (.I0(\dp.rf.rf[6][26] ),
    .I1(_04707_),
    .S(_04782_),
    .Z(_00917_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10108_ (.I0(\dp.rf.rf[6][27] ),
    .I1(_04709_),
    .S(_04782_),
    .Z(_00918_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10109_ (.I0(\dp.rf.rf[6][28] ),
    .I1(_04710_),
    .S(_04782_),
    .Z(_00919_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10110_ (.I0(\dp.rf.rf[6][29] ),
    .I1(_04711_),
    .S(_04782_),
    .Z(_00920_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10111_ (.I0(\dp.rf.rf[6][2] ),
    .I1(_04712_),
    .S(_04782_),
    .Z(_00921_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10112_ (.I0(\dp.rf.rf[6][30] ),
    .I1(_04713_),
    .S(_04782_),
    .Z(_00922_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10113_ (.A1(_04678_),
    .A2(_04780_),
    .Z(_04783_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10114_ (.A1(\dp.rf.rf[6][31] ),
    .A2(_04780_),
    .ZN(_04784_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10115_ (.A1(_04603_),
    .A2(_04783_),
    .B(_04784_),
    .ZN(_00923_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10116_ (.I0(\dp.rf.rf[6][3] ),
    .I1(_04716_),
    .S(_04782_),
    .Z(_00924_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10117_ (.I0(\dp.rf.rf[6][4] ),
    .I1(_04717_),
    .S(_04782_),
    .Z(_00925_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10118_ (.I0(\dp.rf.rf[6][5] ),
    .I1(_04718_),
    .S(_04782_),
    .Z(_00926_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10119_ (.I0(\dp.rf.rf[6][6] ),
    .I1(_04719_),
    .S(_04782_),
    .Z(_00927_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10120_ (.I0(\dp.rf.rf[6][7] ),
    .I1(_04720_),
    .S(_04779_),
    .Z(_00928_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10121_ (.I0(\dp.rf.rf[6][8] ),
    .I1(_04721_),
    .S(_04779_),
    .Z(_00929_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10122_ (.I0(\dp.rf.rf[6][9] ),
    .I1(_04722_),
    .S(_04779_),
    .Z(_00930_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10123_ (.A1(_04545_),
    .A2(_04766_),
    .Z(_04785_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _10124_ (.I(_04785_),
    .Z(_04786_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10125_ (.I0(\dp.rf.rf[7][0] ),
    .I1(_04686_),
    .S(_04786_),
    .Z(_00931_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10126_ (.I0(\dp.rf.rf[7][10] ),
    .I1(_04689_),
    .S(_04786_),
    .Z(_00932_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10127_ (.I0(\dp.rf.rf[7][11] ),
    .I1(_04690_),
    .S(_04786_),
    .Z(_00933_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10128_ (.I0(\dp.rf.rf[7][12] ),
    .I1(_04691_),
    .S(_04786_),
    .Z(_00934_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10129_ (.I0(\dp.rf.rf[7][13] ),
    .I1(_04692_),
    .S(_04786_),
    .Z(_00935_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10130_ (.I0(\dp.rf.rf[7][14] ),
    .I1(_04693_),
    .S(_04786_),
    .Z(_00936_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10131_ (.I0(\dp.rf.rf[7][15] ),
    .I1(_04694_),
    .S(_04786_),
    .Z(_00937_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10132_ (.I0(\dp.rf.rf[7][16] ),
    .I1(_04695_),
    .S(_04786_),
    .Z(_00938_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _10133_ (.I(_04785_),
    .Z(_04787_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10134_ (.I0(\dp.rf.rf[7][17] ),
    .I1(_04696_),
    .S(_04787_),
    .Z(_00939_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10135_ (.I0(\dp.rf.rf[7][18] ),
    .I1(_04698_),
    .S(_04787_),
    .Z(_00940_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10136_ (.I0(\dp.rf.rf[7][19] ),
    .I1(_04699_),
    .S(_04787_),
    .Z(_00941_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10137_ (.I0(\dp.rf.rf[7][1] ),
    .I1(_04700_),
    .S(_04787_),
    .Z(_00942_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10138_ (.I0(\dp.rf.rf[7][20] ),
    .I1(_04701_),
    .S(_04787_),
    .Z(_00943_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10139_ (.I0(\dp.rf.rf[7][21] ),
    .I1(_04702_),
    .S(_04787_),
    .Z(_00944_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10140_ (.I0(\dp.rf.rf[7][22] ),
    .I1(_04703_),
    .S(_04787_),
    .Z(_00945_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10141_ (.I0(\dp.rf.rf[7][23] ),
    .I1(_04704_),
    .S(_04787_),
    .Z(_00946_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10142_ (.I0(\dp.rf.rf[7][24] ),
    .I1(_04705_),
    .S(_04787_),
    .Z(_00947_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10143_ (.I0(\dp.rf.rf[7][25] ),
    .I1(_04706_),
    .S(_04787_),
    .Z(_00948_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _10144_ (.I(_04785_),
    .Z(_04788_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10145_ (.I0(\dp.rf.rf[7][26] ),
    .I1(_04707_),
    .S(_04788_),
    .Z(_00949_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10146_ (.I0(\dp.rf.rf[7][27] ),
    .I1(_04709_),
    .S(_04788_),
    .Z(_00950_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10147_ (.I0(\dp.rf.rf[7][28] ),
    .I1(_04710_),
    .S(_04788_),
    .Z(_00951_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10148_ (.I0(\dp.rf.rf[7][29] ),
    .I1(_04711_),
    .S(_04788_),
    .Z(_00952_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10149_ (.I0(\dp.rf.rf[7][2] ),
    .I1(_04712_),
    .S(_04788_),
    .Z(_00953_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10150_ (.I0(\dp.rf.rf[7][30] ),
    .I1(_04713_),
    .S(_04788_),
    .Z(_00954_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10151_ (.A1(_04482_),
    .A2(_04786_),
    .Z(_04789_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10152_ (.A1(\dp.rf.rf[7][31] ),
    .A2(_04786_),
    .ZN(_04790_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10153_ (.A1(_04603_),
    .A2(_04789_),
    .B(_04790_),
    .ZN(_00955_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10154_ (.I0(\dp.rf.rf[7][3] ),
    .I1(_04716_),
    .S(_04788_),
    .Z(_00956_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10155_ (.I0(\dp.rf.rf[7][4] ),
    .I1(_04717_),
    .S(_04788_),
    .Z(_00957_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10156_ (.I0(\dp.rf.rf[7][5] ),
    .I1(_04718_),
    .S(_04788_),
    .Z(_00958_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10157_ (.I0(\dp.rf.rf[7][6] ),
    .I1(_04719_),
    .S(_04788_),
    .Z(_00959_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10158_ (.I0(\dp.rf.rf[7][7] ),
    .I1(_04720_),
    .S(_04785_),
    .Z(_00960_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10159_ (.I0(\dp.rf.rf[7][8] ),
    .I1(_04721_),
    .S(_04785_),
    .Z(_00961_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10160_ (.I0(\dp.rf.rf[7][9] ),
    .I1(_04722_),
    .S(_04785_),
    .Z(_00962_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10161_ (.A1(_04075_),
    .A2(_04558_),
    .Z(_04791_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _10162_ (.I(_04791_),
    .Z(_04792_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10163_ (.I0(\dp.rf.rf[8][0] ),
    .I1(_04072_),
    .S(_04792_),
    .Z(_00963_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10164_ (.I0(\dp.rf.rf[8][10] ),
    .I1(_04119_),
    .S(_04792_),
    .Z(_00964_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10165_ (.I0(\dp.rf.rf[8][11] ),
    .I1(_04149_),
    .S(_04792_),
    .Z(_00965_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10166_ (.I0(\dp.rf.rf[8][12] ),
    .I1(_04163_),
    .S(_04792_),
    .Z(_00966_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10167_ (.I0(\dp.rf.rf[8][13] ),
    .I1(_04177_),
    .S(_04792_),
    .Z(_00967_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10168_ (.I0(\dp.rf.rf[8][14] ),
    .I1(_04195_),
    .S(_04792_),
    .Z(_00968_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10169_ (.I0(\dp.rf.rf[8][15] ),
    .I1(_04208_),
    .S(_04792_),
    .Z(_00969_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10170_ (.I0(\dp.rf.rf[8][16] ),
    .I1(_04226_),
    .S(_04792_),
    .Z(_00970_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _10171_ (.I(_04791_),
    .Z(_04793_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10172_ (.I0(\dp.rf.rf[8][17] ),
    .I1(_04243_),
    .S(_04793_),
    .Z(_00971_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10173_ (.I0(\dp.rf.rf[8][18] ),
    .I1(_04258_),
    .S(_04793_),
    .Z(_00972_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10174_ (.I0(\dp.rf.rf[8][19] ),
    .I1(_04269_),
    .S(_04793_),
    .Z(_00973_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10175_ (.I0(\dp.rf.rf[8][1] ),
    .I1(_04274_),
    .S(_04793_),
    .Z(_00974_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10176_ (.I0(\dp.rf.rf[8][20] ),
    .I1(_04291_),
    .S(_04793_),
    .Z(_00975_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10177_ (.I0(\dp.rf.rf[8][21] ),
    .I1(_04312_),
    .S(_04793_),
    .Z(_00976_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10178_ (.I0(\dp.rf.rf[8][22] ),
    .I1(_04327_),
    .S(_04793_),
    .Z(_00977_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10179_ (.I0(\dp.rf.rf[8][23] ),
    .I1(_04341_),
    .S(_04793_),
    .Z(_00978_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10180_ (.I0(\dp.rf.rf[8][24] ),
    .I1(_04358_),
    .S(_04793_),
    .Z(_00979_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10181_ (.I0(\dp.rf.rf[8][25] ),
    .I1(_04380_),
    .S(_04793_),
    .Z(_00980_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _10182_ (.I(_04791_),
    .Z(_04794_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10183_ (.I0(\dp.rf.rf[8][26] ),
    .I1(_04394_),
    .S(_04794_),
    .Z(_00981_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10184_ (.I0(\dp.rf.rf[8][27] ),
    .I1(_04408_),
    .S(_04794_),
    .Z(_00982_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10185_ (.I0(\dp.rf.rf[8][28] ),
    .I1(_04420_),
    .S(_04794_),
    .Z(_00983_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10186_ (.I0(\dp.rf.rf[8][29] ),
    .I1(_04438_),
    .S(_04794_),
    .Z(_00984_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10187_ (.I0(\dp.rf.rf[8][2] ),
    .I1(_04445_),
    .S(_04794_),
    .Z(_00985_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10188_ (.I0(\dp.rf.rf[8][30] ),
    .I1(_04461_),
    .S(_04794_),
    .Z(_00986_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10189_ (.A1(_04482_),
    .A2(_04792_),
    .Z(_04795_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10190_ (.A1(\dp.rf.rf[8][31] ),
    .A2(_04792_),
    .ZN(_04796_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10191_ (.A1(_04603_),
    .A2(_04795_),
    .B(_04796_),
    .ZN(_00987_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10192_ (.I0(\dp.rf.rf[8][3] ),
    .I1(_04487_),
    .S(_04794_),
    .Z(_00988_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10193_ (.I0(\dp.rf.rf[8][4] ),
    .I1(_04495_),
    .S(_04794_),
    .Z(_00989_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10194_ (.I0(\dp.rf.rf[8][5] ),
    .I1(_04503_),
    .S(_04794_),
    .Z(_00990_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10195_ (.I0(\dp.rf.rf[8][6] ),
    .I1(_04511_),
    .S(_04794_),
    .Z(_00991_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10196_ (.I0(\dp.rf.rf[8][7] ),
    .I1(_04522_),
    .S(_04791_),
    .Z(_00992_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10197_ (.I0(\dp.rf.rf[8][8] ),
    .I1(_04533_),
    .S(_04791_),
    .Z(_00993_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10198_ (.I0(\dp.rf.rf[8][9] ),
    .I1(_04543_),
    .S(_04791_),
    .Z(_00994_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10199_ (.A1(_04075_),
    .A2(_04595_),
    .ZN(_04797_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _10200_ (.I(_04797_),
    .Z(_04798_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10201_ (.I0(_04073_),
    .I1(\dp.rf.rf[9][0] ),
    .S(_04798_),
    .Z(_00995_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10202_ (.I0(_04120_),
    .I1(\dp.rf.rf[9][10] ),
    .S(_04798_),
    .Z(_00996_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10203_ (.I0(_04150_),
    .I1(\dp.rf.rf[9][11] ),
    .S(_04798_),
    .Z(_00997_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10204_ (.I0(_04164_),
    .I1(\dp.rf.rf[9][12] ),
    .S(_04798_),
    .Z(_00998_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10205_ (.I0(_04178_),
    .I1(\dp.rf.rf[9][13] ),
    .S(_04798_),
    .Z(_00999_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10206_ (.I0(_04196_),
    .I1(\dp.rf.rf[9][14] ),
    .S(_04798_),
    .Z(_01000_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10207_ (.I0(_04209_),
    .I1(\dp.rf.rf[9][15] ),
    .S(_04798_),
    .Z(_01001_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10208_ (.I0(_04227_),
    .I1(\dp.rf.rf[9][16] ),
    .S(_04798_),
    .Z(_01002_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10209_ (.I0(_04244_),
    .I1(\dp.rf.rf[9][17] ),
    .S(_04798_),
    .Z(_01003_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _10210_ (.I(_04797_),
    .Z(_04799_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10211_ (.I0(_04259_),
    .I1(\dp.rf.rf[9][18] ),
    .S(_04799_),
    .Z(_01004_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10212_ (.I0(_04270_),
    .I1(\dp.rf.rf[9][19] ),
    .S(_04799_),
    .Z(_01005_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10213_ (.I0(_04275_),
    .I1(\dp.rf.rf[9][1] ),
    .S(_04799_),
    .Z(_01006_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10214_ (.I0(_04292_),
    .I1(\dp.rf.rf[9][20] ),
    .S(_04799_),
    .Z(_01007_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10215_ (.I0(_04313_),
    .I1(\dp.rf.rf[9][21] ),
    .S(_04799_),
    .Z(_01008_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10216_ (.I0(_04328_),
    .I1(\dp.rf.rf[9][22] ),
    .S(_04799_),
    .Z(_01009_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10217_ (.I0(_04342_),
    .I1(\dp.rf.rf[9][23] ),
    .S(_04799_),
    .Z(_01010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10218_ (.I0(_04359_),
    .I1(\dp.rf.rf[9][24] ),
    .S(_04799_),
    .Z(_01011_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10219_ (.I0(_04381_),
    .I1(\dp.rf.rf[9][25] ),
    .S(_04799_),
    .Z(_01012_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10220_ (.I0(_04395_),
    .I1(\dp.rf.rf[9][26] ),
    .S(_04799_),
    .Z(_01013_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _10221_ (.I(_04797_),
    .Z(_04800_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10222_ (.I0(_04409_),
    .I1(\dp.rf.rf[9][27] ),
    .S(_04800_),
    .Z(_01014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10223_ (.I0(_04421_),
    .I1(\dp.rf.rf[9][28] ),
    .S(_04800_),
    .Z(_01015_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10224_ (.I0(_04439_),
    .I1(\dp.rf.rf[9][29] ),
    .S(_04800_),
    .Z(_01016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10225_ (.I0(_04446_),
    .I1(\dp.rf.rf[9][2] ),
    .S(_04800_),
    .Z(_01017_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10226_ (.I0(_04462_),
    .I1(\dp.rf.rf[9][30] ),
    .S(_04800_),
    .Z(_01018_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10227_ (.I(\dp.rf.rf[9][31] ),
    .ZN(_04801_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10228_ (.A1(_04075_),
    .A2(_04481_),
    .A3(_04601_),
    .Z(_04802_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10229_ (.A1(_04801_),
    .A2(_04798_),
    .B1(_04802_),
    .B2(_04471_),
    .ZN(_01019_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10230_ (.I0(_04488_),
    .I1(\dp.rf.rf[9][3] ),
    .S(_04800_),
    .Z(_01020_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10231_ (.I0(_04496_),
    .I1(\dp.rf.rf[9][4] ),
    .S(_04800_),
    .Z(_01021_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10232_ (.I0(_04504_),
    .I1(\dp.rf.rf[9][5] ),
    .S(_04800_),
    .Z(_01022_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10233_ (.I0(_04512_),
    .I1(\dp.rf.rf[9][6] ),
    .S(_04800_),
    .Z(_01023_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10234_ (.I0(_04523_),
    .I1(\dp.rf.rf[9][7] ),
    .S(_04800_),
    .Z(_01024_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10235_ (.I0(_04534_),
    .I1(\dp.rf.rf[9][8] ),
    .S(_04797_),
    .Z(_01025_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10236_ (.I0(_04544_),
    .I1(\dp.rf.rf[9][9] ),
    .S(_04797_),
    .Z(_01026_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _10237_ (.A1(_04161_),
    .A2(_04059_),
    .ZN(_04803_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _10238_ (.I(_04803_),
    .Z(_04804_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10239_ (.I0(_04112_),
    .I1(_04117_),
    .S(_04804_),
    .Z(\dp.ISRmux.d0[10] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10240_ (.I0(_04142_),
    .I1(_04147_),
    .S(_04804_),
    .Z(\dp.ISRmux.d0[11] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10241_ (.I0(_04158_),
    .I1(_04160_),
    .S(_04804_),
    .Z(\dp.ISRmux.d0[12] ));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10242_ (.A1(_04182_),
    .A2(_04059_),
    .A3(_04175_),
    .Z(_04805_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10243_ (.A1(_04804_),
    .A2(_04173_),
    .B(_04805_),
    .ZN(\dp.ISRmux.d0[13] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10244_ (.I0(_04185_),
    .I1(_04193_),
    .S(_04061_),
    .Z(\dp.ISRmux.d0[14] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10245_ (.I0(_04200_),
    .I1(_04203_),
    .S(_04804_),
    .Z(\dp.ISRmux.d0[15] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10246_ (.I0(_04220_),
    .I1(_04224_),
    .S(_04061_),
    .Z(\dp.ISRmux.d0[16] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10247_ (.I0(_04234_),
    .I1(_04241_),
    .S(_04061_),
    .Z(\dp.ISRmux.d0[17] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10248_ (.I0(_04251_),
    .I1(_04256_),
    .S(_04061_),
    .Z(\dp.ISRmux.d0[18] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10249_ (.I0(_04264_),
    .I1(_04267_),
    .S(_04061_),
    .Z(\dp.ISRmux.d0[19] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10250_ (.I0(_04286_),
    .I1(_04289_),
    .S(_04804_),
    .Z(\dp.ISRmux.d0[20] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10251_ (.I0(_04307_),
    .I1(_04310_),
    .S(_04804_),
    .Z(\dp.ISRmux.d0[21] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10252_ (.I0(_04323_),
    .I1(_04325_),
    .S(_04804_),
    .Z(\dp.ISRmux.d0[22] ));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10253_ (.A1(_04182_),
    .A2(_04059_),
    .A3(_04340_),
    .Z(_04806_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10254_ (.A1(_04804_),
    .A2(_04333_),
    .B(_04806_),
    .ZN(\dp.ISRmux.d0[23] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10255_ (.I0(_04350_),
    .I1(_04356_),
    .S(_04061_),
    .Z(\dp.ISRmux.d0[24] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10256_ (.I0(_04365_),
    .I1(_04378_),
    .S(_04060_),
    .Z(\dp.ISRmux.d0[25] ));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10257_ (.A1(_04182_),
    .A2(_04059_),
    .A3(_04390_),
    .Z(_04807_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10258_ (.A1(_04804_),
    .A2(_04388_),
    .B(_04807_),
    .ZN(\dp.ISRmux.d0[26] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10259_ (.I0(_04404_),
    .I1(_04406_),
    .S(_04803_),
    .Z(\dp.ISRmux.d0[27] ));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _10260_ (.A1(_04182_),
    .A2(_04059_),
    .A3(_04415_),
    .ZN(_04808_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10261_ (.A1(_04061_),
    .A2(_04412_),
    .B(_04808_),
    .ZN(\dp.ISRmux.d0[28] ));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10262_ (.A1(_05196_),
    .A2(_04428_),
    .Z(_04809_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10263_ (.I0(_04432_),
    .I1(_04809_),
    .S(_04060_),
    .Z(\dp.ISRmux.d0[29] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10264_ (.I0(_04442_),
    .I1(_04443_),
    .S(_04060_),
    .Z(\dp.ISRmux.d0[2] ));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _10265_ (.A1(_04182_),
    .A2(_04059_),
    .A3(_04459_),
    .ZN(_04810_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10266_ (.A1(_04061_),
    .A2(_04453_),
    .B(_04810_),
    .ZN(\dp.ISRmux.d0[30] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10267_ (.I0(_04470_),
    .I1(_04474_),
    .S(_04803_),
    .Z(\dp.ISRmux.d0[31] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10268_ (.I0(_05092_),
    .I1(_04485_),
    .S(_04060_),
    .Z(\dp.ISRmux.d0[3] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10269_ (.I0(_04492_),
    .I1(_04493_),
    .S(_04060_),
    .Z(\dp.ISRmux.d0[4] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10270_ (.I0(_04499_),
    .I1(_04501_),
    .S(_04803_),
    .Z(\dp.ISRmux.d0[5] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10271_ (.I0(_04505_),
    .I1(_04507_),
    .S(_04803_),
    .Z(\dp.ISRmux.d0[6] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10272_ (.I0(_04519_),
    .I1(_04516_),
    .S(_04060_),
    .Z(\dp.ISRmux.d0[7] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10273_ (.I0(_04529_),
    .I1(_04531_),
    .S(_04803_),
    .Z(\dp.ISRmux.d0[8] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10274_ (.I0(_04539_),
    .I1(_04541_),
    .S(_04803_),
    .Z(\dp.ISRmux.d0[9] ));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10275_ (.A1(net22),
    .A2(_01079_),
    .A3(_01081_),
    .Z(net127));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10276_ (.A1(net94),
    .A2(_03015_),
    .ZN(_04811_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10277_ (.A1(net275),
    .A2(_04811_),
    .Z(net129));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10278_ (.A1(_02375_),
    .A2(_04811_),
    .Z(net130));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10279_ (.A1(net94),
    .A2(_03015_),
    .B(_02336_),
    .ZN(net131));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10280_ (.A1(_03876_),
    .A2(_04811_),
    .Z(net132));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10281_ (.A1(_02244_),
    .A2(_04811_),
    .Z(net133));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10282_ (.A1(_03940_),
    .A2(_04811_),
    .Z(net134));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10283_ (.A1(_01068_),
    .A2(net94),
    .Z(_04812_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _10284_ (.I(_04812_),
    .Z(_04813_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10285_ (.A1(net255),
    .A2(_04813_),
    .ZN(net135));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10286_ (.A1(_02095_),
    .A2(_04813_),
    .ZN(net136));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10287_ (.A1(_02050_),
    .A2(_04813_),
    .ZN(net137));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10288_ (.A1(_01989_),
    .A2(_04813_),
    .ZN(net138));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10289_ (.A1(_01938_),
    .A2(_04813_),
    .ZN(net140));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10290_ (.A1(_01886_),
    .A2(_04813_),
    .ZN(net141));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10291_ (.A1(_01841_),
    .A2(_04813_),
    .ZN(net142));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10292_ (.A1(_01785_),
    .A2(_04813_),
    .ZN(net143));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10293_ (.A1(_03995_),
    .A2(_04813_),
    .ZN(net144));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10294_ (.A1(_01683_),
    .A2(_04813_),
    .ZN(net145));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10295_ (.A1(_01621_),
    .A2(_04812_),
    .ZN(net146));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10296_ (.A1(_01565_),
    .A2(_04812_),
    .ZN(net147));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10297_ (.A1(_01489_),
    .A2(_04812_),
    .ZN(net148));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10298_ (.A1(_01412_),
    .A2(_04812_),
    .ZN(net149));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10299_ (.A1(_01321_),
    .A2(_04812_),
    .ZN(net151));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10300_ (.A1(_01284_),
    .A2(_04812_),
    .ZN(net152));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10301_ (.A1(_02516_),
    .A2(_04811_),
    .Z(net158));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10302_ (.A1(_02477_),
    .A2(_04811_),
    .Z(net159));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _10303_ (.A(_04814_),
    .B(_04815_),
    .CI(_04816_),
    .CO(_04817_),
    .S(_04818_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _10304_ (.A(_04819_),
    .B(_04820_),
    .CI(_04821_),
    .CO(_04822_),
    .S(_04823_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10305_ (.A(net169),
    .B(_04825_),
    .CO(_04826_),
    .S(_04827_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10306_ (.A(_04828_),
    .B(_04829_),
    .CO(_04830_),
    .S(_04831_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10307_ (.A(_04832_),
    .B(_04833_),
    .CO(_04834_),
    .S(_04835_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10308_ (.A(_04836_),
    .B(_04837_),
    .CO(_04838_),
    .S(_04839_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10309_ (.A(_04840_),
    .B(_04841_),
    .CO(_04842_),
    .S(_04843_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10310_ (.A(_04844_),
    .B(_04845_),
    .CO(_04846_),
    .S(_04847_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10311_ (.A(_04848_),
    .B(_04849_),
    .CO(_04850_),
    .S(_04851_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10312_ (.A(_04852_),
    .B(_04853_),
    .CO(_04854_),
    .S(_04855_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10313_ (.A(_04856_),
    .B(_04857_),
    .CO(_04858_),
    .S(_04859_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10314_ (.A(_04860_),
    .B(_04861_),
    .CO(_04862_),
    .S(_04863_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10315_ (.A(_04864_),
    .B(_04865_),
    .CO(_04866_),
    .S(_04867_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10316_ (.A(_04868_),
    .B(_04869_),
    .CO(_04870_),
    .S(_04871_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10317_ (.A(_04872_),
    .B(_04873_),
    .CO(_04874_),
    .S(_04875_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10318_ (.A(_04876_),
    .B(_04877_),
    .CO(_04878_),
    .S(_04879_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10319_ (.A(_04880_),
    .B(_04881_),
    .CO(_04882_),
    .S(_04883_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10320_ (.A(_04884_),
    .B(_04885_),
    .CO(_04886_),
    .S(_04887_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10321_ (.A(_04888_),
    .B(_04889_),
    .CO(_04890_),
    .S(_04891_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10322_ (.A(_04892_),
    .B(_04893_),
    .CO(_04894_),
    .S(_04895_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10323_ (.A(_04896_),
    .B(_04897_),
    .CO(_04898_),
    .S(_04899_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10324_ (.A(_04900_),
    .B(_04901_),
    .CO(_04902_),
    .S(_04903_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10325_ (.A(_04904_),
    .B(_04905_),
    .CO(_04906_),
    .S(_04907_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10326_ (.A(_04908_),
    .B(_04909_),
    .CO(_04910_),
    .S(_04911_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10327_ (.A(_04912_),
    .B(_04913_),
    .CO(_04914_),
    .S(_04915_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10328_ (.A(_04916_),
    .B(_04917_),
    .CO(_04918_),
    .S(_04919_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10329_ (.A(_04920_),
    .B(_04921_),
    .CO(_04922_),
    .S(_04923_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10330_ (.A(_04924_),
    .B(_04925_),
    .CO(_04926_),
    .S(_04927_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10331_ (.A(_04928_),
    .B(_04929_),
    .CO(_04930_),
    .S(_04931_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10332_ (.A(_04932_),
    .B(_04933_),
    .CO(_04934_),
    .S(_04935_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10333_ (.A(_04936_),
    .B(_04937_),
    .CO(_04938_),
    .S(_04939_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10334_ (.A(_04940_),
    .B(_04941_),
    .CO(_04942_),
    .S(_04943_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10335_ (.A(_04944_),
    .B(_04945_),
    .CO(_04946_),
    .S(_04947_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10336_ (.A(_04948_),
    .B(_04949_),
    .CO(_04950_),
    .S(_04951_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10337_ (.A(_04952_),
    .B(_04953_),
    .CO(_04954_),
    .S(_04955_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10338_ (.A(_04956_),
    .B(_04957_),
    .CO(_04958_),
    .S(_04959_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10339_ (.A(_04960_),
    .B(_04961_),
    .CO(_04962_),
    .S(_04963_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10340_ (.A(_04964_),
    .B(_04965_),
    .CO(_04966_),
    .S(_04967_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10341_ (.A(_04968_),
    .B(_04969_),
    .CO(_04970_),
    .S(_04971_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10342_ (.A(_04972_),
    .B(_04973_),
    .CO(_04974_),
    .S(_04975_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10343_ (.A(_04976_),
    .B(_04977_),
    .CO(_04978_),
    .S(_04979_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10344_ (.A(_04980_),
    .B(_04981_),
    .CO(_04982_),
    .S(_04983_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10345_ (.A(_04984_),
    .B(_04985_),
    .CO(_04986_),
    .S(_04987_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10346_ (.A(_04988_),
    .B(_04989_),
    .CO(_04990_),
    .S(_04991_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10347_ (.A(_04992_),
    .B(_04993_),
    .CO(_04994_),
    .S(_04995_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10348_ (.A(_04996_),
    .B(_04997_),
    .CO(_04998_),
    .S(_04999_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10349_ (.A(_05000_),
    .B(_05001_),
    .CO(_05002_),
    .S(_05003_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10350_ (.A(_05004_),
    .B(_05005_),
    .CO(_05006_),
    .S(_05007_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10351_ (.A(net181),
    .B(_05009_),
    .CO(_05010_),
    .S(_05011_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10352_ (.A(_05012_),
    .B(_05013_),
    .CO(_05014_),
    .S(_05015_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10353_ (.A(_05017_),
    .B(net170),
    .CO(_05018_),
    .S(_05019_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10354_ (.A(_05020_),
    .B(_05021_),
    .CO(_05022_),
    .S(_05023_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10355_ (.A(_05024_),
    .B(_05025_),
    .CO(_05026_),
    .S(_05027_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10356_ (.A(_05028_),
    .B(_05029_),
    .CO(_05030_),
    .S(_05031_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10357_ (.A(_05032_),
    .B(_05033_),
    .CO(_05034_),
    .S(_05035_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10358_ (.A(_05036_),
    .B(_05037_),
    .CO(_05038_),
    .S(_05039_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10359_ (.A(_05040_),
    .B(_05041_),
    .CO(_05042_),
    .S(_05043_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10360_ (.A(_05044_),
    .B(_05045_),
    .CO(_05046_),
    .S(_05047_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10361_ (.A(_05048_),
    .B(_05049_),
    .CO(_05050_),
    .S(_05051_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10362_ (.A(_05052_),
    .B(_05053_),
    .CO(_05054_),
    .S(_05055_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10363_ (.A(_05056_),
    .B(_05057_),
    .CO(_05058_),
    .S(_05059_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10364_ (.A(_05060_),
    .B(_05061_),
    .CO(_05062_),
    .S(_05063_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10365_ (.A(_05065_),
    .B(net266),
    .CO(_05066_),
    .S(_05067_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10366_ (.A(_05068_),
    .B(_05069_),
    .CO(_05070_),
    .S(_05071_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10367_ (.A(_04815_),
    .B(_04816_),
    .CO(_05072_),
    .S(_05073_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10368_ (.A(_05074_),
    .B(_05075_),
    .CO(_05076_),
    .S(_05077_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10369_ (.A(_05078_),
    .B(_05079_),
    .CO(_04819_),
    .S(_05080_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10370_ (.A(_04820_),
    .B(_04821_),
    .CO(_05081_),
    .S(_05082_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10371_ (.A(_05083_),
    .B(_05084_),
    .CO(_05085_),
    .S(_05086_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10372_ (.A(_05087_),
    .B(_05088_),
    .CO(_05089_),
    .S(_05090_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10373_ (.A(net117),
    .B(net120),
    .CO(_05091_),
    .S(_05092_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10374_ (.A(_05093_),
    .B(_05094_),
    .CO(_05095_),
    .S(_05096_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10375_ (.A(_05097_),
    .B(_05098_),
    .CO(_05099_),
    .S(_05100_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10376_ (.A(_05101_),
    .B(_05102_),
    .CO(_05103_),
    .S(_05104_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10377_ (.A(_05105_),
    .B(_05106_),
    .CO(_05107_),
    .S(_05108_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10378_ (.A(_05109_),
    .B(_05110_),
    .CO(_05111_),
    .S(_05112_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10379_ (.A(_05113_),
    .B(_05114_),
    .CO(_05115_),
    .S(_05116_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10380_ (.A(_05117_),
    .B(_05118_),
    .CO(_05119_),
    .S(_05120_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10381_ (.A(_05121_),
    .B(_05122_),
    .CO(_05123_),
    .S(_05124_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10382_ (.A(_05125_),
    .B(_05126_),
    .CO(_05127_),
    .S(_05128_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10383_ (.A(_05129_),
    .B(_05130_),
    .CO(_05131_),
    .S(_05132_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10384_ (.A(_05133_),
    .B(_05134_),
    .CO(_05135_),
    .S(_05136_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10385_ (.A(_05137_),
    .B(_05138_),
    .CO(_05139_),
    .S(_05140_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10386_ (.A(_05141_),
    .B(_05142_),
    .CO(_05143_),
    .S(_05144_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10387_ (.A(_05145_),
    .B(_05146_),
    .CO(_05147_),
    .S(_05148_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10388_ (.A(_05149_),
    .B(_05150_),
    .CO(_05151_),
    .S(_05152_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10389_ (.A(_05153_),
    .B(_05154_),
    .CO(_05155_),
    .S(_05156_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10390_ (.A(_05157_),
    .B(_05158_),
    .CO(_05159_),
    .S(_05160_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10391_ (.A(_05161_),
    .B(_05162_),
    .CO(_05163_),
    .S(_05164_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10392_ (.A(_05165_),
    .B(_05166_),
    .CO(_05167_),
    .S(_05168_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10393_ (.A(_05169_),
    .B(_05170_),
    .CO(_05171_),
    .S(_05172_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10394_ (.A(_05173_),
    .B(_05174_),
    .CO(_05175_),
    .S(_05176_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10395_ (.A(_05177_),
    .B(_05178_),
    .CO(_05179_),
    .S(_05180_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10396_ (.A(_05181_),
    .B(_05182_),
    .CO(_05183_),
    .S(_05184_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10397_ (.A(_05185_),
    .B(_05186_),
    .CO(_05187_),
    .S(_05188_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10398_ (.A(_05189_),
    .B(_05190_),
    .CO(_05191_),
    .S(_05192_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10399_ (.A(_05193_),
    .B(_05194_),
    .CO(_05195_),
    .S(_05196_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _10400_ (.A(_05197_),
    .B(_05198_),
    .CO(_05199_),
    .S(_05200_));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[0]$_DFFE_PP0P_  (.D(_00001_),
    .RN(_00000_),
    .CLK(clknet_leaf_25_clk),
    .Q(net95));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[10]$_DFF_PP0_  (.D(\dp.ISRmux.d0[10] ),
    .RN(_00000_),
    .CLK(clknet_leaf_22_clk),
    .Q(net96));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[11]$_DFF_PP0_  (.D(\dp.ISRmux.d0[11] ),
    .RN(_00000_),
    .CLK(clknet_leaf_22_clk),
    .Q(net97));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[12]$_DFF_PP0_  (.D(\dp.ISRmux.d0[12] ),
    .RN(_00000_),
    .CLK(clknet_leaf_22_clk),
    .Q(net98));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[13]$_DFF_PP0_  (.D(\dp.ISRmux.d0[13] ),
    .RN(_00000_),
    .CLK(clknet_leaf_22_clk),
    .Q(net99));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[14]$_DFF_PP0_  (.D(\dp.ISRmux.d0[14] ),
    .RN(_00000_),
    .CLK(clknet_leaf_22_clk),
    .Q(net100));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[15]$_DFF_PP0_  (.D(\dp.ISRmux.d0[15] ),
    .RN(_00000_),
    .CLK(clknet_leaf_22_clk),
    .Q(net101));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[16]$_DFF_PP0_  (.D(\dp.ISRmux.d0[16] ),
    .RN(_00000_),
    .CLK(clknet_leaf_22_clk),
    .Q(net102));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[17]$_DFF_PP0_  (.D(\dp.ISRmux.d0[17] ),
    .RN(_00000_),
    .CLK(clknet_leaf_22_clk),
    .Q(net103));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[18]$_DFF_PP0_  (.D(\dp.ISRmux.d0[18] ),
    .RN(_00000_),
    .CLK(clknet_leaf_22_clk),
    .Q(net104));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[19]$_DFF_PP0_  (.D(\dp.ISRmux.d0[19] ),
    .RN(_00000_),
    .CLK(clknet_leaf_22_clk),
    .Q(net105));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[1]$_DFFE_PP0P_  (.D(_00002_),
    .RN(_00000_),
    .CLK(clknet_leaf_25_clk),
    .Q(net106));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[20]$_DFF_PP0_  (.D(\dp.ISRmux.d0[20] ),
    .RN(_00000_),
    .CLK(clknet_leaf_22_clk),
    .Q(net107));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[21]$_DFF_PP0_  (.D(\dp.ISRmux.d0[21] ),
    .RN(_00000_),
    .CLK(clknet_leaf_22_clk),
    .Q(net108));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[22]$_DFF_PP0_  (.D(\dp.ISRmux.d0[22] ),
    .RN(_00000_),
    .CLK(clknet_leaf_22_clk),
    .Q(net109));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[23]$_DFF_PP0_  (.D(\dp.ISRmux.d0[23] ),
    .RN(_00000_),
    .CLK(clknet_leaf_22_clk),
    .Q(net110));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[24]$_DFF_PP0_  (.D(\dp.ISRmux.d0[24] ),
    .RN(_00000_),
    .CLK(clknet_leaf_22_clk),
    .Q(net111));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[25]$_DFF_PP0_  (.D(\dp.ISRmux.d0[25] ),
    .RN(_00000_),
    .CLK(clknet_leaf_23_clk),
    .Q(net112));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[26]$_DFF_PP0_  (.D(\dp.ISRmux.d0[26] ),
    .RN(_00000_),
    .CLK(clknet_leaf_23_clk),
    .Q(net113));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[27]$_DFF_PP0_  (.D(\dp.ISRmux.d0[27] ),
    .RN(_00000_),
    .CLK(clknet_leaf_23_clk),
    .Q(net114));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[28]$_DFF_PP0_  (.D(\dp.ISRmux.d0[28] ),
    .RN(_00000_),
    .CLK(clknet_leaf_23_clk),
    .Q(net115));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[29]$_DFF_PP0_  (.D(\dp.ISRmux.d0[29] ),
    .RN(_00000_),
    .CLK(clknet_leaf_23_clk),
    .Q(net116));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[2]$_DFF_PP0_  (.D(\dp.ISRmux.d0[2] ),
    .RN(_00000_),
    .CLK(clknet_leaf_25_clk),
    .Q(net117));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[30]$_DFF_PP0_  (.D(\dp.ISRmux.d0[30] ),
    .RN(_00000_),
    .CLK(clknet_leaf_23_clk),
    .Q(net118));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[31]$_DFF_PP0_  (.D(\dp.ISRmux.d0[31] ),
    .RN(_00000_),
    .CLK(clknet_leaf_25_clk),
    .Q(net119));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[3]$_DFF_PP0_  (.D(\dp.ISRmux.d0[3] ),
    .RN(_00000_),
    .CLK(clknet_leaf_25_clk),
    .Q(net120));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[4]$_DFF_PP0_  (.D(\dp.ISRmux.d0[4] ),
    .RN(_00000_),
    .CLK(clknet_leaf_25_clk),
    .Q(net121));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[5]$_DFF_PP0_  (.D(\dp.ISRmux.d0[5] ),
    .RN(_00000_),
    .CLK(clknet_leaf_25_clk),
    .Q(net122));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[6]$_DFF_PP0_  (.D(\dp.ISRmux.d0[6] ),
    .RN(_00000_),
    .CLK(clknet_leaf_25_clk),
    .Q(net123));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[7]$_DFF_PP0_  (.D(\dp.ISRmux.d0[7] ),
    .RN(_00000_),
    .CLK(clknet_leaf_25_clk),
    .Q(net124));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[8]$_DFF_PP0_  (.D(\dp.ISRmux.d0[8] ),
    .RN(_00000_),
    .CLK(clknet_leaf_25_clk),
    .Q(net125));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[9]$_DFF_PP0_  (.D(\dp.ISRmux.d0[9] ),
    .RN(_00000_),
    .CLK(clknet_leaf_25_clk),
    .Q(net126));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][0]$_DFFE_PP_  (.D(_00003_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[0][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][10]$_DFFE_PP_  (.D(_00004_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[0][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][11]$_DFFE_PP_  (.D(_00005_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[0][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][12]$_DFFE_PP_  (.D(_00006_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[0][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][13]$_DFFE_PP_  (.D(_00007_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[0][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][14]$_DFFE_PP_  (.D(_00008_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[0][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][15]$_DFFE_PP_  (.D(_00009_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[0][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][16]$_DFFE_PP_  (.D(_00010_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[0][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][17]$_DFFE_PP_  (.D(_00011_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[0][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][18]$_DFFE_PP_  (.D(_00012_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[0][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][19]$_DFFE_PP_  (.D(_00013_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[0][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][1]$_DFFE_PP_  (.D(_00014_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[0][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][20]$_DFFE_PP_  (.D(_00015_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[0][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][21]$_DFFE_PP_  (.D(_00016_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[0][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][22]$_DFFE_PP_  (.D(_00017_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[0][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][23]$_DFFE_PP_  (.D(_00018_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[0][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][24]$_DFFE_PP_  (.D(_00019_),
    .CLK(clknet_leaf_23_clk),
    .Q(\dp.rf.rf[0][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][25]$_DFFE_PP_  (.D(_00020_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[0][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][26]$_DFFE_PP_  (.D(_00021_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[0][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][27]$_DFFE_PP_  (.D(_00022_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[0][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][28]$_DFFE_PP_  (.D(_00023_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[0][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][29]$_DFFE_PP_  (.D(_00024_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[0][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][2]$_DFFE_PP_  (.D(_00025_),
    .CLK(clknet_leaf_3_clk),
    .Q(\dp.rf.rf[0][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][30]$_DFFE_PP_  (.D(_00026_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[0][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][31]$_DFFE_PP_  (.D(_00027_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[0][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][3]$_DFFE_PP_  (.D(_00028_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[0][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][4]$_DFFE_PP_  (.D(_00029_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[0][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][5]$_DFFE_PP_  (.D(_00030_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[0][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][6]$_DFFE_PP_  (.D(_00031_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[0][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][7]$_DFFE_PP_  (.D(_00032_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[0][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][8]$_DFFE_PP_  (.D(_00033_),
    .CLK(clknet_leaf_3_clk),
    .Q(\dp.rf.rf[0][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][9]$_DFFE_PP_  (.D(_00034_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[0][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][0]$_DFFE_PP_  (.D(_00035_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[10][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][10]$_DFFE_PP_  (.D(_00036_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[10][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][11]$_DFFE_PP_  (.D(_00037_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[10][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][12]$_DFFE_PP_  (.D(_00038_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[10][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][13]$_DFFE_PP_  (.D(_00039_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[10][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][14]$_DFFE_PP_  (.D(_00040_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[10][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][15]$_DFFE_PP_  (.D(_00041_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[10][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][16]$_DFFE_PP_  (.D(_00042_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[10][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][17]$_DFFE_PP_  (.D(_00043_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[10][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][18]$_DFFE_PP_  (.D(_00044_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[10][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][19]$_DFFE_PP_  (.D(_00045_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[10][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][1]$_DFFE_PP_  (.D(_00046_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[10][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][20]$_DFFE_PP_  (.D(_00047_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[10][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][21]$_DFFE_PP_  (.D(_00048_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[10][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][22]$_DFFE_PP_  (.D(_00049_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[10][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][23]$_DFFE_PP_  (.D(_00050_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[10][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][24]$_DFFE_PP_  (.D(_00051_),
    .CLK(clknet_leaf_23_clk),
    .Q(\dp.rf.rf[10][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][25]$_DFFE_PP_  (.D(_00052_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[10][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][26]$_DFFE_PP_  (.D(_00053_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[10][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][27]$_DFFE_PP_  (.D(_00054_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[10][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][28]$_DFFE_PP_  (.D(_00055_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[10][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][29]$_DFFE_PP_  (.D(_00056_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[10][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][2]$_DFFE_PP_  (.D(_00057_),
    .CLK(clknet_leaf_3_clk),
    .Q(\dp.rf.rf[10][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][30]$_DFFE_PP_  (.D(_00058_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[10][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][31]$_DFFE_PP_  (.D(_00059_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[10][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][3]$_DFFE_PP_  (.D(_00060_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[10][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][4]$_DFFE_PP_  (.D(_00061_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[10][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][5]$_DFFE_PP_  (.D(_00062_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[10][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][6]$_DFFE_PP_  (.D(_00063_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[10][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][7]$_DFFE_PP_  (.D(_00064_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[10][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][8]$_DFFE_PP_  (.D(_00065_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[10][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][9]$_DFFE_PP_  (.D(_00066_),
    .CLK(clknet_leaf_3_clk),
    .Q(\dp.rf.rf[10][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][0]$_DFFE_PP_  (.D(_00067_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[11][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][10]$_DFFE_PP_  (.D(_00068_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[11][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][11]$_DFFE_PP_  (.D(_00069_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[11][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][12]$_DFFE_PP_  (.D(_00070_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[11][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][13]$_DFFE_PP_  (.D(_00071_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[11][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][14]$_DFFE_PP_  (.D(_00072_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[11][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][15]$_DFFE_PP_  (.D(_00073_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[11][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][16]$_DFFE_PP_  (.D(_00074_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[11][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][17]$_DFFE_PP_  (.D(_00075_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[11][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][18]$_DFFE_PP_  (.D(_00076_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[11][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][19]$_DFFE_PP_  (.D(_00077_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[11][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][1]$_DFFE_PP_  (.D(_00078_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[11][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][20]$_DFFE_PP_  (.D(_00079_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[11][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][21]$_DFFE_PP_  (.D(_00080_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[11][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][22]$_DFFE_PP_  (.D(_00081_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[11][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][23]$_DFFE_PP_  (.D(_00082_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[11][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][24]$_DFFE_PP_  (.D(_00083_),
    .CLK(clknet_leaf_24_clk),
    .Q(\dp.rf.rf[11][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][25]$_DFFE_PP_  (.D(_00084_),
    .CLK(clknet_leaf_22_clk),
    .Q(\dp.rf.rf[11][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][26]$_DFFE_PP_  (.D(_00085_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[11][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][27]$_DFFE_PP_  (.D(_00086_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[11][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][28]$_DFFE_PP_  (.D(_00087_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[11][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][29]$_DFFE_PP_  (.D(_00088_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[11][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][2]$_DFFE_PP_  (.D(_00089_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[11][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][30]$_DFFE_PP_  (.D(_00090_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[11][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][31]$_DFFE_PP_  (.D(_00091_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[11][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][3]$_DFFE_PP_  (.D(_00092_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[11][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][4]$_DFFE_PP_  (.D(_00093_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[11][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][5]$_DFFE_PP_  (.D(_00094_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[11][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][6]$_DFFE_PP_  (.D(_00095_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[11][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][7]$_DFFE_PP_  (.D(_00096_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[11][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][8]$_DFFE_PP_  (.D(_00097_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[11][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][9]$_DFFE_PP_  (.D(_00098_),
    .CLK(clknet_leaf_3_clk),
    .Q(\dp.rf.rf[11][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][0]$_DFFE_PP_  (.D(_00099_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[12][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][10]$_DFFE_PP_  (.D(_00100_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[12][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][11]$_DFFE_PP_  (.D(_00101_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[12][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][12]$_DFFE_PP_  (.D(_00102_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[12][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][13]$_DFFE_PP_  (.D(_00103_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[12][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][14]$_DFFE_PP_  (.D(_00104_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[12][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][15]$_DFFE_PP_  (.D(_00105_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[12][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][16]$_DFFE_PP_  (.D(_00106_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[12][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][17]$_DFFE_PP_  (.D(_00107_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[12][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][18]$_DFFE_PP_  (.D(_00108_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[12][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][19]$_DFFE_PP_  (.D(_00109_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[12][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][1]$_DFFE_PP_  (.D(_00110_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[12][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][20]$_DFFE_PP_  (.D(_00111_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[12][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][21]$_DFFE_PP_  (.D(_00112_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[12][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][22]$_DFFE_PP_  (.D(_00113_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[12][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][23]$_DFFE_PP_  (.D(_00114_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[12][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][24]$_DFFE_PP_  (.D(_00115_),
    .CLK(clknet_leaf_23_clk),
    .Q(\dp.rf.rf[12][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][25]$_DFFE_PP_  (.D(_00116_),
    .CLK(clknet_leaf_22_clk),
    .Q(\dp.rf.rf[12][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][26]$_DFFE_PP_  (.D(_00117_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[12][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][27]$_DFFE_PP_  (.D(_00118_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[12][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][28]$_DFFE_PP_  (.D(_00119_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[12][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][29]$_DFFE_PP_  (.D(_00120_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[12][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][2]$_DFFE_PP_  (.D(_00121_),
    .CLK(clknet_leaf_3_clk),
    .Q(\dp.rf.rf[12][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][30]$_DFFE_PP_  (.D(_00122_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[12][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][31]$_DFFE_PP_  (.D(_00123_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[12][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][3]$_DFFE_PP_  (.D(_00124_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[12][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][4]$_DFFE_PP_  (.D(_00125_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[12][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][5]$_DFFE_PP_  (.D(_00126_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[12][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][6]$_DFFE_PP_  (.D(_00127_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[12][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][7]$_DFFE_PP_  (.D(_00128_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[12][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][8]$_DFFE_PP_  (.D(_00129_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[12][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][9]$_DFFE_PP_  (.D(_00130_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[12][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][0]$_DFFE_PP_  (.D(_00131_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[13][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][10]$_DFFE_PP_  (.D(_00132_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[13][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][11]$_DFFE_PP_  (.D(_00133_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[13][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][12]$_DFFE_PP_  (.D(_00134_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[13][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][13]$_DFFE_PP_  (.D(_00135_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[13][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][14]$_DFFE_PP_  (.D(_00136_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[13][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][15]$_DFFE_PP_  (.D(_00137_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[13][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][16]$_DFFE_PP_  (.D(_00138_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[13][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][17]$_DFFE_PP_  (.D(_00139_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[13][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][18]$_DFFE_PP_  (.D(_00140_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[13][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][19]$_DFFE_PP_  (.D(_00141_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[13][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][1]$_DFFE_PP_  (.D(_00142_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[13][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][20]$_DFFE_PP_  (.D(_00143_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[13][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][21]$_DFFE_PP_  (.D(_00144_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[13][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][22]$_DFFE_PP_  (.D(_00145_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[13][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][23]$_DFFE_PP_  (.D(_00146_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[13][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][24]$_DFFE_PP_  (.D(_00147_),
    .CLK(clknet_leaf_23_clk),
    .Q(\dp.rf.rf[13][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][25]$_DFFE_PP_  (.D(_00148_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[13][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][26]$_DFFE_PP_  (.D(_00149_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[13][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][27]$_DFFE_PP_  (.D(_00150_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[13][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][28]$_DFFE_PP_  (.D(_00151_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[13][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][29]$_DFFE_PP_  (.D(_00152_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[13][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][2]$_DFFE_PP_  (.D(_00153_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[13][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][30]$_DFFE_PP_  (.D(_00154_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[13][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][31]$_DFFE_PP_  (.D(_00155_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[13][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][3]$_DFFE_PP_  (.D(_00156_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[13][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][4]$_DFFE_PP_  (.D(_00157_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[13][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][5]$_DFFE_PP_  (.D(_00158_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[13][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][6]$_DFFE_PP_  (.D(_00159_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[13][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][7]$_DFFE_PP_  (.D(_00160_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[13][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][8]$_DFFE_PP_  (.D(_00161_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[13][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][9]$_DFFE_PP_  (.D(_00162_),
    .CLK(clknet_leaf_3_clk),
    .Q(\dp.rf.rf[13][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][0]$_DFFE_PP_  (.D(_00163_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[14][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][10]$_DFFE_PP_  (.D(_00164_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[14][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][11]$_DFFE_PP_  (.D(_00165_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[14][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][12]$_DFFE_PP_  (.D(_00166_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[14][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][13]$_DFFE_PP_  (.D(_00167_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[14][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][14]$_DFFE_PP_  (.D(_00168_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[14][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][15]$_DFFE_PP_  (.D(_00169_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[14][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][16]$_DFFE_PP_  (.D(_00170_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[14][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][17]$_DFFE_PP_  (.D(_00171_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[14][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][18]$_DFFE_PP_  (.D(_00172_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[14][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][19]$_DFFE_PP_  (.D(_00173_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[14][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][1]$_DFFE_PP_  (.D(_00174_),
    .CLK(clknet_leaf_24_clk),
    .Q(\dp.rf.rf[14][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][20]$_DFFE_PP_  (.D(_00175_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[14][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][21]$_DFFE_PP_  (.D(_00176_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[14][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][22]$_DFFE_PP_  (.D(_00177_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[14][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][23]$_DFFE_PP_  (.D(_00178_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[14][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][24]$_DFFE_PP_  (.D(_00179_),
    .CLK(clknet_leaf_24_clk),
    .Q(\dp.rf.rf[14][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][25]$_DFFE_PP_  (.D(_00180_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[14][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][26]$_DFFE_PP_  (.D(_00181_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[14][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][27]$_DFFE_PP_  (.D(_00182_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[14][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][28]$_DFFE_PP_  (.D(_00183_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[14][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][29]$_DFFE_PP_  (.D(_00184_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[14][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][2]$_DFFE_PP_  (.D(_00185_),
    .CLK(clknet_leaf_3_clk),
    .Q(\dp.rf.rf[14][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][30]$_DFFE_PP_  (.D(_00186_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[14][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][31]$_DFFE_PP_  (.D(_00187_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[14][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][3]$_DFFE_PP_  (.D(_00188_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[14][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][4]$_DFFE_PP_  (.D(_00189_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[14][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][5]$_DFFE_PP_  (.D(_00190_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[14][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][6]$_DFFE_PP_  (.D(_00191_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[14][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][7]$_DFFE_PP_  (.D(_00192_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[14][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][8]$_DFFE_PP_  (.D(_00193_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[14][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][9]$_DFFE_PP_  (.D(_00194_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[14][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][0]$_DFFE_PP_  (.D(_00195_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[15][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][10]$_DFFE_PP_  (.D(_00196_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[15][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][11]$_DFFE_PP_  (.D(_00197_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[15][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][12]$_DFFE_PP_  (.D(_00198_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[15][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][13]$_DFFE_PP_  (.D(_00199_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[15][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][14]$_DFFE_PP_  (.D(_00200_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[15][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][15]$_DFFE_PP_  (.D(_00201_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[15][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][16]$_DFFE_PP_  (.D(_00202_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[15][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][17]$_DFFE_PP_  (.D(_00203_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[15][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][18]$_DFFE_PP_  (.D(_00204_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[15][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][19]$_DFFE_PP_  (.D(_00205_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[15][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][1]$_DFFE_PP_  (.D(_00206_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[15][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][20]$_DFFE_PP_  (.D(_00207_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[15][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][21]$_DFFE_PP_  (.D(_00208_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[15][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][22]$_DFFE_PP_  (.D(_00209_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[15][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][23]$_DFFE_PP_  (.D(_00210_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[15][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][24]$_DFFE_PP_  (.D(_00211_),
    .CLK(clknet_leaf_24_clk),
    .Q(\dp.rf.rf[15][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][25]$_DFFE_PP_  (.D(_00212_),
    .CLK(clknet_leaf_22_clk),
    .Q(\dp.rf.rf[15][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][26]$_DFFE_PP_  (.D(_00213_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[15][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][27]$_DFFE_PP_  (.D(_00214_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[15][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][28]$_DFFE_PP_  (.D(_00215_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[15][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][29]$_DFFE_PP_  (.D(_00216_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[15][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][2]$_DFFE_PP_  (.D(_00217_),
    .CLK(clknet_leaf_3_clk),
    .Q(\dp.rf.rf[15][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][30]$_DFFE_PP_  (.D(_00218_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[15][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][31]$_DFFE_PP_  (.D(_00219_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[15][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][3]$_DFFE_PP_  (.D(_00220_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[15][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][4]$_DFFE_PP_  (.D(_00221_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[15][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][5]$_DFFE_PP_  (.D(_00222_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[15][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][6]$_DFFE_PP_  (.D(_00223_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[15][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][7]$_DFFE_PP_  (.D(_00224_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[15][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][8]$_DFFE_PP_  (.D(_00225_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[15][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][9]$_DFFE_PP_  (.D(_00226_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[15][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][0]$_DFFE_PP_  (.D(_00227_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[16][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][10]$_DFFE_PP_  (.D(_00228_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[16][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][11]$_DFFE_PP_  (.D(_00229_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[16][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][12]$_DFFE_PP_  (.D(_00230_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[16][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][13]$_DFFE_PP_  (.D(_00231_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[16][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][14]$_DFFE_PP_  (.D(_00232_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[16][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][15]$_DFFE_PP_  (.D(_00233_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[16][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][16]$_DFFE_PP_  (.D(_00234_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[16][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][17]$_DFFE_PP_  (.D(_00235_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[16][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][18]$_DFFE_PP_  (.D(_00236_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[16][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][19]$_DFFE_PP_  (.D(_00237_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[16][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][1]$_DFFE_PP_  (.D(_00238_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[16][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][20]$_DFFE_PP_  (.D(_00239_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[16][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][21]$_DFFE_PP_  (.D(_00240_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[16][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][22]$_DFFE_PP_  (.D(_00241_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[16][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][23]$_DFFE_PP_  (.D(_00242_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[16][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][24]$_DFFE_PP_  (.D(_00243_),
    .CLK(clknet_leaf_23_clk),
    .Q(\dp.rf.rf[16][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][25]$_DFFE_PP_  (.D(_00244_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[16][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][26]$_DFFE_PP_  (.D(_00245_),
    .CLK(clknet_leaf_24_clk),
    .Q(\dp.rf.rf[16][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][27]$_DFFE_PP_  (.D(_00246_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[16][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][28]$_DFFE_PP_  (.D(_00247_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[16][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][29]$_DFFE_PP_  (.D(_00248_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[16][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][2]$_DFFE_PP_  (.D(_00249_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[16][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][30]$_DFFE_PP_  (.D(_00250_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[16][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][31]$_DFFE_PP_  (.D(_00251_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[16][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][3]$_DFFE_PP_  (.D(_00252_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[16][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][4]$_DFFE_PP_  (.D(_00253_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[16][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][5]$_DFFE_PP_  (.D(_00254_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[16][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][6]$_DFFE_PP_  (.D(_00255_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[16][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][7]$_DFFE_PP_  (.D(_00256_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[16][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][8]$_DFFE_PP_  (.D(_00257_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[16][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][9]$_DFFE_PP_  (.D(_00258_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[16][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][0]$_DFFE_PP_  (.D(_00259_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[17][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][10]$_DFFE_PP_  (.D(_00260_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[17][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][11]$_DFFE_PP_  (.D(_00261_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[17][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][12]$_DFFE_PP_  (.D(_00262_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[17][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][13]$_DFFE_PP_  (.D(_00263_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[17][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][14]$_DFFE_PP_  (.D(_00264_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[17][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][15]$_DFFE_PP_  (.D(_00265_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[17][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][16]$_DFFE_PP_  (.D(_00266_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[17][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][17]$_DFFE_PP_  (.D(_00267_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[17][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][18]$_DFFE_PP_  (.D(_00268_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[17][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][19]$_DFFE_PP_  (.D(_00269_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[17][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][1]$_DFFE_PP_  (.D(_00270_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[17][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][20]$_DFFE_PP_  (.D(_00271_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[17][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][21]$_DFFE_PP_  (.D(_00272_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[17][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][22]$_DFFE_PP_  (.D(_00273_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[17][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][23]$_DFFE_PP_  (.D(_00274_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[17][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][24]$_DFFE_PP_  (.D(_00275_),
    .CLK(clknet_leaf_23_clk),
    .Q(\dp.rf.rf[17][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][25]$_DFFE_PP_  (.D(_00276_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[17][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][26]$_DFFE_PP_  (.D(_00277_),
    .CLK(clknet_leaf_24_clk),
    .Q(\dp.rf.rf[17][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][27]$_DFFE_PP_  (.D(_00278_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[17][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][28]$_DFFE_PP_  (.D(_00279_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[17][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][29]$_DFFE_PP_  (.D(_00280_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[17][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][2]$_DFFE_PP_  (.D(_00281_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[17][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][30]$_DFFE_PP_  (.D(_00282_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[17][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][31]$_DFFE_PP_  (.D(_00283_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[17][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][3]$_DFFE_PP_  (.D(_00284_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[17][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][4]$_DFFE_PP_  (.D(_00285_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[17][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][5]$_DFFE_PP_  (.D(_00286_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[17][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][6]$_DFFE_PP_  (.D(_00287_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[17][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][7]$_DFFE_PP_  (.D(_00288_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[17][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][8]$_DFFE_PP_  (.D(_00289_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[17][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][9]$_DFFE_PP_  (.D(_00290_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[17][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][0]$_DFFE_PP_  (.D(_00291_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[18][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][10]$_DFFE_PP_  (.D(_00292_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[18][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][11]$_DFFE_PP_  (.D(_00293_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[18][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][12]$_DFFE_PP_  (.D(_00294_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[18][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][13]$_DFFE_PP_  (.D(_00295_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[18][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][14]$_DFFE_PP_  (.D(_00296_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[18][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][15]$_DFFE_PP_  (.D(_00297_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[18][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][16]$_DFFE_PP_  (.D(_00298_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[18][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][17]$_DFFE_PP_  (.D(_00299_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[18][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][18]$_DFFE_PP_  (.D(_00300_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[18][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][19]$_DFFE_PP_  (.D(_00301_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[18][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][1]$_DFFE_PP_  (.D(_00302_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[18][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][20]$_DFFE_PP_  (.D(_00303_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[18][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][21]$_DFFE_PP_  (.D(_00304_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[18][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][22]$_DFFE_PP_  (.D(_00305_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[18][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][23]$_DFFE_PP_  (.D(_00306_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[18][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][24]$_DFFE_PP_  (.D(_00307_),
    .CLK(clknet_leaf_23_clk),
    .Q(\dp.rf.rf[18][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][25]$_DFFE_PP_  (.D(_00308_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[18][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][26]$_DFFE_PP_  (.D(_00309_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[18][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][27]$_DFFE_PP_  (.D(_00310_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[18][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][28]$_DFFE_PP_  (.D(_00311_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[18][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][29]$_DFFE_PP_  (.D(_00312_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[18][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][2]$_DFFE_PP_  (.D(_00313_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[18][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][30]$_DFFE_PP_  (.D(_00314_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[18][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][31]$_DFFE_PP_  (.D(_00315_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[18][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][3]$_DFFE_PP_  (.D(_00316_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[18][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][4]$_DFFE_PP_  (.D(_00317_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[18][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][5]$_DFFE_PP_  (.D(_00318_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[18][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][6]$_DFFE_PP_  (.D(_00319_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[18][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][7]$_DFFE_PP_  (.D(_00320_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[18][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][8]$_DFFE_PP_  (.D(_00321_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[18][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][9]$_DFFE_PP_  (.D(_00322_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[18][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][0]$_DFFE_PP_  (.D(_00323_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[19][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][10]$_DFFE_PP_  (.D(_00324_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[19][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][11]$_DFFE_PP_  (.D(_00325_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[19][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][12]$_DFFE_PP_  (.D(_00326_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[19][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][13]$_DFFE_PP_  (.D(_00327_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[19][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][14]$_DFFE_PP_  (.D(_00328_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[19][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][15]$_DFFE_PP_  (.D(_00329_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[19][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][16]$_DFFE_PP_  (.D(_00330_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[19][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][17]$_DFFE_PP_  (.D(_00331_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[19][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][18]$_DFFE_PP_  (.D(_00332_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[19][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][19]$_DFFE_PP_  (.D(_00333_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[19][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][1]$_DFFE_PP_  (.D(_00334_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[19][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][20]$_DFFE_PP_  (.D(_00335_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[19][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][21]$_DFFE_PP_  (.D(_00336_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[19][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][22]$_DFFE_PP_  (.D(_00337_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[19][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][23]$_DFFE_PP_  (.D(_00338_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[19][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][24]$_DFFE_PP_  (.D(_00339_),
    .CLK(clknet_leaf_23_clk),
    .Q(\dp.rf.rf[19][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][25]$_DFFE_PP_  (.D(_00340_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[19][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][26]$_DFFE_PP_  (.D(_00341_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[19][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][27]$_DFFE_PP_  (.D(_00342_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[19][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][28]$_DFFE_PP_  (.D(_00343_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[19][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][29]$_DFFE_PP_  (.D(_00344_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[19][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][2]$_DFFE_PP_  (.D(_00345_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[19][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][30]$_DFFE_PP_  (.D(_00346_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[19][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][31]$_DFFE_PP_  (.D(_00347_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[19][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][3]$_DFFE_PP_  (.D(_00348_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[19][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][4]$_DFFE_PP_  (.D(_00349_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[19][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][5]$_DFFE_PP_  (.D(_00350_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[19][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][6]$_DFFE_PP_  (.D(_00351_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[19][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][7]$_DFFE_PP_  (.D(_00352_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[19][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][8]$_DFFE_PP_  (.D(_00353_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[19][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][9]$_DFFE_PP_  (.D(_00354_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[19][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][0]$_DFFE_PP_  (.D(_00355_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[1][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][10]$_DFFE_PP_  (.D(_00356_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[1][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][11]$_DFFE_PP_  (.D(_00357_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[1][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][12]$_DFFE_PP_  (.D(_00358_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[1][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][13]$_DFFE_PP_  (.D(_00359_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[1][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][14]$_DFFE_PP_  (.D(_00360_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[1][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][15]$_DFFE_PP_  (.D(_00361_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[1][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][16]$_DFFE_PP_  (.D(_00362_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[1][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][17]$_DFFE_PP_  (.D(_00363_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[1][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][18]$_DFFE_PP_  (.D(_00364_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[1][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][19]$_DFFE_PP_  (.D(_00365_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[1][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][1]$_DFFE_PP_  (.D(_00366_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[1][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][20]$_DFFE_PP_  (.D(_00367_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[1][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][21]$_DFFE_PP_  (.D(_00368_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[1][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][22]$_DFFE_PP_  (.D(_00369_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[1][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][23]$_DFFE_PP_  (.D(_00370_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[1][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][24]$_DFFE_PP_  (.D(_00371_),
    .CLK(clknet_leaf_23_clk),
    .Q(\dp.rf.rf[1][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][25]$_DFFE_PP_  (.D(_00372_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[1][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][26]$_DFFE_PP_  (.D(_00373_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[1][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][27]$_DFFE_PP_  (.D(_00374_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[1][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][28]$_DFFE_PP_  (.D(_00375_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[1][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][29]$_DFFE_PP_  (.D(_00376_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[1][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][2]$_DFFE_PP_  (.D(_00377_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[1][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][30]$_DFFE_PP_  (.D(_00378_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[1][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][31]$_DFFE_PP_  (.D(_00379_),
    .CLK(clknet_leaf_3_clk),
    .Q(\dp.rf.rf[1][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][3]$_DFFE_PP_  (.D(_00380_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[1][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][4]$_DFFE_PP_  (.D(_00381_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[1][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][5]$_DFFE_PP_  (.D(_00382_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[1][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][6]$_DFFE_PP_  (.D(_00383_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[1][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][7]$_DFFE_PP_  (.D(_00384_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[1][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][8]$_DFFE_PP_  (.D(_00385_),
    .CLK(clknet_leaf_3_clk),
    .Q(\dp.rf.rf[1][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][9]$_DFFE_PP_  (.D(_00386_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[1][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][0]$_DFFE_PP_  (.D(_00387_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[20][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][10]$_DFFE_PP_  (.D(_00388_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[20][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][11]$_DFFE_PP_  (.D(_00389_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[20][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][12]$_DFFE_PP_  (.D(_00390_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[20][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][13]$_DFFE_PP_  (.D(_00391_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[20][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][14]$_DFFE_PP_  (.D(_00392_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[20][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][15]$_DFFE_PP_  (.D(_00393_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[20][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][16]$_DFFE_PP_  (.D(_00394_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[20][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][17]$_DFFE_PP_  (.D(_00395_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[20][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][18]$_DFFE_PP_  (.D(_00396_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[20][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][19]$_DFFE_PP_  (.D(_00397_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[20][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][1]$_DFFE_PP_  (.D(_00398_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[20][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][20]$_DFFE_PP_  (.D(_00399_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[20][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][21]$_DFFE_PP_  (.D(_00400_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[20][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][22]$_DFFE_PP_  (.D(_00401_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[20][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][23]$_DFFE_PP_  (.D(_00402_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[20][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][24]$_DFFE_PP_  (.D(_00403_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[20][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][25]$_DFFE_PP_  (.D(_00404_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[20][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][26]$_DFFE_PP_  (.D(_00405_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[20][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][27]$_DFFE_PP_  (.D(_00406_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[20][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][28]$_DFFE_PP_  (.D(_00407_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[20][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][29]$_DFFE_PP_  (.D(_00408_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[20][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][2]$_DFFE_PP_  (.D(_00409_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[20][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][30]$_DFFE_PP_  (.D(_00410_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[20][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][31]$_DFFE_PP_  (.D(_00411_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[20][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][3]$_DFFE_PP_  (.D(_00412_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[20][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][4]$_DFFE_PP_  (.D(_00413_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[20][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][5]$_DFFE_PP_  (.D(_00414_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[20][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][6]$_DFFE_PP_  (.D(_00415_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[20][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][7]$_DFFE_PP_  (.D(_00416_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[20][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][8]$_DFFE_PP_  (.D(_00417_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[20][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][9]$_DFFE_PP_  (.D(_00418_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[20][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][0]$_DFFE_PP_  (.D(_00419_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[21][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][10]$_DFFE_PP_  (.D(_00420_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[21][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][11]$_DFFE_PP_  (.D(_00421_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[21][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][12]$_DFFE_PP_  (.D(_00422_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[21][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][13]$_DFFE_PP_  (.D(_00423_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[21][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][14]$_DFFE_PP_  (.D(_00424_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[21][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][15]$_DFFE_PP_  (.D(_00425_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[21][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][16]$_DFFE_PP_  (.D(_00426_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[21][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][17]$_DFFE_PP_  (.D(_00427_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[21][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][18]$_DFFE_PP_  (.D(_00428_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[21][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][19]$_DFFE_PP_  (.D(_00429_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[21][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][1]$_DFFE_PP_  (.D(_00430_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[21][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][20]$_DFFE_PP_  (.D(_00431_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[21][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][21]$_DFFE_PP_  (.D(_00432_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[21][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][22]$_DFFE_PP_  (.D(_00433_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[21][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][23]$_DFFE_PP_  (.D(_00434_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[21][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][24]$_DFFE_PP_  (.D(_00435_),
    .CLK(clknet_leaf_24_clk),
    .Q(\dp.rf.rf[21][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][25]$_DFFE_PP_  (.D(_00436_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[21][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][26]$_DFFE_PP_  (.D(_00437_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[21][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][27]$_DFFE_PP_  (.D(_00438_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[21][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][28]$_DFFE_PP_  (.D(_00439_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[21][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][29]$_DFFE_PP_  (.D(_00440_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[21][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][2]$_DFFE_PP_  (.D(_00441_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[21][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][30]$_DFFE_PP_  (.D(_00442_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[21][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][31]$_DFFE_PP_  (.D(_00443_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[21][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][3]$_DFFE_PP_  (.D(_00444_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[21][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][4]$_DFFE_PP_  (.D(_00445_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[21][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][5]$_DFFE_PP_  (.D(_00446_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[21][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][6]$_DFFE_PP_  (.D(_00447_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[21][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][7]$_DFFE_PP_  (.D(_00448_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[21][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][8]$_DFFE_PP_  (.D(_00449_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[21][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][9]$_DFFE_PP_  (.D(_00450_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[21][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][0]$_DFFE_PP_  (.D(_00451_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[22][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][10]$_DFFE_PP_  (.D(_00452_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[22][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][11]$_DFFE_PP_  (.D(_00453_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[22][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][12]$_DFFE_PP_  (.D(_00454_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[22][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][13]$_DFFE_PP_  (.D(_00455_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[22][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][14]$_DFFE_PP_  (.D(_00456_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[22][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][15]$_DFFE_PP_  (.D(_00457_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[22][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][16]$_DFFE_PP_  (.D(_00458_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[22][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][17]$_DFFE_PP_  (.D(_00459_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[22][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][18]$_DFFE_PP_  (.D(_00460_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[22][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][19]$_DFFE_PP_  (.D(_00461_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[22][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][1]$_DFFE_PP_  (.D(_00462_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[22][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][20]$_DFFE_PP_  (.D(_00463_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[22][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][21]$_DFFE_PP_  (.D(_00464_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[22][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][22]$_DFFE_PP_  (.D(_00465_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[22][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][23]$_DFFE_PP_  (.D(_00466_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[22][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][24]$_DFFE_PP_  (.D(_00467_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[22][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][25]$_DFFE_PP_  (.D(_00468_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[22][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][26]$_DFFE_PP_  (.D(_00469_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[22][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][27]$_DFFE_PP_  (.D(_00470_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[22][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][28]$_DFFE_PP_  (.D(_00471_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[22][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][29]$_DFFE_PP_  (.D(_00472_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[22][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][2]$_DFFE_PP_  (.D(_00473_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[22][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][30]$_DFFE_PP_  (.D(_00474_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[22][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][31]$_DFFE_PP_  (.D(_00475_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[22][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][3]$_DFFE_PP_  (.D(_00476_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[22][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][4]$_DFFE_PP_  (.D(_00477_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[22][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][5]$_DFFE_PP_  (.D(_00478_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[22][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][6]$_DFFE_PP_  (.D(_00479_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[22][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][7]$_DFFE_PP_  (.D(_00480_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[22][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][8]$_DFFE_PP_  (.D(_00481_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[22][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][9]$_DFFE_PP_  (.D(_00482_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[22][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][0]$_DFFE_PP_  (.D(_00483_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[23][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][10]$_DFFE_PP_  (.D(_00484_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[23][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][11]$_DFFE_PP_  (.D(_00485_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[23][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][12]$_DFFE_PP_  (.D(_00486_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[23][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][13]$_DFFE_PP_  (.D(_00487_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[23][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][14]$_DFFE_PP_  (.D(_00488_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[23][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][15]$_DFFE_PP_  (.D(_00489_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[23][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][16]$_DFFE_PP_  (.D(_00490_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[23][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][17]$_DFFE_PP_  (.D(_00491_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[23][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][18]$_DFFE_PP_  (.D(_00492_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[23][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][19]$_DFFE_PP_  (.D(_00493_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[23][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][1]$_DFFE_PP_  (.D(_00494_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[23][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][20]$_DFFE_PP_  (.D(_00495_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[23][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][21]$_DFFE_PP_  (.D(_00496_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[23][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][22]$_DFFE_PP_  (.D(_00497_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[23][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][23]$_DFFE_PP_  (.D(_00498_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[23][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][24]$_DFFE_PP_  (.D(_00499_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[23][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][25]$_DFFE_PP_  (.D(_00500_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[23][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][26]$_DFFE_PP_  (.D(_00501_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[23][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][27]$_DFFE_PP_  (.D(_00502_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[23][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][28]$_DFFE_PP_  (.D(_00503_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[23][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][29]$_DFFE_PP_  (.D(_00504_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[23][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][2]$_DFFE_PP_  (.D(_00505_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[23][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][30]$_DFFE_PP_  (.D(_00506_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[23][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][31]$_DFFE_PP_  (.D(_00507_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[23][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][3]$_DFFE_PP_  (.D(_00508_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[23][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][4]$_DFFE_PP_  (.D(_00509_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[23][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][5]$_DFFE_PP_  (.D(_00510_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[23][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][6]$_DFFE_PP_  (.D(_00511_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[23][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][7]$_DFFE_PP_  (.D(_00512_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[23][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][8]$_DFFE_PP_  (.D(_00513_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[23][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][9]$_DFFE_PP_  (.D(_00514_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[23][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][0]$_DFFE_PP_  (.D(_00515_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[24][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][10]$_DFFE_PP_  (.D(_00516_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[24][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][11]$_DFFE_PP_  (.D(_00517_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[24][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][12]$_DFFE_PP_  (.D(_00518_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[24][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][13]$_DFFE_PP_  (.D(_00519_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[24][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][14]$_DFFE_PP_  (.D(_00520_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[24][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][15]$_DFFE_PP_  (.D(_00521_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[24][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][16]$_DFFE_PP_  (.D(_00522_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[24][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][17]$_DFFE_PP_  (.D(_00523_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[24][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][18]$_DFFE_PP_  (.D(_00524_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[24][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][19]$_DFFE_PP_  (.D(_00525_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[24][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][1]$_DFFE_PP_  (.D(_00526_),
    .CLK(clknet_leaf_24_clk),
    .Q(\dp.rf.rf[24][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][20]$_DFFE_PP_  (.D(_00527_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[24][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][21]$_DFFE_PP_  (.D(_00528_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[24][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][22]$_DFFE_PP_  (.D(_00529_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[24][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][23]$_DFFE_PP_  (.D(_00530_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[24][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][24]$_DFFE_PP_  (.D(_00531_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[24][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][25]$_DFFE_PP_  (.D(_00532_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[24][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][26]$_DFFE_PP_  (.D(_00533_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[24][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][27]$_DFFE_PP_  (.D(_00534_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[24][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][28]$_DFFE_PP_  (.D(_00535_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[24][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][29]$_DFFE_PP_  (.D(_00536_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[24][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][2]$_DFFE_PP_  (.D(_00537_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[24][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][30]$_DFFE_PP_  (.D(_00538_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[24][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][31]$_DFFE_PP_  (.D(_00539_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[24][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][3]$_DFFE_PP_  (.D(_00540_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[24][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][4]$_DFFE_PP_  (.D(_00541_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[24][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][5]$_DFFE_PP_  (.D(_00542_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[24][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][6]$_DFFE_PP_  (.D(_00543_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[24][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][7]$_DFFE_PP_  (.D(_00544_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[24][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][8]$_DFFE_PP_  (.D(_00545_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[24][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][9]$_DFFE_PP_  (.D(_00546_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[24][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][0]$_DFFE_PP_  (.D(_00547_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[25][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][10]$_DFFE_PP_  (.D(_00548_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[25][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][11]$_DFFE_PP_  (.D(_00549_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[25][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][12]$_DFFE_PP_  (.D(_00550_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[25][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][13]$_DFFE_PP_  (.D(_00551_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[25][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][14]$_DFFE_PP_  (.D(_00552_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[25][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][15]$_DFFE_PP_  (.D(_00553_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[25][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][16]$_DFFE_PP_  (.D(_00554_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[25][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][17]$_DFFE_PP_  (.D(_00555_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[25][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][18]$_DFFE_PP_  (.D(_00556_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[25][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][19]$_DFFE_PP_  (.D(_00557_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[25][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][1]$_DFFE_PP_  (.D(_00558_),
    .CLK(clknet_leaf_23_clk),
    .Q(\dp.rf.rf[25][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][20]$_DFFE_PP_  (.D(_00559_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[25][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][21]$_DFFE_PP_  (.D(_00560_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[25][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][22]$_DFFE_PP_  (.D(_00561_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[25][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][23]$_DFFE_PP_  (.D(_00562_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[25][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][24]$_DFFE_PP_  (.D(_00563_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[25][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][25]$_DFFE_PP_  (.D(_00564_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[25][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][26]$_DFFE_PP_  (.D(_00565_),
    .CLK(clknet_leaf_24_clk),
    .Q(\dp.rf.rf[25][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][27]$_DFFE_PP_  (.D(_00566_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[25][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][28]$_DFFE_PP_  (.D(_00567_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[25][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][29]$_DFFE_PP_  (.D(_00568_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[25][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][2]$_DFFE_PP_  (.D(_00569_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[25][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][30]$_DFFE_PP_  (.D(_00570_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[25][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][31]$_DFFE_PP_  (.D(_00571_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[25][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][3]$_DFFE_PP_  (.D(_00572_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[25][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][4]$_DFFE_PP_  (.D(_00573_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[25][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][5]$_DFFE_PP_  (.D(_00574_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[25][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][6]$_DFFE_PP_  (.D(_00575_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[25][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][7]$_DFFE_PP_  (.D(_00576_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[25][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][8]$_DFFE_PP_  (.D(_00577_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[25][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][9]$_DFFE_PP_  (.D(_00578_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[25][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][0]$_DFFE_PP_  (.D(_00579_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[26][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][10]$_DFFE_PP_  (.D(_00580_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[26][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][11]$_DFFE_PP_  (.D(_00581_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[26][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][12]$_DFFE_PP_  (.D(_00582_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[26][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][13]$_DFFE_PP_  (.D(_00583_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[26][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][14]$_DFFE_PP_  (.D(_00584_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[26][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][15]$_DFFE_PP_  (.D(_00585_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[26][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][16]$_DFFE_PP_  (.D(_00586_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[26][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][17]$_DFFE_PP_  (.D(_00587_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[26][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][18]$_DFFE_PP_  (.D(_00588_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[26][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][19]$_DFFE_PP_  (.D(_00589_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[26][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][1]$_DFFE_PP_  (.D(_00590_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[26][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][20]$_DFFE_PP_  (.D(_00591_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[26][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][21]$_DFFE_PP_  (.D(_00592_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[26][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][22]$_DFFE_PP_  (.D(_00593_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[26][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][23]$_DFFE_PP_  (.D(_00594_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[26][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][24]$_DFFE_PP_  (.D(_00595_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[26][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][25]$_DFFE_PP_  (.D(_00596_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[26][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][26]$_DFFE_PP_  (.D(_00597_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[26][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][27]$_DFFE_PP_  (.D(_00598_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[26][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][28]$_DFFE_PP_  (.D(_00599_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[26][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][29]$_DFFE_PP_  (.D(_00600_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[26][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][2]$_DFFE_PP_  (.D(_00601_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[26][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][30]$_DFFE_PP_  (.D(_00602_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[26][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][31]$_DFFE_PP_  (.D(_00603_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[26][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][3]$_DFFE_PP_  (.D(_00604_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[26][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][4]$_DFFE_PP_  (.D(_00605_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[26][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][5]$_DFFE_PP_  (.D(_00606_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[26][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][6]$_DFFE_PP_  (.D(_00607_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[26][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][7]$_DFFE_PP_  (.D(_00608_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[26][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][8]$_DFFE_PP_  (.D(_00609_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[26][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][9]$_DFFE_PP_  (.D(_00610_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[26][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][0]$_DFFE_PP_  (.D(_00611_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[27][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][10]$_DFFE_PP_  (.D(_00612_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[27][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][11]$_DFFE_PP_  (.D(_00613_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[27][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][12]$_DFFE_PP_  (.D(_00614_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[27][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][13]$_DFFE_PP_  (.D(_00615_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[27][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][14]$_DFFE_PP_  (.D(_00616_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[27][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][15]$_DFFE_PP_  (.D(_00617_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[27][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][16]$_DFFE_PP_  (.D(_00618_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[27][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][17]$_DFFE_PP_  (.D(_00619_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[27][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][18]$_DFFE_PP_  (.D(_00620_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[27][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][19]$_DFFE_PP_  (.D(_00621_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[27][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][1]$_DFFE_PP_  (.D(_00622_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[27][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][20]$_DFFE_PP_  (.D(_00623_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[27][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][21]$_DFFE_PP_  (.D(_00624_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[27][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][22]$_DFFE_PP_  (.D(_00625_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[27][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][23]$_DFFE_PP_  (.D(_00626_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[27][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][24]$_DFFE_PP_  (.D(_00627_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[27][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][25]$_DFFE_PP_  (.D(_00628_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[27][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][26]$_DFFE_PP_  (.D(_00629_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[27][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][27]$_DFFE_PP_  (.D(_00630_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[27][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][28]$_DFFE_PP_  (.D(_00631_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[27][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][29]$_DFFE_PP_  (.D(_00632_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[27][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][2]$_DFFE_PP_  (.D(_00633_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[27][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][30]$_DFFE_PP_  (.D(_00634_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[27][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][31]$_DFFE_PP_  (.D(_00635_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[27][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][3]$_DFFE_PP_  (.D(_00636_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[27][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][4]$_DFFE_PP_  (.D(_00637_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[27][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][5]$_DFFE_PP_  (.D(_00638_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[27][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][6]$_DFFE_PP_  (.D(_00639_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[27][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][7]$_DFFE_PP_  (.D(_00640_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[27][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][8]$_DFFE_PP_  (.D(_00641_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[27][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][9]$_DFFE_PP_  (.D(_00642_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[27][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][0]$_DFFE_PP_  (.D(_00643_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[28][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][10]$_DFFE_PP_  (.D(_00644_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[28][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][11]$_DFFE_PP_  (.D(_00645_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[28][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][12]$_DFFE_PP_  (.D(_00646_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[28][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][13]$_DFFE_PP_  (.D(_00647_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[28][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][14]$_DFFE_PP_  (.D(_00648_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[28][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][15]$_DFFE_PP_  (.D(_00649_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[28][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][16]$_DFFE_PP_  (.D(_00650_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[28][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][17]$_DFFE_PP_  (.D(_00651_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[28][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][18]$_DFFE_PP_  (.D(_00652_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[28][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][19]$_DFFE_PP_  (.D(_00653_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[28][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][1]$_DFFE_PP_  (.D(_00654_),
    .CLK(clknet_leaf_24_clk),
    .Q(\dp.rf.rf[28][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][20]$_DFFE_PP_  (.D(_00655_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[28][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][21]$_DFFE_PP_  (.D(_00656_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[28][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][22]$_DFFE_PP_  (.D(_00657_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[28][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][23]$_DFFE_PP_  (.D(_00658_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[28][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][24]$_DFFE_PP_  (.D(_00659_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[28][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][25]$_DFFE_PP_  (.D(_00660_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[28][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][26]$_DFFE_PP_  (.D(_00661_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[28][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][27]$_DFFE_PP_  (.D(_00662_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[28][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][28]$_DFFE_PP_  (.D(_00663_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[28][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][29]$_DFFE_PP_  (.D(_00664_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[28][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][2]$_DFFE_PP_  (.D(_00665_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[28][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][30]$_DFFE_PP_  (.D(_00666_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[28][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][31]$_DFFE_PP_  (.D(_00667_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[28][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][3]$_DFFE_PP_  (.D(_00668_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[28][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][4]$_DFFE_PP_  (.D(_00669_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[28][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][5]$_DFFE_PP_  (.D(_00670_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[28][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][6]$_DFFE_PP_  (.D(_00671_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[28][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][7]$_DFFE_PP_  (.D(_00672_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[28][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][8]$_DFFE_PP_  (.D(_00673_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[28][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][9]$_DFFE_PP_  (.D(_00674_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[28][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][0]$_DFFE_PP_  (.D(_00675_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[29][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][10]$_DFFE_PP_  (.D(_00676_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[29][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][11]$_DFFE_PP_  (.D(_00677_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[29][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][12]$_DFFE_PP_  (.D(_00678_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[29][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][13]$_DFFE_PP_  (.D(_00679_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[29][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][14]$_DFFE_PP_  (.D(_00680_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[29][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][15]$_DFFE_PP_  (.D(_00681_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[29][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][16]$_DFFE_PP_  (.D(_00682_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[29][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][17]$_DFFE_PP_  (.D(_00683_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[29][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][18]$_DFFE_PP_  (.D(_00684_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[29][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][19]$_DFFE_PP_  (.D(_00685_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[29][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][1]$_DFFE_PP_  (.D(_00686_),
    .CLK(clknet_leaf_24_clk),
    .Q(\dp.rf.rf[29][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][20]$_DFFE_PP_  (.D(_00687_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[29][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][21]$_DFFE_PP_  (.D(_00688_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[29][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][22]$_DFFE_PP_  (.D(_00689_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[29][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][23]$_DFFE_PP_  (.D(_00690_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[29][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][24]$_DFFE_PP_  (.D(_00691_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[29][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][25]$_DFFE_PP_  (.D(_00692_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[29][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][26]$_DFFE_PP_  (.D(_00693_),
    .CLK(clknet_leaf_24_clk),
    .Q(\dp.rf.rf[29][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][27]$_DFFE_PP_  (.D(_00694_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[29][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][28]$_DFFE_PP_  (.D(_00695_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[29][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][29]$_DFFE_PP_  (.D(_00696_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[29][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][2]$_DFFE_PP_  (.D(_00697_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[29][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][30]$_DFFE_PP_  (.D(_00698_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[29][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][31]$_DFFE_PP_  (.D(_00699_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[29][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][3]$_DFFE_PP_  (.D(_00700_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[29][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][4]$_DFFE_PP_  (.D(_00701_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[29][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][5]$_DFFE_PP_  (.D(_00702_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[29][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][6]$_DFFE_PP_  (.D(_00703_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[29][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][7]$_DFFE_PP_  (.D(_00704_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[29][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][8]$_DFFE_PP_  (.D(_00705_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[29][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][9]$_DFFE_PP_  (.D(_00706_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[29][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][0]$_DFFE_PP_  (.D(_00707_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[2][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][10]$_DFFE_PP_  (.D(_00708_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[2][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][11]$_DFFE_PP_  (.D(_00709_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[2][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][12]$_DFFE_PP_  (.D(_00710_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[2][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][13]$_DFFE_PP_  (.D(_00711_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[2][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][14]$_DFFE_PP_  (.D(_00712_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[2][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][15]$_DFFE_PP_  (.D(_00713_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[2][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][16]$_DFFE_PP_  (.D(_00714_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[2][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][17]$_DFFE_PP_  (.D(_00715_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[2][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][18]$_DFFE_PP_  (.D(_00716_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[2][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][19]$_DFFE_PP_  (.D(_00717_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[2][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][1]$_DFFE_PP_  (.D(_00718_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[2][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][20]$_DFFE_PP_  (.D(_00719_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[2][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][21]$_DFFE_PP_  (.D(_00720_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[2][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][22]$_DFFE_PP_  (.D(_00721_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[2][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][23]$_DFFE_PP_  (.D(_00722_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[2][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][24]$_DFFE_PP_  (.D(_00723_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[2][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][25]$_DFFE_PP_  (.D(_00724_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[2][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][26]$_DFFE_PP_  (.D(_00725_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[2][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][27]$_DFFE_PP_  (.D(_00726_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[2][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][28]$_DFFE_PP_  (.D(_00727_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[2][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][29]$_DFFE_PP_  (.D(_00728_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[2][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][2]$_DFFE_PP_  (.D(_00729_),
    .CLK(clknet_leaf_3_clk),
    .Q(\dp.rf.rf[2][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][30]$_DFFE_PP_  (.D(_00730_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[2][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][31]$_DFFE_PP_  (.D(_00731_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[2][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][3]$_DFFE_PP_  (.D(_00732_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[2][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][4]$_DFFE_PP_  (.D(_00733_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[2][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][5]$_DFFE_PP_  (.D(_00734_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[2][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][6]$_DFFE_PP_  (.D(_00735_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[2][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][7]$_DFFE_PP_  (.D(_00736_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[2][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][8]$_DFFE_PP_  (.D(_00737_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[2][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][9]$_DFFE_PP_  (.D(_00738_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[2][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][0]$_DFFE_PP_  (.D(_00739_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[30][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][10]$_DFFE_PP_  (.D(_00740_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[30][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][11]$_DFFE_PP_  (.D(_00741_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[30][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][12]$_DFFE_PP_  (.D(_00742_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[30][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][13]$_DFFE_PP_  (.D(_00743_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[30][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][14]$_DFFE_PP_  (.D(_00744_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[30][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][15]$_DFFE_PP_  (.D(_00745_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[30][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][16]$_DFFE_PP_  (.D(_00746_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[30][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][17]$_DFFE_PP_  (.D(_00747_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[30][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][18]$_DFFE_PP_  (.D(_00748_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[30][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][19]$_DFFE_PP_  (.D(_00749_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[30][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][1]$_DFFE_PP_  (.D(_00750_),
    .CLK(clknet_leaf_24_clk),
    .Q(\dp.rf.rf[30][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][20]$_DFFE_PP_  (.D(_00751_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[30][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][21]$_DFFE_PP_  (.D(_00752_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[30][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][22]$_DFFE_PP_  (.D(_00753_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[30][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][23]$_DFFE_PP_  (.D(_00754_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[30][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][24]$_DFFE_PP_  (.D(_00755_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[30][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][25]$_DFFE_PP_  (.D(_00756_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[30][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][26]$_DFFE_PP_  (.D(_00757_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[30][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][27]$_DFFE_PP_  (.D(_00758_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[30][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][28]$_DFFE_PP_  (.D(_00759_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[30][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][29]$_DFFE_PP_  (.D(_00760_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[30][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][2]$_DFFE_PP_  (.D(_00761_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[30][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][30]$_DFFE_PP_  (.D(_00762_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[30][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][31]$_DFFE_PP_  (.D(_00763_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[30][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][3]$_DFFE_PP_  (.D(_00764_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[30][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][4]$_DFFE_PP_  (.D(_00765_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[30][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][5]$_DFFE_PP_  (.D(_00766_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[30][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][6]$_DFFE_PP_  (.D(_00767_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[30][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][7]$_DFFE_PP_  (.D(_00768_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[30][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][8]$_DFFE_PP_  (.D(_00769_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[30][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][9]$_DFFE_PP_  (.D(_00770_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[30][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][0]$_DFFE_PP_  (.D(_00771_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[31][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][10]$_DFFE_PP_  (.D(_00772_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[31][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][11]$_DFFE_PP_  (.D(_00773_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[31][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][12]$_DFFE_PP_  (.D(_00774_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[31][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][13]$_DFFE_PP_  (.D(_00775_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[31][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][14]$_DFFE_PP_  (.D(_00776_),
    .CLK(clknet_leaf_7_clk),
    .Q(\dp.rf.rf[31][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][15]$_DFFE_PP_  (.D(_00777_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[31][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][16]$_DFFE_PP_  (.D(_00778_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[31][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][17]$_DFFE_PP_  (.D(_00779_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[31][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][18]$_DFFE_PP_  (.D(_00780_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[31][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][19]$_DFFE_PP_  (.D(_00781_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[31][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][1]$_DFFE_PP_  (.D(_00782_),
    .CLK(clknet_leaf_24_clk),
    .Q(\dp.rf.rf[31][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][20]$_DFFE_PP_  (.D(_00783_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[31][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][21]$_DFFE_PP_  (.D(_00784_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[31][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][22]$_DFFE_PP_  (.D(_00785_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[31][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][23]$_DFFE_PP_  (.D(_00786_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[31][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][24]$_DFFE_PP_  (.D(_00787_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[31][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][25]$_DFFE_PP_  (.D(_00788_),
    .CLK(clknet_leaf_21_clk),
    .Q(\dp.rf.rf[31][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][26]$_DFFE_PP_  (.D(_00789_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[31][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][27]$_DFFE_PP_  (.D(_00790_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[31][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][28]$_DFFE_PP_  (.D(_00791_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[31][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][29]$_DFFE_PP_  (.D(_00792_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[31][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][2]$_DFFE_PP_  (.D(_00793_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[31][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][30]$_DFFE_PP_  (.D(_00794_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[31][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][31]$_DFFE_PP_  (.D(_00795_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[31][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][3]$_DFFE_PP_  (.D(_00796_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[31][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][4]$_DFFE_PP_  (.D(_00797_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[31][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][5]$_DFFE_PP_  (.D(_00798_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[31][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][6]$_DFFE_PP_  (.D(_00799_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[31][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][7]$_DFFE_PP_  (.D(_00800_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[31][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][8]$_DFFE_PP_  (.D(_00801_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[31][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][9]$_DFFE_PP_  (.D(_00802_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[31][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][0]$_DFFE_PP_  (.D(_00803_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[3][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][10]$_DFFE_PP_  (.D(_00804_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[3][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][11]$_DFFE_PP_  (.D(_00805_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[3][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][12]$_DFFE_PP_  (.D(_00806_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[3][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][13]$_DFFE_PP_  (.D(_00807_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[3][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][14]$_DFFE_PP_  (.D(_00808_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[3][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][15]$_DFFE_PP_  (.D(_00809_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[3][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][16]$_DFFE_PP_  (.D(_00810_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[3][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][17]$_DFFE_PP_  (.D(_00811_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[3][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][18]$_DFFE_PP_  (.D(_00812_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[3][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][19]$_DFFE_PP_  (.D(_00813_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[3][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][1]$_DFFE_PP_  (.D(_00814_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[3][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][20]$_DFFE_PP_  (.D(_00815_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[3][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][21]$_DFFE_PP_  (.D(_00816_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[3][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][22]$_DFFE_PP_  (.D(_00817_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[3][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][23]$_DFFE_PP_  (.D(_00818_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[3][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][24]$_DFFE_PP_  (.D(_00819_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[3][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][25]$_DFFE_PP_  (.D(_00820_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[3][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][26]$_DFFE_PP_  (.D(_00821_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[3][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][27]$_DFFE_PP_  (.D(_00822_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[3][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][28]$_DFFE_PP_  (.D(_00823_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[3][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][29]$_DFFE_PP_  (.D(_00824_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[3][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][2]$_DFFE_PP_  (.D(_00825_),
    .CLK(clknet_leaf_3_clk),
    .Q(\dp.rf.rf[3][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][30]$_DFFE_PP_  (.D(_00826_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[3][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][31]$_DFFE_PP_  (.D(_00827_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[3][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][3]$_DFFE_PP_  (.D(_00828_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[3][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][4]$_DFFE_PP_  (.D(_00829_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[3][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][5]$_DFFE_PP_  (.D(_00830_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[3][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][6]$_DFFE_PP_  (.D(_00831_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[3][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][7]$_DFFE_PP_  (.D(_00832_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[3][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][8]$_DFFE_PP_  (.D(_00833_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[3][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][9]$_DFFE_PP_  (.D(_00834_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[3][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][0]$_DFFE_PP_  (.D(_00835_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[4][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][10]$_DFFE_PP_  (.D(_00836_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[4][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][11]$_DFFE_PP_  (.D(_00837_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[4][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][12]$_DFFE_PP_  (.D(_00838_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[4][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][13]$_DFFE_PP_  (.D(_00839_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[4][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][14]$_DFFE_PP_  (.D(_00840_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[4][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][15]$_DFFE_PP_  (.D(_00841_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[4][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][16]$_DFFE_PP_  (.D(_00842_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[4][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][17]$_DFFE_PP_  (.D(_00843_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[4][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][18]$_DFFE_PP_  (.D(_00844_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[4][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][19]$_DFFE_PP_  (.D(_00845_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[4][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][1]$_DFFE_PP_  (.D(_00846_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[4][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][20]$_DFFE_PP_  (.D(_00847_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[4][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][21]$_DFFE_PP_  (.D(_00848_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[4][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][22]$_DFFE_PP_  (.D(_00849_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[4][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][23]$_DFFE_PP_  (.D(_00850_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[4][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][24]$_DFFE_PP_  (.D(_00851_),
    .CLK(clknet_leaf_23_clk),
    .Q(\dp.rf.rf[4][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][25]$_DFFE_PP_  (.D(_00852_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[4][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][26]$_DFFE_PP_  (.D(_00853_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[4][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][27]$_DFFE_PP_  (.D(_00854_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[4][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][28]$_DFFE_PP_  (.D(_00855_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[4][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][29]$_DFFE_PP_  (.D(_00856_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[4][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][2]$_DFFE_PP_  (.D(_00857_),
    .CLK(clknet_leaf_3_clk),
    .Q(\dp.rf.rf[4][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][30]$_DFFE_PP_  (.D(_00858_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[4][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][31]$_DFFE_PP_  (.D(_00859_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[4][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][3]$_DFFE_PP_  (.D(_00860_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[4][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][4]$_DFFE_PP_  (.D(_00861_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[4][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][5]$_DFFE_PP_  (.D(_00862_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[4][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][6]$_DFFE_PP_  (.D(_00863_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[4][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][7]$_DFFE_PP_  (.D(_00864_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[4][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][8]$_DFFE_PP_  (.D(_00865_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[4][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][9]$_DFFE_PP_  (.D(_00866_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[4][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][0]$_DFFE_PP_  (.D(_00867_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[5][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][10]$_DFFE_PP_  (.D(_00868_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[5][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][11]$_DFFE_PP_  (.D(_00869_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[5][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][12]$_DFFE_PP_  (.D(_00870_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[5][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][13]$_DFFE_PP_  (.D(_00871_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[5][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][14]$_DFFE_PP_  (.D(_00872_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[5][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][15]$_DFFE_PP_  (.D(_00873_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[5][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][16]$_DFFE_PP_  (.D(_00874_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[5][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][17]$_DFFE_PP_  (.D(_00875_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[5][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][18]$_DFFE_PP_  (.D(_00876_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[5][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][19]$_DFFE_PP_  (.D(_00877_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[5][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][1]$_DFFE_PP_  (.D(_00878_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[5][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][20]$_DFFE_PP_  (.D(_00879_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[5][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][21]$_DFFE_PP_  (.D(_00880_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[5][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][22]$_DFFE_PP_  (.D(_00881_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[5][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][23]$_DFFE_PP_  (.D(_00882_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[5][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][24]$_DFFE_PP_  (.D(_00883_),
    .CLK(clknet_leaf_23_clk),
    .Q(\dp.rf.rf[5][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][25]$_DFFE_PP_  (.D(_00884_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[5][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][26]$_DFFE_PP_  (.D(_00885_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[5][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][27]$_DFFE_PP_  (.D(_00886_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[5][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][28]$_DFFE_PP_  (.D(_00887_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[5][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][29]$_DFFE_PP_  (.D(_00888_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[5][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][2]$_DFFE_PP_  (.D(_00889_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[5][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][30]$_DFFE_PP_  (.D(_00890_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[5][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][31]$_DFFE_PP_  (.D(_00891_),
    .CLK(clknet_leaf_3_clk),
    .Q(\dp.rf.rf[5][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][3]$_DFFE_PP_  (.D(_00892_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[5][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][4]$_DFFE_PP_  (.D(_00893_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[5][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][5]$_DFFE_PP_  (.D(_00894_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[5][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][6]$_DFFE_PP_  (.D(_00895_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[5][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][7]$_DFFE_PP_  (.D(_00896_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[5][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][8]$_DFFE_PP_  (.D(_00897_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[5][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][9]$_DFFE_PP_  (.D(_00898_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[5][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][0]$_DFFE_PP_  (.D(_00899_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[6][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][10]$_DFFE_PP_  (.D(_00900_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[6][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][11]$_DFFE_PP_  (.D(_00901_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[6][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][12]$_DFFE_PP_  (.D(_00902_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[6][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][13]$_DFFE_PP_  (.D(_00903_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[6][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][14]$_DFFE_PP_  (.D(_00904_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[6][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][15]$_DFFE_PP_  (.D(_00905_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[6][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][16]$_DFFE_PP_  (.D(_00906_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[6][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][17]$_DFFE_PP_  (.D(_00907_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[6][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][18]$_DFFE_PP_  (.D(_00908_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[6][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][19]$_DFFE_PP_  (.D(_00909_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[6][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][1]$_DFFE_PP_  (.D(_00910_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[6][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][20]$_DFFE_PP_  (.D(_00911_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[6][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][21]$_DFFE_PP_  (.D(_00912_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[6][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][22]$_DFFE_PP_  (.D(_00913_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[6][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][23]$_DFFE_PP_  (.D(_00914_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[6][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][24]$_DFFE_PP_  (.D(_00915_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[6][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][25]$_DFFE_PP_  (.D(_00916_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[6][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][26]$_DFFE_PP_  (.D(_00917_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[6][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][27]$_DFFE_PP_  (.D(_00918_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[6][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][28]$_DFFE_PP_  (.D(_00919_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[6][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][29]$_DFFE_PP_  (.D(_00920_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[6][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][2]$_DFFE_PP_  (.D(_00921_),
    .CLK(clknet_leaf_3_clk),
    .Q(\dp.rf.rf[6][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][30]$_DFFE_PP_  (.D(_00922_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[6][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][31]$_DFFE_PP_  (.D(_00923_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[6][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][3]$_DFFE_PP_  (.D(_00924_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[6][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][4]$_DFFE_PP_  (.D(_00925_),
    .CLK(clknet_leaf_32_clk),
    .Q(\dp.rf.rf[6][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][5]$_DFFE_PP_  (.D(_00926_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[6][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][6]$_DFFE_PP_  (.D(_00927_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[6][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][7]$_DFFE_PP_  (.D(_00928_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[6][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][8]$_DFFE_PP_  (.D(_00929_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[6][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][9]$_DFFE_PP_  (.D(_00930_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[6][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][0]$_DFFE_PP_  (.D(_00931_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[7][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][10]$_DFFE_PP_  (.D(_00932_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[7][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][11]$_DFFE_PP_  (.D(_00933_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[7][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][12]$_DFFE_PP_  (.D(_00934_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[7][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][13]$_DFFE_PP_  (.D(_00935_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[7][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][14]$_DFFE_PP_  (.D(_00936_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[7][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][15]$_DFFE_PP_  (.D(_00937_),
    .CLK(clknet_leaf_5_clk),
    .Q(\dp.rf.rf[7][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][16]$_DFFE_PP_  (.D(_00938_),
    .CLK(clknet_leaf_8_clk),
    .Q(\dp.rf.rf[7][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][17]$_DFFE_PP_  (.D(_00939_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[7][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][18]$_DFFE_PP_  (.D(_00940_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[7][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][19]$_DFFE_PP_  (.D(_00941_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[7][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][1]$_DFFE_PP_  (.D(_00942_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[7][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][20]$_DFFE_PP_  (.D(_00943_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[7][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][21]$_DFFE_PP_  (.D(_00944_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[7][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][22]$_DFFE_PP_  (.D(_00945_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[7][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][23]$_DFFE_PP_  (.D(_00946_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[7][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][24]$_DFFE_PP_  (.D(_00947_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[7][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][25]$_DFFE_PP_  (.D(_00948_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[7][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][26]$_DFFE_PP_  (.D(_00949_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[7][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][27]$_DFFE_PP_  (.D(_00950_),
    .CLK(clknet_leaf_29_clk),
    .Q(\dp.rf.rf[7][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][28]$_DFFE_PP_  (.D(_00951_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[7][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][29]$_DFFE_PP_  (.D(_00952_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[7][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][2]$_DFFE_PP_  (.D(_00953_),
    .CLK(clknet_leaf_3_clk),
    .Q(\dp.rf.rf[7][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][30]$_DFFE_PP_  (.D(_00954_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[7][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][31]$_DFFE_PP_  (.D(_00955_),
    .CLK(clknet_leaf_3_clk),
    .Q(\dp.rf.rf[7][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][3]$_DFFE_PP_  (.D(_00956_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[7][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][4]$_DFFE_PP_  (.D(_00957_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[7][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][5]$_DFFE_PP_  (.D(_00958_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[7][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][6]$_DFFE_PP_  (.D(_00959_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[7][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][7]$_DFFE_PP_  (.D(_00960_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[7][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][8]$_DFFE_PP_  (.D(_00961_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[7][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][9]$_DFFE_PP_  (.D(_00962_),
    .CLK(clknet_leaf_38_clk),
    .Q(\dp.rf.rf[7][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][0]$_DFFE_PP_  (.D(_00963_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[8][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][10]$_DFFE_PP_  (.D(_00964_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[8][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][11]$_DFFE_PP_  (.D(_00965_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[8][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][12]$_DFFE_PP_  (.D(_00966_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[8][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][13]$_DFFE_PP_  (.D(_00967_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[8][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][14]$_DFFE_PP_  (.D(_00968_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[8][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][15]$_DFFE_PP_  (.D(_00969_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[8][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][16]$_DFFE_PP_  (.D(_00970_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[8][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][17]$_DFFE_PP_  (.D(_00971_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[8][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][18]$_DFFE_PP_  (.D(_00972_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[8][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][19]$_DFFE_PP_  (.D(_00973_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[8][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][1]$_DFFE_PP_  (.D(_00974_),
    .CLK(clknet_leaf_24_clk),
    .Q(\dp.rf.rf[8][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][20]$_DFFE_PP_  (.D(_00975_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[8][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][21]$_DFFE_PP_  (.D(_00976_),
    .CLK(clknet_leaf_16_clk),
    .Q(\dp.rf.rf[8][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][22]$_DFFE_PP_  (.D(_00977_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[8][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][23]$_DFFE_PP_  (.D(_00978_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[8][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][24]$_DFFE_PP_  (.D(_00979_),
    .CLK(clknet_leaf_23_clk),
    .Q(\dp.rf.rf[8][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][25]$_DFFE_PP_  (.D(_00980_),
    .CLK(clknet_leaf_22_clk),
    .Q(\dp.rf.rf[8][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][26]$_DFFE_PP_  (.D(_00981_),
    .CLK(clknet_leaf_24_clk),
    .Q(\dp.rf.rf[8][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][27]$_DFFE_PP_  (.D(_00982_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[8][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][28]$_DFFE_PP_  (.D(_00983_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[8][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][29]$_DFFE_PP_  (.D(_00984_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[8][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][2]$_DFFE_PP_  (.D(_00985_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[8][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][30]$_DFFE_PP_  (.D(_00986_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[8][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][31]$_DFFE_PP_  (.D(_00987_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[8][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][3]$_DFFE_PP_  (.D(_00988_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[8][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][4]$_DFFE_PP_  (.D(_00989_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[8][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][5]$_DFFE_PP_  (.D(_00990_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[8][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][6]$_DFFE_PP_  (.D(_00991_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[8][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][7]$_DFFE_PP_  (.D(_00992_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[8][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][8]$_DFFE_PP_  (.D(_00993_),
    .CLK(clknet_leaf_3_clk),
    .Q(\dp.rf.rf[8][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][9]$_DFFE_PP_  (.D(_00994_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[8][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][0]$_DFFE_PP_  (.D(_00995_),
    .CLK(clknet_leaf_1_clk),
    .Q(\dp.rf.rf[9][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][10]$_DFFE_PP_  (.D(_00996_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[9][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][11]$_DFFE_PP_  (.D(_00997_),
    .CLK(clknet_leaf_9_clk),
    .Q(\dp.rf.rf[9][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][12]$_DFFE_PP_  (.D(_00998_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[9][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][13]$_DFFE_PP_  (.D(_00999_),
    .CLK(clknet_leaf_10_clk),
    .Q(\dp.rf.rf[9][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][14]$_DFFE_PP_  (.D(_01000_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[9][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][15]$_DFFE_PP_  (.D(_01001_),
    .CLK(clknet_leaf_15_clk),
    .Q(\dp.rf.rf[9][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][16]$_DFFE_PP_  (.D(_01002_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[9][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][17]$_DFFE_PP_  (.D(_01003_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[9][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][18]$_DFFE_PP_  (.D(_01004_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[9][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][19]$_DFFE_PP_  (.D(_01005_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[9][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][1]$_DFFE_PP_  (.D(_01006_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[9][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][20]$_DFFE_PP_  (.D(_01007_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[9][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][21]$_DFFE_PP_  (.D(_01008_),
    .CLK(clknet_leaf_17_clk),
    .Q(\dp.rf.rf[9][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][22]$_DFFE_PP_  (.D(_01009_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[9][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][23]$_DFFE_PP_  (.D(_01010_),
    .CLK(clknet_leaf_19_clk),
    .Q(\dp.rf.rf[9][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][24]$_DFFE_PP_  (.D(_01011_),
    .CLK(clknet_leaf_23_clk),
    .Q(\dp.rf.rf[9][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][25]$_DFFE_PP_  (.D(_01012_),
    .CLK(clknet_leaf_22_clk),
    .Q(\dp.rf.rf[9][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][26]$_DFFE_PP_  (.D(_01013_),
    .CLK(clknet_leaf_31_clk),
    .Q(\dp.rf.rf[9][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][27]$_DFFE_PP_  (.D(_01014_),
    .CLK(clknet_leaf_30_clk),
    .Q(\dp.rf.rf[9][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][28]$_DFFE_PP_  (.D(_01015_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[9][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][29]$_DFFE_PP_  (.D(_01016_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[9][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][2]$_DFFE_PP_  (.D(_01017_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[9][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][30]$_DFFE_PP_  (.D(_01018_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[9][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][31]$_DFFE_PP_  (.D(_01019_),
    .CLK(clknet_leaf_4_clk),
    .Q(\dp.rf.rf[9][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][3]$_DFFE_PP_  (.D(_01020_),
    .CLK(clknet_leaf_35_clk),
    .Q(\dp.rf.rf[9][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][4]$_DFFE_PP_  (.D(_01021_),
    .CLK(clknet_leaf_34_clk),
    .Q(\dp.rf.rf[9][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][5]$_DFFE_PP_  (.D(_01022_),
    .CLK(clknet_leaf_36_clk),
    .Q(\dp.rf.rf[9][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][6]$_DFFE_PP_  (.D(_01023_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[9][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][7]$_DFFE_PP_  (.D(_01024_),
    .CLK(clknet_leaf_37_clk),
    .Q(\dp.rf.rf[9][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][8]$_DFFE_PP_  (.D(_01025_),
    .CLK(clknet_leaf_3_clk),
    .Q(\dp.rf.rf[9][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][9]$_DFFE_PP_  (.D(_01026_),
    .CLK(clknet_leaf_33_clk),
    .Q(\dp.rf.rf[9][9] ));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Right_145 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Right_146 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Right_147 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Right_148 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Right_149 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Right_150 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Right_151 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Right_152 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Right_153 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Right_154 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Right_155 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Right_156 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Right_157 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Right_158 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_159_Right_159 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_160_Right_160 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_161_Right_161 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_162_Right_162 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_163 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_164 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_165 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_166 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_167 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_168 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_169 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_170 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_171 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_172 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_173 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_174 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_175 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_176 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_177 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_178 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_179 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_180 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_181 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_182 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_183 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_184 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_185 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_186 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_187 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_188 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_189 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_190 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_191 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_192 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_193 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_194 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_195 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_196 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_197 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_198 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_199 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_200 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_201 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_202 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_203 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_204 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_205 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Left_206 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Left_207 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Left_208 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Left_209 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Left_210 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Left_211 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Left_212 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Left_213 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Left_214 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Left_215 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Left_216 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Left_217 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Left_218 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Left_219 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Left_220 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Left_221 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Left_222 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Left_223 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Left_224 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Left_225 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Left_226 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Left_227 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Left_228 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Left_229 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Left_230 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Left_231 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Left_232 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Left_233 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Left_234 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Left_235 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Left_236 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Left_237 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Left_238 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Left_239 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Left_240 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Left_241 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Left_242 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Left_243 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Left_244 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Left_245 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Left_246 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Left_247 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Left_248 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Left_249 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Left_250 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Left_251 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Left_252 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Left_253 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Left_254 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Left_255 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Left_256 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Left_257 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Left_258 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Left_259 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Left_260 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Left_261 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Left_262 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Left_263 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Left_264 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Left_265 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Left_266 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Left_267 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Left_268 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Left_269 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Left_270 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Left_271 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Left_272 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Left_273 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Left_274 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Left_275 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Left_276 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Left_277 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Left_278 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Left_279 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Left_280 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Left_281 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Left_282 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Left_283 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Left_284 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Left_285 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Left_286 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Left_287 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Left_288 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Left_289 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Left_290 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Left_291 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Left_292 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Left_293 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Left_294 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Left_295 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Left_296 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Left_297 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Left_298 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Left_299 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Left_300 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Left_301 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Left_302 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Left_303 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Left_304 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Left_305 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Left_306 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Left_307 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Left_308 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Left_309 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Left_310 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Left_311 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Left_312 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Left_313 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Left_314 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Left_315 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Left_316 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Left_317 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Left_318 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Left_319 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Left_320 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Left_321 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_159_Left_322 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_160_Left_323 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_161_Left_324 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_162_Left_325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_359 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_360 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_361 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_362 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_363 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_364 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_365 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_366 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_367 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_368 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_369 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_370 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_375 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_376 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_377 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_378 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_379 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_380 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_381 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_382 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_383 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_384 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_385 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_386 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_387 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_388 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_467 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_468 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_961 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_962 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_963 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_964 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_965 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_966 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_967 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_968 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_969 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_970 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_971 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_972 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_973 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_974 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_975 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_976 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_977 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_978 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_979 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_980 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_981 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_982 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_983 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_984 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_985 ();
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 input1 (.I(instr[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input2 (.I(instr[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input3 (.I(instr[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input4 (.I(instr[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input5 (.I(instr[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input6 (.I(instr[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input7 (.I(instr[16]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input8 (.I(instr[18]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input9 (.I(instr[19]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 input10 (.I(instr[1]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input11 (.I(instr[22]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input12 (.I(instr[23]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input13 (.I(instr[24]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input14 (.I(instr[25]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input15 (.I(instr[26]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input16 (.I(instr[27]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input17 (.I(instr[28]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input18 (.I(instr[29]),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input19 (.I(instr[30]),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input20 (.I(instr[31]),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 input21 (.I(instr[3]),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 input22 (.I(instr[4]),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input23 (.I(instr[5]),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 input24 (.I(instr[6]),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input25 (.I(instr[7]),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input26 (.I(instr[8]),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input27 (.I(instr[9]),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input28 (.I(readdata[0]),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input29 (.I(readdata[10]),
    .Z(net29));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input30 (.I(readdata[11]),
    .Z(net30));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input31 (.I(readdata[12]),
    .Z(net31));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input32 (.I(readdata[13]),
    .Z(net32));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input33 (.I(readdata[14]),
    .Z(net33));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input34 (.I(readdata[15]),
    .Z(net34));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input35 (.I(readdata[16]),
    .Z(net35));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input36 (.I(readdata[17]),
    .Z(net36));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input37 (.I(readdata[18]),
    .Z(net37));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input38 (.I(readdata[19]),
    .Z(net38));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input39 (.I(readdata[1]),
    .Z(net39));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input40 (.I(readdata[20]),
    .Z(net40));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input41 (.I(readdata[21]),
    .Z(net41));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input42 (.I(readdata[22]),
    .Z(net42));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input43 (.I(readdata[23]),
    .Z(net43));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input44 (.I(readdata[24]),
    .Z(net44));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input45 (.I(readdata[25]),
    .Z(net45));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input46 (.I(readdata[26]),
    .Z(net46));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input47 (.I(readdata[27]),
    .Z(net47));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input48 (.I(readdata[28]),
    .Z(net48));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input49 (.I(readdata[29]),
    .Z(net49));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input50 (.I(readdata[2]),
    .Z(net50));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input51 (.I(readdata[30]),
    .Z(net51));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input52 (.I(readdata[31]),
    .Z(net52));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input53 (.I(readdata[3]),
    .Z(net53));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input54 (.I(readdata[4]),
    .Z(net54));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input55 (.I(readdata[5]),
    .Z(net55));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input56 (.I(readdata[6]),
    .Z(net56));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input57 (.I(readdata[7]),
    .Z(net57));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input58 (.I(readdata[8]),
    .Z(net58));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input59 (.I(readdata[9]),
    .Z(net59));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input60 (.I(reset),
    .Z(net60));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output61 (.I(net61),
    .Z(aluout[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output62 (.I(net62),
    .Z(aluout[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output63 (.I(net63),
    .Z(aluout[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output64 (.I(net64),
    .Z(aluout[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output65 (.I(net65),
    .Z(aluout[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output66 (.I(net66),
    .Z(aluout[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output67 (.I(net67),
    .Z(aluout[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output68 (.I(net68),
    .Z(aluout[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output69 (.I(net69),
    .Z(aluout[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output70 (.I(net70),
    .Z(aluout[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output71 (.I(net71),
    .Z(aluout[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output72 (.I(net72),
    .Z(aluout[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output73 (.I(net73),
    .Z(aluout[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output74 (.I(net74),
    .Z(aluout[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output75 (.I(net75),
    .Z(aluout[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output76 (.I(net76),
    .Z(aluout[23]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output77 (.I(net77),
    .Z(aluout[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output78 (.I(net78),
    .Z(aluout[25]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output79 (.I(net79),
    .Z(aluout[26]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output80 (.I(net80),
    .Z(aluout[27]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output81 (.I(net81),
    .Z(aluout[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output82 (.I(net82),
    .Z(aluout[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output83 (.I(net83),
    .Z(aluout[2]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output84 (.I(net84),
    .Z(aluout[30]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output85 (.I(net85),
    .Z(aluout[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output86 (.I(net86),
    .Z(aluout[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output87 (.I(net87),
    .Z(aluout[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output88 (.I(net88),
    .Z(aluout[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output89 (.I(net89),
    .Z(aluout[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output90 (.I(net90),
    .Z(aluout[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output91 (.I(net91),
    .Z(aluout[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output92 (.I(net92),
    .Z(aluout[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output93 (.I(net93),
    .Z(memread));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output94 (.I(net94),
    .Z(memwrite));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output95 (.I(net95),
    .Z(pc[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output96 (.I(net96),
    .Z(pc[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output97 (.I(net97),
    .Z(pc[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output98 (.I(net98),
    .Z(pc[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output99 (.I(net99),
    .Z(pc[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output100 (.I(net100),
    .Z(pc[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output101 (.I(net101),
    .Z(pc[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output102 (.I(net102),
    .Z(pc[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output103 (.I(net103),
    .Z(pc[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output104 (.I(net104),
    .Z(pc[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output105 (.I(net105),
    .Z(pc[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output106 (.I(net106),
    .Z(pc[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output107 (.I(net107),
    .Z(pc[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output108 (.I(net108),
    .Z(pc[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output109 (.I(net109),
    .Z(pc[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output110 (.I(net110),
    .Z(pc[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output111 (.I(net111),
    .Z(pc[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output112 (.I(net112),
    .Z(pc[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output113 (.I(net113),
    .Z(pc[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output114 (.I(net114),
    .Z(pc[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output115 (.I(net115),
    .Z(pc[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output116 (.I(net116),
    .Z(pc[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output117 (.I(net117),
    .Z(pc[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output118 (.I(net118),
    .Z(pc[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output119 (.I(net119),
    .Z(pc[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output120 (.I(net120),
    .Z(pc[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output121 (.I(net121),
    .Z(pc[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output122 (.I(net122),
    .Z(pc[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output123 (.I(net123),
    .Z(pc[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output124 (.I(net124),
    .Z(pc[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output125 (.I(net125),
    .Z(pc[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output126 (.I(net126),
    .Z(pc[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output127 (.I(net127),
    .Z(suspend));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output128 (.I(net128),
    .Z(writedata[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output129 (.I(net129),
    .Z(writedata[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output130 (.I(net130),
    .Z(writedata[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output131 (.I(net131),
    .Z(writedata[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output132 (.I(net132),
    .Z(writedata[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output133 (.I(net133),
    .Z(writedata[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output134 (.I(net134),
    .Z(writedata[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output135 (.I(net135),
    .Z(writedata[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output136 (.I(net136),
    .Z(writedata[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output137 (.I(net137),
    .Z(writedata[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output138 (.I(net138),
    .Z(writedata[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output139 (.I(net139),
    .Z(writedata[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output140 (.I(net140),
    .Z(writedata[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output141 (.I(net141),
    .Z(writedata[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output142 (.I(net142),
    .Z(writedata[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output143 (.I(net143),
    .Z(writedata[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output144 (.I(net144),
    .Z(writedata[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output145 (.I(net145),
    .Z(writedata[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output146 (.I(net146),
    .Z(writedata[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output147 (.I(net147),
    .Z(writedata[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output148 (.I(net148),
    .Z(writedata[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output149 (.I(net149),
    .Z(writedata[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output150 (.I(net150),
    .Z(writedata[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output151 (.I(net151),
    .Z(writedata[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output152 (.I(net152),
    .Z(writedata[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output153 (.I(net153),
    .Z(writedata[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output154 (.I(net154),
    .Z(writedata[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output155 (.I(net155),
    .Z(writedata[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output156 (.I(net156),
    .Z(writedata[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output157 (.I(net157),
    .Z(writedata[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output158 (.I(net158),
    .Z(writedata[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output159 (.I(net159),
    .Z(writedata[9]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_0_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_1_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_2_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_3_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_4_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_5_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_6_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_7_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_8_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_9_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_10_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_11_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_12_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_13_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_14_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_15_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_16_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_16_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_17_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_18_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_19_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_20_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_21_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_22_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_23_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_24_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_25_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_26_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_27_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_28_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_29_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_29_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_30_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_31_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_32_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_33_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_34_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_35_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_35_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_36_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_37_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_38_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_2_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_2_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_2_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_2_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_20 clkload0 (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload1 (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload2 (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload3 (.I(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload4 (.I(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 clkload5 (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload6 (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload7 (.I(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload8 (.I(clknet_leaf_35_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload9 (.I(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload10 (.I(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 clkload11 (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload12 (.I(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload13 (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload14 (.I(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 clkload15 (.I(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload16 (.I(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload17 (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload18 (.I(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload19 (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload20 (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload21 (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload22 (.I(clknet_leaf_16_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 clkload23 (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload24 (.I(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload25 (.I(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload26 (.I(clknet_leaf_29_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload27 (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload28 (.I(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload29 (.I(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkload30 (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkload31 (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 clkload32 (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 rebuffer1 (.I(_01076_),
    .Z(net160));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2 (.I(net160),
    .Z(net161));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer3 (.I(net160),
    .Z(net162));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 split4 (.I(_02814_),
    .Z(net163));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer6 (.I(net164),
    .Z(net165));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer7 (.I(_02747_),
    .Z(net166));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 split10 (.I(_04824_),
    .Z(net169));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer11 (.I(_05016_),
    .Z(net170));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer12 (.I(net170),
    .Z(net171));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer13 (.I(net170),
    .Z(net172));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer14 (.I(net170),
    .Z(net173));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer15 (.I(net173),
    .Z(net174));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer17 (.I(net181),
    .Z(net176));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer18 (.I(_01206_),
    .Z(net177));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 split19 (.I(_02750_),
    .Z(net178));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 split20 (.I(_02816_),
    .Z(net179));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 split21 (.I(_01073_),
    .Z(net180));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer23 (.I(net181),
    .Z(net182));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer24 (.I(net181),
    .Z(net183));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer25 (.I(net181),
    .Z(net184));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer26 (.I(net181),
    .Z(net185));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer27 (.I(_01076_),
    .Z(net186));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer29 (.I(_01588_),
    .Z(net188));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer30 (.I(_01588_),
    .Z(net189));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer31 (.I(net189),
    .Z(net190));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer32 (.I(_01588_),
    .Z(net191));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 split33 (.I(_01608_),
    .Z(net192));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer34 (.I(_02811_),
    .Z(net193));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer35 (.I(_01047_),
    .Z(net194));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer36 (.I(_01047_),
    .Z(net195));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer37 (.I(net195),
    .Z(net196));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer38 (.I(_01056_),
    .Z(net197));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer39 (.I(_01097_),
    .Z(net198));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer40 (.I(net198),
    .Z(net199));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer41 (.I(_01342_),
    .Z(net200));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer42 (.I(net200),
    .Z(net201));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer43 (.I(_01342_),
    .Z(net202));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer44 (.I(net202),
    .Z(net203));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer45 (.I(net202),
    .Z(net204));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 split46 (.I(_01207_),
    .Z(net205));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 split47 (.I(_01078_),
    .Z(net206));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer48 (.I(_01358_),
    .Z(net207));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer49 (.I(net207),
    .Z(net208));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer50 (.I(net207),
    .Z(net209));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer51 (.I(_01358_),
    .Z(net210));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer52 (.I(net210),
    .Z(net211));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer53 (.I(_01048_),
    .Z(net212));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer54 (.I(_01778_),
    .Z(net213));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer55 (.I(net213),
    .Z(net214));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer56 (.I(net213),
    .Z(net215));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer57 (.I(_01075_),
    .Z(net216));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer58 (.I(net269),
    .Z(net217));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer59 (.I(net269),
    .Z(net218));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer60 (.I(_05056_),
    .Z(net219));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer61 (.I(net219),
    .Z(net220));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 split63 (.I(_02750_),
    .Z(net222));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer71 (.I(_01032_),
    .Z(net230));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer72 (.I(net230),
    .Z(net231));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer73 (.I(net230),
    .Z(net232));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer74 (.I(net232),
    .Z(net233));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer78 (.I(_04992_),
    .Z(net237));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer79 (.I(net237),
    .Z(net238));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer92 (.I(_01073_),
    .Z(net251));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer93 (.I(_03350_),
    .Z(net252));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer4 (.I(_01677_),
    .Z(net223));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer9 (.I(net223),
    .Z(net224));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer10 (.I(net224),
    .Z(net225));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 split11 (.I(_01547_),
    .Z(net226));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer16 (.I(_01349_),
    .Z(net227));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer19 (.I(_01349_),
    .Z(net228));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer20 (.I(net228),
    .Z(net229));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer21 (.I(net228),
    .Z(net234));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer28 (.I(net234),
    .Z(net235));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer33 (.I(_02030_),
    .Z(net236));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer46 (.I(net236),
    .Z(net239));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer47 (.I(net239),
    .Z(net240));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 rebuffer62 (.I(net240),
    .Z(net241));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 split64 (.I(_04815_),
    .Z(net242));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer65 (.I(_02228_),
    .Z(net243));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer66 (.I(_02814_),
    .Z(net244));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer67 (.I(_01085_),
    .Z(net245));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer68 (.I(net245),
    .Z(net246));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer69 (.I(net245),
    .Z(net247));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer70 (.I(net247),
    .Z(net248));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 split71 (.I(_01548_),
    .Z(net249));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer75 (.I(_02697_),
    .Z(net250));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer76 (.I(_02697_),
    .Z(net253));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer77 (.I(net253),
    .Z(net254));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer80 (.I(_02139_),
    .Z(net255));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer81 (.I(_01553_),
    .Z(net256));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 split82 (.I(_01324_),
    .Z(net257));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer83 (.I(_05064_),
    .Z(net258));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer84 (.I(net266),
    .Z(net259));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer85 (.I(_05064_),
    .Z(net260));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer86 (.I(_01547_),
    .Z(net261));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer87 (.I(_01049_),
    .Z(net262));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 split88 (.I(_04952_),
    .Z(net263));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer90 (.I(_03649_),
    .Z(net265));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer91 (.I(_05064_),
    .Z(net266));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer94 (.I(_01142_),
    .Z(net267));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer95 (.I(_02971_),
    .Z(net268));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer96 (.I(_01075_),
    .Z(net269));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer97 (.I(_01062_),
    .Z(net270));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 split98 (.I(_02892_),
    .Z(net271));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer99 (.I(_01150_),
    .Z(net272));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer100 (.I(net272),
    .Z(net273));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer101 (.I(net273),
    .Z(net274));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_1 (.I(_01588_));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_2 (.I(net157));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_3 (.I(net153));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_11 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1477 ();
endmodule
