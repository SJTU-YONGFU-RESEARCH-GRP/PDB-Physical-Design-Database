module leading_zero_counter (valid_input,
    data_in,
    zero_count);
 output valid_input;
 input [31:0] data_in;
 output [5:0] zero_count;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;

 sky130_fd_sc_hd__nor4_1 _058_ (.A(net32),
    .B(net31),
    .C(net3),
    .D(net2),
    .Y(_003_));
 sky130_fd_sc_hd__nor4_1 _059_ (.A(net5),
    .B(net4),
    .C(net7),
    .D(net6),
    .Y(_004_));
 sky130_fd_sc_hd__nor4_1 _060_ (.A(net26),
    .B(net23),
    .C(net30),
    .D(net29),
    .Y(_005_));
 sky130_fd_sc_hd__nor2_1 _061_ (.A(net12),
    .B(net1),
    .Y(_006_));
 sky130_fd_sc_hd__nor2_1 _062_ (.A(net28),
    .B(net27),
    .Y(_007_));
 sky130_fd_sc_hd__and3_1 _063_ (.A(_005_),
    .B(_006_),
    .C(_007_),
    .X(_008_));
 sky130_fd_sc_hd__nand3_1 _064_ (.A(_003_),
    .B(_004_),
    .C(_008_),
    .Y(net38));
 sky130_fd_sc_hd__or4_1 _065_ (.A(net9),
    .B(net8),
    .C(net11),
    .D(net10),
    .X(_009_));
 sky130_fd_sc_hd__or4_1 _066_ (.A(net14),
    .B(net13),
    .C(net16),
    .D(net15),
    .X(_010_));
 sky130_fd_sc_hd__nor2_1 _067_ (.A(_009_),
    .B(_010_),
    .Y(_011_));
 sky130_fd_sc_hd__nor4_1 _068_ (.A(net18),
    .B(net17),
    .C(net20),
    .D(net19),
    .Y(_012_));
 sky130_fd_sc_hd__nor2_1 _069_ (.A(net22),
    .B(net21),
    .Y(_013_));
 sky130_fd_sc_hd__nor2_1 _070_ (.A(net25),
    .B(net24),
    .Y(_014_));
 sky130_fd_sc_hd__nand4_1 _071_ (.A(_011_),
    .B(_012_),
    .C(_013_),
    .D(_014_),
    .Y(_015_));
 sky130_fd_sc_hd__nor2_1 _072_ (.A(net38),
    .B(_015_),
    .Y(net39));
 sky130_fd_sc_hd__or2_0 _073_ (.A(net38),
    .B(_015_),
    .X(net33));
 sky130_fd_sc_hd__inv_1 _074_ (.A(net29),
    .Y(_016_));
 sky130_fd_sc_hd__nand2b_1 _075_ (.A_N(net30),
    .B(net31),
    .Y(_017_));
 sky130_fd_sc_hd__a21oi_1 _076_ (.A1(_016_),
    .A2(_017_),
    .B1(net28),
    .Y(_018_));
 sky130_fd_sc_hd__nor3_1 _077_ (.A(net1),
    .B(net23),
    .C(net27),
    .Y(_019_));
 sky130_fd_sc_hd__nor2b_1 _078_ (.A(_018_),
    .B_N(_019_),
    .Y(_020_));
 sky130_fd_sc_hd__inv_1 _079_ (.A(net4),
    .Y(_021_));
 sky130_fd_sc_hd__a21oi_1 _080_ (.A1(net5),
    .A2(_021_),
    .B1(net3),
    .Y(_022_));
 sky130_fd_sc_hd__nor3_1 _081_ (.A(net28),
    .B(net30),
    .C(net32),
    .Y(_023_));
 sky130_fd_sc_hd__o21ai_0 _082_ (.A1(net2),
    .A2(_022_),
    .B1(_023_),
    .Y(_024_));
 sky130_fd_sc_hd__inv_1 _083_ (.A(net19),
    .Y(_025_));
 sky130_fd_sc_hd__nand2b_1 _084_ (.A_N(net22),
    .B(net24),
    .Y(_026_));
 sky130_fd_sc_hd__nor2_1 _085_ (.A(net19),
    .B(net21),
    .Y(_027_));
 sky130_fd_sc_hd__a221oi_1 _086_ (.A1(net20),
    .A2(_025_),
    .B1(_026_),
    .B2(_027_),
    .C1(net18),
    .Y(_028_));
 sky130_fd_sc_hd__or3_1 _087_ (.A(net13),
    .B(net15),
    .C(net17),
    .X(_029_));
 sky130_fd_sc_hd__inv_1 _088_ (.A(net13),
    .Y(_030_));
 sky130_fd_sc_hd__nor2_1 _089_ (.A(net13),
    .B(net15),
    .Y(_031_));
 sky130_fd_sc_hd__or3_1 _090_ (.A(net7),
    .B(net9),
    .C(net11),
    .X(_032_));
 sky130_fd_sc_hd__a221oi_1 _091_ (.A1(net14),
    .A2(_030_),
    .B1(net16),
    .B2(_031_),
    .C1(_032_),
    .Y(_033_));
 sky130_fd_sc_hd__o21ai_1 _092_ (.A1(_028_),
    .A2(_029_),
    .B1(_033_),
    .Y(_034_));
 sky130_fd_sc_hd__and2b_1 _093_ (.A_N(net9),
    .B(net10),
    .X(_035_));
 sky130_fd_sc_hd__o21bai_1 _094_ (.A1(net8),
    .A2(_035_),
    .B1_N(net7),
    .Y(_036_));
 sky130_fd_sc_hd__nor3_1 _095_ (.A(net2),
    .B(net4),
    .C(net6),
    .Y(_037_));
 sky130_fd_sc_hd__and4b_1 _096_ (.A_N(_018_),
    .B(_019_),
    .C(_036_),
    .D(_037_),
    .X(_038_));
 sky130_fd_sc_hd__inv_1 _097_ (.A(net23),
    .Y(_039_));
 sky130_fd_sc_hd__a21oi_1 _098_ (.A1(net26),
    .A2(_039_),
    .B1(net12),
    .Y(_040_));
 sky130_fd_sc_hd__nor2_1 _099_ (.A(net1),
    .B(_040_),
    .Y(_041_));
 sky130_fd_sc_hd__a221oi_1 _100_ (.A1(_020_),
    .A2(_024_),
    .B1(_034_),
    .B2(_038_),
    .C1(_041_),
    .Y(net34));
 sky130_fd_sc_hd__nor2_1 _101_ (.A(net11),
    .B(net10),
    .Y(_042_));
 sky130_fd_sc_hd__nor2_1 _102_ (.A(net18),
    .B(net17),
    .Y(_043_));
 sky130_fd_sc_hd__nor2_1 _103_ (.A(net14),
    .B(net13),
    .Y(_044_));
 sky130_fd_sc_hd__o311ai_2 _104_ (.A1(net20),
    .A2(net19),
    .A3(_013_),
    .B1(_043_),
    .C1(_044_),
    .Y(_045_));
 sky130_fd_sc_hd__o21ai_0 _105_ (.A1(net16),
    .A2(net15),
    .B1(_044_),
    .Y(_046_));
 sky130_fd_sc_hd__or4_1 _106_ (.A(net5),
    .B(net4),
    .C(net9),
    .D(net8),
    .X(_047_));
 sky130_fd_sc_hd__a31oi_1 _107_ (.A1(_042_),
    .A2(_045_),
    .A3(_046_),
    .B1(_047_),
    .Y(_048_));
 sky130_fd_sc_hd__nor2_1 _108_ (.A(net7),
    .B(net6),
    .Y(_049_));
 sky130_fd_sc_hd__nor2_1 _109_ (.A(net3),
    .B(net2),
    .Y(_050_));
 sky130_fd_sc_hd__o311ai_0 _110_ (.A1(net5),
    .A2(net4),
    .A3(_049_),
    .B1(_005_),
    .C1(_050_),
    .Y(_051_));
 sky130_fd_sc_hd__nor2_1 _111_ (.A(net26),
    .B(net23),
    .Y(_052_));
 sky130_fd_sc_hd__nor2_1 _112_ (.A(net32),
    .B(net31),
    .Y(_053_));
 sky130_fd_sc_hd__o31ai_1 _113_ (.A1(net30),
    .A2(net29),
    .A3(_053_),
    .B1(_007_),
    .Y(_054_));
 sky130_fd_sc_hd__a21boi_0 _114_ (.A1(_052_),
    .A2(_054_),
    .B1_N(_006_),
    .Y(_055_));
 sky130_fd_sc_hd__o21ai_0 _115_ (.A1(_048_),
    .A2(_051_),
    .B1(_055_),
    .Y(net35));
 sky130_fd_sc_hd__nor2_1 _116_ (.A(net30),
    .B(net29),
    .Y(_056_));
 sky130_fd_sc_hd__nand2_1 _117_ (.A(_056_),
    .B(_007_),
    .Y(_057_));
 sky130_fd_sc_hd__o21bai_1 _118_ (.A1(_010_),
    .A2(_012_),
    .B1_N(_009_),
    .Y(_000_));
 sky130_fd_sc_hd__a21boi_0 _119_ (.A1(_004_),
    .A2(_000_),
    .B1_N(_003_),
    .Y(_001_));
 sky130_fd_sc_hd__o211ai_1 _120_ (.A1(_057_),
    .A2(_001_),
    .B1(_052_),
    .C1(_006_),
    .Y(net36));
 sky130_fd_sc_hd__nand2_1 _121_ (.A(_003_),
    .B(_004_),
    .Y(_002_));
 sky130_fd_sc_hd__o21ai_0 _122_ (.A1(_002_),
    .A2(_011_),
    .B1(_008_),
    .Y(net37));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_45 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(data_in[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(data_in[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(data_in[11]),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(data_in[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(data_in[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(data_in[14]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(data_in[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(data_in[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(data_in[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(data_in[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(data_in[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(data_in[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(data_in[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(data_in[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(data_in[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(data_in[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(data_in[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(data_in[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(data_in[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(data_in[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(data_in[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(data_in[29]),
    .X(net22));
 sky130_fd_sc_hd__dlymetal6s2s_1 input23 (.A(data_in[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(data_in[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(data_in[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(data_in[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(data_in[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(data_in[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(data_in[6]),
    .X(net29));
 sky130_fd_sc_hd__dlymetal6s2s_1 input30 (.A(data_in[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(data_in[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(data_in[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 output33 (.A(net33),
    .X(valid_input));
 sky130_fd_sc_hd__clkbuf_1 output34 (.A(net34),
    .X(zero_count[0]));
 sky130_fd_sc_hd__clkbuf_1 output35 (.A(net35),
    .X(zero_count[1]));
 sky130_fd_sc_hd__clkbuf_1 output36 (.A(net36),
    .X(zero_count[2]));
 sky130_fd_sc_hd__clkbuf_1 output37 (.A(net37),
    .X(zero_count[3]));
 sky130_fd_sc_hd__clkbuf_1 output38 (.A(net38),
    .X(zero_count[4]));
 sky130_fd_sc_hd__clkbuf_1 output39 (.A(net39),
    .X(zero_count[5]));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_70 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_92 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_87 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_129 ();
endmodule
