module configurable_sync_fifo (almost_empty,
    almost_full,
    clk,
    empty,
    full,
    rd_en,
    rst_n,
    wr_en,
    data_in,
    data_out,
    fill_level);
 output almost_empty;
 output almost_full;
 input clk;
 output empty;
 output full;
 input rd_en;
 input rst_n;
 input wr_en;
 input [7:0] data_in;
 output [7:0] data_out;
 output [4:0] fill_level;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire \memory[0][0] ;
 wire \memory[0][1] ;
 wire \memory[0][2] ;
 wire \memory[0][3] ;
 wire \memory[0][4] ;
 wire \memory[0][5] ;
 wire \memory[0][6] ;
 wire \memory[0][7] ;
 wire \memory[10][0] ;
 wire \memory[10][1] ;
 wire \memory[10][2] ;
 wire \memory[10][3] ;
 wire \memory[10][4] ;
 wire \memory[10][5] ;
 wire \memory[10][6] ;
 wire \memory[10][7] ;
 wire \memory[11][0] ;
 wire \memory[11][1] ;
 wire \memory[11][2] ;
 wire \memory[11][3] ;
 wire \memory[11][4] ;
 wire \memory[11][5] ;
 wire \memory[11][6] ;
 wire \memory[11][7] ;
 wire \memory[12][0] ;
 wire \memory[12][1] ;
 wire \memory[12][2] ;
 wire \memory[12][3] ;
 wire \memory[12][4] ;
 wire \memory[12][5] ;
 wire \memory[12][6] ;
 wire \memory[12][7] ;
 wire \memory[13][0] ;
 wire \memory[13][1] ;
 wire \memory[13][2] ;
 wire \memory[13][3] ;
 wire \memory[13][4] ;
 wire \memory[13][5] ;
 wire \memory[13][6] ;
 wire \memory[13][7] ;
 wire \memory[14][0] ;
 wire \memory[14][1] ;
 wire \memory[14][2] ;
 wire \memory[14][3] ;
 wire \memory[14][4] ;
 wire \memory[14][5] ;
 wire \memory[14][6] ;
 wire \memory[14][7] ;
 wire \memory[15][0] ;
 wire \memory[15][1] ;
 wire \memory[15][2] ;
 wire \memory[15][3] ;
 wire \memory[15][4] ;
 wire \memory[15][5] ;
 wire \memory[15][6] ;
 wire \memory[15][7] ;
 wire \memory[1][0] ;
 wire \memory[1][1] ;
 wire \memory[1][2] ;
 wire \memory[1][3] ;
 wire \memory[1][4] ;
 wire \memory[1][5] ;
 wire \memory[1][6] ;
 wire \memory[1][7] ;
 wire \memory[2][0] ;
 wire \memory[2][1] ;
 wire \memory[2][2] ;
 wire \memory[2][3] ;
 wire \memory[2][4] ;
 wire \memory[2][5] ;
 wire \memory[2][6] ;
 wire \memory[2][7] ;
 wire \memory[3][0] ;
 wire \memory[3][1] ;
 wire \memory[3][2] ;
 wire \memory[3][3] ;
 wire \memory[3][4] ;
 wire \memory[3][5] ;
 wire \memory[3][6] ;
 wire \memory[3][7] ;
 wire \memory[4][0] ;
 wire \memory[4][1] ;
 wire \memory[4][2] ;
 wire \memory[4][3] ;
 wire \memory[4][4] ;
 wire \memory[4][5] ;
 wire \memory[4][6] ;
 wire \memory[4][7] ;
 wire \memory[5][0] ;
 wire \memory[5][1] ;
 wire \memory[5][2] ;
 wire \memory[5][3] ;
 wire \memory[5][4] ;
 wire \memory[5][5] ;
 wire \memory[5][6] ;
 wire \memory[5][7] ;
 wire \memory[6][0] ;
 wire \memory[6][1] ;
 wire \memory[6][2] ;
 wire \memory[6][3] ;
 wire \memory[6][4] ;
 wire \memory[6][5] ;
 wire \memory[6][6] ;
 wire \memory[6][7] ;
 wire \memory[7][0] ;
 wire \memory[7][1] ;
 wire \memory[7][2] ;
 wire \memory[7][3] ;
 wire \memory[7][4] ;
 wire \memory[7][5] ;
 wire \memory[7][6] ;
 wire \memory[7][7] ;
 wire \memory[8][0] ;
 wire \memory[8][1] ;
 wire \memory[8][2] ;
 wire \memory[8][3] ;
 wire \memory[8][4] ;
 wire \memory[8][5] ;
 wire \memory[8][6] ;
 wire \memory[8][7] ;
 wire \memory[9][0] ;
 wire \memory[9][1] ;
 wire \memory[9][2] ;
 wire \memory[9][3] ;
 wire \memory[9][4] ;
 wire \memory[9][5] ;
 wire \memory[9][6] ;
 wire \memory[9][7] ;
 wire \rd_ptr[0] ;
 wire \rd_ptr[1] ;
 wire \rd_ptr[2] ;
 wire \rd_ptr[3] ;
 wire \wr_ptr[0] ;
 wire \wr_ptr[1] ;
 wire \wr_ptr[2] ;
 wire \wr_ptr[3] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 CLKBUF_X2 _0581_ (.A(net18),
    .Z(_0152_));
 BUF_X4 _0582_ (.A(net16),
    .Z(_0153_));
 NOR4_X4 _0583_ (.A1(net15),
    .A2(net14),
    .A3(net17),
    .A4(_0153_),
    .ZN(_0154_));
 AND2_X1 _0584_ (.A1(_0152_),
    .A2(_0154_),
    .ZN(net19));
 INV_X1 _0585_ (.A(net2),
    .ZN(_0155_));
 AOI21_X4 _0586_ (.A(_0155_),
    .B1(_0152_),
    .B2(_0154_),
    .ZN(_0156_));
 BUF_X4 _0587_ (.A(_0156_),
    .Z(_0557_));
 NOR2_X1 _0588_ (.A1(net15),
    .A2(net14),
    .ZN(_0157_));
 NOR2_X1 _0589_ (.A1(net17),
    .A2(_0153_),
    .ZN(_0158_));
 NAND3_X2 _0590_ (.A1(_0000_),
    .A2(_0157_),
    .A3(_0158_),
    .ZN(_0159_));
 INV_X2 _0591_ (.A(_0159_),
    .ZN(net13));
 NAND2_X1 _0592_ (.A1(net1),
    .A2(_0159_),
    .ZN(_0160_));
 CLKBUF_X3 _0593_ (.A(_0160_),
    .Z(_0558_));
 INV_X2 _0594_ (.A(_0554_),
    .ZN(_0572_));
 BUF_X1 _0595_ (.A(data_in[0]),
    .Z(_0161_));
 BUF_X2 _0596_ (.A(_0161_),
    .Z(_0162_));
 BUF_X4 _0597_ (.A(\wr_ptr[3] ),
    .Z(_0163_));
 BUF_X4 _0598_ (.A(\wr_ptr[2] ),
    .Z(_0164_));
 CLKBUF_X3 _0599_ (.A(_0562_),
    .Z(_0165_));
 BUF_X1 _0600_ (.A(rst_n),
    .Z(_0166_));
 BUF_X4 _0601_ (.A(_0166_),
    .Z(_0167_));
 NAND3_X1 _0602_ (.A1(_0165_),
    .A2(_0167_),
    .A3(_0156_),
    .ZN(_0168_));
 NOR3_X4 _0603_ (.A1(_0163_),
    .A2(_0164_),
    .A3(_0168_),
    .ZN(_0169_));
 MUX2_X1 _0604_ (.A(\memory[0][0] ),
    .B(_0162_),
    .S(_0169_),
    .Z(_0016_));
 CLKBUF_X2 _0605_ (.A(data_in[1]),
    .Z(_0170_));
 BUF_X2 _0606_ (.A(_0170_),
    .Z(_0171_));
 MUX2_X1 _0607_ (.A(\memory[0][1] ),
    .B(_0171_),
    .S(_0169_),
    .Z(_0017_));
 CLKBUF_X2 _0608_ (.A(data_in[2]),
    .Z(_0172_));
 BUF_X2 _0609_ (.A(_0172_),
    .Z(_0173_));
 MUX2_X1 _0610_ (.A(\memory[0][2] ),
    .B(_0173_),
    .S(_0169_),
    .Z(_0018_));
 CLKBUF_X2 _0611_ (.A(data_in[3]),
    .Z(_0174_));
 BUF_X2 _0612_ (.A(_0174_),
    .Z(_0175_));
 MUX2_X1 _0613_ (.A(\memory[0][3] ),
    .B(_0175_),
    .S(_0169_),
    .Z(_0019_));
 CLKBUF_X2 _0614_ (.A(data_in[4]),
    .Z(_0176_));
 BUF_X2 _0615_ (.A(_0176_),
    .Z(_0177_));
 MUX2_X1 _0616_ (.A(\memory[0][4] ),
    .B(_0177_),
    .S(_0169_),
    .Z(_0020_));
 CLKBUF_X2 _0617_ (.A(data_in[5]),
    .Z(_0178_));
 BUF_X2 _0618_ (.A(_0178_),
    .Z(_0179_));
 MUX2_X1 _0619_ (.A(\memory[0][5] ),
    .B(_0179_),
    .S(_0169_),
    .Z(_0021_));
 CLKBUF_X2 _0620_ (.A(data_in[6]),
    .Z(_0180_));
 BUF_X2 _0621_ (.A(_0180_),
    .Z(_0181_));
 MUX2_X1 _0622_ (.A(\memory[0][6] ),
    .B(_0181_),
    .S(_0169_),
    .Z(_0022_));
 CLKBUF_X2 _0623_ (.A(data_in[7]),
    .Z(_0182_));
 BUF_X2 _0624_ (.A(_0182_),
    .Z(_0183_));
 MUX2_X1 _0625_ (.A(\memory[0][7] ),
    .B(_0183_),
    .S(_0169_),
    .Z(_0023_));
 BUF_X8 _0626_ (.A(_0167_),
    .Z(_0184_));
 CLKBUF_X3 _0627_ (.A(_0564_),
    .Z(_0185_));
 INV_X2 _0628_ (.A(_0164_),
    .ZN(_0186_));
 AND3_X1 _0629_ (.A1(_0163_),
    .A2(_0186_),
    .A3(_0156_),
    .ZN(_0187_));
 BUF_X4 _0630_ (.A(_0187_),
    .Z(_0188_));
 NAND3_X4 _0631_ (.A1(_0184_),
    .A2(_0185_),
    .A3(_0188_),
    .ZN(_0189_));
 MUX2_X1 _0632_ (.A(_0162_),
    .B(\memory[10][0] ),
    .S(_0189_),
    .Z(_0024_));
 MUX2_X1 _0633_ (.A(_0171_),
    .B(\memory[10][1] ),
    .S(_0189_),
    .Z(_0025_));
 MUX2_X1 _0634_ (.A(_0173_),
    .B(\memory[10][2] ),
    .S(_0189_),
    .Z(_0026_));
 MUX2_X1 _0635_ (.A(_0175_),
    .B(\memory[10][3] ),
    .S(_0189_),
    .Z(_0027_));
 MUX2_X1 _0636_ (.A(_0177_),
    .B(\memory[10][4] ),
    .S(_0189_),
    .Z(_0028_));
 MUX2_X1 _0637_ (.A(_0179_),
    .B(\memory[10][5] ),
    .S(_0189_),
    .Z(_0029_));
 MUX2_X1 _0638_ (.A(_0181_),
    .B(\memory[10][6] ),
    .S(_0189_),
    .Z(_0030_));
 MUX2_X1 _0639_ (.A(_0183_),
    .B(\memory[10][7] ),
    .S(_0189_),
    .Z(_0031_));
 BUF_X4 _0640_ (.A(_0568_),
    .Z(_0190_));
 NAND3_X4 _0641_ (.A1(_0190_),
    .A2(_0184_),
    .A3(_0188_),
    .ZN(_0191_));
 MUX2_X1 _0642_ (.A(_0162_),
    .B(\memory[11][0] ),
    .S(_0191_),
    .Z(_0032_));
 MUX2_X1 _0643_ (.A(_0171_),
    .B(\memory[11][1] ),
    .S(_0191_),
    .Z(_0033_));
 MUX2_X1 _0644_ (.A(_0173_),
    .B(\memory[11][2] ),
    .S(_0191_),
    .Z(_0034_));
 MUX2_X1 _0645_ (.A(_0175_),
    .B(\memory[11][3] ),
    .S(_0191_),
    .Z(_0035_));
 MUX2_X1 _0646_ (.A(_0177_),
    .B(\memory[11][4] ),
    .S(_0191_),
    .Z(_0036_));
 MUX2_X1 _0647_ (.A(_0179_),
    .B(\memory[11][5] ),
    .S(_0191_),
    .Z(_0037_));
 MUX2_X1 _0648_ (.A(_0181_),
    .B(\memory[11][6] ),
    .S(_0191_),
    .Z(_0038_));
 MUX2_X1 _0649_ (.A(_0183_),
    .B(\memory[11][7] ),
    .S(_0191_),
    .Z(_0039_));
 INV_X2 _0650_ (.A(_0163_),
    .ZN(_0192_));
 NOR2_X4 _0651_ (.A1(_0192_),
    .A2(_0186_),
    .ZN(_0193_));
 NAND4_X4 _0652_ (.A1(_0165_),
    .A2(_0167_),
    .A3(_0557_),
    .A4(_0193_),
    .ZN(_0194_));
 MUX2_X1 _0653_ (.A(_0162_),
    .B(\memory[12][0] ),
    .S(_0194_),
    .Z(_0040_));
 MUX2_X1 _0654_ (.A(_0171_),
    .B(\memory[12][1] ),
    .S(_0194_),
    .Z(_0041_));
 MUX2_X1 _0655_ (.A(_0173_),
    .B(\memory[12][2] ),
    .S(_0194_),
    .Z(_0042_));
 MUX2_X1 _0656_ (.A(_0175_),
    .B(\memory[12][3] ),
    .S(_0194_),
    .Z(_0043_));
 MUX2_X1 _0657_ (.A(_0177_),
    .B(\memory[12][4] ),
    .S(_0194_),
    .Z(_0044_));
 MUX2_X1 _0658_ (.A(_0179_),
    .B(\memory[12][5] ),
    .S(_0194_),
    .Z(_0045_));
 MUX2_X1 _0659_ (.A(_0181_),
    .B(\memory[12][6] ),
    .S(_0194_),
    .Z(_0046_));
 MUX2_X1 _0660_ (.A(_0183_),
    .B(\memory[12][7] ),
    .S(_0194_),
    .Z(_0047_));
 CLKBUF_X3 _0661_ (.A(_0566_),
    .Z(_0195_));
 NAND4_X4 _0662_ (.A1(_0167_),
    .A2(_0195_),
    .A3(_0557_),
    .A4(_0193_),
    .ZN(_0196_));
 MUX2_X1 _0663_ (.A(_0162_),
    .B(\memory[13][0] ),
    .S(_0196_),
    .Z(_0048_));
 MUX2_X1 _0664_ (.A(_0171_),
    .B(\memory[13][1] ),
    .S(_0196_),
    .Z(_0049_));
 MUX2_X1 _0665_ (.A(_0173_),
    .B(\memory[13][2] ),
    .S(_0196_),
    .Z(_0050_));
 MUX2_X1 _0666_ (.A(_0175_),
    .B(\memory[13][3] ),
    .S(_0196_),
    .Z(_0051_));
 MUX2_X1 _0667_ (.A(_0177_),
    .B(\memory[13][4] ),
    .S(_0196_),
    .Z(_0052_));
 MUX2_X1 _0668_ (.A(_0179_),
    .B(\memory[13][5] ),
    .S(_0196_),
    .Z(_0053_));
 MUX2_X1 _0669_ (.A(_0181_),
    .B(\memory[13][6] ),
    .S(_0196_),
    .Z(_0054_));
 MUX2_X1 _0670_ (.A(_0183_),
    .B(\memory[13][7] ),
    .S(_0196_),
    .Z(_0055_));
 NAND4_X4 _0671_ (.A1(_0167_),
    .A2(_0185_),
    .A3(_0557_),
    .A4(_0193_),
    .ZN(_0197_));
 MUX2_X1 _0672_ (.A(_0162_),
    .B(\memory[14][0] ),
    .S(_0197_),
    .Z(_0056_));
 MUX2_X1 _0673_ (.A(_0171_),
    .B(\memory[14][1] ),
    .S(_0197_),
    .Z(_0057_));
 MUX2_X1 _0674_ (.A(_0173_),
    .B(\memory[14][2] ),
    .S(_0197_),
    .Z(_0058_));
 MUX2_X1 _0675_ (.A(_0175_),
    .B(\memory[14][3] ),
    .S(_0197_),
    .Z(_0059_));
 MUX2_X1 _0676_ (.A(_0177_),
    .B(\memory[14][4] ),
    .S(_0197_),
    .Z(_0060_));
 MUX2_X1 _0677_ (.A(_0179_),
    .B(\memory[14][5] ),
    .S(_0197_),
    .Z(_0061_));
 MUX2_X1 _0678_ (.A(_0181_),
    .B(\memory[14][6] ),
    .S(_0197_),
    .Z(_0062_));
 MUX2_X1 _0679_ (.A(_0183_),
    .B(\memory[14][7] ),
    .S(_0197_),
    .Z(_0063_));
 NAND4_X4 _0680_ (.A1(_0190_),
    .A2(_0167_),
    .A3(_0557_),
    .A4(_0193_),
    .ZN(_0198_));
 MUX2_X1 _0681_ (.A(_0162_),
    .B(\memory[15][0] ),
    .S(_0198_),
    .Z(_0064_));
 MUX2_X1 _0682_ (.A(_0171_),
    .B(\memory[15][1] ),
    .S(_0198_),
    .Z(_0065_));
 MUX2_X1 _0683_ (.A(_0173_),
    .B(\memory[15][2] ),
    .S(_0198_),
    .Z(_0066_));
 MUX2_X1 _0684_ (.A(_0175_),
    .B(\memory[15][3] ),
    .S(_0198_),
    .Z(_0067_));
 MUX2_X1 _0685_ (.A(_0177_),
    .B(\memory[15][4] ),
    .S(_0198_),
    .Z(_0068_));
 MUX2_X1 _0686_ (.A(_0179_),
    .B(\memory[15][5] ),
    .S(_0198_),
    .Z(_0069_));
 MUX2_X1 _0687_ (.A(_0181_),
    .B(\memory[15][6] ),
    .S(_0198_),
    .Z(_0070_));
 MUX2_X1 _0688_ (.A(_0183_),
    .B(\memory[15][7] ),
    .S(_0198_),
    .Z(_0071_));
 NAND3_X1 _0689_ (.A1(_0167_),
    .A2(_0195_),
    .A3(_0156_),
    .ZN(_0199_));
 NOR3_X4 _0690_ (.A1(_0163_),
    .A2(_0164_),
    .A3(_0199_),
    .ZN(_0200_));
 MUX2_X1 _0691_ (.A(\memory[1][0] ),
    .B(_0162_),
    .S(_0200_),
    .Z(_0072_));
 MUX2_X1 _0692_ (.A(\memory[1][1] ),
    .B(_0171_),
    .S(_0200_),
    .Z(_0073_));
 MUX2_X1 _0693_ (.A(\memory[1][2] ),
    .B(_0173_),
    .S(_0200_),
    .Z(_0074_));
 MUX2_X1 _0694_ (.A(\memory[1][3] ),
    .B(_0175_),
    .S(_0200_),
    .Z(_0075_));
 MUX2_X1 _0695_ (.A(\memory[1][4] ),
    .B(_0177_),
    .S(_0200_),
    .Z(_0076_));
 MUX2_X1 _0696_ (.A(\memory[1][5] ),
    .B(_0179_),
    .S(_0200_),
    .Z(_0077_));
 MUX2_X1 _0697_ (.A(\memory[1][6] ),
    .B(_0181_),
    .S(_0200_),
    .Z(_0078_));
 MUX2_X1 _0698_ (.A(\memory[1][7] ),
    .B(_0183_),
    .S(_0200_),
    .Z(_0079_));
 NAND3_X1 _0699_ (.A1(_0167_),
    .A2(_0185_),
    .A3(_0156_),
    .ZN(_0201_));
 NOR3_X4 _0700_ (.A1(_0163_),
    .A2(_0164_),
    .A3(_0201_),
    .ZN(_0202_));
 MUX2_X1 _0701_ (.A(\memory[2][0] ),
    .B(_0162_),
    .S(_0202_),
    .Z(_0080_));
 MUX2_X1 _0702_ (.A(\memory[2][1] ),
    .B(_0171_),
    .S(_0202_),
    .Z(_0081_));
 MUX2_X1 _0703_ (.A(\memory[2][2] ),
    .B(_0173_),
    .S(_0202_),
    .Z(_0082_));
 MUX2_X1 _0704_ (.A(\memory[2][3] ),
    .B(_0175_),
    .S(_0202_),
    .Z(_0083_));
 MUX2_X1 _0705_ (.A(\memory[2][4] ),
    .B(_0177_),
    .S(_0202_),
    .Z(_0084_));
 MUX2_X1 _0706_ (.A(\memory[2][5] ),
    .B(_0179_),
    .S(_0202_),
    .Z(_0085_));
 MUX2_X1 _0707_ (.A(\memory[2][6] ),
    .B(_0181_),
    .S(_0202_),
    .Z(_0086_));
 MUX2_X1 _0708_ (.A(\memory[2][7] ),
    .B(_0183_),
    .S(_0202_),
    .Z(_0087_));
 NAND3_X1 _0709_ (.A1(_0190_),
    .A2(_0167_),
    .A3(_0156_),
    .ZN(_0203_));
 NOR3_X4 _0710_ (.A1(_0163_),
    .A2(_0164_),
    .A3(_0203_),
    .ZN(_0204_));
 MUX2_X1 _0711_ (.A(\memory[3][0] ),
    .B(_0162_),
    .S(_0204_),
    .Z(_0088_));
 MUX2_X1 _0712_ (.A(\memory[3][1] ),
    .B(_0171_),
    .S(_0204_),
    .Z(_0089_));
 MUX2_X1 _0713_ (.A(\memory[3][2] ),
    .B(_0173_),
    .S(_0204_),
    .Z(_0090_));
 MUX2_X1 _0714_ (.A(\memory[3][3] ),
    .B(_0175_),
    .S(_0204_),
    .Z(_0091_));
 MUX2_X1 _0715_ (.A(\memory[3][4] ),
    .B(_0177_),
    .S(_0204_),
    .Z(_0092_));
 MUX2_X1 _0716_ (.A(\memory[3][5] ),
    .B(_0179_),
    .S(_0204_),
    .Z(_0093_));
 MUX2_X1 _0717_ (.A(\memory[3][6] ),
    .B(_0181_),
    .S(_0204_),
    .Z(_0094_));
 MUX2_X1 _0718_ (.A(\memory[3][7] ),
    .B(_0183_),
    .S(_0204_),
    .Z(_0095_));
 AND3_X1 _0719_ (.A1(_0192_),
    .A2(_0164_),
    .A3(_0156_),
    .ZN(_0205_));
 BUF_X4 _0720_ (.A(_0205_),
    .Z(_0206_));
 NAND3_X4 _0721_ (.A1(_0165_),
    .A2(_0184_),
    .A3(_0206_),
    .ZN(_0207_));
 MUX2_X1 _0722_ (.A(_0161_),
    .B(\memory[4][0] ),
    .S(_0207_),
    .Z(_0096_));
 MUX2_X1 _0723_ (.A(_0170_),
    .B(\memory[4][1] ),
    .S(_0207_),
    .Z(_0097_));
 MUX2_X1 _0724_ (.A(_0172_),
    .B(\memory[4][2] ),
    .S(_0207_),
    .Z(_0098_));
 MUX2_X1 _0725_ (.A(_0174_),
    .B(\memory[4][3] ),
    .S(_0207_),
    .Z(_0099_));
 MUX2_X1 _0726_ (.A(_0176_),
    .B(\memory[4][4] ),
    .S(_0207_),
    .Z(_0100_));
 MUX2_X1 _0727_ (.A(_0178_),
    .B(\memory[4][5] ),
    .S(_0207_),
    .Z(_0101_));
 MUX2_X1 _0728_ (.A(_0180_),
    .B(\memory[4][6] ),
    .S(_0207_),
    .Z(_0102_));
 MUX2_X1 _0729_ (.A(_0182_),
    .B(\memory[4][7] ),
    .S(_0207_),
    .Z(_0103_));
 NAND3_X4 _0730_ (.A1(_0184_),
    .A2(_0195_),
    .A3(_0206_),
    .ZN(_0208_));
 MUX2_X1 _0731_ (.A(_0161_),
    .B(\memory[5][0] ),
    .S(_0208_),
    .Z(_0104_));
 MUX2_X1 _0732_ (.A(_0170_),
    .B(\memory[5][1] ),
    .S(_0208_),
    .Z(_0105_));
 MUX2_X1 _0733_ (.A(_0172_),
    .B(\memory[5][2] ),
    .S(_0208_),
    .Z(_0106_));
 MUX2_X1 _0734_ (.A(_0174_),
    .B(\memory[5][3] ),
    .S(_0208_),
    .Z(_0107_));
 MUX2_X1 _0735_ (.A(_0176_),
    .B(\memory[5][4] ),
    .S(_0208_),
    .Z(_0108_));
 MUX2_X1 _0736_ (.A(_0178_),
    .B(\memory[5][5] ),
    .S(_0208_),
    .Z(_0109_));
 MUX2_X1 _0737_ (.A(_0180_),
    .B(\memory[5][6] ),
    .S(_0208_),
    .Z(_0110_));
 MUX2_X1 _0738_ (.A(_0182_),
    .B(\memory[5][7] ),
    .S(_0208_),
    .Z(_0111_));
 NAND3_X4 _0739_ (.A1(_0184_),
    .A2(_0185_),
    .A3(_0206_),
    .ZN(_0209_));
 MUX2_X1 _0740_ (.A(_0161_),
    .B(\memory[6][0] ),
    .S(_0209_),
    .Z(_0112_));
 MUX2_X1 _0741_ (.A(_0170_),
    .B(\memory[6][1] ),
    .S(_0209_),
    .Z(_0113_));
 MUX2_X1 _0742_ (.A(_0172_),
    .B(\memory[6][2] ),
    .S(_0209_),
    .Z(_0114_));
 MUX2_X1 _0743_ (.A(_0174_),
    .B(\memory[6][3] ),
    .S(_0209_),
    .Z(_0115_));
 MUX2_X1 _0744_ (.A(_0176_),
    .B(\memory[6][4] ),
    .S(_0209_),
    .Z(_0116_));
 MUX2_X1 _0745_ (.A(_0178_),
    .B(\memory[6][5] ),
    .S(_0209_),
    .Z(_0117_));
 MUX2_X1 _0746_ (.A(_0180_),
    .B(\memory[6][6] ),
    .S(_0209_),
    .Z(_0118_));
 MUX2_X1 _0747_ (.A(_0182_),
    .B(\memory[6][7] ),
    .S(_0209_),
    .Z(_0119_));
 NAND3_X4 _0748_ (.A1(_0190_),
    .A2(_0184_),
    .A3(_0206_),
    .ZN(_0210_));
 MUX2_X1 _0749_ (.A(_0161_),
    .B(\memory[7][0] ),
    .S(_0210_),
    .Z(_0120_));
 MUX2_X1 _0750_ (.A(_0170_),
    .B(\memory[7][1] ),
    .S(_0210_),
    .Z(_0121_));
 MUX2_X1 _0751_ (.A(_0172_),
    .B(\memory[7][2] ),
    .S(_0210_),
    .Z(_0122_));
 MUX2_X1 _0752_ (.A(_0174_),
    .B(\memory[7][3] ),
    .S(_0210_),
    .Z(_0123_));
 MUX2_X1 _0753_ (.A(_0176_),
    .B(\memory[7][4] ),
    .S(_0210_),
    .Z(_0124_));
 MUX2_X1 _0754_ (.A(_0178_),
    .B(\memory[7][5] ),
    .S(_0210_),
    .Z(_0125_));
 MUX2_X1 _0755_ (.A(_0180_),
    .B(\memory[7][6] ),
    .S(_0210_),
    .Z(_0126_));
 MUX2_X1 _0756_ (.A(_0182_),
    .B(\memory[7][7] ),
    .S(_0210_),
    .Z(_0127_));
 NAND3_X4 _0757_ (.A1(_0165_),
    .A2(_0167_),
    .A3(_0188_),
    .ZN(_0211_));
 MUX2_X1 _0758_ (.A(_0161_),
    .B(\memory[8][0] ),
    .S(_0211_),
    .Z(_0128_));
 MUX2_X1 _0759_ (.A(_0170_),
    .B(\memory[8][1] ),
    .S(_0211_),
    .Z(_0129_));
 MUX2_X1 _0760_ (.A(_0172_),
    .B(\memory[8][2] ),
    .S(_0211_),
    .Z(_0130_));
 MUX2_X1 _0761_ (.A(_0174_),
    .B(\memory[8][3] ),
    .S(_0211_),
    .Z(_0131_));
 MUX2_X1 _0762_ (.A(_0176_),
    .B(\memory[8][4] ),
    .S(_0211_),
    .Z(_0132_));
 MUX2_X1 _0763_ (.A(_0178_),
    .B(\memory[8][5] ),
    .S(_0211_),
    .Z(_0133_));
 MUX2_X1 _0764_ (.A(_0180_),
    .B(\memory[8][6] ),
    .S(_0211_),
    .Z(_0134_));
 MUX2_X1 _0765_ (.A(_0182_),
    .B(\memory[8][7] ),
    .S(_0211_),
    .Z(_0135_));
 NAND3_X4 _0766_ (.A1(_0184_),
    .A2(_0195_),
    .A3(_0188_),
    .ZN(_0212_));
 MUX2_X1 _0767_ (.A(_0161_),
    .B(\memory[9][0] ),
    .S(_0212_),
    .Z(_0136_));
 MUX2_X1 _0768_ (.A(_0170_),
    .B(\memory[9][1] ),
    .S(_0212_),
    .Z(_0137_));
 MUX2_X1 _0769_ (.A(_0172_),
    .B(\memory[9][2] ),
    .S(_0212_),
    .Z(_0138_));
 MUX2_X1 _0770_ (.A(_0174_),
    .B(\memory[9][3] ),
    .S(_0212_),
    .Z(_0139_));
 MUX2_X1 _0771_ (.A(_0176_),
    .B(\memory[9][4] ),
    .S(_0212_),
    .Z(_0140_));
 MUX2_X1 _0772_ (.A(_0178_),
    .B(\memory[9][5] ),
    .S(_0212_),
    .Z(_0141_));
 MUX2_X1 _0773_ (.A(_0180_),
    .B(\memory[9][6] ),
    .S(_0212_),
    .Z(_0142_));
 MUX2_X1 _0774_ (.A(_0182_),
    .B(\memory[9][7] ),
    .S(_0212_),
    .Z(_0143_));
 BUF_X2 _0775_ (.A(_0184_),
    .Z(_0213_));
 BUF_X2 _0776_ (.A(_0559_),
    .Z(_0214_));
 MUX2_X1 _0777_ (.A(_0002_),
    .B(net14),
    .S(_0214_),
    .Z(_0215_));
 AND2_X1 _0778_ (.A1(_0213_),
    .A2(_0215_),
    .ZN(_0003_));
 INV_X2 _0779_ (.A(_0166_),
    .ZN(_0216_));
 CLKBUF_X3 _0780_ (.A(_0216_),
    .Z(_0217_));
 NOR2_X1 _0781_ (.A1(_0556_),
    .A2(_0214_),
    .ZN(_0218_));
 AOI21_X1 _0782_ (.A(_0218_),
    .B1(_0214_),
    .B2(net15),
    .ZN(_0219_));
 NOR2_X1 _0783_ (.A1(_0217_),
    .A2(_0219_),
    .ZN(_0004_));
 XOR2_X1 _0784_ (.A(_0576_),
    .B(_0555_),
    .Z(_0220_));
 NOR2_X1 _0785_ (.A1(_0214_),
    .A2(_0220_),
    .ZN(_0221_));
 AOI21_X1 _0786_ (.A(_0221_),
    .B1(_0214_),
    .B2(_0153_),
    .ZN(_0222_));
 NOR2_X1 _0787_ (.A1(_0217_),
    .A2(_0222_),
    .ZN(_0005_));
 AND2_X1 _0788_ (.A1(net14),
    .A2(_0574_),
    .ZN(_0223_));
 AOI221_X2 _0789_ (.A(_0575_),
    .B1(_0223_),
    .B2(_0580_),
    .C1(_0573_),
    .C2(_0576_),
    .ZN(_0224_));
 XOR2_X1 _0790_ (.A(_0578_),
    .B(_0224_),
    .Z(_0225_));
 INV_X1 _0791_ (.A(net17),
    .ZN(_0226_));
 MUX2_X1 _0792_ (.A(_0225_),
    .B(_0226_),
    .S(_0214_),
    .Z(_0227_));
 NOR2_X1 _0793_ (.A1(_0217_),
    .A2(_0227_),
    .ZN(_0006_));
 INV_X1 _0794_ (.A(_0152_),
    .ZN(_0228_));
 NOR2_X1 _0795_ (.A1(_0228_),
    .A2(_0217_),
    .ZN(_0229_));
 NOR2_X1 _0796_ (.A1(_0152_),
    .A2(_0217_),
    .ZN(_0230_));
 NOR2_X1 _0797_ (.A1(_0572_),
    .A2(_0214_),
    .ZN(_0231_));
 NOR2_X1 _0798_ (.A1(_0554_),
    .A2(_0214_),
    .ZN(_0232_));
 INV_X1 _0799_ (.A(_0575_),
    .ZN(_0233_));
 INV_X1 _0800_ (.A(_0580_),
    .ZN(_0234_));
 OAI21_X1 _0801_ (.A(_0233_),
    .B1(_0234_),
    .B2(_0555_),
    .ZN(_0235_));
 AOI21_X1 _0802_ (.A(_0577_),
    .B1(_0578_),
    .B2(_0235_),
    .ZN(_0236_));
 MUX2_X1 _0803_ (.A(_0231_),
    .B(_0232_),
    .S(_0236_),
    .Z(_0237_));
 MUX2_X1 _0804_ (.A(_0229_),
    .B(_0230_),
    .S(_0237_),
    .Z(_0007_));
 BUF_X4 _0805_ (.A(\rd_ptr[3] ),
    .Z(_0238_));
 BUF_X16 _0806_ (.A(_0238_),
    .Z(_0239_));
 BUF_X8 _0807_ (.A(_0239_),
    .Z(_0240_));
 MUX2_X1 _0808_ (.A(\memory[0][0] ),
    .B(\memory[8][0] ),
    .S(_0240_),
    .Z(_0241_));
 MUX2_X1 _0809_ (.A(\memory[4][0] ),
    .B(\memory[12][0] ),
    .S(_0240_),
    .Z(_0242_));
 CLKBUF_X3 _0810_ (.A(\rd_ptr[2] ),
    .Z(_0243_));
 BUF_X4 _0811_ (.A(_0243_),
    .Z(_0244_));
 MUX2_X1 _0812_ (.A(_0241_),
    .B(_0242_),
    .S(_0244_),
    .Z(_0245_));
 MUX2_X1 _0813_ (.A(\memory[2][0] ),
    .B(\memory[10][0] ),
    .S(_0240_),
    .Z(_0246_));
 MUX2_X1 _0814_ (.A(\memory[6][0] ),
    .B(\memory[14][0] ),
    .S(_0240_),
    .Z(_0247_));
 MUX2_X1 _0815_ (.A(_0246_),
    .B(_0247_),
    .S(_0244_),
    .Z(_0248_));
 BUF_X4 _0816_ (.A(\rd_ptr[1] ),
    .Z(_0249_));
 CLKBUF_X3 _0817_ (.A(_0249_),
    .Z(_0250_));
 MUX2_X1 _0818_ (.A(_0245_),
    .B(_0248_),
    .S(_0250_),
    .Z(_0251_));
 INV_X2 _0819_ (.A(net1),
    .ZN(_0252_));
 CLKBUF_X2 _0820_ (.A(\rd_ptr[0] ),
    .Z(_0253_));
 NOR4_X4 _0821_ (.A1(_0252_),
    .A2(_0253_),
    .A3(_0216_),
    .A4(net13),
    .ZN(_0254_));
 INV_X1 _0822_ (.A(_0253_),
    .ZN(_0255_));
 NOR4_X4 _0823_ (.A1(_0252_),
    .A2(_0255_),
    .A3(_0216_),
    .A4(net13),
    .ZN(_0256_));
 MUX2_X1 _0824_ (.A(\memory[1][0] ),
    .B(\memory[9][0] ),
    .S(_0239_),
    .Z(_0257_));
 MUX2_X1 _0825_ (.A(\memory[5][0] ),
    .B(\memory[13][0] ),
    .S(_0239_),
    .Z(_0258_));
 MUX2_X1 _0826_ (.A(_0257_),
    .B(_0258_),
    .S(_0243_),
    .Z(_0259_));
 MUX2_X1 _0827_ (.A(\memory[3][0] ),
    .B(\memory[11][0] ),
    .S(_0239_),
    .Z(_0260_));
 MUX2_X1 _0828_ (.A(\memory[7][0] ),
    .B(\memory[15][0] ),
    .S(_0239_),
    .Z(_0261_));
 MUX2_X1 _0829_ (.A(_0260_),
    .B(_0261_),
    .S(_0243_),
    .Z(_0262_));
 MUX2_X1 _0830_ (.A(_0259_),
    .B(_0262_),
    .S(_0249_),
    .Z(_0263_));
 AOI22_X1 _0831_ (.A1(_0251_),
    .A2(_0254_),
    .B1(_0256_),
    .B2(_0263_),
    .ZN(_0264_));
 NAND3_X1 _0832_ (.A1(_0213_),
    .A2(net5),
    .A3(_0558_),
    .ZN(_0265_));
 NAND2_X1 _0833_ (.A1(_0264_),
    .A2(_0265_),
    .ZN(_0008_));
 BUF_X8 _0834_ (.A(_0239_),
    .Z(_0266_));
 MUX2_X1 _0835_ (.A(\memory[0][1] ),
    .B(\memory[8][1] ),
    .S(_0266_),
    .Z(_0267_));
 MUX2_X1 _0836_ (.A(\memory[4][1] ),
    .B(\memory[12][1] ),
    .S(_0266_),
    .Z(_0268_));
 BUF_X4 _0837_ (.A(_0243_),
    .Z(_0269_));
 MUX2_X1 _0838_ (.A(_0267_),
    .B(_0268_),
    .S(_0269_),
    .Z(_0270_));
 BUF_X8 _0839_ (.A(_0239_),
    .Z(_0271_));
 MUX2_X1 _0840_ (.A(\memory[2][1] ),
    .B(\memory[10][1] ),
    .S(_0271_),
    .Z(_0272_));
 MUX2_X1 _0841_ (.A(\memory[6][1] ),
    .B(\memory[14][1] ),
    .S(_0240_),
    .Z(_0273_));
 MUX2_X1 _0842_ (.A(_0272_),
    .B(_0273_),
    .S(_0244_),
    .Z(_0274_));
 MUX2_X1 _0843_ (.A(_0270_),
    .B(_0274_),
    .S(_0250_),
    .Z(_0275_));
 BUF_X4 _0844_ (.A(_0238_),
    .Z(_0276_));
 MUX2_X1 _0845_ (.A(\memory[1][1] ),
    .B(\memory[9][1] ),
    .S(_0276_),
    .Z(_0277_));
 BUF_X4 _0846_ (.A(_0238_),
    .Z(_0278_));
 MUX2_X1 _0847_ (.A(\memory[5][1] ),
    .B(\memory[13][1] ),
    .S(_0278_),
    .Z(_0279_));
 CLKBUF_X3 _0848_ (.A(_0243_),
    .Z(_0280_));
 MUX2_X1 _0849_ (.A(_0277_),
    .B(_0279_),
    .S(_0280_),
    .Z(_0281_));
 MUX2_X1 _0850_ (.A(\memory[3][1] ),
    .B(\memory[11][1] ),
    .S(_0278_),
    .Z(_0282_));
 BUF_X4 _0851_ (.A(_0238_),
    .Z(_0283_));
 MUX2_X1 _0852_ (.A(\memory[7][1] ),
    .B(\memory[15][1] ),
    .S(_0283_),
    .Z(_0284_));
 MUX2_X1 _0853_ (.A(_0282_),
    .B(_0284_),
    .S(_0269_),
    .Z(_0285_));
 MUX2_X1 _0854_ (.A(_0281_),
    .B(_0285_),
    .S(_0249_),
    .Z(_0286_));
 AOI22_X1 _0855_ (.A1(_0254_),
    .A2(_0275_),
    .B1(_0286_),
    .B2(_0256_),
    .ZN(_0287_));
 NAND3_X1 _0856_ (.A1(_0213_),
    .A2(net6),
    .A3(_0558_),
    .ZN(_0288_));
 NAND2_X1 _0857_ (.A1(_0287_),
    .A2(_0288_),
    .ZN(_0009_));
 MUX2_X1 _0858_ (.A(\memory[0][2] ),
    .B(\memory[8][2] ),
    .S(_0266_),
    .Z(_0289_));
 MUX2_X1 _0859_ (.A(\memory[4][2] ),
    .B(\memory[12][2] ),
    .S(_0266_),
    .Z(_0290_));
 MUX2_X1 _0860_ (.A(_0289_),
    .B(_0290_),
    .S(_0269_),
    .Z(_0291_));
 MUX2_X1 _0861_ (.A(\memory[2][2] ),
    .B(\memory[10][2] ),
    .S(_0271_),
    .Z(_0292_));
 MUX2_X1 _0862_ (.A(\memory[6][2] ),
    .B(\memory[14][2] ),
    .S(_0240_),
    .Z(_0293_));
 MUX2_X1 _0863_ (.A(_0292_),
    .B(_0293_),
    .S(_0244_),
    .Z(_0294_));
 MUX2_X1 _0864_ (.A(_0291_),
    .B(_0294_),
    .S(_0250_),
    .Z(_0295_));
 MUX2_X1 _0865_ (.A(\memory[1][2] ),
    .B(\memory[9][2] ),
    .S(_0276_),
    .Z(_0296_));
 MUX2_X1 _0866_ (.A(\memory[5][2] ),
    .B(\memory[13][2] ),
    .S(_0276_),
    .Z(_0297_));
 MUX2_X1 _0867_ (.A(_0296_),
    .B(_0297_),
    .S(_0280_),
    .Z(_0298_));
 MUX2_X1 _0868_ (.A(\memory[3][2] ),
    .B(\memory[11][2] ),
    .S(_0278_),
    .Z(_0299_));
 MUX2_X1 _0869_ (.A(\memory[7][2] ),
    .B(\memory[15][2] ),
    .S(_0283_),
    .Z(_0300_));
 MUX2_X1 _0870_ (.A(_0299_),
    .B(_0300_),
    .S(_0280_),
    .Z(_0301_));
 MUX2_X1 _0871_ (.A(_0298_),
    .B(_0301_),
    .S(_0249_),
    .Z(_0302_));
 AOI22_X2 _0872_ (.A1(_0254_),
    .A2(_0295_),
    .B1(_0302_),
    .B2(_0256_),
    .ZN(_0303_));
 NAND3_X1 _0873_ (.A1(_0213_),
    .A2(net7),
    .A3(_0558_),
    .ZN(_0304_));
 NAND2_X1 _0874_ (.A1(_0303_),
    .A2(_0304_),
    .ZN(_0010_));
 MUX2_X1 _0875_ (.A(\memory[0][3] ),
    .B(\memory[8][3] ),
    .S(_0283_),
    .Z(_0305_));
 MUX2_X1 _0876_ (.A(\memory[4][3] ),
    .B(\memory[12][3] ),
    .S(_0266_),
    .Z(_0306_));
 MUX2_X1 _0877_ (.A(_0305_),
    .B(_0306_),
    .S(_0269_),
    .Z(_0307_));
 MUX2_X1 _0878_ (.A(\memory[2][3] ),
    .B(\memory[10][3] ),
    .S(_0271_),
    .Z(_0308_));
 MUX2_X1 _0879_ (.A(\memory[6][3] ),
    .B(\memory[14][3] ),
    .S(_0240_),
    .Z(_0309_));
 MUX2_X1 _0880_ (.A(_0308_),
    .B(_0309_),
    .S(_0244_),
    .Z(_0310_));
 MUX2_X1 _0881_ (.A(_0307_),
    .B(_0310_),
    .S(_0250_),
    .Z(_0311_));
 MUX2_X1 _0882_ (.A(\memory[1][3] ),
    .B(\memory[9][3] ),
    .S(_0276_),
    .Z(_0312_));
 MUX2_X1 _0883_ (.A(\memory[5][3] ),
    .B(\memory[13][3] ),
    .S(_0276_),
    .Z(_0313_));
 MUX2_X1 _0884_ (.A(_0312_),
    .B(_0313_),
    .S(_0280_),
    .Z(_0314_));
 MUX2_X1 _0885_ (.A(\memory[3][3] ),
    .B(\memory[11][3] ),
    .S(_0278_),
    .Z(_0315_));
 MUX2_X1 _0886_ (.A(\memory[7][3] ),
    .B(\memory[15][3] ),
    .S(_0283_),
    .Z(_0316_));
 MUX2_X1 _0887_ (.A(_0315_),
    .B(_0316_),
    .S(_0280_),
    .Z(_0317_));
 MUX2_X1 _0888_ (.A(_0314_),
    .B(_0317_),
    .S(_0249_),
    .Z(_0318_));
 AOI22_X2 _0889_ (.A1(_0254_),
    .A2(_0311_),
    .B1(_0318_),
    .B2(_0256_),
    .ZN(_0319_));
 NAND3_X1 _0890_ (.A1(_0213_),
    .A2(net8),
    .A3(_0558_),
    .ZN(_0320_));
 NAND2_X1 _0891_ (.A1(_0319_),
    .A2(_0320_),
    .ZN(_0011_));
 MUX2_X1 _0892_ (.A(\memory[0][4] ),
    .B(\memory[8][4] ),
    .S(_0283_),
    .Z(_0321_));
 MUX2_X1 _0893_ (.A(\memory[4][4] ),
    .B(\memory[12][4] ),
    .S(_0266_),
    .Z(_0322_));
 MUX2_X1 _0894_ (.A(_0321_),
    .B(_0322_),
    .S(_0269_),
    .Z(_0323_));
 MUX2_X1 _0895_ (.A(\memory[2][4] ),
    .B(\memory[10][4] ),
    .S(_0271_),
    .Z(_0324_));
 MUX2_X1 _0896_ (.A(\memory[6][4] ),
    .B(\memory[14][4] ),
    .S(_0271_),
    .Z(_0325_));
 MUX2_X1 _0897_ (.A(_0324_),
    .B(_0325_),
    .S(_0244_),
    .Z(_0326_));
 MUX2_X1 _0898_ (.A(_0323_),
    .B(_0326_),
    .S(_0250_),
    .Z(_0327_));
 MUX2_X1 _0899_ (.A(\memory[1][4] ),
    .B(\memory[9][4] ),
    .S(_0276_),
    .Z(_0328_));
 MUX2_X1 _0900_ (.A(\memory[5][4] ),
    .B(\memory[13][4] ),
    .S(_0276_),
    .Z(_0329_));
 MUX2_X1 _0901_ (.A(_0328_),
    .B(_0329_),
    .S(_0280_),
    .Z(_0330_));
 MUX2_X1 _0902_ (.A(\memory[3][4] ),
    .B(\memory[11][4] ),
    .S(_0278_),
    .Z(_0331_));
 MUX2_X1 _0903_ (.A(\memory[7][4] ),
    .B(\memory[15][4] ),
    .S(_0283_),
    .Z(_0332_));
 MUX2_X1 _0904_ (.A(_0331_),
    .B(_0332_),
    .S(_0280_),
    .Z(_0333_));
 MUX2_X1 _0905_ (.A(_0330_),
    .B(_0333_),
    .S(_0249_),
    .Z(_0334_));
 AOI22_X2 _0906_ (.A1(_0254_),
    .A2(_0327_),
    .B1(_0334_),
    .B2(_0256_),
    .ZN(_0335_));
 NAND3_X1 _0907_ (.A1(_0213_),
    .A2(net9),
    .A3(_0558_),
    .ZN(_0336_));
 NAND2_X1 _0908_ (.A1(_0335_),
    .A2(_0336_),
    .ZN(_0012_));
 MUX2_X1 _0909_ (.A(\memory[0][5] ),
    .B(\memory[8][5] ),
    .S(_0283_),
    .Z(_0337_));
 MUX2_X1 _0910_ (.A(\memory[4][5] ),
    .B(\memory[12][5] ),
    .S(_0266_),
    .Z(_0338_));
 MUX2_X1 _0911_ (.A(_0337_),
    .B(_0338_),
    .S(_0269_),
    .Z(_0339_));
 MUX2_X1 _0912_ (.A(\memory[2][5] ),
    .B(\memory[10][5] ),
    .S(_0271_),
    .Z(_0340_));
 MUX2_X1 _0913_ (.A(\memory[6][5] ),
    .B(\memory[14][5] ),
    .S(_0271_),
    .Z(_0341_));
 MUX2_X1 _0914_ (.A(_0340_),
    .B(_0341_),
    .S(_0244_),
    .Z(_0342_));
 MUX2_X1 _0915_ (.A(_0339_),
    .B(_0342_),
    .S(_0250_),
    .Z(_0343_));
 MUX2_X1 _0916_ (.A(\memory[1][5] ),
    .B(\memory[9][5] ),
    .S(_0239_),
    .Z(_0344_));
 MUX2_X1 _0917_ (.A(\memory[5][5] ),
    .B(\memory[13][5] ),
    .S(_0276_),
    .Z(_0345_));
 MUX2_X1 _0918_ (.A(_0344_),
    .B(_0345_),
    .S(_0243_),
    .Z(_0346_));
 MUX2_X1 _0919_ (.A(\memory[3][5] ),
    .B(\memory[11][5] ),
    .S(_0278_),
    .Z(_0347_));
 MUX2_X1 _0920_ (.A(\memory[7][5] ),
    .B(\memory[15][5] ),
    .S(_0283_),
    .Z(_0348_));
 MUX2_X1 _0921_ (.A(_0347_),
    .B(_0348_),
    .S(_0280_),
    .Z(_0349_));
 MUX2_X1 _0922_ (.A(_0346_),
    .B(_0349_),
    .S(_0249_),
    .Z(_0350_));
 AOI22_X1 _0923_ (.A1(_0254_),
    .A2(_0343_),
    .B1(_0350_),
    .B2(_0256_),
    .ZN(_0351_));
 NAND3_X1 _0924_ (.A1(_0213_),
    .A2(net10),
    .A3(_0558_),
    .ZN(_0352_));
 NAND2_X1 _0925_ (.A1(_0351_),
    .A2(_0352_),
    .ZN(_0013_));
 MUX2_X1 _0926_ (.A(\memory[0][6] ),
    .B(\memory[8][6] ),
    .S(_0283_),
    .Z(_0353_));
 MUX2_X1 _0927_ (.A(\memory[4][6] ),
    .B(\memory[12][6] ),
    .S(_0266_),
    .Z(_0354_));
 MUX2_X1 _0928_ (.A(_0353_),
    .B(_0354_),
    .S(_0269_),
    .Z(_0355_));
 MUX2_X1 _0929_ (.A(\memory[2][6] ),
    .B(\memory[10][6] ),
    .S(_0271_),
    .Z(_0356_));
 MUX2_X1 _0930_ (.A(\memory[6][6] ),
    .B(\memory[14][6] ),
    .S(_0271_),
    .Z(_0357_));
 MUX2_X1 _0931_ (.A(_0356_),
    .B(_0357_),
    .S(_0269_),
    .Z(_0358_));
 MUX2_X1 _0932_ (.A(_0355_),
    .B(_0358_),
    .S(_0250_),
    .Z(_0359_));
 MUX2_X1 _0933_ (.A(\memory[1][6] ),
    .B(\memory[9][6] ),
    .S(_0239_),
    .Z(_0360_));
 MUX2_X1 _0934_ (.A(\memory[5][6] ),
    .B(\memory[13][6] ),
    .S(_0276_),
    .Z(_0361_));
 MUX2_X1 _0935_ (.A(_0360_),
    .B(_0361_),
    .S(_0243_),
    .Z(_0362_));
 MUX2_X1 _0936_ (.A(\memory[3][6] ),
    .B(\memory[11][6] ),
    .S(_0278_),
    .Z(_0363_));
 MUX2_X1 _0937_ (.A(\memory[7][6] ),
    .B(\memory[15][6] ),
    .S(_0278_),
    .Z(_0364_));
 MUX2_X1 _0938_ (.A(_0363_),
    .B(_0364_),
    .S(_0280_),
    .Z(_0365_));
 MUX2_X1 _0939_ (.A(_0362_),
    .B(_0365_),
    .S(_0249_),
    .Z(_0366_));
 AOI22_X2 _0940_ (.A1(_0254_),
    .A2(_0359_),
    .B1(_0366_),
    .B2(_0256_),
    .ZN(_0367_));
 NAND3_X1 _0941_ (.A1(_0184_),
    .A2(net11),
    .A3(_0558_),
    .ZN(_0368_));
 NAND2_X1 _0942_ (.A1(_0367_),
    .A2(_0368_),
    .ZN(_0014_));
 MUX2_X1 _0943_ (.A(\memory[0][7] ),
    .B(\memory[8][7] ),
    .S(_0283_),
    .Z(_0369_));
 MUX2_X1 _0944_ (.A(\memory[4][7] ),
    .B(\memory[12][7] ),
    .S(_0266_),
    .Z(_0370_));
 MUX2_X1 _0945_ (.A(_0369_),
    .B(_0370_),
    .S(_0269_),
    .Z(_0371_));
 MUX2_X1 _0946_ (.A(\memory[2][7] ),
    .B(\memory[10][7] ),
    .S(_0266_),
    .Z(_0372_));
 MUX2_X1 _0947_ (.A(\memory[6][7] ),
    .B(\memory[14][7] ),
    .S(_0271_),
    .Z(_0373_));
 MUX2_X1 _0948_ (.A(_0372_),
    .B(_0373_),
    .S(_0269_),
    .Z(_0374_));
 MUX2_X1 _0949_ (.A(_0371_),
    .B(_0374_),
    .S(_0249_),
    .Z(_0375_));
 MUX2_X1 _0950_ (.A(\memory[1][7] ),
    .B(\memory[9][7] ),
    .S(_0239_),
    .Z(_0376_));
 MUX2_X1 _0951_ (.A(\memory[5][7] ),
    .B(\memory[13][7] ),
    .S(_0276_),
    .Z(_0377_));
 MUX2_X1 _0952_ (.A(_0376_),
    .B(_0377_),
    .S(_0243_),
    .Z(_0378_));
 MUX2_X1 _0953_ (.A(\memory[3][7] ),
    .B(\memory[11][7] ),
    .S(_0278_),
    .Z(_0379_));
 MUX2_X1 _0954_ (.A(\memory[7][7] ),
    .B(\memory[15][7] ),
    .S(_0278_),
    .Z(_0380_));
 MUX2_X1 _0955_ (.A(_0379_),
    .B(_0380_),
    .S(_0280_),
    .Z(_0381_));
 MUX2_X1 _0956_ (.A(_0378_),
    .B(_0381_),
    .S(_0249_),
    .Z(_0382_));
 AOI22_X2 _0957_ (.A1(_0254_),
    .A2(_0375_),
    .B1(_0382_),
    .B2(_0256_),
    .ZN(_0383_));
 NAND3_X1 _0958_ (.A1(_0184_),
    .A2(net12),
    .A3(_0558_),
    .ZN(_0384_));
 NAND2_X1 _0959_ (.A1(_0383_),
    .A2(_0384_),
    .ZN(_0015_));
 NAND3_X1 _0960_ (.A1(_0244_),
    .A2(_0240_),
    .A3(_0570_),
    .ZN(_0385_));
 NAND2_X1 _0961_ (.A1(_0255_),
    .A2(_0385_),
    .ZN(_0386_));
 MUX2_X1 _0962_ (.A(_0386_),
    .B(_0255_),
    .S(_0558_),
    .Z(_0387_));
 NOR2_X1 _0963_ (.A1(_0217_),
    .A2(_0387_),
    .ZN(_0144_));
 MUX2_X1 _0964_ (.A(_0571_),
    .B(_0250_),
    .S(_0160_),
    .Z(_0388_));
 AND2_X1 _0965_ (.A1(_0213_),
    .A2(_0388_),
    .ZN(_0145_));
 NAND3_X1 _0966_ (.A1(net1),
    .A2(_0570_),
    .A3(_0159_),
    .ZN(_0389_));
 XOR2_X1 _0967_ (.A(_0244_),
    .B(_0389_),
    .Z(_0390_));
 NOR2_X1 _0968_ (.A1(_0217_),
    .A2(_0390_),
    .ZN(_0146_));
 NAND3_X1 _0969_ (.A1(net1),
    .A2(_0244_),
    .A3(_0159_),
    .ZN(_0391_));
 AOI21_X1 _0970_ (.A(_0570_),
    .B1(_0250_),
    .B2(_0253_),
    .ZN(_0392_));
 OAI21_X1 _0971_ (.A(_0240_),
    .B1(_0391_),
    .B2(_0392_),
    .ZN(_0393_));
 NAND2_X1 _0972_ (.A1(_0253_),
    .A2(_0250_),
    .ZN(_0394_));
 OR3_X1 _0973_ (.A1(_0240_),
    .A2(_0394_),
    .A3(_0391_),
    .ZN(_0395_));
 AOI21_X1 _0974_ (.A(_0217_),
    .B1(_0393_),
    .B2(_0395_),
    .ZN(_0147_));
 AOI21_X1 _0975_ (.A(\wr_ptr[0] ),
    .B1(_0193_),
    .B2(_0190_),
    .ZN(_0396_));
 MUX2_X1 _0976_ (.A(\wr_ptr[0] ),
    .B(_0396_),
    .S(_0557_),
    .Z(_0397_));
 AND2_X1 _0977_ (.A1(_0213_),
    .A2(_0397_),
    .ZN(_0148_));
 MUX2_X1 _0978_ (.A(\wr_ptr[1] ),
    .B(_0563_),
    .S(_0557_),
    .Z(_0398_));
 AND2_X1 _0979_ (.A1(_0213_),
    .A2(_0398_),
    .ZN(_0149_));
 NAND2_X1 _0980_ (.A1(_0190_),
    .A2(_0557_),
    .ZN(_0399_));
 XNOR2_X1 _0981_ (.A(_0186_),
    .B(_0399_),
    .ZN(_0400_));
 NOR2_X1 _0982_ (.A1(_0217_),
    .A2(_0400_),
    .ZN(_0150_));
 AOI21_X1 _0983_ (.A(_0190_),
    .B1(\wr_ptr[0] ),
    .B2(\wr_ptr[1] ),
    .ZN(_0401_));
 NOR3_X1 _0984_ (.A1(_0192_),
    .A2(_0186_),
    .A3(_0401_),
    .ZN(_0402_));
 NAND4_X1 _0985_ (.A1(_0164_),
    .A2(\wr_ptr[0] ),
    .A3(\wr_ptr[1] ),
    .A4(_0557_),
    .ZN(_0403_));
 AOI221_X1 _0986_ (.A(_0217_),
    .B1(_0557_),
    .B2(_0402_),
    .C1(_0403_),
    .C2(_0192_),
    .ZN(_0151_));
 INV_X1 _0987_ (.A(_0001_),
    .ZN(_0404_));
 NAND2_X1 _0988_ (.A1(_0153_),
    .A2(_0002_),
    .ZN(_0405_));
 OAI21_X1 _0989_ (.A(_0404_),
    .B1(_0405_),
    .B2(net15),
    .ZN(_0406_));
 NAND2_X1 _0990_ (.A1(_0228_),
    .A2(_0406_),
    .ZN(_0407_));
 NAND3_X1 _0991_ (.A1(_0153_),
    .A2(_0000_),
    .A3(_0157_),
    .ZN(_0408_));
 AOI21_X1 _0992_ (.A(net17),
    .B1(_0407_),
    .B2(_0408_),
    .ZN(net3));
 AND3_X1 _0993_ (.A1(_0228_),
    .A2(_0406_),
    .A3(_0408_),
    .ZN(_0409_));
 AOI21_X1 _0994_ (.A(_0409_),
    .B1(_0228_),
    .B2(_0226_),
    .ZN(net4));
 FA_X1 _0995_ (.A(_0002_),
    .B(_0553_),
    .CI(_0554_),
    .CO(_0555_),
    .S(_0556_));
 HA_X1 _0996_ (.A(_0557_),
    .B(_0558_),
    .CO(_0554_),
    .S(_0559_));
 HA_X1 _0997_ (.A(_0560_),
    .B(_0561_),
    .CO(_0562_),
    .S(_0563_));
 HA_X1 _0998_ (.A(_0560_),
    .B(\wr_ptr[1] ),
    .CO(_0564_),
    .S(_0565_));
 HA_X1 _0999_ (.A(\wr_ptr[0] ),
    .B(_0561_),
    .CO(_0566_),
    .S(_0567_));
 HA_X1 _1000_ (.A(\wr_ptr[0] ),
    .B(\wr_ptr[1] ),
    .CO(_0568_),
    .S(_0569_));
 HA_X1 _1001_ (.A(\rd_ptr[0] ),
    .B(\rd_ptr[1] ),
    .CO(_0570_),
    .S(_0571_));
 HA_X1 _1002_ (.A(net15),
    .B(_0572_),
    .CO(_0573_),
    .S(_0574_));
 HA_X1 _1003_ (.A(net16),
    .B(_0572_),
    .CO(_0575_),
    .S(_0576_));
 HA_X1 _1004_ (.A(net17),
    .B(_0572_),
    .CO(_0577_),
    .S(_0578_));
 HA_X1 _1005_ (.A(net16),
    .B(_0572_),
    .CO(_0579_),
    .S(_0580_));
 DFF_X2 \count[0]$_SDFFE_PN0P_  (.D(_0003_),
    .CK(clknet_4_5_0_clk),
    .Q(net14),
    .QN(_0002_));
 DFF_X2 \count[1]$_SDFFE_PN0P_  (.D(_0004_),
    .CK(clknet_4_5_0_clk),
    .Q(net15),
    .QN(_0553_));
 DFF_X2 \count[2]$_SDFFE_PN0P_  (.D(_0005_),
    .CK(clknet_4_5_0_clk),
    .Q(net16),
    .QN(_0001_));
 DFF_X2 \count[3]$_SDFFE_PN0P_  (.D(_0006_),
    .CK(clknet_4_5_0_clk),
    .Q(net17),
    .QN(_0552_));
 DFF_X1 \count[4]$_SDFFE_PN0P_  (.D(_0007_),
    .CK(clknet_4_5_0_clk),
    .Q(net18),
    .QN(_0000_));
 DFF_X1 \data_out[0]$_SDFFE_PN0P_  (.D(_0008_),
    .CK(clknet_4_13_0_clk),
    .Q(net5),
    .QN(_0551_));
 DFF_X1 \data_out[1]$_SDFFE_PN0P_  (.D(_0009_),
    .CK(clknet_4_7_0_clk),
    .Q(net6),
    .QN(_0550_));
 DFF_X1 \data_out[2]$_SDFFE_PN0P_  (.D(_0010_),
    .CK(clknet_4_13_0_clk),
    .Q(net7),
    .QN(_0549_));
 DFF_X1 \data_out[3]$_SDFFE_PN0P_  (.D(_0011_),
    .CK(clknet_4_13_0_clk),
    .Q(net8),
    .QN(_0548_));
 DFF_X1 \data_out[4]$_SDFFE_PN0P_  (.D(_0012_),
    .CK(clknet_4_7_0_clk),
    .Q(net9),
    .QN(_0547_));
 DFF_X1 \data_out[5]$_SDFFE_PN0P_  (.D(_0013_),
    .CK(clknet_4_13_0_clk),
    .Q(net10),
    .QN(_0546_));
 DFF_X1 \data_out[6]$_SDFFE_PN0P_  (.D(_0014_),
    .CK(clknet_4_13_0_clk),
    .Q(net11),
    .QN(_0545_));
 DFF_X1 \data_out[7]$_SDFFE_PN0P_  (.D(_0015_),
    .CK(clknet_4_13_0_clk),
    .Q(net12),
    .QN(_0544_));
 DFF_X1 \memory[0][0]$_DFFE_PP_  (.D(_0016_),
    .CK(clknet_4_15_0_clk),
    .Q(\memory[0][0] ),
    .QN(_0543_));
 DFF_X1 \memory[0][1]$_DFFE_PP_  (.D(_0017_),
    .CK(clknet_4_4_0_clk),
    .Q(\memory[0][1] ),
    .QN(_0542_));
 DFF_X1 \memory[0][2]$_DFFE_PP_  (.D(_0018_),
    .CK(clknet_4_14_0_clk),
    .Q(\memory[0][2] ),
    .QN(_0541_));
 DFF_X1 \memory[0][3]$_DFFE_PP_  (.D(_0019_),
    .CK(clknet_4_9_0_clk),
    .Q(\memory[0][3] ),
    .QN(_0540_));
 DFF_X1 \memory[0][4]$_DFFE_PP_  (.D(_0020_),
    .CK(clknet_4_1_0_clk),
    .Q(\memory[0][4] ),
    .QN(_0539_));
 DFF_X1 \memory[0][5]$_DFFE_PP_  (.D(_0021_),
    .CK(clknet_4_14_0_clk),
    .Q(\memory[0][5] ),
    .QN(_0538_));
 DFF_X1 \memory[0][6]$_DFFE_PP_  (.D(_0022_),
    .CK(clknet_4_3_0_clk),
    .Q(\memory[0][6] ),
    .QN(_0537_));
 DFF_X1 \memory[0][7]$_DFFE_PP_  (.D(_0023_),
    .CK(clknet_4_11_0_clk),
    .Q(\memory[0][7] ),
    .QN(_0536_));
 DFF_X1 \memory[10][0]$_DFFE_PP_  (.D(_0024_),
    .CK(clknet_4_12_0_clk),
    .Q(\memory[10][0] ),
    .QN(_0535_));
 DFF_X1 \memory[10][1]$_DFFE_PP_  (.D(_0025_),
    .CK(clknet_4_7_0_clk),
    .Q(\memory[10][1] ),
    .QN(_0534_));
 DFF_X1 \memory[10][2]$_DFFE_PP_  (.D(_0026_),
    .CK(clknet_4_12_0_clk),
    .Q(\memory[10][2] ),
    .QN(_0533_));
 DFF_X1 \memory[10][3]$_DFFE_PP_  (.D(_0027_),
    .CK(clknet_4_12_0_clk),
    .Q(\memory[10][3] ),
    .QN(_0532_));
 DFF_X1 \memory[10][4]$_DFFE_PP_  (.D(_0028_),
    .CK(clknet_4_4_0_clk),
    .Q(\memory[10][4] ),
    .QN(_0531_));
 DFF_X1 \memory[10][5]$_DFFE_PP_  (.D(_0029_),
    .CK(clknet_4_12_0_clk),
    .Q(\memory[10][5] ),
    .QN(_0530_));
 DFF_X1 \memory[10][6]$_DFFE_PP_  (.D(_0030_),
    .CK(clknet_4_7_0_clk),
    .Q(\memory[10][6] ),
    .QN(_0529_));
 DFF_X1 \memory[10][7]$_DFFE_PP_  (.D(_0031_),
    .CK(clknet_4_9_0_clk),
    .Q(\memory[10][7] ),
    .QN(_0528_));
 DFF_X1 \memory[11][0]$_DFFE_PP_  (.D(_0032_),
    .CK(clknet_4_13_0_clk),
    .Q(\memory[11][0] ),
    .QN(_0527_));
 DFF_X1 \memory[11][1]$_DFFE_PP_  (.D(_0033_),
    .CK(clknet_4_0_0_clk),
    .Q(\memory[11][1] ),
    .QN(_0526_));
 DFF_X1 \memory[11][2]$_DFFE_PP_  (.D(_0034_),
    .CK(clknet_4_8_0_clk),
    .Q(\memory[11][2] ),
    .QN(_0525_));
 DFF_X1 \memory[11][3]$_DFFE_PP_  (.D(_0035_),
    .CK(clknet_4_8_0_clk),
    .Q(\memory[11][3] ),
    .QN(_0524_));
 DFF_X1 \memory[11][4]$_DFFE_PP_  (.D(_0036_),
    .CK(clknet_4_0_0_clk),
    .Q(\memory[11][4] ),
    .QN(_0523_));
 DFF_X1 \memory[11][5]$_DFFE_PP_  (.D(_0037_),
    .CK(clknet_4_9_0_clk),
    .Q(\memory[11][5] ),
    .QN(_0522_));
 DFF_X1 \memory[11][6]$_DFFE_PP_  (.D(_0038_),
    .CK(clknet_4_2_0_clk),
    .Q(\memory[11][6] ),
    .QN(_0521_));
 DFF_X1 \memory[11][7]$_DFFE_PP_  (.D(_0039_),
    .CK(clknet_4_8_0_clk),
    .Q(\memory[11][7] ),
    .QN(_0520_));
 DFF_X1 \memory[12][0]$_DFFE_PP_  (.D(_0040_),
    .CK(clknet_4_15_0_clk),
    .Q(\memory[12][0] ),
    .QN(_0519_));
 DFF_X1 \memory[12][1]$_DFFE_PP_  (.D(_0041_),
    .CK(clknet_4_5_0_clk),
    .Q(\memory[12][1] ),
    .QN(_0518_));
 DFF_X1 \memory[12][2]$_DFFE_PP_  (.D(_0042_),
    .CK(clknet_4_14_0_clk),
    .Q(\memory[12][2] ),
    .QN(_0517_));
 DFF_X1 \memory[12][3]$_DFFE_PP_  (.D(_0043_),
    .CK(clknet_4_9_0_clk),
    .Q(\memory[12][3] ),
    .QN(_0516_));
 DFF_X1 \memory[12][4]$_DFFE_PP_  (.D(_0044_),
    .CK(clknet_4_4_0_clk),
    .Q(\memory[12][4] ),
    .QN(_0515_));
 DFF_X1 \memory[12][5]$_DFFE_PP_  (.D(_0045_),
    .CK(clknet_4_14_0_clk),
    .Q(\memory[12][5] ),
    .QN(_0514_));
 DFF_X1 \memory[12][6]$_DFFE_PP_  (.D(_0046_),
    .CK(clknet_4_6_0_clk),
    .Q(\memory[12][6] ),
    .QN(_0513_));
 DFF_X1 \memory[12][7]$_DFFE_PP_  (.D(_0047_),
    .CK(clknet_4_11_0_clk),
    .Q(\memory[12][7] ),
    .QN(_0512_));
 DFF_X1 \memory[13][0]$_DFFE_PP_  (.D(_0048_),
    .CK(clknet_4_15_0_clk),
    .Q(\memory[13][0] ),
    .QN(_0511_));
 DFF_X1 \memory[13][1]$_DFFE_PP_  (.D(_0049_),
    .CK(clknet_4_1_0_clk),
    .Q(\memory[13][1] ),
    .QN(_0510_));
 DFF_X1 \memory[13][2]$_DFFE_PP_  (.D(_0050_),
    .CK(clknet_4_10_0_clk),
    .Q(\memory[13][2] ),
    .QN(_0509_));
 DFF_X1 \memory[13][3]$_DFFE_PP_  (.D(_0051_),
    .CK(clknet_4_2_0_clk),
    .Q(\memory[13][3] ),
    .QN(_0508_));
 DFF_X1 \memory[13][4]$_DFFE_PP_  (.D(_0052_),
    .CK(clknet_4_0_0_clk),
    .Q(\memory[13][4] ),
    .QN(_0507_));
 DFF_X1 \memory[13][5]$_DFFE_PP_  (.D(_0053_),
    .CK(clknet_4_11_0_clk),
    .Q(\memory[13][5] ),
    .QN(_0506_));
 DFF_X1 \memory[13][6]$_DFFE_PP_  (.D(_0054_),
    .CK(clknet_4_2_0_clk),
    .Q(\memory[13][6] ),
    .QN(_0505_));
 DFF_X1 \memory[13][7]$_DFFE_PP_  (.D(_0055_),
    .CK(clknet_4_10_0_clk),
    .Q(\memory[13][7] ),
    .QN(_0504_));
 DFF_X1 \memory[14][0]$_DFFE_PP_  (.D(_0056_),
    .CK(clknet_4_15_0_clk),
    .Q(\memory[14][0] ),
    .QN(_0503_));
 DFF_X1 \memory[14][1]$_DFFE_PP_  (.D(_0057_),
    .CK(clknet_4_4_0_clk),
    .Q(\memory[14][1] ),
    .QN(_0502_));
 DFF_X1 \memory[14][2]$_DFFE_PP_  (.D(_0058_),
    .CK(clknet_4_14_0_clk),
    .Q(\memory[14][2] ),
    .QN(_0501_));
 DFF_X1 \memory[14][3]$_DFFE_PP_  (.D(_0059_),
    .CK(clknet_4_12_0_clk),
    .Q(\memory[14][3] ),
    .QN(_0500_));
 DFF_X1 \memory[14][4]$_DFFE_PP_  (.D(_0060_),
    .CK(clknet_4_4_0_clk),
    .Q(\memory[14][4] ),
    .QN(_0499_));
 DFF_X1 \memory[14][5]$_DFFE_PP_  (.D(_0061_),
    .CK(clknet_4_15_0_clk),
    .Q(\memory[14][5] ),
    .QN(_0498_));
 DFF_X1 \memory[14][6]$_DFFE_PP_  (.D(_0062_),
    .CK(clknet_4_6_0_clk),
    .Q(\memory[14][6] ),
    .QN(_0497_));
 DFF_X1 \memory[14][7]$_DFFE_PP_  (.D(_0063_),
    .CK(clknet_4_11_0_clk),
    .Q(\memory[14][7] ),
    .QN(_0496_));
 DFF_X1 \memory[15][0]$_DFFE_PP_  (.D(_0064_),
    .CK(clknet_4_15_0_clk),
    .Q(\memory[15][0] ),
    .QN(_0495_));
 DFF_X1 \memory[15][1]$_DFFE_PP_  (.D(_0065_),
    .CK(clknet_4_1_0_clk),
    .Q(\memory[15][1] ),
    .QN(_0494_));
 DFF_X1 \memory[15][2]$_DFFE_PP_  (.D(_0066_),
    .CK(clknet_4_10_0_clk),
    .Q(\memory[15][2] ),
    .QN(_0493_));
 DFF_X1 \memory[15][3]$_DFFE_PP_  (.D(_0067_),
    .CK(clknet_4_3_0_clk),
    .Q(\memory[15][3] ),
    .QN(_0492_));
 DFF_X1 \memory[15][4]$_DFFE_PP_  (.D(_0068_),
    .CK(clknet_4_0_0_clk),
    .Q(\memory[15][4] ),
    .QN(_0491_));
 DFF_X1 \memory[15][5]$_DFFE_PP_  (.D(_0069_),
    .CK(clknet_4_9_0_clk),
    .Q(\memory[15][5] ),
    .QN(_0490_));
 DFF_X1 \memory[15][6]$_DFFE_PP_  (.D(_0070_),
    .CK(clknet_4_2_0_clk),
    .Q(\memory[15][6] ),
    .QN(_0489_));
 DFF_X1 \memory[15][7]$_DFFE_PP_  (.D(_0071_),
    .CK(clknet_4_10_0_clk),
    .Q(\memory[15][7] ),
    .QN(_0488_));
 DFF_X1 \memory[1][0]$_DFFE_PP_  (.D(_0072_),
    .CK(clknet_4_15_0_clk),
    .Q(\memory[1][0] ),
    .QN(_0487_));
 DFF_X1 \memory[1][1]$_DFFE_PP_  (.D(_0073_),
    .CK(clknet_4_0_0_clk),
    .Q(\memory[1][1] ),
    .QN(_0486_));
 DFF_X1 \memory[1][2]$_DFFE_PP_  (.D(_0074_),
    .CK(clknet_4_10_0_clk),
    .Q(\memory[1][2] ),
    .QN(_0485_));
 DFF_X1 \memory[1][3]$_DFFE_PP_  (.D(_0075_),
    .CK(clknet_4_2_0_clk),
    .Q(\memory[1][3] ),
    .QN(_0484_));
 DFF_X1 \memory[1][4]$_DFFE_PP_  (.D(_0076_),
    .CK(clknet_4_0_0_clk),
    .Q(\memory[1][4] ),
    .QN(_0483_));
 DFF_X1 \memory[1][5]$_DFFE_PP_  (.D(_0077_),
    .CK(clknet_4_15_0_clk),
    .Q(\memory[1][5] ),
    .QN(_0482_));
 DFF_X1 \memory[1][6]$_DFFE_PP_  (.D(_0078_),
    .CK(clknet_4_3_0_clk),
    .Q(\memory[1][6] ),
    .QN(_0481_));
 DFF_X1 \memory[1][7]$_DFFE_PP_  (.D(_0079_),
    .CK(clknet_4_10_0_clk),
    .Q(\memory[1][7] ),
    .QN(_0480_));
 DFF_X1 \memory[2][0]$_DFFE_PP_  (.D(_0080_),
    .CK(clknet_4_13_0_clk),
    .Q(\memory[2][0] ),
    .QN(_0479_));
 DFF_X1 \memory[2][1]$_DFFE_PP_  (.D(_0081_),
    .CK(clknet_4_6_0_clk),
    .Q(\memory[2][1] ),
    .QN(_0478_));
 DFF_X1 \memory[2][2]$_DFFE_PP_  (.D(_0082_),
    .CK(clknet_4_12_0_clk),
    .Q(\memory[2][2] ),
    .QN(_0477_));
 DFF_X1 \memory[2][3]$_DFFE_PP_  (.D(_0083_),
    .CK(clknet_4_12_0_clk),
    .Q(\memory[2][3] ),
    .QN(_0476_));
 DFF_X1 \memory[2][4]$_DFFE_PP_  (.D(_0084_),
    .CK(clknet_4_1_0_clk),
    .Q(\memory[2][4] ),
    .QN(_0475_));
 DFF_X1 \memory[2][5]$_DFFE_PP_  (.D(_0085_),
    .CK(clknet_4_14_0_clk),
    .Q(\memory[2][5] ),
    .QN(_0474_));
 DFF_X1 \memory[2][6]$_DFFE_PP_  (.D(_0086_),
    .CK(clknet_4_7_0_clk),
    .Q(\memory[2][6] ),
    .QN(_0473_));
 DFF_X1 \memory[2][7]$_DFFE_PP_  (.D(_0087_),
    .CK(clknet_4_9_0_clk),
    .Q(\memory[2][7] ),
    .QN(_0472_));
 DFF_X1 \memory[3][0]$_DFFE_PP_  (.D(_0088_),
    .CK(clknet_4_13_0_clk),
    .Q(\memory[3][0] ),
    .QN(_0471_));
 DFF_X1 \memory[3][1]$_DFFE_PP_  (.D(_0089_),
    .CK(clknet_4_0_0_clk),
    .Q(\memory[3][1] ),
    .QN(_0470_));
 DFF_X1 \memory[3][2]$_DFFE_PP_  (.D(_0090_),
    .CK(clknet_4_8_0_clk),
    .Q(\memory[3][2] ),
    .QN(_0469_));
 DFF_X1 \memory[3][3]$_DFFE_PP_  (.D(_0091_),
    .CK(clknet_4_8_0_clk),
    .Q(\memory[3][3] ),
    .QN(_0468_));
 DFF_X1 \memory[3][4]$_DFFE_PP_  (.D(_0092_),
    .CK(clknet_4_0_0_clk),
    .Q(\memory[3][4] ),
    .QN(_0467_));
 DFF_X1 \memory[3][5]$_DFFE_PP_  (.D(_0093_),
    .CK(clknet_4_8_0_clk),
    .Q(\memory[3][5] ),
    .QN(_0466_));
 DFF_X1 \memory[3][6]$_DFFE_PP_  (.D(_0094_),
    .CK(clknet_4_2_0_clk),
    .Q(\memory[3][6] ),
    .QN(_0465_));
 DFF_X1 \memory[3][7]$_DFFE_PP_  (.D(_0095_),
    .CK(clknet_4_8_0_clk),
    .Q(\memory[3][7] ),
    .QN(_0464_));
 DFF_X1 \memory[4][0]$_DFFE_PP_  (.D(_0096_),
    .CK(clknet_4_15_0_clk),
    .Q(\memory[4][0] ),
    .QN(_0463_));
 DFF_X1 \memory[4][1]$_DFFE_PP_  (.D(_0097_),
    .CK(clknet_4_4_0_clk),
    .Q(\memory[4][1] ),
    .QN(_0462_));
 DFF_X1 \memory[4][2]$_DFFE_PP_  (.D(_0098_),
    .CK(clknet_4_14_0_clk),
    .Q(\memory[4][2] ),
    .QN(_0461_));
 DFF_X1 \memory[4][3]$_DFFE_PP_  (.D(_0099_),
    .CK(clknet_4_6_0_clk),
    .Q(\memory[4][3] ),
    .QN(_0460_));
 DFF_X1 \memory[4][4]$_DFFE_PP_  (.D(_0100_),
    .CK(clknet_4_4_0_clk),
    .Q(\memory[4][4] ),
    .QN(_0459_));
 DFF_X1 \memory[4][5]$_DFFE_PP_  (.D(_0101_),
    .CK(clknet_4_14_0_clk),
    .Q(\memory[4][5] ),
    .QN(_0458_));
 DFF_X1 \memory[4][6]$_DFFE_PP_  (.D(_0102_),
    .CK(clknet_4_3_0_clk),
    .Q(\memory[4][6] ),
    .QN(_0457_));
 DFF_X1 \memory[4][7]$_DFFE_PP_  (.D(_0103_),
    .CK(clknet_4_11_0_clk),
    .Q(\memory[4][7] ),
    .QN(_0456_));
 DFF_X1 \memory[5][0]$_DFFE_PP_  (.D(_0104_),
    .CK(clknet_4_15_0_clk),
    .Q(\memory[5][0] ),
    .QN(_0455_));
 DFF_X1 \memory[5][1]$_DFFE_PP_  (.D(_0105_),
    .CK(clknet_4_3_0_clk),
    .Q(\memory[5][1] ),
    .QN(_0454_));
 DFF_X1 \memory[5][2]$_DFFE_PP_  (.D(_0106_),
    .CK(clknet_4_10_0_clk),
    .Q(\memory[5][2] ),
    .QN(_0453_));
 DFF_X1 \memory[5][3]$_DFFE_PP_  (.D(_0107_),
    .CK(clknet_4_2_0_clk),
    .Q(\memory[5][3] ),
    .QN(_0452_));
 DFF_X1 \memory[5][4]$_DFFE_PP_  (.D(_0108_),
    .CK(clknet_4_0_0_clk),
    .Q(\memory[5][4] ),
    .QN(_0451_));
 DFF_X1 \memory[5][5]$_DFFE_PP_  (.D(_0109_),
    .CK(clknet_4_11_0_clk),
    .Q(\memory[5][5] ),
    .QN(_0450_));
 DFF_X1 \memory[5][6]$_DFFE_PP_  (.D(_0110_),
    .CK(clknet_4_2_0_clk),
    .Q(\memory[5][6] ),
    .QN(_0449_));
 DFF_X1 \memory[5][7]$_DFFE_PP_  (.D(_0111_),
    .CK(clknet_4_10_0_clk),
    .Q(\memory[5][7] ),
    .QN(_0448_));
 DFF_X1 \memory[6][0]$_DFFE_PP_  (.D(_0112_),
    .CK(clknet_4_15_0_clk),
    .Q(\memory[6][0] ),
    .QN(_0447_));
 DFF_X1 \memory[6][1]$_DFFE_PP_  (.D(_0113_),
    .CK(clknet_4_4_0_clk),
    .Q(\memory[6][1] ),
    .QN(_0446_));
 DFF_X1 \memory[6][2]$_DFFE_PP_  (.D(_0114_),
    .CK(clknet_4_14_0_clk),
    .Q(\memory[6][2] ),
    .QN(_0445_));
 DFF_X1 \memory[6][3]$_DFFE_PP_  (.D(_0115_),
    .CK(clknet_4_12_0_clk),
    .Q(\memory[6][3] ),
    .QN(_0444_));
 DFF_X1 \memory[6][4]$_DFFE_PP_  (.D(_0116_),
    .CK(clknet_4_1_0_clk),
    .Q(\memory[6][4] ),
    .QN(_0443_));
 DFF_X1 \memory[6][5]$_DFFE_PP_  (.D(_0117_),
    .CK(clknet_4_15_0_clk),
    .Q(\memory[6][5] ),
    .QN(_0442_));
 DFF_X1 \memory[6][6]$_DFFE_PP_  (.D(_0118_),
    .CK(clknet_4_6_0_clk),
    .Q(\memory[6][6] ),
    .QN(_0441_));
 DFF_X1 \memory[6][7]$_DFFE_PP_  (.D(_0119_),
    .CK(clknet_4_11_0_clk),
    .Q(\memory[6][7] ),
    .QN(_0440_));
 DFF_X1 \memory[7][0]$_DFFE_PP_  (.D(_0120_),
    .CK(clknet_4_15_0_clk),
    .Q(\memory[7][0] ),
    .QN(_0439_));
 DFF_X1 \memory[7][1]$_DFFE_PP_  (.D(_0121_),
    .CK(clknet_4_1_0_clk),
    .Q(\memory[7][1] ),
    .QN(_0438_));
 DFF_X1 \memory[7][2]$_DFFE_PP_  (.D(_0122_),
    .CK(clknet_4_10_0_clk),
    .Q(\memory[7][2] ),
    .QN(_0437_));
 DFF_X1 \memory[7][3]$_DFFE_PP_  (.D(_0123_),
    .CK(clknet_4_8_0_clk),
    .Q(\memory[7][3] ),
    .QN(_0436_));
 DFF_X1 \memory[7][4]$_DFFE_PP_  (.D(_0124_),
    .CK(clknet_4_0_0_clk),
    .Q(\memory[7][4] ),
    .QN(_0435_));
 DFF_X1 \memory[7][5]$_DFFE_PP_  (.D(_0125_),
    .CK(clknet_4_10_0_clk),
    .Q(\memory[7][5] ),
    .QN(_0434_));
 DFF_X1 \memory[7][6]$_DFFE_PP_  (.D(_0126_),
    .CK(clknet_4_2_0_clk),
    .Q(\memory[7][6] ),
    .QN(_0433_));
 DFF_X1 \memory[7][7]$_DFFE_PP_  (.D(_0127_),
    .CK(clknet_4_10_0_clk),
    .Q(\memory[7][7] ),
    .QN(_0432_));
 DFF_X1 \memory[8][0]$_DFFE_PP_  (.D(_0128_),
    .CK(clknet_4_15_0_clk),
    .Q(\memory[8][0] ),
    .QN(_0431_));
 DFF_X1 \memory[8][1]$_DFFE_PP_  (.D(_0129_),
    .CK(clknet_4_5_0_clk),
    .Q(\memory[8][1] ),
    .QN(_0430_));
 DFF_X1 \memory[8][2]$_DFFE_PP_  (.D(_0130_),
    .CK(clknet_4_14_0_clk),
    .Q(\memory[8][2] ),
    .QN(_0429_));
 DFF_X1 \memory[8][3]$_DFFE_PP_  (.D(_0131_),
    .CK(clknet_4_3_0_clk),
    .Q(\memory[8][3] ),
    .QN(_0428_));
 DFF_X1 \memory[8][4]$_DFFE_PP_  (.D(_0132_),
    .CK(clknet_4_1_0_clk),
    .Q(\memory[8][4] ),
    .QN(_0427_));
 DFF_X1 \memory[8][5]$_DFFE_PP_  (.D(_0133_),
    .CK(clknet_4_14_0_clk),
    .Q(\memory[8][5] ),
    .QN(_0426_));
 DFF_X1 \memory[8][6]$_DFFE_PP_  (.D(_0134_),
    .CK(clknet_4_1_0_clk),
    .Q(\memory[8][6] ),
    .QN(_0425_));
 DFF_X1 \memory[8][7]$_DFFE_PP_  (.D(_0135_),
    .CK(clknet_4_11_0_clk),
    .Q(\memory[8][7] ),
    .QN(_0424_));
 DFF_X1 \memory[9][0]$_DFFE_PP_  (.D(_0136_),
    .CK(clknet_4_15_0_clk),
    .Q(\memory[9][0] ),
    .QN(_0423_));
 DFF_X1 \memory[9][1]$_DFFE_PP_  (.D(_0137_),
    .CK(clknet_4_0_0_clk),
    .Q(\memory[9][1] ),
    .QN(_0422_));
 DFF_X1 \memory[9][2]$_DFFE_PP_  (.D(_0138_),
    .CK(clknet_4_10_0_clk),
    .Q(\memory[9][2] ),
    .QN(_0421_));
 DFF_X1 \memory[9][3]$_DFFE_PP_  (.D(_0139_),
    .CK(clknet_4_2_0_clk),
    .Q(\memory[9][3] ),
    .QN(_0420_));
 DFF_X1 \memory[9][4]$_DFFE_PP_  (.D(_0140_),
    .CK(clknet_4_0_0_clk),
    .Q(\memory[9][4] ),
    .QN(_0419_));
 DFF_X1 \memory[9][5]$_DFFE_PP_  (.D(_0141_),
    .CK(clknet_4_15_0_clk),
    .Q(\memory[9][5] ),
    .QN(_0418_));
 DFF_X1 \memory[9][6]$_DFFE_PP_  (.D(_0142_),
    .CK(clknet_4_2_0_clk),
    .Q(\memory[9][6] ),
    .QN(_0417_));
 DFF_X1 \memory[9][7]$_DFFE_PP_  (.D(_0143_),
    .CK(clknet_4_10_0_clk),
    .Q(\memory[9][7] ),
    .QN(_0416_));
 DFF_X1 \rd_ptr[0]$_SDFFE_PN0P_  (.D(_0144_),
    .CK(clknet_4_13_0_clk),
    .Q(\rd_ptr[0] ),
    .QN(_0415_));
 DFF_X1 \rd_ptr[1]$_SDFFE_PN0P_  (.D(_0145_),
    .CK(clknet_4_13_0_clk),
    .Q(\rd_ptr[1] ),
    .QN(_0414_));
 DFF_X1 \rd_ptr[2]$_SDFFE_PN0P_  (.D(_0146_),
    .CK(clknet_4_7_0_clk),
    .Q(\rd_ptr[2] ),
    .QN(_0413_));
 DFF_X1 \rd_ptr[3]$_SDFFE_PN0P_  (.D(_0147_),
    .CK(clknet_4_7_0_clk),
    .Q(\rd_ptr[3] ),
    .QN(_0412_));
 DFF_X2 \wr_ptr[0]$_SDFFE_PN0P_  (.D(_0148_),
    .CK(clknet_4_5_0_clk),
    .Q(\wr_ptr[0] ),
    .QN(_0560_));
 DFF_X2 \wr_ptr[1]$_SDFFE_PN0P_  (.D(_0149_),
    .CK(clknet_4_5_0_clk),
    .Q(\wr_ptr[1] ),
    .QN(_0561_));
 DFF_X1 \wr_ptr[2]$_SDFFE_PN0P_  (.D(_0150_),
    .CK(clknet_4_5_0_clk),
    .Q(\wr_ptr[2] ),
    .QN(_0411_));
 DFF_X1 \wr_ptr[3]$_SDFFE_PN0P_  (.D(_0151_),
    .CK(clknet_4_5_0_clk),
    .Q(\wr_ptr[3] ),
    .QN(_0410_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_73 ();
 BUF_X1 input1 (.A(rd_en),
    .Z(net1));
 BUF_X1 input2 (.A(wr_en),
    .Z(net2));
 BUF_X1 output3 (.A(net3),
    .Z(almost_empty));
 BUF_X1 output4 (.A(net4),
    .Z(almost_full));
 BUF_X1 output5 (.A(net5),
    .Z(data_out[0]));
 BUF_X1 output6 (.A(net6),
    .Z(data_out[1]));
 BUF_X1 output7 (.A(net7),
    .Z(data_out[2]));
 BUF_X1 output8 (.A(net8),
    .Z(data_out[3]));
 BUF_X1 output9 (.A(net9),
    .Z(data_out[4]));
 BUF_X1 output10 (.A(net10),
    .Z(data_out[5]));
 BUF_X1 output11 (.A(net11),
    .Z(data_out[6]));
 BUF_X1 output12 (.A(net12),
    .Z(data_out[7]));
 BUF_X1 output13 (.A(net13),
    .Z(empty));
 BUF_X1 output14 (.A(net14),
    .Z(fill_level[0]));
 BUF_X1 output15 (.A(net15),
    .Z(fill_level[1]));
 BUF_X1 output16 (.A(net16),
    .Z(fill_level[2]));
 BUF_X1 output17 (.A(net17),
    .Z(fill_level[3]));
 BUF_X1 output18 (.A(net18),
    .Z(fill_level[4]));
 BUF_X1 output19 (.A(net19),
    .Z(full));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 CLKBUF_X3 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 CLKBUF_X3 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 CLKBUF_X3 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 CLKBUF_X3 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 CLKBUF_X3 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 CLKBUF_X3 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 CLKBUF_X3 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 CLKBUF_X3 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 CLKBUF_X3 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 CLKBUF_X3 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 CLKBUF_X3 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 CLKBUF_X3 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 CLKBUF_X3 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 CLKBUF_X3 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 CLKBUF_X3 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 INV_X2 clkload0 (.A(clknet_4_0_0_clk));
 INV_X4 clkload1 (.A(clknet_4_1_0_clk));
 INV_X2 clkload2 (.A(clknet_4_2_0_clk));
 INV_X8 clkload3 (.A(clknet_4_3_0_clk));
 INV_X4 clkload4 (.A(clknet_4_4_0_clk));
 INV_X4 clkload5 (.A(clknet_4_5_0_clk));
 INV_X8 clkload6 (.A(clknet_4_6_0_clk));
 INV_X4 clkload7 (.A(clknet_4_7_0_clk));
 INV_X4 clkload8 (.A(clknet_4_8_0_clk));
 INV_X8 clkload9 (.A(clknet_4_9_0_clk));
 INV_X2 clkload10 (.A(clknet_4_10_0_clk));
 INV_X4 clkload11 (.A(clknet_4_11_0_clk));
 INV_X4 clkload12 (.A(clknet_4_12_0_clk));
 INV_X2 clkload13 (.A(clknet_4_13_0_clk));
 INV_X2 clkload14 (.A(clknet_4_14_0_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X8 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_77 ();
 FILLCELL_X32 FILLER_0_109 ();
 FILLCELL_X32 FILLER_0_141 ();
 FILLCELL_X8 FILLER_0_173 ();
 FILLCELL_X1 FILLER_0_181 ();
 FILLCELL_X32 FILLER_0_201 ();
 FILLCELL_X32 FILLER_0_233 ();
 FILLCELL_X8 FILLER_0_265 ();
 FILLCELL_X4 FILLER_0_273 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X16 FILLER_1_161 ();
 FILLCELL_X4 FILLER_1_177 ();
 FILLCELL_X8 FILLER_1_210 ();
 FILLCELL_X4 FILLER_1_218 ();
 FILLCELL_X1 FILLER_1_222 ();
 FILLCELL_X4 FILLER_1_242 ();
 FILLCELL_X2 FILLER_1_246 ();
 FILLCELL_X1 FILLER_1_248 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X8 FILLER_2_129 ();
 FILLCELL_X4 FILLER_2_137 ();
 FILLCELL_X1 FILLER_2_141 ();
 FILLCELL_X32 FILLER_2_149 ();
 FILLCELL_X2 FILLER_2_181 ();
 FILLCELL_X1 FILLER_2_183 ();
 FILLCELL_X1 FILLER_2_208 ();
 FILLCELL_X4 FILLER_2_214 ();
 FILLCELL_X2 FILLER_2_218 ();
 FILLCELL_X2 FILLER_2_274 ();
 FILLCELL_X1 FILLER_2_276 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X8 FILLER_3_97 ();
 FILLCELL_X4 FILLER_3_105 ();
 FILLCELL_X1 FILLER_3_109 ();
 FILLCELL_X1 FILLER_3_117 ();
 FILLCELL_X16 FILLER_3_152 ();
 FILLCELL_X1 FILLER_3_168 ();
 FILLCELL_X2 FILLER_3_200 ();
 FILLCELL_X2 FILLER_3_209 ();
 FILLCELL_X1 FILLER_3_211 ();
 FILLCELL_X8 FILLER_3_217 ();
 FILLCELL_X2 FILLER_3_225 ();
 FILLCELL_X1 FILLER_3_243 ();
 FILLCELL_X1 FILLER_3_250 ();
 FILLCELL_X1 FILLER_3_273 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X8 FILLER_4_65 ();
 FILLCELL_X2 FILLER_4_73 ();
 FILLCELL_X1 FILLER_4_75 ();
 FILLCELL_X8 FILLER_4_93 ();
 FILLCELL_X2 FILLER_4_101 ();
 FILLCELL_X1 FILLER_4_103 ();
 FILLCELL_X16 FILLER_4_108 ();
 FILLCELL_X4 FILLER_4_124 ();
 FILLCELL_X2 FILLER_4_128 ();
 FILLCELL_X1 FILLER_4_130 ();
 FILLCELL_X16 FILLER_4_138 ();
 FILLCELL_X1 FILLER_4_154 ();
 FILLCELL_X4 FILLER_4_179 ();
 FILLCELL_X2 FILLER_4_183 ();
 FILLCELL_X1 FILLER_4_192 ();
 FILLCELL_X4 FILLER_4_210 ();
 FILLCELL_X1 FILLER_4_214 ();
 FILLCELL_X4 FILLER_4_220 ();
 FILLCELL_X1 FILLER_4_224 ();
 FILLCELL_X4 FILLER_4_228 ();
 FILLCELL_X2 FILLER_4_232 ();
 FILLCELL_X2 FILLER_4_241 ();
 FILLCELL_X1 FILLER_4_276 ();
 FILLCELL_X8 FILLER_5_1 ();
 FILLCELL_X4 FILLER_5_9 ();
 FILLCELL_X1 FILLER_5_13 ();
 FILLCELL_X2 FILLER_5_48 ();
 FILLCELL_X1 FILLER_5_50 ();
 FILLCELL_X4 FILLER_5_55 ();
 FILLCELL_X8 FILLER_5_93 ();
 FILLCELL_X1 FILLER_5_101 ();
 FILLCELL_X4 FILLER_5_119 ();
 FILLCELL_X1 FILLER_5_123 ();
 FILLCELL_X8 FILLER_5_148 ();
 FILLCELL_X1 FILLER_5_156 ();
 FILLCELL_X16 FILLER_5_164 ();
 FILLCELL_X8 FILLER_5_180 ();
 FILLCELL_X16 FILLER_5_210 ();
 FILLCELL_X8 FILLER_5_226 ();
 FILLCELL_X2 FILLER_5_244 ();
 FILLCELL_X1 FILLER_5_250 ();
 FILLCELL_X2 FILLER_5_257 ();
 FILLCELL_X4 FILLER_5_269 ();
 FILLCELL_X1 FILLER_5_273 ();
 FILLCELL_X8 FILLER_6_1 ();
 FILLCELL_X1 FILLER_6_9 ();
 FILLCELL_X2 FILLER_6_27 ();
 FILLCELL_X2 FILLER_6_36 ();
 FILLCELL_X1 FILLER_6_38 ();
 FILLCELL_X2 FILLER_6_56 ();
 FILLCELL_X4 FILLER_6_75 ();
 FILLCELL_X1 FILLER_6_86 ();
 FILLCELL_X1 FILLER_6_118 ();
 FILLCELL_X4 FILLER_6_133 ();
 FILLCELL_X2 FILLER_6_137 ();
 FILLCELL_X1 FILLER_6_163 ();
 FILLCELL_X1 FILLER_6_188 ();
 FILLCELL_X1 FILLER_6_199 ();
 FILLCELL_X1 FILLER_6_209 ();
 FILLCELL_X4 FILLER_6_228 ();
 FILLCELL_X2 FILLER_6_232 ();
 FILLCELL_X2 FILLER_6_251 ();
 FILLCELL_X1 FILLER_6_253 ();
 FILLCELL_X4 FILLER_6_270 ();
 FILLCELL_X2 FILLER_6_274 ();
 FILLCELL_X1 FILLER_6_276 ();
 FILLCELL_X8 FILLER_7_1 ();
 FILLCELL_X1 FILLER_7_9 ();
 FILLCELL_X4 FILLER_7_31 ();
 FILLCELL_X2 FILLER_7_35 ();
 FILLCELL_X4 FILLER_7_51 ();
 FILLCELL_X2 FILLER_7_55 ();
 FILLCELL_X2 FILLER_7_78 ();
 FILLCELL_X2 FILLER_7_87 ();
 FILLCELL_X1 FILLER_7_89 ();
 FILLCELL_X4 FILLER_7_97 ();
 FILLCELL_X2 FILLER_7_101 ();
 FILLCELL_X16 FILLER_7_110 ();
 FILLCELL_X4 FILLER_7_133 ();
 FILLCELL_X2 FILLER_7_137 ();
 FILLCELL_X1 FILLER_7_139 ();
 FILLCELL_X8 FILLER_7_171 ();
 FILLCELL_X4 FILLER_7_179 ();
 FILLCELL_X2 FILLER_7_183 ();
 FILLCELL_X1 FILLER_7_185 ();
 FILLCELL_X1 FILLER_7_193 ();
 FILLCELL_X1 FILLER_7_197 ();
 FILLCELL_X1 FILLER_7_230 ();
 FILLCELL_X4 FILLER_7_249 ();
 FILLCELL_X1 FILLER_7_253 ();
 FILLCELL_X1 FILLER_7_276 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X8 FILLER_8_33 ();
 FILLCELL_X4 FILLER_8_41 ();
 FILLCELL_X1 FILLER_8_45 ();
 FILLCELL_X32 FILLER_8_53 ();
 FILLCELL_X32 FILLER_8_85 ();
 FILLCELL_X4 FILLER_8_117 ();
 FILLCELL_X2 FILLER_8_121 ();
 FILLCELL_X16 FILLER_8_140 ();
 FILLCELL_X2 FILLER_8_156 ();
 FILLCELL_X1 FILLER_8_158 ();
 FILLCELL_X8 FILLER_8_176 ();
 FILLCELL_X2 FILLER_8_184 ();
 FILLCELL_X1 FILLER_8_186 ();
 FILLCELL_X1 FILLER_8_213 ();
 FILLCELL_X4 FILLER_8_239 ();
 FILLCELL_X8 FILLER_9_1 ();
 FILLCELL_X4 FILLER_9_9 ();
 FILLCELL_X8 FILLER_9_17 ();
 FILLCELL_X2 FILLER_9_25 ();
 FILLCELL_X1 FILLER_9_27 ();
 FILLCELL_X8 FILLER_9_45 ();
 FILLCELL_X4 FILLER_9_53 ();
 FILLCELL_X1 FILLER_9_74 ();
 FILLCELL_X4 FILLER_9_82 ();
 FILLCELL_X32 FILLER_9_93 ();
 FILLCELL_X16 FILLER_9_125 ();
 FILLCELL_X2 FILLER_9_141 ();
 FILLCELL_X1 FILLER_9_143 ();
 FILLCELL_X8 FILLER_9_149 ();
 FILLCELL_X2 FILLER_9_164 ();
 FILLCELL_X1 FILLER_9_166 ();
 FILLCELL_X4 FILLER_9_174 ();
 FILLCELL_X2 FILLER_9_178 ();
 FILLCELL_X1 FILLER_9_180 ();
 FILLCELL_X2 FILLER_9_186 ();
 FILLCELL_X2 FILLER_9_202 ();
 FILLCELL_X16 FILLER_9_221 ();
 FILLCELL_X8 FILLER_9_237 ();
 FILLCELL_X2 FILLER_10_1 ();
 FILLCELL_X1 FILLER_10_3 ();
 FILLCELL_X1 FILLER_10_21 ();
 FILLCELL_X1 FILLER_10_29 ();
 FILLCELL_X1 FILLER_10_37 ();
 FILLCELL_X2 FILLER_10_55 ();
 FILLCELL_X2 FILLER_10_81 ();
 FILLCELL_X4 FILLER_10_107 ();
 FILLCELL_X4 FILLER_10_128 ();
 FILLCELL_X2 FILLER_10_132 ();
 FILLCELL_X2 FILLER_10_141 ();
 FILLCELL_X1 FILLER_10_143 ();
 FILLCELL_X1 FILLER_10_156 ();
 FILLCELL_X4 FILLER_10_186 ();
 FILLCELL_X1 FILLER_10_204 ();
 FILLCELL_X2 FILLER_10_232 ();
 FILLCELL_X2 FILLER_10_251 ();
 FILLCELL_X2 FILLER_10_265 ();
 FILLCELL_X1 FILLER_10_267 ();
 FILLCELL_X16 FILLER_11_1 ();
 FILLCELL_X4 FILLER_11_28 ();
 FILLCELL_X16 FILLER_11_46 ();
 FILLCELL_X1 FILLER_11_62 ();
 FILLCELL_X4 FILLER_11_78 ();
 FILLCELL_X2 FILLER_11_82 ();
 FILLCELL_X4 FILLER_11_91 ();
 FILLCELL_X1 FILLER_11_95 ();
 FILLCELL_X2 FILLER_11_147 ();
 FILLCELL_X1 FILLER_11_149 ();
 FILLCELL_X4 FILLER_11_167 ();
 FILLCELL_X2 FILLER_11_171 ();
 FILLCELL_X4 FILLER_11_197 ();
 FILLCELL_X1 FILLER_11_201 ();
 FILLCELL_X2 FILLER_11_215 ();
 FILLCELL_X1 FILLER_11_217 ();
 FILLCELL_X4 FILLER_11_231 ();
 FILLCELL_X1 FILLER_11_235 ();
 FILLCELL_X8 FILLER_11_256 ();
 FILLCELL_X2 FILLER_11_274 ();
 FILLCELL_X1 FILLER_11_276 ();
 FILLCELL_X1 FILLER_12_1 ();
 FILLCELL_X8 FILLER_12_33 ();
 FILLCELL_X4 FILLER_12_41 ();
 FILLCELL_X2 FILLER_12_45 ();
 FILLCELL_X1 FILLER_12_47 ();
 FILLCELL_X8 FILLER_12_55 ();
 FILLCELL_X2 FILLER_12_63 ();
 FILLCELL_X2 FILLER_12_89 ();
 FILLCELL_X8 FILLER_12_98 ();
 FILLCELL_X4 FILLER_12_106 ();
 FILLCELL_X1 FILLER_12_110 ();
 FILLCELL_X1 FILLER_12_125 ();
 FILLCELL_X1 FILLER_12_133 ();
 FILLCELL_X2 FILLER_12_141 ();
 FILLCELL_X2 FILLER_12_150 ();
 FILLCELL_X2 FILLER_12_161 ();
 FILLCELL_X1 FILLER_12_163 ();
 FILLCELL_X16 FILLER_12_178 ();
 FILLCELL_X8 FILLER_12_194 ();
 FILLCELL_X2 FILLER_12_202 ();
 FILLCELL_X1 FILLER_12_204 ();
 FILLCELL_X16 FILLER_12_231 ();
 FILLCELL_X2 FILLER_12_247 ();
 FILLCELL_X1 FILLER_12_252 ();
 FILLCELL_X2 FILLER_12_256 ();
 FILLCELL_X1 FILLER_12_258 ();
 FILLCELL_X8 FILLER_12_262 ();
 FILLCELL_X4 FILLER_12_270 ();
 FILLCELL_X2 FILLER_12_274 ();
 FILLCELL_X1 FILLER_12_276 ();
 FILLCELL_X16 FILLER_13_1 ();
 FILLCELL_X8 FILLER_13_17 ();
 FILLCELL_X4 FILLER_13_25 ();
 FILLCELL_X2 FILLER_13_53 ();
 FILLCELL_X16 FILLER_13_72 ();
 FILLCELL_X4 FILLER_13_88 ();
 FILLCELL_X2 FILLER_13_92 ();
 FILLCELL_X1 FILLER_13_94 ();
 FILLCELL_X32 FILLER_13_119 ();
 FILLCELL_X16 FILLER_13_151 ();
 FILLCELL_X2 FILLER_13_167 ();
 FILLCELL_X16 FILLER_13_181 ();
 FILLCELL_X4 FILLER_13_197 ();
 FILLCELL_X2 FILLER_13_201 ();
 FILLCELL_X1 FILLER_13_203 ();
 FILLCELL_X8 FILLER_13_230 ();
 FILLCELL_X1 FILLER_13_256 ();
 FILLCELL_X2 FILLER_13_274 ();
 FILLCELL_X1 FILLER_13_276 ();
 FILLCELL_X4 FILLER_14_1 ();
 FILLCELL_X2 FILLER_14_5 ();
 FILLCELL_X1 FILLER_14_7 ();
 FILLCELL_X4 FILLER_14_25 ();
 FILLCELL_X2 FILLER_14_29 ();
 FILLCELL_X4 FILLER_14_35 ();
 FILLCELL_X2 FILLER_14_39 ();
 FILLCELL_X2 FILLER_14_48 ();
 FILLCELL_X1 FILLER_14_50 ();
 FILLCELL_X8 FILLER_14_82 ();
 FILLCELL_X4 FILLER_14_90 ();
 FILLCELL_X1 FILLER_14_94 ();
 FILLCELL_X8 FILLER_14_112 ();
 FILLCELL_X8 FILLER_14_137 ();
 FILLCELL_X4 FILLER_14_145 ();
 FILLCELL_X2 FILLER_14_149 ();
 FILLCELL_X1 FILLER_14_151 ();
 FILLCELL_X4 FILLER_14_190 ();
 FILLCELL_X1 FILLER_14_204 ();
 FILLCELL_X16 FILLER_14_218 ();
 FILLCELL_X2 FILLER_14_234 ();
 FILLCELL_X1 FILLER_14_236 ();
 FILLCELL_X2 FILLER_14_255 ();
 FILLCELL_X4 FILLER_15_1 ();
 FILLCELL_X1 FILLER_15_5 ();
 FILLCELL_X1 FILLER_15_54 ();
 FILLCELL_X1 FILLER_15_79 ();
 FILLCELL_X2 FILLER_15_87 ();
 FILLCELL_X1 FILLER_15_103 ();
 FILLCELL_X4 FILLER_15_118 ();
 FILLCELL_X1 FILLER_15_122 ();
 FILLCELL_X1 FILLER_15_130 ();
 FILLCELL_X16 FILLER_15_176 ();
 FILLCELL_X8 FILLER_15_192 ();
 FILLCELL_X4 FILLER_15_200 ();
 FILLCELL_X8 FILLER_15_226 ();
 FILLCELL_X4 FILLER_15_234 ();
 FILLCELL_X1 FILLER_15_243 ();
 FILLCELL_X1 FILLER_15_248 ();
 FILLCELL_X2 FILLER_15_257 ();
 FILLCELL_X1 FILLER_15_259 ();
 FILLCELL_X2 FILLER_15_271 ();
 FILLCELL_X1 FILLER_15_273 ();
 FILLCELL_X8 FILLER_16_1 ();
 FILLCELL_X4 FILLER_16_9 ();
 FILLCELL_X2 FILLER_16_13 ();
 FILLCELL_X16 FILLER_16_29 ();
 FILLCELL_X4 FILLER_16_45 ();
 FILLCELL_X1 FILLER_16_56 ();
 FILLCELL_X2 FILLER_16_93 ();
 FILLCELL_X1 FILLER_16_95 ();
 FILLCELL_X1 FILLER_16_103 ();
 FILLCELL_X2 FILLER_16_135 ();
 FILLCELL_X16 FILLER_16_185 ();
 FILLCELL_X8 FILLER_16_201 ();
 FILLCELL_X2 FILLER_16_209 ();
 FILLCELL_X8 FILLER_16_214 ();
 FILLCELL_X2 FILLER_16_222 ();
 FILLCELL_X1 FILLER_16_245 ();
 FILLCELL_X2 FILLER_16_253 ();
 FILLCELL_X8 FILLER_16_259 ();
 FILLCELL_X4 FILLER_16_270 ();
 FILLCELL_X16 FILLER_17_1 ();
 FILLCELL_X8 FILLER_17_17 ();
 FILLCELL_X4 FILLER_17_25 ();
 FILLCELL_X1 FILLER_17_29 ();
 FILLCELL_X8 FILLER_17_47 ();
 FILLCELL_X2 FILLER_17_55 ();
 FILLCELL_X4 FILLER_17_60 ();
 FILLCELL_X2 FILLER_17_64 ();
 FILLCELL_X1 FILLER_17_66 ();
 FILLCELL_X2 FILLER_17_74 ();
 FILLCELL_X8 FILLER_17_83 ();
 FILLCELL_X1 FILLER_17_91 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X16 FILLER_17_129 ();
 FILLCELL_X8 FILLER_17_145 ();
 FILLCELL_X1 FILLER_17_153 ();
 FILLCELL_X32 FILLER_17_170 ();
 FILLCELL_X4 FILLER_17_202 ();
 FILLCELL_X2 FILLER_17_206 ();
 FILLCELL_X4 FILLER_17_228 ();
 FILLCELL_X2 FILLER_17_232 ();
 FILLCELL_X2 FILLER_17_253 ();
 FILLCELL_X1 FILLER_17_255 ();
 FILLCELL_X8 FILLER_17_263 ();
 FILLCELL_X2 FILLER_17_271 ();
 FILLCELL_X1 FILLER_17_273 ();
 FILLCELL_X2 FILLER_18_1 ();
 FILLCELL_X1 FILLER_18_3 ();
 FILLCELL_X4 FILLER_18_28 ();
 FILLCELL_X1 FILLER_18_32 ();
 FILLCELL_X16 FILLER_18_50 ();
 FILLCELL_X8 FILLER_18_66 ();
 FILLCELL_X2 FILLER_18_74 ();
 FILLCELL_X1 FILLER_18_76 ();
 FILLCELL_X2 FILLER_18_84 ();
 FILLCELL_X1 FILLER_18_86 ();
 FILLCELL_X1 FILLER_18_94 ();
 FILLCELL_X8 FILLER_18_102 ();
 FILLCELL_X4 FILLER_18_110 ();
 FILLCELL_X1 FILLER_18_114 ();
 FILLCELL_X1 FILLER_18_122 ();
 FILLCELL_X8 FILLER_18_145 ();
 FILLCELL_X32 FILLER_18_166 ();
 FILLCELL_X8 FILLER_18_198 ();
 FILLCELL_X4 FILLER_18_206 ();
 FILLCELL_X1 FILLER_18_210 ();
 FILLCELL_X4 FILLER_18_218 ();
 FILLCELL_X2 FILLER_18_246 ();
 FILLCELL_X4 FILLER_18_253 ();
 FILLCELL_X2 FILLER_18_274 ();
 FILLCELL_X1 FILLER_18_276 ();
 FILLCELL_X2 FILLER_19_1 ();
 FILLCELL_X1 FILLER_19_3 ();
 FILLCELL_X1 FILLER_19_28 ();
 FILLCELL_X16 FILLER_19_50 ();
 FILLCELL_X4 FILLER_19_66 ();
 FILLCELL_X2 FILLER_19_70 ();
 FILLCELL_X2 FILLER_19_96 ();
 FILLCELL_X1 FILLER_19_98 ();
 FILLCELL_X1 FILLER_19_123 ();
 FILLCELL_X2 FILLER_19_131 ();
 FILLCELL_X4 FILLER_19_140 ();
 FILLCELL_X2 FILLER_19_151 ();
 FILLCELL_X4 FILLER_19_162 ();
 FILLCELL_X1 FILLER_19_173 ();
 FILLCELL_X4 FILLER_19_223 ();
 FILLCELL_X2 FILLER_19_227 ();
 FILLCELL_X1 FILLER_19_229 ();
 FILLCELL_X4 FILLER_19_234 ();
 FILLCELL_X4 FILLER_19_252 ();
 FILLCELL_X2 FILLER_19_256 ();
 FILLCELL_X1 FILLER_19_258 ();
 FILLCELL_X2 FILLER_19_262 ();
 FILLCELL_X1 FILLER_19_264 ();
 FILLCELL_X4 FILLER_19_269 ();
 FILLCELL_X1 FILLER_19_273 ();
 FILLCELL_X8 FILLER_20_1 ();
 FILLCELL_X2 FILLER_20_9 ();
 FILLCELL_X8 FILLER_20_22 ();
 FILLCELL_X2 FILLER_20_30 ();
 FILLCELL_X1 FILLER_20_32 ();
 FILLCELL_X8 FILLER_20_37 ();
 FILLCELL_X1 FILLER_20_45 ();
 FILLCELL_X16 FILLER_20_77 ();
 FILLCELL_X4 FILLER_20_93 ();
 FILLCELL_X1 FILLER_20_97 ();
 FILLCELL_X8 FILLER_20_105 ();
 FILLCELL_X2 FILLER_20_113 ();
 FILLCELL_X1 FILLER_20_122 ();
 FILLCELL_X4 FILLER_20_140 ();
 FILLCELL_X2 FILLER_20_178 ();
 FILLCELL_X1 FILLER_20_180 ();
 FILLCELL_X16 FILLER_20_188 ();
 FILLCELL_X2 FILLER_20_204 ();
 FILLCELL_X8 FILLER_20_213 ();
 FILLCELL_X4 FILLER_20_221 ();
 FILLCELL_X1 FILLER_20_225 ();
 FILLCELL_X2 FILLER_20_250 ();
 FILLCELL_X1 FILLER_20_276 ();
 FILLCELL_X16 FILLER_21_1 ();
 FILLCELL_X2 FILLER_21_24 ();
 FILLCELL_X1 FILLER_21_26 ();
 FILLCELL_X4 FILLER_21_34 ();
 FILLCELL_X2 FILLER_21_38 ();
 FILLCELL_X2 FILLER_21_47 ();
 FILLCELL_X1 FILLER_21_49 ();
 FILLCELL_X4 FILLER_21_57 ();
 FILLCELL_X2 FILLER_21_61 ();
 FILLCELL_X16 FILLER_21_77 ();
 FILLCELL_X4 FILLER_21_93 ();
 FILLCELL_X8 FILLER_21_114 ();
 FILLCELL_X4 FILLER_21_122 ();
 FILLCELL_X1 FILLER_21_126 ();
 FILLCELL_X8 FILLER_21_141 ();
 FILLCELL_X4 FILLER_21_149 ();
 FILLCELL_X1 FILLER_21_153 ();
 FILLCELL_X4 FILLER_21_175 ();
 FILLCELL_X1 FILLER_21_179 ();
 FILLCELL_X32 FILLER_21_204 ();
 FILLCELL_X8 FILLER_21_236 ();
 FILLCELL_X1 FILLER_21_244 ();
 FILLCELL_X1 FILLER_21_250 ();
 FILLCELL_X2 FILLER_21_274 ();
 FILLCELL_X1 FILLER_21_276 ();
 FILLCELL_X8 FILLER_22_1 ();
 FILLCELL_X2 FILLER_22_9 ();
 FILLCELL_X1 FILLER_22_11 ();
 FILLCELL_X16 FILLER_22_46 ();
 FILLCELL_X2 FILLER_22_62 ();
 FILLCELL_X1 FILLER_22_64 ();
 FILLCELL_X32 FILLER_22_82 ();
 FILLCELL_X32 FILLER_22_114 ();
 FILLCELL_X32 FILLER_22_146 ();
 FILLCELL_X16 FILLER_22_178 ();
 FILLCELL_X8 FILLER_22_194 ();
 FILLCELL_X4 FILLER_22_202 ();
 FILLCELL_X1 FILLER_22_206 ();
 FILLCELL_X16 FILLER_22_224 ();
 FILLCELL_X8 FILLER_22_240 ();
 FILLCELL_X2 FILLER_22_248 ();
 FILLCELL_X1 FILLER_22_250 ();
 FILLCELL_X8 FILLER_22_263 ();
 FILLCELL_X16 FILLER_23_1 ();
 FILLCELL_X16 FILLER_23_31 ();
 FILLCELL_X4 FILLER_23_47 ();
 FILLCELL_X1 FILLER_23_51 ();
 FILLCELL_X2 FILLER_23_76 ();
 FILLCELL_X2 FILLER_23_85 ();
 FILLCELL_X4 FILLER_23_94 ();
 FILLCELL_X2 FILLER_23_98 ();
 FILLCELL_X16 FILLER_23_134 ();
 FILLCELL_X1 FILLER_23_150 ();
 FILLCELL_X1 FILLER_23_182 ();
 FILLCELL_X8 FILLER_23_200 ();
 FILLCELL_X2 FILLER_23_208 ();
 FILLCELL_X1 FILLER_23_210 ();
 FILLCELL_X8 FILLER_23_235 ();
 FILLCELL_X4 FILLER_23_243 ();
 FILLCELL_X2 FILLER_23_247 ();
 FILLCELL_X8 FILLER_23_269 ();
 FILLCELL_X2 FILLER_24_1 ();
 FILLCELL_X16 FILLER_24_37 ();
 FILLCELL_X4 FILLER_24_53 ();
 FILLCELL_X2 FILLER_24_57 ();
 FILLCELL_X1 FILLER_24_59 ();
 FILLCELL_X4 FILLER_24_79 ();
 FILLCELL_X2 FILLER_24_107 ();
 FILLCELL_X2 FILLER_24_118 ();
 FILLCELL_X1 FILLER_24_120 ();
 FILLCELL_X8 FILLER_24_135 ();
 FILLCELL_X2 FILLER_24_143 ();
 FILLCELL_X1 FILLER_24_145 ();
 FILLCELL_X1 FILLER_24_163 ();
 FILLCELL_X1 FILLER_24_171 ();
 FILLCELL_X1 FILLER_24_189 ();
 FILLCELL_X1 FILLER_24_197 ();
 FILLCELL_X1 FILLER_24_205 ();
 FILLCELL_X8 FILLER_24_242 ();
 FILLCELL_X1 FILLER_24_250 ();
 FILLCELL_X4 FILLER_24_271 ();
 FILLCELL_X2 FILLER_24_275 ();
 FILLCELL_X16 FILLER_25_1 ();
 FILLCELL_X8 FILLER_25_17 ();
 FILLCELL_X4 FILLER_25_25 ();
 FILLCELL_X16 FILLER_25_36 ();
 FILLCELL_X8 FILLER_25_52 ();
 FILLCELL_X16 FILLER_25_82 ();
 FILLCELL_X8 FILLER_25_98 ();
 FILLCELL_X2 FILLER_25_106 ();
 FILLCELL_X1 FILLER_25_108 ();
 FILLCELL_X16 FILLER_25_121 ();
 FILLCELL_X8 FILLER_25_137 ();
 FILLCELL_X4 FILLER_25_145 ();
 FILLCELL_X4 FILLER_25_158 ();
 FILLCELL_X2 FILLER_25_162 ();
 FILLCELL_X2 FILLER_25_190 ();
 FILLCELL_X4 FILLER_25_204 ();
 FILLCELL_X2 FILLER_25_242 ();
 FILLCELL_X4 FILLER_25_249 ();
 FILLCELL_X1 FILLER_25_253 ();
 FILLCELL_X2 FILLER_25_274 ();
 FILLCELL_X1 FILLER_25_276 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X2 FILLER_26_33 ();
 FILLCELL_X1 FILLER_26_35 ();
 FILLCELL_X4 FILLER_26_57 ();
 FILLCELL_X1 FILLER_26_61 ();
 FILLCELL_X2 FILLER_26_83 ();
 FILLCELL_X2 FILLER_26_92 ();
 FILLCELL_X4 FILLER_26_101 ();
 FILLCELL_X2 FILLER_26_112 ();
 FILLCELL_X4 FILLER_26_131 ();
 FILLCELL_X8 FILLER_26_149 ();
 FILLCELL_X2 FILLER_26_157 ();
 FILLCELL_X1 FILLER_26_159 ();
 FILLCELL_X8 FILLER_26_174 ();
 FILLCELL_X2 FILLER_26_182 ();
 FILLCELL_X1 FILLER_26_184 ();
 FILLCELL_X2 FILLER_26_192 ();
 FILLCELL_X1 FILLER_26_194 ();
 FILLCELL_X16 FILLER_26_202 ();
 FILLCELL_X2 FILLER_26_218 ();
 FILLCELL_X1 FILLER_26_220 ();
 FILLCELL_X2 FILLER_26_228 ();
 FILLCELL_X4 FILLER_26_237 ();
 FILLCELL_X16 FILLER_26_255 ();
 FILLCELL_X4 FILLER_26_271 ();
 FILLCELL_X2 FILLER_26_275 ();
 FILLCELL_X8 FILLER_27_1 ();
 FILLCELL_X2 FILLER_27_33 ();
 FILLCELL_X8 FILLER_27_69 ();
 FILLCELL_X4 FILLER_27_106 ();
 FILLCELL_X1 FILLER_27_110 ();
 FILLCELL_X8 FILLER_27_118 ();
 FILLCELL_X2 FILLER_27_133 ();
 FILLCELL_X8 FILLER_27_142 ();
 FILLCELL_X1 FILLER_27_150 ();
 FILLCELL_X2 FILLER_27_175 ();
 FILLCELL_X1 FILLER_27_177 ();
 FILLCELL_X4 FILLER_27_209 ();
 FILLCELL_X2 FILLER_27_213 ();
 FILLCELL_X4 FILLER_27_222 ();
 FILLCELL_X16 FILLER_27_233 ();
 FILLCELL_X4 FILLER_27_249 ();
 FILLCELL_X2 FILLER_27_253 ();
 FILLCELL_X8 FILLER_27_262 ();
 FILLCELL_X4 FILLER_27_270 ();
 FILLCELL_X2 FILLER_27_274 ();
 FILLCELL_X1 FILLER_27_276 ();
 FILLCELL_X8 FILLER_28_1 ();
 FILLCELL_X4 FILLER_28_9 ();
 FILLCELL_X1 FILLER_28_13 ();
 FILLCELL_X2 FILLER_28_21 ();
 FILLCELL_X1 FILLER_28_23 ();
 FILLCELL_X2 FILLER_28_31 ();
 FILLCELL_X4 FILLER_28_40 ();
 FILLCELL_X2 FILLER_28_44 ();
 FILLCELL_X8 FILLER_28_60 ();
 FILLCELL_X2 FILLER_28_68 ();
 FILLCELL_X4 FILLER_28_77 ();
 FILLCELL_X1 FILLER_28_81 ();
 FILLCELL_X2 FILLER_28_109 ();
 FILLCELL_X1 FILLER_28_111 ();
 FILLCELL_X4 FILLER_28_117 ();
 FILLCELL_X2 FILLER_28_121 ();
 FILLCELL_X4 FILLER_28_140 ();
 FILLCELL_X2 FILLER_28_200 ();
 FILLCELL_X4 FILLER_28_207 ();
 FILLCELL_X2 FILLER_28_211 ();
 FILLCELL_X4 FILLER_28_237 ();
 FILLCELL_X2 FILLER_28_241 ();
 FILLCELL_X2 FILLER_28_257 ();
 FILLCELL_X1 FILLER_28_259 ();
 FILLCELL_X8 FILLER_29_1 ();
 FILLCELL_X4 FILLER_29_9 ();
 FILLCELL_X2 FILLER_29_13 ();
 FILLCELL_X1 FILLER_29_15 ();
 FILLCELL_X2 FILLER_29_33 ();
 FILLCELL_X1 FILLER_29_35 ();
 FILLCELL_X2 FILLER_29_53 ();
 FILLCELL_X1 FILLER_29_55 ();
 FILLCELL_X16 FILLER_29_73 ();
 FILLCELL_X1 FILLER_29_89 ();
 FILLCELL_X8 FILLER_29_97 ();
 FILLCELL_X1 FILLER_29_105 ();
 FILLCELL_X16 FILLER_29_132 ();
 FILLCELL_X8 FILLER_29_148 ();
 FILLCELL_X4 FILLER_29_156 ();
 FILLCELL_X2 FILLER_29_160 ();
 FILLCELL_X8 FILLER_29_169 ();
 FILLCELL_X1 FILLER_29_177 ();
 FILLCELL_X16 FILLER_29_185 ();
 FILLCELL_X4 FILLER_29_201 ();
 FILLCELL_X2 FILLER_29_205 ();
 FILLCELL_X8 FILLER_29_231 ();
 FILLCELL_X4 FILLER_29_239 ();
 FILLCELL_X16 FILLER_29_260 ();
 FILLCELL_X1 FILLER_29_276 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X4 FILLER_30_65 ();
 FILLCELL_X2 FILLER_30_69 ();
 FILLCELL_X8 FILLER_30_88 ();
 FILLCELL_X1 FILLER_30_96 ();
 FILLCELL_X4 FILLER_30_101 ();
 FILLCELL_X2 FILLER_30_105 ();
 FILLCELL_X1 FILLER_30_107 ();
 FILLCELL_X16 FILLER_30_125 ();
 FILLCELL_X4 FILLER_30_165 ();
 FILLCELL_X1 FILLER_30_169 ();
 FILLCELL_X1 FILLER_30_177 ();
 FILLCELL_X32 FILLER_30_185 ();
 FILLCELL_X16 FILLER_30_217 ();
 FILLCELL_X8 FILLER_30_233 ();
 FILLCELL_X2 FILLER_30_241 ();
 FILLCELL_X16 FILLER_30_257 ();
 FILLCELL_X4 FILLER_30_273 ();
 FILLCELL_X16 FILLER_31_1 ();
 FILLCELL_X8 FILLER_31_17 ();
 FILLCELL_X1 FILLER_31_25 ();
 FILLCELL_X16 FILLER_31_50 ();
 FILLCELL_X4 FILLER_31_66 ();
 FILLCELL_X2 FILLER_31_70 ();
 FILLCELL_X1 FILLER_31_72 ();
 FILLCELL_X8 FILLER_31_87 ();
 FILLCELL_X4 FILLER_31_95 ();
 FILLCELL_X1 FILLER_31_99 ();
 FILLCELL_X2 FILLER_31_107 ();
 FILLCELL_X4 FILLER_31_126 ();
 FILLCELL_X2 FILLER_31_130 ();
 FILLCELL_X1 FILLER_31_132 ();
 FILLCELL_X4 FILLER_31_164 ();
 FILLCELL_X1 FILLER_31_168 ();
 FILLCELL_X32 FILLER_31_186 ();
 FILLCELL_X1 FILLER_31_218 ();
 FILLCELL_X1 FILLER_31_233 ();
 FILLCELL_X16 FILLER_31_258 ();
 FILLCELL_X2 FILLER_31_274 ();
 FILLCELL_X1 FILLER_31_276 ();
 FILLCELL_X16 FILLER_32_1 ();
 FILLCELL_X4 FILLER_32_17 ();
 FILLCELL_X2 FILLER_32_21 ();
 FILLCELL_X4 FILLER_32_54 ();
 FILLCELL_X2 FILLER_32_58 ();
 FILLCELL_X1 FILLER_32_60 ();
 FILLCELL_X2 FILLER_32_65 ();
 FILLCELL_X4 FILLER_32_74 ();
 FILLCELL_X1 FILLER_32_78 ();
 FILLCELL_X1 FILLER_32_86 ();
 FILLCELL_X8 FILLER_32_101 ();
 FILLCELL_X2 FILLER_32_109 ();
 FILLCELL_X8 FILLER_32_118 ();
 FILLCELL_X16 FILLER_32_130 ();
 FILLCELL_X8 FILLER_32_146 ();
 FILLCELL_X4 FILLER_32_154 ();
 FILLCELL_X2 FILLER_32_158 ();
 FILLCELL_X4 FILLER_32_167 ();
 FILLCELL_X16 FILLER_32_202 ();
 FILLCELL_X4 FILLER_32_270 ();
 FILLCELL_X2 FILLER_32_274 ();
 FILLCELL_X1 FILLER_32_276 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X16 FILLER_33_33 ();
 FILLCELL_X4 FILLER_33_49 ();
 FILLCELL_X2 FILLER_33_53 ();
 FILLCELL_X1 FILLER_33_55 ();
 FILLCELL_X2 FILLER_33_63 ();
 FILLCELL_X1 FILLER_33_65 ();
 FILLCELL_X16 FILLER_33_100 ();
 FILLCELL_X1 FILLER_33_116 ();
 FILLCELL_X8 FILLER_33_124 ();
 FILLCELL_X1 FILLER_33_132 ();
 FILLCELL_X1 FILLER_33_153 ();
 FILLCELL_X4 FILLER_33_178 ();
 FILLCELL_X2 FILLER_33_182 ();
 FILLCELL_X1 FILLER_33_184 ();
 FILLCELL_X4 FILLER_33_199 ();
 FILLCELL_X2 FILLER_33_203 ();
 FILLCELL_X1 FILLER_33_212 ();
 FILLCELL_X8 FILLER_33_237 ();
 FILLCELL_X2 FILLER_33_245 ();
 FILLCELL_X1 FILLER_33_247 ();
 FILLCELL_X8 FILLER_33_262 ();
 FILLCELL_X4 FILLER_33_270 ();
 FILLCELL_X2 FILLER_33_274 ();
 FILLCELL_X1 FILLER_33_276 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X16 FILLER_34_33 ();
 FILLCELL_X8 FILLER_34_49 ();
 FILLCELL_X2 FILLER_34_57 ();
 FILLCELL_X1 FILLER_34_59 ();
 FILLCELL_X4 FILLER_34_84 ();
 FILLCELL_X2 FILLER_34_88 ();
 FILLCELL_X16 FILLER_34_97 ();
 FILLCELL_X4 FILLER_34_130 ();
 FILLCELL_X1 FILLER_34_134 ();
 FILLCELL_X2 FILLER_34_142 ();
 FILLCELL_X4 FILLER_34_161 ();
 FILLCELL_X2 FILLER_34_182 ();
 FILLCELL_X4 FILLER_34_201 ();
 FILLCELL_X2 FILLER_34_229 ();
 FILLCELL_X4 FILLER_34_251 ();
 FILLCELL_X2 FILLER_34_255 ();
 FILLCELL_X2 FILLER_34_274 ();
 FILLCELL_X1 FILLER_34_276 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X4 FILLER_35_65 ();
 FILLCELL_X1 FILLER_35_69 ();
 FILLCELL_X4 FILLER_35_77 ();
 FILLCELL_X2 FILLER_35_81 ();
 FILLCELL_X8 FILLER_35_100 ();
 FILLCELL_X2 FILLER_35_108 ();
 FILLCELL_X1 FILLER_35_110 ();
 FILLCELL_X4 FILLER_35_118 ();
 FILLCELL_X1 FILLER_35_122 ();
 FILLCELL_X8 FILLER_35_130 ();
 FILLCELL_X1 FILLER_35_138 ();
 FILLCELL_X8 FILLER_35_156 ();
 FILLCELL_X1 FILLER_35_164 ();
 FILLCELL_X4 FILLER_35_172 ();
 FILLCELL_X1 FILLER_35_176 ();
 FILLCELL_X4 FILLER_35_201 ();
 FILLCELL_X2 FILLER_35_205 ();
 FILLCELL_X16 FILLER_35_231 ();
 FILLCELL_X8 FILLER_35_264 ();
 FILLCELL_X4 FILLER_35_272 ();
 FILLCELL_X1 FILLER_35_276 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X2 FILLER_36_33 ();
 FILLCELL_X16 FILLER_36_39 ();
 FILLCELL_X8 FILLER_36_55 ();
 FILLCELL_X2 FILLER_36_63 ();
 FILLCELL_X16 FILLER_36_86 ();
 FILLCELL_X4 FILLER_36_102 ();
 FILLCELL_X2 FILLER_36_106 ();
 FILLCELL_X1 FILLER_36_108 ();
 FILLCELL_X32 FILLER_36_130 ();
 FILLCELL_X32 FILLER_36_162 ();
 FILLCELL_X32 FILLER_36_194 ();
 FILLCELL_X2 FILLER_36_226 ();
 FILLCELL_X1 FILLER_36_228 ();
 FILLCELL_X32 FILLER_36_232 ();
 FILLCELL_X8 FILLER_36_264 ();
 FILLCELL_X4 FILLER_36_272 ();
 FILLCELL_X1 FILLER_36_276 ();
endmodule
