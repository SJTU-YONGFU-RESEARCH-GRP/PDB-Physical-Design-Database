module showahead_fifo (almost_empty,
    almost_full,
    clk,
    empty,
    full,
    peek_en,
    rd_en,
    rst_n,
    valid,
    wr_en,
    data_count,
    rd_data,
    wr_data);
 output almost_empty;
 output almost_full;
 input clk;
 output empty;
 output full;
 input peek_en;
 input rd_en;
 input rst_n;
 output valid;
 input wr_en;
 output [4:0] data_count;
 output [7:0] rd_data;
 input [7:0] wr_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire _433_;
 wire _434_;
 wire _435_;
 wire _436_;
 wire _437_;
 wire _438_;
 wire _439_;
 wire _440_;
 wire _441_;
 wire _442_;
 wire _443_;
 wire _444_;
 wire _445_;
 wire _446_;
 wire _447_;
 wire _448_;
 wire _449_;
 wire _450_;
 wire _451_;
 wire _452_;
 wire _453_;
 wire _454_;
 wire _455_;
 wire _456_;
 wire _457_;
 wire _458_;
 wire _459_;
 wire _460_;
 wire _461_;
 wire _462_;
 wire _463_;
 wire _464_;
 wire _465_;
 wire _466_;
 wire _467_;
 wire _468_;
 wire _469_;
 wire _470_;
 wire _471_;
 wire _472_;
 wire _473_;
 wire _474_;
 wire _475_;
 wire _476_;
 wire _477_;
 wire _478_;
 wire _479_;
 wire _480_;
 wire _481_;
 wire _482_;
 wire _483_;
 wire _484_;
 wire _485_;
 wire _486_;
 wire _487_;
 wire _488_;
 wire _489_;
 wire _490_;
 wire _491_;
 wire _492_;
 wire _493_;
 wire _494_;
 wire _495_;
 wire _496_;
 wire _497_;
 wire _498_;
 wire _499_;
 wire _500_;
 wire _501_;
 wire _502_;
 wire _503_;
 wire _504_;
 wire _505_;
 wire _506_;
 wire _507_;
 wire _508_;
 wire _509_;
 wire _510_;
 wire _511_;
 wire _512_;
 wire _513_;
 wire _514_;
 wire _515_;
 wire _516_;
 wire _517_;
 wire _518_;
 wire _519_;
 wire _520_;
 wire _521_;
 wire _522_;
 wire _523_;
 wire _524_;
 wire _525_;
 wire _526_;
 wire _527_;
 wire _528_;
 wire _529_;
 wire _530_;
 wire _531_;
 wire _532_;
 wire _533_;
 wire _534_;
 wire _535_;
 wire _536_;
 wire _537_;
 wire _538_;
 wire _539_;
 wire _540_;
 wire _541_;
 wire _542_;
 wire _543_;
 wire _544_;
 wire _545_;
 wire _546_;
 wire _547_;
 wire _548_;
 wire _549_;
 wire _550_;
 wire _551_;
 wire _552_;
 wire _553_;
 wire _554_;
 wire _555_;
 wire _556_;
 wire _557_;
 wire \mem[0][0] ;
 wire \mem[0][1] ;
 wire \mem[0][2] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[10][0] ;
 wire \mem[10][1] ;
 wire \mem[10][2] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[11][0] ;
 wire \mem[11][1] ;
 wire \mem[11][2] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[12][0] ;
 wire \mem[12][1] ;
 wire \mem[12][2] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[13][0] ;
 wire \mem[13][1] ;
 wire \mem[13][2] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[14][0] ;
 wire \mem[14][1] ;
 wire \mem[14][2] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[15][0] ;
 wire \mem[15][1] ;
 wire \mem[15][2] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[1][0] ;
 wire \mem[1][1] ;
 wire \mem[1][2] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[2][0] ;
 wire \mem[2][1] ;
 wire \mem[2][2] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[3][0] ;
 wire \mem[3][1] ;
 wire \mem[3][2] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[4][0] ;
 wire \mem[4][1] ;
 wire \mem[4][2] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[5][0] ;
 wire \mem[5][1] ;
 wire \mem[5][2] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[6][0] ;
 wire \mem[6][1] ;
 wire \mem[6][2] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[7][0] ;
 wire \mem[7][1] ;
 wire \mem[7][2] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[8][0] ;
 wire \mem[8][1] ;
 wire \mem[8][2] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[9][0] ;
 wire \mem[9][1] ;
 wire \mem[9][2] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \rd_ptr[0] ;
 wire \rd_ptr[1] ;
 wire \rd_ptr[2] ;
 wire \rd_ptr[3] ;
 wire \rd_ptr[4] ;
 wire \wr_ptr[0] ;
 wire \wr_ptr[1] ;
 wire \wr_ptr[2] ;
 wire \wr_ptr[3] ;
 wire \wr_ptr[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 CLKBUF_X2 _558_ (.A(_557_),
    .Z(_275_));
 INV_X2 _559_ (.A(_275_),
    .ZN(net5));
 BUF_X4 _560_ (.A(_541_),
    .Z(_276_));
 AND2_X1 _561_ (.A1(_546_),
    .A2(_543_),
    .ZN(_277_));
 INV_X1 _562_ (.A(_556_),
    .ZN(_537_));
 AOI221_X2 _563_ (.A(_545_),
    .B1(_277_),
    .B2(_537_),
    .C1(_542_),
    .C2(_546_),
    .ZN(_278_));
 XNOR2_X2 _564_ (.A(_276_),
    .B(_278_),
    .ZN(net8));
 XNOR2_X2 _565_ (.A(_546_),
    .B(_538_),
    .ZN(_279_));
 INV_X4 _566_ (.A(_279_),
    .ZN(net7));
 AND2_X1 _567_ (.A1(_276_),
    .A2(_546_),
    .ZN(_280_));
 AOI221_X2 _568_ (.A(_540_),
    .B1(_545_),
    .B2(_276_),
    .C1(_280_),
    .C2(_538_),
    .ZN(_281_));
 XNOR2_X1 _569_ (.A(\wr_ptr[4] ),
    .B(\rd_ptr[4] ),
    .ZN(_282_));
 XOR2_X2 _570_ (.A(_281_),
    .B(_282_),
    .Z(_283_));
 BUF_X8 _571_ (.A(_283_),
    .Z(_284_));
 INV_X8 _572_ (.A(_284_),
    .ZN(net9));
 BUF_X8 _573_ (.A(_283_),
    .Z(_285_));
 BUF_X2 _574_ (.A(net6),
    .Z(_286_));
 INV_X1 _575_ (.A(_286_),
    .ZN(_287_));
 NAND4_X1 _576_ (.A1(_276_),
    .A2(_275_),
    .A3(_287_),
    .A4(_279_),
    .ZN(_288_));
 INV_X1 _577_ (.A(_276_),
    .ZN(_289_));
 NAND4_X1 _578_ (.A1(_289_),
    .A2(_275_),
    .A3(_287_),
    .A4(_279_),
    .ZN(_290_));
 MUX2_X1 _579_ (.A(_288_),
    .B(_290_),
    .S(_278_),
    .Z(_291_));
 BUF_X8 _580_ (.A(_291_),
    .Z(_292_));
 BUF_X16 _581_ (.A(_292_),
    .Z(_293_));
 NOR2_X4 _582_ (.A1(_285_),
    .A2(_293_),
    .ZN(net11));
 NOR2_X4 _583_ (.A1(net9),
    .A2(_293_),
    .ZN(net10));
 BUF_X2 _584_ (.A(wr_data[0]),
    .Z(_294_));
 BUF_X2 _585_ (.A(_294_),
    .Z(_295_));
 INV_X2 _586_ (.A(\wr_ptr[3] ),
    .ZN(_296_));
 INV_X2 _587_ (.A(\wr_ptr[2] ),
    .ZN(_297_));
 NAND2_X2 _588_ (.A1(_296_),
    .A2(_297_),
    .ZN(_298_));
 CLKBUF_X3 _589_ (.A(wr_en),
    .Z(_299_));
 NAND2_X1 _590_ (.A1(_299_),
    .A2(_549_),
    .ZN(_300_));
 NOR2_X1 _591_ (.A1(_298_),
    .A2(_300_),
    .ZN(_301_));
 OAI21_X4 _592_ (.A(_301_),
    .B1(_293_),
    .B2(_285_),
    .ZN(_302_));
 MUX2_X1 _593_ (.A(_295_),
    .B(\mem[0][0] ),
    .S(_302_),
    .Z(_140_));
 CLKBUF_X2 _594_ (.A(wr_data[1]),
    .Z(_303_));
 BUF_X2 _595_ (.A(_303_),
    .Z(_304_));
 MUX2_X1 _596_ (.A(_304_),
    .B(\mem[0][1] ),
    .S(_302_),
    .Z(_141_));
 BUF_X2 _597_ (.A(wr_data[2]),
    .Z(_305_));
 BUF_X2 _598_ (.A(_305_),
    .Z(_306_));
 MUX2_X1 _599_ (.A(_306_),
    .B(\mem[0][2] ),
    .S(_302_),
    .Z(_142_));
 CLKBUF_X2 _600_ (.A(wr_data[3]),
    .Z(_307_));
 BUF_X2 _601_ (.A(_307_),
    .Z(_308_));
 MUX2_X1 _602_ (.A(_308_),
    .B(\mem[0][3] ),
    .S(_302_),
    .Z(_143_));
 CLKBUF_X2 _603_ (.A(wr_data[4]),
    .Z(_309_));
 BUF_X2 _604_ (.A(_309_),
    .Z(_310_));
 MUX2_X1 _605_ (.A(_310_),
    .B(\mem[0][4] ),
    .S(_302_),
    .Z(_144_));
 CLKBUF_X2 _606_ (.A(wr_data[5]),
    .Z(_311_));
 BUF_X2 _607_ (.A(_311_),
    .Z(_312_));
 MUX2_X1 _608_ (.A(_312_),
    .B(\mem[0][5] ),
    .S(_302_),
    .Z(_145_));
 CLKBUF_X2 _609_ (.A(wr_data[6]),
    .Z(_313_));
 BUF_X2 _610_ (.A(_313_),
    .Z(_314_));
 MUX2_X1 _611_ (.A(_314_),
    .B(\mem[0][6] ),
    .S(_302_),
    .Z(_146_));
 CLKBUF_X2 _612_ (.A(wr_data[7]),
    .Z(_315_));
 BUF_X2 _613_ (.A(_315_),
    .Z(_316_));
 MUX2_X1 _614_ (.A(_316_),
    .B(\mem[0][7] ),
    .S(_302_),
    .Z(_147_));
 NAND2_X2 _615_ (.A1(\wr_ptr[3] ),
    .A2(_297_),
    .ZN(_317_));
 NAND2_X1 _616_ (.A1(_299_),
    .A2(_550_),
    .ZN(_318_));
 NOR2_X1 _617_ (.A1(_317_),
    .A2(_318_),
    .ZN(_319_));
 OAI21_X4 _618_ (.A(_319_),
    .B1(_293_),
    .B2(_285_),
    .ZN(_320_));
 MUX2_X1 _619_ (.A(_295_),
    .B(\mem[10][0] ),
    .S(_320_),
    .Z(_148_));
 MUX2_X1 _620_ (.A(_304_),
    .B(\mem[10][1] ),
    .S(_320_),
    .Z(_149_));
 MUX2_X1 _621_ (.A(_306_),
    .B(\mem[10][2] ),
    .S(_320_),
    .Z(_150_));
 MUX2_X1 _622_ (.A(_308_),
    .B(\mem[10][3] ),
    .S(_320_),
    .Z(_151_));
 MUX2_X1 _623_ (.A(_310_),
    .B(\mem[10][4] ),
    .S(_320_),
    .Z(_152_));
 MUX2_X1 _624_ (.A(_312_),
    .B(\mem[10][5] ),
    .S(_320_),
    .Z(_153_));
 MUX2_X1 _625_ (.A(_314_),
    .B(\mem[10][6] ),
    .S(_320_),
    .Z(_154_));
 MUX2_X1 _626_ (.A(_316_),
    .B(\mem[10][7] ),
    .S(_320_),
    .Z(_155_));
 NAND2_X1 _627_ (.A1(_299_),
    .A2(_554_),
    .ZN(_321_));
 NOR2_X1 _628_ (.A1(_317_),
    .A2(_321_),
    .ZN(_322_));
 OAI21_X4 _629_ (.A(_322_),
    .B1(_293_),
    .B2(_285_),
    .ZN(_323_));
 MUX2_X1 _630_ (.A(_295_),
    .B(\mem[11][0] ),
    .S(_323_),
    .Z(_156_));
 MUX2_X1 _631_ (.A(_304_),
    .B(\mem[11][1] ),
    .S(_323_),
    .Z(_157_));
 MUX2_X1 _632_ (.A(_306_),
    .B(\mem[11][2] ),
    .S(_323_),
    .Z(_158_));
 MUX2_X1 _633_ (.A(_308_),
    .B(\mem[11][3] ),
    .S(_323_),
    .Z(_159_));
 MUX2_X1 _634_ (.A(_310_),
    .B(\mem[11][4] ),
    .S(_323_),
    .Z(_160_));
 MUX2_X1 _635_ (.A(_312_),
    .B(\mem[11][5] ),
    .S(_323_),
    .Z(_161_));
 MUX2_X1 _636_ (.A(_314_),
    .B(\mem[11][6] ),
    .S(_323_),
    .Z(_162_));
 MUX2_X1 _637_ (.A(_316_),
    .B(\mem[11][7] ),
    .S(_323_),
    .Z(_163_));
 NOR2_X2 _638_ (.A1(_296_),
    .A2(_297_),
    .ZN(_324_));
 NAND3_X1 _639_ (.A1(_299_),
    .A2(_549_),
    .A3(_324_),
    .ZN(_325_));
 NOR4_X1 _640_ (.A1(_289_),
    .A2(net5),
    .A3(_286_),
    .A4(net7),
    .ZN(_326_));
 NOR4_X1 _641_ (.A1(_276_),
    .A2(net5),
    .A3(_286_),
    .A4(net7),
    .ZN(_327_));
 MUX2_X1 _642_ (.A(_326_),
    .B(_327_),
    .S(_278_),
    .Z(_328_));
 BUF_X8 _643_ (.A(_328_),
    .Z(_329_));
 AOI21_X4 _644_ (.A(_325_),
    .B1(_329_),
    .B2(net9),
    .ZN(_330_));
 MUX2_X1 _645_ (.A(\mem[12][0] ),
    .B(_295_),
    .S(_330_),
    .Z(_164_));
 MUX2_X1 _646_ (.A(\mem[12][1] ),
    .B(_304_),
    .S(_330_),
    .Z(_165_));
 MUX2_X1 _647_ (.A(\mem[12][2] ),
    .B(_306_),
    .S(_330_),
    .Z(_166_));
 MUX2_X1 _648_ (.A(\mem[12][3] ),
    .B(_308_),
    .S(_330_),
    .Z(_167_));
 MUX2_X1 _649_ (.A(\mem[12][4] ),
    .B(_310_),
    .S(_330_),
    .Z(_168_));
 MUX2_X1 _650_ (.A(\mem[12][5] ),
    .B(_312_),
    .S(_330_),
    .Z(_169_));
 MUX2_X1 _651_ (.A(\mem[12][6] ),
    .B(_314_),
    .S(_330_),
    .Z(_170_));
 MUX2_X1 _652_ (.A(\mem[12][7] ),
    .B(_316_),
    .S(_330_),
    .Z(_171_));
 NAND3_X1 _653_ (.A1(_299_),
    .A2(_552_),
    .A3(_324_),
    .ZN(_331_));
 AOI21_X4 _654_ (.A(_331_),
    .B1(_329_),
    .B2(net9),
    .ZN(_332_));
 MUX2_X1 _655_ (.A(\mem[13][0] ),
    .B(_295_),
    .S(_332_),
    .Z(_172_));
 MUX2_X1 _656_ (.A(\mem[13][1] ),
    .B(_304_),
    .S(_332_),
    .Z(_173_));
 MUX2_X1 _657_ (.A(\mem[13][2] ),
    .B(_306_),
    .S(_332_),
    .Z(_174_));
 MUX2_X1 _658_ (.A(\mem[13][3] ),
    .B(_308_),
    .S(_332_),
    .Z(_175_));
 MUX2_X1 _659_ (.A(\mem[13][4] ),
    .B(_310_),
    .S(_332_),
    .Z(_176_));
 MUX2_X1 _660_ (.A(\mem[13][5] ),
    .B(_312_),
    .S(_332_),
    .Z(_177_));
 MUX2_X1 _661_ (.A(\mem[13][6] ),
    .B(_314_),
    .S(_332_),
    .Z(_178_));
 MUX2_X1 _662_ (.A(\mem[13][7] ),
    .B(_316_),
    .S(_332_),
    .Z(_179_));
 NAND3_X2 _663_ (.A1(_299_),
    .A2(_550_),
    .A3(_324_),
    .ZN(_333_));
 AOI21_X4 _664_ (.A(_333_),
    .B1(_329_),
    .B2(net9),
    .ZN(_334_));
 MUX2_X1 _665_ (.A(\mem[14][0] ),
    .B(_295_),
    .S(_334_),
    .Z(_180_));
 MUX2_X1 _666_ (.A(\mem[14][1] ),
    .B(_304_),
    .S(_334_),
    .Z(_181_));
 MUX2_X1 _667_ (.A(\mem[14][2] ),
    .B(_306_),
    .S(_334_),
    .Z(_182_));
 MUX2_X1 _668_ (.A(\mem[14][3] ),
    .B(_308_),
    .S(_334_),
    .Z(_183_));
 MUX2_X1 _669_ (.A(\mem[14][4] ),
    .B(_310_),
    .S(_334_),
    .Z(_184_));
 MUX2_X1 _670_ (.A(\mem[14][5] ),
    .B(_312_),
    .S(_334_),
    .Z(_185_));
 MUX2_X1 _671_ (.A(\mem[14][6] ),
    .B(_314_),
    .S(_334_),
    .Z(_186_));
 MUX2_X1 _672_ (.A(\mem[14][7] ),
    .B(_316_),
    .S(_334_),
    .Z(_187_));
 NAND3_X2 _673_ (.A1(_299_),
    .A2(_554_),
    .A3(_324_),
    .ZN(_335_));
 AOI21_X4 _674_ (.A(_335_),
    .B1(_329_),
    .B2(net9),
    .ZN(_336_));
 MUX2_X1 _675_ (.A(\mem[15][0] ),
    .B(_295_),
    .S(_336_),
    .Z(_188_));
 MUX2_X1 _676_ (.A(\mem[15][1] ),
    .B(_304_),
    .S(_336_),
    .Z(_189_));
 MUX2_X1 _677_ (.A(\mem[15][2] ),
    .B(_306_),
    .S(_336_),
    .Z(_190_));
 MUX2_X1 _678_ (.A(\mem[15][3] ),
    .B(_308_),
    .S(_336_),
    .Z(_191_));
 MUX2_X1 _679_ (.A(\mem[15][4] ),
    .B(_310_),
    .S(_336_),
    .Z(_192_));
 MUX2_X1 _680_ (.A(\mem[15][5] ),
    .B(_312_),
    .S(_336_),
    .Z(_193_));
 MUX2_X1 _681_ (.A(\mem[15][6] ),
    .B(_314_),
    .S(_336_),
    .Z(_194_));
 MUX2_X1 _682_ (.A(\mem[15][7] ),
    .B(_316_),
    .S(_336_),
    .Z(_195_));
 NAND2_X1 _683_ (.A1(_299_),
    .A2(_552_),
    .ZN(_337_));
 NOR2_X1 _684_ (.A1(_298_),
    .A2(_337_),
    .ZN(_338_));
 OAI21_X4 _685_ (.A(_338_),
    .B1(_293_),
    .B2(_284_),
    .ZN(_339_));
 MUX2_X1 _686_ (.A(_295_),
    .B(\mem[1][0] ),
    .S(_339_),
    .Z(_196_));
 MUX2_X1 _687_ (.A(_304_),
    .B(\mem[1][1] ),
    .S(_339_),
    .Z(_197_));
 MUX2_X1 _688_ (.A(_306_),
    .B(\mem[1][2] ),
    .S(_339_),
    .Z(_198_));
 MUX2_X1 _689_ (.A(_308_),
    .B(\mem[1][3] ),
    .S(_339_),
    .Z(_199_));
 MUX2_X1 _690_ (.A(_310_),
    .B(\mem[1][4] ),
    .S(_339_),
    .Z(_200_));
 MUX2_X1 _691_ (.A(_312_),
    .B(\mem[1][5] ),
    .S(_339_),
    .Z(_201_));
 MUX2_X1 _692_ (.A(_314_),
    .B(\mem[1][6] ),
    .S(_339_),
    .Z(_202_));
 MUX2_X1 _693_ (.A(_316_),
    .B(\mem[1][7] ),
    .S(_339_),
    .Z(_203_));
 NOR2_X1 _694_ (.A1(_298_),
    .A2(_318_),
    .ZN(_340_));
 OAI21_X4 _695_ (.A(_340_),
    .B1(_293_),
    .B2(_284_),
    .ZN(_341_));
 MUX2_X1 _696_ (.A(_295_),
    .B(\mem[2][0] ),
    .S(_341_),
    .Z(_204_));
 MUX2_X1 _697_ (.A(_304_),
    .B(\mem[2][1] ),
    .S(_341_),
    .Z(_205_));
 MUX2_X1 _698_ (.A(_306_),
    .B(\mem[2][2] ),
    .S(_341_),
    .Z(_206_));
 MUX2_X1 _699_ (.A(_308_),
    .B(\mem[2][3] ),
    .S(_341_),
    .Z(_207_));
 MUX2_X1 _700_ (.A(_310_),
    .B(\mem[2][4] ),
    .S(_341_),
    .Z(_208_));
 MUX2_X1 _701_ (.A(_312_),
    .B(\mem[2][5] ),
    .S(_341_),
    .Z(_209_));
 MUX2_X1 _702_ (.A(_314_),
    .B(\mem[2][6] ),
    .S(_341_),
    .Z(_210_));
 MUX2_X1 _703_ (.A(_316_),
    .B(\mem[2][7] ),
    .S(_341_),
    .Z(_211_));
 NOR2_X1 _704_ (.A1(_298_),
    .A2(_321_),
    .ZN(_342_));
 OAI21_X4 _705_ (.A(_342_),
    .B1(_293_),
    .B2(_284_),
    .ZN(_343_));
 MUX2_X1 _706_ (.A(_295_),
    .B(\mem[3][0] ),
    .S(_343_),
    .Z(_212_));
 MUX2_X1 _707_ (.A(_304_),
    .B(\mem[3][1] ),
    .S(_343_),
    .Z(_213_));
 MUX2_X1 _708_ (.A(_306_),
    .B(\mem[3][2] ),
    .S(_343_),
    .Z(_214_));
 MUX2_X1 _709_ (.A(_308_),
    .B(\mem[3][3] ),
    .S(_343_),
    .Z(_215_));
 MUX2_X1 _710_ (.A(_310_),
    .B(\mem[3][4] ),
    .S(_343_),
    .Z(_216_));
 MUX2_X1 _711_ (.A(_312_),
    .B(\mem[3][5] ),
    .S(_343_),
    .Z(_217_));
 MUX2_X1 _712_ (.A(_314_),
    .B(\mem[3][6] ),
    .S(_343_),
    .Z(_218_));
 MUX2_X1 _713_ (.A(_316_),
    .B(\mem[3][7] ),
    .S(_343_),
    .Z(_219_));
 NAND2_X2 _714_ (.A1(_296_),
    .A2(\wr_ptr[2] ),
    .ZN(_344_));
 NOR2_X1 _715_ (.A1(_300_),
    .A2(_344_),
    .ZN(_345_));
 OAI21_X4 _716_ (.A(_345_),
    .B1(_293_),
    .B2(_284_),
    .ZN(_346_));
 MUX2_X1 _717_ (.A(_294_),
    .B(\mem[4][0] ),
    .S(_346_),
    .Z(_220_));
 MUX2_X1 _718_ (.A(_303_),
    .B(\mem[4][1] ),
    .S(_346_),
    .Z(_221_));
 MUX2_X1 _719_ (.A(_305_),
    .B(\mem[4][2] ),
    .S(_346_),
    .Z(_222_));
 MUX2_X1 _720_ (.A(_307_),
    .B(\mem[4][3] ),
    .S(_346_),
    .Z(_223_));
 MUX2_X1 _721_ (.A(_309_),
    .B(\mem[4][4] ),
    .S(_346_),
    .Z(_224_));
 MUX2_X1 _722_ (.A(_311_),
    .B(\mem[4][5] ),
    .S(_346_),
    .Z(_225_));
 MUX2_X1 _723_ (.A(_313_),
    .B(\mem[4][6] ),
    .S(_346_),
    .Z(_226_));
 MUX2_X1 _724_ (.A(_315_),
    .B(\mem[4][7] ),
    .S(_346_),
    .Z(_227_));
 NOR2_X1 _725_ (.A1(_337_),
    .A2(_344_),
    .ZN(_347_));
 OAI21_X4 _726_ (.A(_347_),
    .B1(_292_),
    .B2(_284_),
    .ZN(_348_));
 MUX2_X1 _727_ (.A(_294_),
    .B(\mem[5][0] ),
    .S(_348_),
    .Z(_228_));
 MUX2_X1 _728_ (.A(_303_),
    .B(\mem[5][1] ),
    .S(_348_),
    .Z(_229_));
 MUX2_X1 _729_ (.A(_305_),
    .B(\mem[5][2] ),
    .S(_348_),
    .Z(_230_));
 MUX2_X1 _730_ (.A(_307_),
    .B(\mem[5][3] ),
    .S(_348_),
    .Z(_231_));
 MUX2_X1 _731_ (.A(_309_),
    .B(\mem[5][4] ),
    .S(_348_),
    .Z(_232_));
 MUX2_X1 _732_ (.A(_311_),
    .B(\mem[5][5] ),
    .S(_348_),
    .Z(_233_));
 MUX2_X1 _733_ (.A(_313_),
    .B(\mem[5][6] ),
    .S(_348_),
    .Z(_234_));
 MUX2_X1 _734_ (.A(_315_),
    .B(\mem[5][7] ),
    .S(_348_),
    .Z(_235_));
 NOR2_X1 _735_ (.A1(_318_),
    .A2(_344_),
    .ZN(_349_));
 OAI21_X4 _736_ (.A(_349_),
    .B1(_292_),
    .B2(_284_),
    .ZN(_350_));
 MUX2_X1 _737_ (.A(_294_),
    .B(\mem[6][0] ),
    .S(_350_),
    .Z(_236_));
 MUX2_X1 _738_ (.A(_303_),
    .B(\mem[6][1] ),
    .S(_350_),
    .Z(_237_));
 MUX2_X1 _739_ (.A(_305_),
    .B(\mem[6][2] ),
    .S(_350_),
    .Z(_238_));
 MUX2_X1 _740_ (.A(_307_),
    .B(\mem[6][3] ),
    .S(_350_),
    .Z(_239_));
 MUX2_X1 _741_ (.A(_309_),
    .B(\mem[6][4] ),
    .S(_350_),
    .Z(_240_));
 MUX2_X1 _742_ (.A(_311_),
    .B(\mem[6][5] ),
    .S(_350_),
    .Z(_241_));
 MUX2_X1 _743_ (.A(_313_),
    .B(\mem[6][6] ),
    .S(_350_),
    .Z(_242_));
 MUX2_X1 _744_ (.A(_315_),
    .B(\mem[6][7] ),
    .S(_350_),
    .Z(_243_));
 NOR2_X1 _745_ (.A1(_321_),
    .A2(_344_),
    .ZN(_351_));
 OAI21_X4 _746_ (.A(_351_),
    .B1(_292_),
    .B2(_284_),
    .ZN(_352_));
 MUX2_X1 _747_ (.A(_294_),
    .B(\mem[7][0] ),
    .S(_352_),
    .Z(_244_));
 MUX2_X1 _748_ (.A(_303_),
    .B(\mem[7][1] ),
    .S(_352_),
    .Z(_245_));
 MUX2_X1 _749_ (.A(_305_),
    .B(\mem[7][2] ),
    .S(_352_),
    .Z(_246_));
 MUX2_X1 _750_ (.A(_307_),
    .B(\mem[7][3] ),
    .S(_352_),
    .Z(_247_));
 MUX2_X1 _751_ (.A(_309_),
    .B(\mem[7][4] ),
    .S(_352_),
    .Z(_248_));
 MUX2_X1 _752_ (.A(_311_),
    .B(\mem[7][5] ),
    .S(_352_),
    .Z(_249_));
 MUX2_X1 _753_ (.A(_313_),
    .B(\mem[7][6] ),
    .S(_352_),
    .Z(_250_));
 MUX2_X1 _754_ (.A(_315_),
    .B(\mem[7][7] ),
    .S(_352_),
    .Z(_251_));
 NOR2_X1 _755_ (.A1(_300_),
    .A2(_317_),
    .ZN(_353_));
 OAI21_X4 _756_ (.A(_353_),
    .B1(_292_),
    .B2(_284_),
    .ZN(_354_));
 MUX2_X1 _757_ (.A(_294_),
    .B(\mem[8][0] ),
    .S(_354_),
    .Z(_252_));
 MUX2_X1 _758_ (.A(_303_),
    .B(\mem[8][1] ),
    .S(_354_),
    .Z(_253_));
 MUX2_X1 _759_ (.A(_305_),
    .B(\mem[8][2] ),
    .S(_354_),
    .Z(_254_));
 MUX2_X1 _760_ (.A(_307_),
    .B(\mem[8][3] ),
    .S(_354_),
    .Z(_255_));
 MUX2_X1 _761_ (.A(_309_),
    .B(\mem[8][4] ),
    .S(_354_),
    .Z(_256_));
 MUX2_X1 _762_ (.A(_311_),
    .B(\mem[8][5] ),
    .S(_354_),
    .Z(_257_));
 MUX2_X1 _763_ (.A(_313_),
    .B(\mem[8][6] ),
    .S(_354_),
    .Z(_258_));
 MUX2_X1 _764_ (.A(_315_),
    .B(\mem[8][7] ),
    .S(_354_),
    .Z(_259_));
 NOR2_X1 _765_ (.A1(_317_),
    .A2(_337_),
    .ZN(_355_));
 OAI21_X4 _766_ (.A(_355_),
    .B1(_292_),
    .B2(_284_),
    .ZN(_356_));
 MUX2_X1 _767_ (.A(_294_),
    .B(\mem[9][0] ),
    .S(_356_),
    .Z(_260_));
 MUX2_X1 _768_ (.A(_303_),
    .B(\mem[9][1] ),
    .S(_356_),
    .Z(_261_));
 MUX2_X1 _769_ (.A(_305_),
    .B(\mem[9][2] ),
    .S(_356_),
    .Z(_262_));
 MUX2_X1 _770_ (.A(_307_),
    .B(\mem[9][3] ),
    .S(_356_),
    .Z(_263_));
 MUX2_X1 _771_ (.A(_309_),
    .B(\mem[9][4] ),
    .S(_356_),
    .Z(_264_));
 MUX2_X1 _772_ (.A(_311_),
    .B(\mem[9][5] ),
    .S(_356_),
    .Z(_265_));
 MUX2_X1 _773_ (.A(_313_),
    .B(\mem[9][6] ),
    .S(_356_),
    .Z(_266_));
 MUX2_X1 _774_ (.A(_315_),
    .B(\mem[9][7] ),
    .S(_356_),
    .Z(_267_));
 AND2_X1 _775_ (.A1(\rd_ptr[0] ),
    .A2(net2),
    .ZN(_357_));
 INV_X2 _776_ (.A(net2),
    .ZN(_358_));
 NOR2_X1 _777_ (.A1(\rd_ptr[0] ),
    .A2(_358_),
    .ZN(_359_));
 INV_X1 _778_ (.A(net1),
    .ZN(_360_));
 AOI21_X2 _779_ (.A(_360_),
    .B1(_285_),
    .B2(_329_),
    .ZN(_361_));
 MUX2_X1 _780_ (.A(_357_),
    .B(_359_),
    .S(_361_),
    .Z(_136_));
 BUF_X2 _781_ (.A(net2),
    .Z(_362_));
 AND2_X1 _782_ (.A1(\rd_ptr[1] ),
    .A2(_362_),
    .ZN(_363_));
 AND2_X1 _783_ (.A1(_135_),
    .A2(_362_),
    .ZN(_364_));
 MUX2_X1 _784_ (.A(_363_),
    .B(_364_),
    .S(_361_),
    .Z(_137_));
 AND2_X1 _785_ (.A1(\rd_ptr[2] ),
    .A2(_362_),
    .ZN(_365_));
 NOR2_X1 _786_ (.A1(\rd_ptr[2] ),
    .A2(_358_),
    .ZN(_366_));
 NAND2_X1 _787_ (.A1(net1),
    .A2(_547_),
    .ZN(_367_));
 AOI21_X1 _788_ (.A(_367_),
    .B1(_329_),
    .B2(_285_),
    .ZN(_368_));
 MUX2_X1 _789_ (.A(_365_),
    .B(_366_),
    .S(_368_),
    .Z(_138_));
 AND2_X1 _790_ (.A1(\rd_ptr[3] ),
    .A2(_362_),
    .ZN(_369_));
 NOR2_X1 _791_ (.A1(\rd_ptr[3] ),
    .A2(_358_),
    .ZN(_370_));
 NAND4_X1 _792_ (.A1(net1),
    .A2(\rd_ptr[0] ),
    .A3(\rd_ptr[2] ),
    .A4(\rd_ptr[1] ),
    .ZN(_371_));
 AOI21_X1 _793_ (.A(_371_),
    .B1(_329_),
    .B2(_285_),
    .ZN(_372_));
 MUX2_X1 _794_ (.A(_369_),
    .B(_370_),
    .S(_372_),
    .Z(_139_));
 AND2_X1 _795_ (.A1(_134_),
    .A2(_362_),
    .ZN(_373_));
 MUX2_X1 _796_ (.A(_357_),
    .B(_373_),
    .S(_361_),
    .Z(_268_));
 AND2_X1 _797_ (.A1(\rd_ptr[4] ),
    .A2(_362_),
    .ZN(_374_));
 NOR2_X1 _798_ (.A1(\rd_ptr[4] ),
    .A2(_358_),
    .ZN(_375_));
 NAND4_X1 _799_ (.A1(net1),
    .A2(_547_),
    .A3(\rd_ptr[2] ),
    .A4(\rd_ptr[3] ),
    .ZN(_376_));
 AOI21_X1 _800_ (.A(_376_),
    .B1(_329_),
    .B2(_285_),
    .ZN(_377_));
 MUX2_X1 _801_ (.A(_374_),
    .B(_375_),
    .S(_377_),
    .Z(_269_));
 AND2_X1 _802_ (.A1(_132_),
    .A2(_362_),
    .ZN(_378_));
 AND2_X1 _803_ (.A1(\wr_ptr[0] ),
    .A2(_362_),
    .ZN(_379_));
 OAI21_X1 _804_ (.A(_299_),
    .B1(_285_),
    .B2(_293_),
    .ZN(_380_));
 MUX2_X1 _805_ (.A(_378_),
    .B(_379_),
    .S(_380_),
    .Z(_270_));
 AND2_X1 _806_ (.A1(_133_),
    .A2(_362_),
    .ZN(_381_));
 AND2_X1 _807_ (.A1(\wr_ptr[1] ),
    .A2(_362_),
    .ZN(_382_));
 MUX2_X1 _808_ (.A(_381_),
    .B(_382_),
    .S(_380_),
    .Z(_271_));
 NOR2_X1 _809_ (.A1(_297_),
    .A2(_358_),
    .ZN(_383_));
 NOR2_X1 _810_ (.A1(\wr_ptr[2] ),
    .A2(_358_),
    .ZN(_384_));
 AOI21_X1 _811_ (.A(_321_),
    .B1(_329_),
    .B2(net9),
    .ZN(_385_));
 MUX2_X1 _812_ (.A(_383_),
    .B(_384_),
    .S(_385_),
    .Z(_272_));
 NOR2_X1 _813_ (.A1(_296_),
    .A2(_358_),
    .ZN(_386_));
 NOR2_X1 _814_ (.A1(\wr_ptr[3] ),
    .A2(_358_),
    .ZN(_387_));
 NAND4_X1 _815_ (.A1(_299_),
    .A2(\wr_ptr[2] ),
    .A3(\wr_ptr[1] ),
    .A4(\wr_ptr[0] ),
    .ZN(_388_));
 AOI21_X1 _816_ (.A(_388_),
    .B1(_329_),
    .B2(net9),
    .ZN(_389_));
 MUX2_X1 _817_ (.A(_386_),
    .B(_387_),
    .S(_389_),
    .Z(_273_));
 AND2_X1 _818_ (.A1(\wr_ptr[4] ),
    .A2(net2),
    .ZN(_390_));
 NOR2_X1 _819_ (.A1(\wr_ptr[4] ),
    .A2(_358_),
    .ZN(_391_));
 MUX2_X1 _820_ (.A(_390_),
    .B(_391_),
    .S(_336_),
    .Z(_274_));
 INV_X1 _821_ (.A(net10),
    .ZN(net20));
 XOR2_X2 _822_ (.A(_275_),
    .B(_286_),
    .Z(_392_));
 NOR4_X1 _823_ (.A1(net8),
    .A2(net7),
    .A3(net9),
    .A4(_392_),
    .ZN(net3));
 NAND3_X2 _824_ (.A1(_286_),
    .A2(net8),
    .A3(net7),
    .ZN(_393_));
 NAND2_X4 _825_ (.A1(_285_),
    .A2(_393_),
    .ZN(net4));
 BUF_X4 _826_ (.A(_002_),
    .Z(_394_));
 BUF_X4 _827_ (.A(_394_),
    .Z(_395_));
 MUX2_X1 _828_ (.A(_004_),
    .B(_008_),
    .S(_395_),
    .Z(_396_));
 BUF_X4 _829_ (.A(_394_),
    .Z(_397_));
 MUX2_X1 _830_ (.A(_005_),
    .B(_009_),
    .S(_397_),
    .Z(_398_));
 CLKBUF_X3 _831_ (.A(_000_),
    .Z(_399_));
 BUF_X4 _832_ (.A(_399_),
    .Z(_400_));
 MUX2_X1 _833_ (.A(_396_),
    .B(_398_),
    .S(_400_),
    .Z(_401_));
 MUX2_X1 _834_ (.A(_012_),
    .B(_016_),
    .S(_397_),
    .Z(_402_));
 BUF_X4 _835_ (.A(_394_),
    .Z(_403_));
 MUX2_X1 _836_ (.A(_013_),
    .B(_017_),
    .S(_403_),
    .Z(_404_));
 BUF_X4 _837_ (.A(_399_),
    .Z(_405_));
 MUX2_X1 _838_ (.A(_402_),
    .B(_404_),
    .S(_405_),
    .Z(_406_));
 CLKBUF_X3 _839_ (.A(_003_),
    .Z(_407_));
 BUF_X4 _840_ (.A(_407_),
    .Z(_408_));
 MUX2_X1 _841_ (.A(_401_),
    .B(_406_),
    .S(_408_),
    .Z(_409_));
 BUF_X4 _842_ (.A(_394_),
    .Z(_410_));
 MUX2_X1 _843_ (.A(_006_),
    .B(_010_),
    .S(_410_),
    .Z(_411_));
 BUF_X4 _844_ (.A(_394_),
    .Z(_412_));
 MUX2_X1 _845_ (.A(_007_),
    .B(_011_),
    .S(_412_),
    .Z(_413_));
 BUF_X4 _846_ (.A(_399_),
    .Z(_414_));
 MUX2_X1 _847_ (.A(_411_),
    .B(_413_),
    .S(_414_),
    .Z(_415_));
 BUF_X4 _848_ (.A(_394_),
    .Z(_416_));
 MUX2_X1 _849_ (.A(_014_),
    .B(_018_),
    .S(_416_),
    .Z(_417_));
 MUX2_X1 _850_ (.A(_015_),
    .B(_019_),
    .S(_412_),
    .Z(_418_));
 MUX2_X1 _851_ (.A(_417_),
    .B(_418_),
    .S(_414_),
    .Z(_419_));
 MUX2_X1 _852_ (.A(_415_),
    .B(_419_),
    .S(_408_),
    .Z(_420_));
 BUF_X4 _853_ (.A(_001_),
    .Z(_421_));
 MUX2_X2 _854_ (.A(_409_),
    .B(_420_),
    .S(_421_),
    .Z(_422_));
 NOR2_X1 _855_ (.A1(net10),
    .A2(_422_),
    .ZN(net12));
 MUX2_X1 _856_ (.A(_020_),
    .B(_024_),
    .S(_395_),
    .Z(_423_));
 MUX2_X1 _857_ (.A(_021_),
    .B(_025_),
    .S(_397_),
    .Z(_424_));
 MUX2_X1 _858_ (.A(_423_),
    .B(_424_),
    .S(_400_),
    .Z(_425_));
 MUX2_X1 _859_ (.A(_028_),
    .B(_032_),
    .S(_397_),
    .Z(_426_));
 MUX2_X1 _860_ (.A(_029_),
    .B(_033_),
    .S(_403_),
    .Z(_427_));
 MUX2_X1 _861_ (.A(_426_),
    .B(_427_),
    .S(_405_),
    .Z(_428_));
 MUX2_X1 _862_ (.A(_425_),
    .B(_428_),
    .S(_408_),
    .Z(_429_));
 MUX2_X1 _863_ (.A(_022_),
    .B(_026_),
    .S(_410_),
    .Z(_430_));
 MUX2_X1 _864_ (.A(_023_),
    .B(_027_),
    .S(_412_),
    .Z(_431_));
 MUX2_X1 _865_ (.A(_430_),
    .B(_431_),
    .S(_414_),
    .Z(_432_));
 MUX2_X1 _866_ (.A(_030_),
    .B(_034_),
    .S(_416_),
    .Z(_433_));
 MUX2_X1 _867_ (.A(_031_),
    .B(_035_),
    .S(_412_),
    .Z(_434_));
 MUX2_X1 _868_ (.A(_433_),
    .B(_434_),
    .S(_414_),
    .Z(_435_));
 MUX2_X1 _869_ (.A(_432_),
    .B(_435_),
    .S(_408_),
    .Z(_436_));
 MUX2_X2 _870_ (.A(_429_),
    .B(_436_),
    .S(_421_),
    .Z(_437_));
 NOR2_X1 _871_ (.A1(net10),
    .A2(_437_),
    .ZN(net13));
 MUX2_X1 _872_ (.A(_036_),
    .B(_040_),
    .S(_395_),
    .Z(_438_));
 MUX2_X1 _873_ (.A(_037_),
    .B(_041_),
    .S(_397_),
    .Z(_439_));
 MUX2_X1 _874_ (.A(_438_),
    .B(_439_),
    .S(_400_),
    .Z(_440_));
 MUX2_X1 _875_ (.A(_044_),
    .B(_048_),
    .S(_397_),
    .Z(_441_));
 MUX2_X1 _876_ (.A(_045_),
    .B(_049_),
    .S(_403_),
    .Z(_442_));
 MUX2_X1 _877_ (.A(_441_),
    .B(_442_),
    .S(_405_),
    .Z(_443_));
 MUX2_X1 _878_ (.A(_440_),
    .B(_443_),
    .S(_407_),
    .Z(_444_));
 MUX2_X1 _879_ (.A(_038_),
    .B(_042_),
    .S(_410_),
    .Z(_445_));
 MUX2_X1 _880_ (.A(_039_),
    .B(_043_),
    .S(_416_),
    .Z(_446_));
 MUX2_X1 _881_ (.A(_445_),
    .B(_446_),
    .S(_405_),
    .Z(_447_));
 MUX2_X1 _882_ (.A(_046_),
    .B(_050_),
    .S(_416_),
    .Z(_448_));
 MUX2_X1 _883_ (.A(_047_),
    .B(_051_),
    .S(_412_),
    .Z(_449_));
 MUX2_X1 _884_ (.A(_448_),
    .B(_449_),
    .S(_414_),
    .Z(_450_));
 MUX2_X1 _885_ (.A(_447_),
    .B(_450_),
    .S(_408_),
    .Z(_451_));
 MUX2_X2 _886_ (.A(_444_),
    .B(_451_),
    .S(_421_),
    .Z(_452_));
 NOR2_X1 _887_ (.A1(net10),
    .A2(_452_),
    .ZN(net14));
 MUX2_X1 _888_ (.A(_052_),
    .B(_056_),
    .S(_395_),
    .Z(_453_));
 MUX2_X1 _889_ (.A(_053_),
    .B(_057_),
    .S(_397_),
    .Z(_454_));
 MUX2_X1 _890_ (.A(_453_),
    .B(_454_),
    .S(_400_),
    .Z(_455_));
 MUX2_X1 _891_ (.A(_060_),
    .B(_064_),
    .S(_397_),
    .Z(_456_));
 MUX2_X1 _892_ (.A(_061_),
    .B(_065_),
    .S(_403_),
    .Z(_457_));
 MUX2_X1 _893_ (.A(_456_),
    .B(_457_),
    .S(_405_),
    .Z(_458_));
 MUX2_X1 _894_ (.A(_455_),
    .B(_458_),
    .S(_407_),
    .Z(_459_));
 MUX2_X1 _895_ (.A(_054_),
    .B(_058_),
    .S(_410_),
    .Z(_460_));
 MUX2_X1 _896_ (.A(_055_),
    .B(_059_),
    .S(_416_),
    .Z(_461_));
 MUX2_X1 _897_ (.A(_460_),
    .B(_461_),
    .S(_405_),
    .Z(_462_));
 MUX2_X1 _898_ (.A(_062_),
    .B(_066_),
    .S(_416_),
    .Z(_463_));
 MUX2_X1 _899_ (.A(_063_),
    .B(_067_),
    .S(_412_),
    .Z(_464_));
 MUX2_X1 _900_ (.A(_463_),
    .B(_464_),
    .S(_414_),
    .Z(_465_));
 MUX2_X1 _901_ (.A(_462_),
    .B(_465_),
    .S(_408_),
    .Z(_466_));
 MUX2_X2 _902_ (.A(_459_),
    .B(_466_),
    .S(_421_),
    .Z(_467_));
 NOR2_X1 _903_ (.A1(net10),
    .A2(_467_),
    .ZN(net15));
 MUX2_X1 _904_ (.A(_068_),
    .B(_072_),
    .S(_394_),
    .Z(_468_));
 MUX2_X1 _905_ (.A(_069_),
    .B(_073_),
    .S(_397_),
    .Z(_469_));
 MUX2_X1 _906_ (.A(_468_),
    .B(_469_),
    .S(_400_),
    .Z(_470_));
 MUX2_X1 _907_ (.A(_076_),
    .B(_080_),
    .S(_397_),
    .Z(_471_));
 MUX2_X1 _908_ (.A(_077_),
    .B(_081_),
    .S(_403_),
    .Z(_472_));
 MUX2_X1 _909_ (.A(_471_),
    .B(_472_),
    .S(_400_),
    .Z(_473_));
 MUX2_X1 _910_ (.A(_470_),
    .B(_473_),
    .S(_407_),
    .Z(_474_));
 MUX2_X1 _911_ (.A(_070_),
    .B(_074_),
    .S(_410_),
    .Z(_475_));
 MUX2_X1 _912_ (.A(_071_),
    .B(_075_),
    .S(_416_),
    .Z(_476_));
 MUX2_X1 _913_ (.A(_475_),
    .B(_476_),
    .S(_405_),
    .Z(_477_));
 MUX2_X1 _914_ (.A(_078_),
    .B(_082_),
    .S(_403_),
    .Z(_478_));
 MUX2_X1 _915_ (.A(_079_),
    .B(_083_),
    .S(_412_),
    .Z(_479_));
 MUX2_X1 _916_ (.A(_478_),
    .B(_479_),
    .S(_414_),
    .Z(_480_));
 MUX2_X1 _917_ (.A(_477_),
    .B(_480_),
    .S(_408_),
    .Z(_481_));
 MUX2_X2 _918_ (.A(_474_),
    .B(_481_),
    .S(_421_),
    .Z(_482_));
 NOR2_X1 _919_ (.A1(net10),
    .A2(_482_),
    .ZN(net16));
 MUX2_X1 _920_ (.A(_084_),
    .B(_088_),
    .S(_394_),
    .Z(_483_));
 MUX2_X1 _921_ (.A(_085_),
    .B(_089_),
    .S(_395_),
    .Z(_484_));
 MUX2_X1 _922_ (.A(_483_),
    .B(_484_),
    .S(_400_),
    .Z(_485_));
 MUX2_X1 _923_ (.A(_092_),
    .B(_096_),
    .S(_395_),
    .Z(_486_));
 MUX2_X1 _924_ (.A(_093_),
    .B(_097_),
    .S(_403_),
    .Z(_487_));
 MUX2_X1 _925_ (.A(_486_),
    .B(_487_),
    .S(_400_),
    .Z(_488_));
 MUX2_X1 _926_ (.A(_485_),
    .B(_488_),
    .S(_407_),
    .Z(_489_));
 MUX2_X1 _927_ (.A(_086_),
    .B(_090_),
    .S(_410_),
    .Z(_490_));
 MUX2_X1 _928_ (.A(_087_),
    .B(_091_),
    .S(_416_),
    .Z(_491_));
 MUX2_X1 _929_ (.A(_490_),
    .B(_491_),
    .S(_405_),
    .Z(_492_));
 MUX2_X1 _930_ (.A(_094_),
    .B(_098_),
    .S(_403_),
    .Z(_493_));
 MUX2_X1 _931_ (.A(_095_),
    .B(_099_),
    .S(_412_),
    .Z(_494_));
 MUX2_X1 _932_ (.A(_493_),
    .B(_494_),
    .S(_414_),
    .Z(_495_));
 MUX2_X1 _933_ (.A(_492_),
    .B(_495_),
    .S(_408_),
    .Z(_496_));
 MUX2_X2 _934_ (.A(_489_),
    .B(_496_),
    .S(_421_),
    .Z(_497_));
 NOR2_X1 _935_ (.A1(net10),
    .A2(_497_),
    .ZN(net17));
 MUX2_X1 _936_ (.A(_100_),
    .B(_104_),
    .S(_394_),
    .Z(_498_));
 MUX2_X1 _937_ (.A(_101_),
    .B(_105_),
    .S(_395_),
    .Z(_499_));
 MUX2_X1 _938_ (.A(_498_),
    .B(_499_),
    .S(_399_),
    .Z(_500_));
 MUX2_X1 _939_ (.A(_108_),
    .B(_112_),
    .S(_395_),
    .Z(_501_));
 MUX2_X1 _940_ (.A(_109_),
    .B(_113_),
    .S(_410_),
    .Z(_502_));
 MUX2_X1 _941_ (.A(_501_),
    .B(_502_),
    .S(_400_),
    .Z(_503_));
 MUX2_X1 _942_ (.A(_500_),
    .B(_503_),
    .S(_407_),
    .Z(_504_));
 MUX2_X1 _943_ (.A(_102_),
    .B(_106_),
    .S(_410_),
    .Z(_505_));
 MUX2_X1 _944_ (.A(_103_),
    .B(_107_),
    .S(_416_),
    .Z(_506_));
 MUX2_X1 _945_ (.A(_505_),
    .B(_506_),
    .S(_405_),
    .Z(_507_));
 MUX2_X1 _946_ (.A(_110_),
    .B(_114_),
    .S(_403_),
    .Z(_508_));
 MUX2_X1 _947_ (.A(_111_),
    .B(_115_),
    .S(_412_),
    .Z(_509_));
 MUX2_X1 _948_ (.A(_508_),
    .B(_509_),
    .S(_414_),
    .Z(_510_));
 MUX2_X1 _949_ (.A(_507_),
    .B(_510_),
    .S(_408_),
    .Z(_511_));
 MUX2_X2 _950_ (.A(_504_),
    .B(_511_),
    .S(_421_),
    .Z(_512_));
 NOR2_X1 _951_ (.A1(net10),
    .A2(_512_),
    .ZN(net18));
 MUX2_X1 _952_ (.A(_116_),
    .B(_120_),
    .S(_394_),
    .Z(_513_));
 MUX2_X1 _953_ (.A(_117_),
    .B(_121_),
    .S(_395_),
    .Z(_514_));
 MUX2_X1 _954_ (.A(_513_),
    .B(_514_),
    .S(_399_),
    .Z(_515_));
 MUX2_X1 _955_ (.A(_124_),
    .B(_128_),
    .S(_395_),
    .Z(_516_));
 MUX2_X1 _956_ (.A(_125_),
    .B(_129_),
    .S(_410_),
    .Z(_517_));
 MUX2_X1 _957_ (.A(_516_),
    .B(_517_),
    .S(_400_),
    .Z(_518_));
 MUX2_X1 _958_ (.A(_515_),
    .B(_518_),
    .S(_407_),
    .Z(_519_));
 MUX2_X1 _959_ (.A(_118_),
    .B(_122_),
    .S(_410_),
    .Z(_520_));
 MUX2_X1 _960_ (.A(_119_),
    .B(_123_),
    .S(_416_),
    .Z(_521_));
 MUX2_X1 _961_ (.A(_520_),
    .B(_521_),
    .S(_405_),
    .Z(_522_));
 MUX2_X1 _962_ (.A(_126_),
    .B(_130_),
    .S(_403_),
    .Z(_523_));
 MUX2_X1 _963_ (.A(_127_),
    .B(_131_),
    .S(_412_),
    .Z(_524_));
 MUX2_X1 _964_ (.A(_523_),
    .B(_524_),
    .S(_414_),
    .Z(_525_));
 MUX2_X1 _965_ (.A(_522_),
    .B(_525_),
    .S(_408_),
    .Z(_526_));
 MUX2_X2 _966_ (.A(_519_),
    .B(_526_),
    .S(_421_),
    .Z(_527_));
 NOR2_X1 _967_ (.A1(net10),
    .A2(_527_),
    .ZN(net19));
 FA_X1 _968_ (.A(_536_),
    .B(\wr_ptr[1] ),
    .CI(_537_),
    .CO(_538_),
    .S(net6));
 HA_X1 _969_ (.A(_539_),
    .B(\wr_ptr[3] ),
    .CO(_540_),
    .S(_541_));
 HA_X1 _970_ (.A(_536_),
    .B(\wr_ptr[1] ),
    .CO(_542_),
    .S(_543_));
 HA_X1 _971_ (.A(_544_),
    .B(\wr_ptr[2] ),
    .CO(_545_),
    .S(_546_));
 HA_X1 _972_ (.A(\rd_ptr[0] ),
    .B(\rd_ptr[1] ),
    .CO(_547_),
    .S(_135_));
 HA_X1 _973_ (.A(_132_),
    .B(_548_),
    .CO(_549_),
    .S(_133_));
 HA_X1 _974_ (.A(_132_),
    .B(\wr_ptr[1] ),
    .CO(_550_),
    .S(_551_));
 HA_X1 _975_ (.A(\wr_ptr[0] ),
    .B(_548_),
    .CO(_552_),
    .S(_553_));
 HA_X1 _976_ (.A(\wr_ptr[0] ),
    .B(\wr_ptr[1] ),
    .CO(_554_),
    .S(_555_));
 HA_X1 _977_ (.A(\rd_ptr[0] ),
    .B(_132_),
    .CO(_556_),
    .S(_557_));
 DFF_X1 _978_ (.D(_136_),
    .CK(clknet_4_4_0_clk),
    .Q(_000_),
    .QN(_535_));
 DFF_X1 _979_ (.D(_137_),
    .CK(clknet_4_1_0_clk),
    .Q(_001_),
    .QN(_534_));
 DFF_X1 _980_ (.D(_138_),
    .CK(clknet_4_4_0_clk),
    .Q(_002_),
    .QN(_533_));
 DFF_X1 _981_ (.D(_139_),
    .CK(clknet_4_4_0_clk),
    .Q(_003_),
    .QN(_532_));
 DFF_X1 \mem[0][0]$_DFFE_PP_  (.D(_140_),
    .CK(clknet_4_13_0_clk),
    .Q(\mem[0][0] ),
    .QN(_004_));
 DFF_X1 \mem[0][1]$_DFFE_PP_  (.D(_141_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[0][1] ),
    .QN(_020_));
 DFF_X1 \mem[0][2]$_DFFE_PP_  (.D(_142_),
    .CK(clknet_4_13_0_clk),
    .Q(\mem[0][2] ),
    .QN(_036_));
 DFF_X1 \mem[0][3]$_DFFE_PP_  (.D(_143_),
    .CK(clknet_4_13_0_clk),
    .Q(\mem[0][3] ),
    .QN(_052_));
 DFF_X1 \mem[0][4]$_DFFE_PP_  (.D(_144_),
    .CK(clknet_4_13_0_clk),
    .Q(\mem[0][4] ),
    .QN(_068_));
 DFF_X1 \mem[0][5]$_DFFE_PP_  (.D(_145_),
    .CK(clknet_4_7_0_clk),
    .Q(\mem[0][5] ),
    .QN(_084_));
 DFF_X1 \mem[0][6]$_DFFE_PP_  (.D(_146_),
    .CK(clknet_4_5_0_clk),
    .Q(\mem[0][6] ),
    .QN(_100_));
 DFF_X1 \mem[0][7]$_DFFE_PP_  (.D(_147_),
    .CK(clknet_4_7_0_clk),
    .Q(\mem[0][7] ),
    .QN(_116_));
 DFF_X1 \mem[10][0]$_DFFE_PP_  (.D(_148_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[10][0] ),
    .QN(_014_));
 DFF_X1 \mem[10][1]$_DFFE_PP_  (.D(_149_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[10][1] ),
    .QN(_030_));
 DFF_X1 \mem[10][2]$_DFFE_PP_  (.D(_150_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[10][2] ),
    .QN(_046_));
 DFF_X1 \mem[10][3]$_DFFE_PP_  (.D(_151_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[10][3] ),
    .QN(_062_));
 DFF_X1 \mem[10][4]$_DFFE_PP_  (.D(_152_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[10][4] ),
    .QN(_078_));
 DFF_X1 \mem[10][5]$_DFFE_PP_  (.D(_153_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[10][5] ),
    .QN(_094_));
 DFF_X1 \mem[10][6]$_DFFE_PP_  (.D(_154_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[10][6] ),
    .QN(_110_));
 DFF_X1 \mem[10][7]$_DFFE_PP_  (.D(_155_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[10][7] ),
    .QN(_126_));
 DFF_X1 \mem[11][0]$_DFFE_PP_  (.D(_156_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[11][0] ),
    .QN(_015_));
 DFF_X1 \mem[11][1]$_DFFE_PP_  (.D(_157_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[11][1] ),
    .QN(_031_));
 DFF_X1 \mem[11][2]$_DFFE_PP_  (.D(_158_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[11][2] ),
    .QN(_047_));
 DFF_X1 \mem[11][3]$_DFFE_PP_  (.D(_159_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[11][3] ),
    .QN(_063_));
 DFF_X1 \mem[11][4]$_DFFE_PP_  (.D(_160_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[11][4] ),
    .QN(_079_));
 DFF_X1 \mem[11][5]$_DFFE_PP_  (.D(_161_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[11][5] ),
    .QN(_095_));
 DFF_X1 \mem[11][6]$_DFFE_PP_  (.D(_162_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[11][6] ),
    .QN(_111_));
 DFF_X1 \mem[11][7]$_DFFE_PP_  (.D(_163_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[11][7] ),
    .QN(_127_));
 DFF_X1 \mem[12][0]$_DFFE_PP_  (.D(_164_),
    .CK(clknet_4_15_0_clk),
    .Q(\mem[12][0] ),
    .QN(_016_));
 DFF_X1 \mem[12][1]$_DFFE_PP_  (.D(_165_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[12][1] ),
    .QN(_032_));
 DFF_X1 \mem[12][2]$_DFFE_PP_  (.D(_166_),
    .CK(clknet_4_15_0_clk),
    .Q(\mem[12][2] ),
    .QN(_048_));
 DFF_X1 \mem[12][3]$_DFFE_PP_  (.D(_167_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[12][3] ),
    .QN(_064_));
 DFF_X1 \mem[12][4]$_DFFE_PP_  (.D(_168_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[12][4] ),
    .QN(_080_));
 DFF_X1 \mem[12][5]$_DFFE_PP_  (.D(_169_),
    .CK(clknet_4_6_0_clk),
    .Q(\mem[12][5] ),
    .QN(_096_));
 DFF_X1 \mem[12][6]$_DFFE_PP_  (.D(_170_),
    .CK(clknet_4_5_0_clk),
    .Q(\mem[12][6] ),
    .QN(_112_));
 DFF_X1 \mem[12][7]$_DFFE_PP_  (.D(_171_),
    .CK(clknet_4_7_0_clk),
    .Q(\mem[12][7] ),
    .QN(_128_));
 DFF_X1 \mem[13][0]$_DFFE_PP_  (.D(_172_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[13][0] ),
    .QN(_017_));
 DFF_X1 \mem[13][1]$_DFFE_PP_  (.D(_173_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[13][1] ),
    .QN(_033_));
 DFF_X1 \mem[13][2]$_DFFE_PP_  (.D(_174_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[13][2] ),
    .QN(_049_));
 DFF_X1 \mem[13][3]$_DFFE_PP_  (.D(_175_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[13][3] ),
    .QN(_065_));
 DFF_X1 \mem[13][4]$_DFFE_PP_  (.D(_176_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[13][4] ),
    .QN(_081_));
 DFF_X1 \mem[13][5]$_DFFE_PP_  (.D(_177_),
    .CK(clknet_4_6_0_clk),
    .Q(\mem[13][5] ),
    .QN(_097_));
 DFF_X1 \mem[13][6]$_DFFE_PP_  (.D(_178_),
    .CK(clknet_4_5_0_clk),
    .Q(\mem[13][6] ),
    .QN(_113_));
 DFF_X1 \mem[13][7]$_DFFE_PP_  (.D(_179_),
    .CK(clknet_4_6_0_clk),
    .Q(\mem[13][7] ),
    .QN(_129_));
 DFF_X1 \mem[14][0]$_DFFE_PP_  (.D(_180_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[14][0] ),
    .QN(_018_));
 DFF_X1 \mem[14][1]$_DFFE_PP_  (.D(_181_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[14][1] ),
    .QN(_034_));
 DFF_X1 \mem[14][2]$_DFFE_PP_  (.D(_182_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[14][2] ),
    .QN(_050_));
 DFF_X1 \mem[14][3]$_DFFE_PP_  (.D(_183_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[14][3] ),
    .QN(_066_));
 DFF_X1 \mem[14][4]$_DFFE_PP_  (.D(_184_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[14][4] ),
    .QN(_082_));
 DFF_X1 \mem[14][5]$_DFFE_PP_  (.D(_185_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[14][5] ),
    .QN(_098_));
 DFF_X1 \mem[14][6]$_DFFE_PP_  (.D(_186_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[14][6] ),
    .QN(_114_));
 DFF_X1 \mem[14][7]$_DFFE_PP_  (.D(_187_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[14][7] ),
    .QN(_130_));
 DFF_X1 \mem[15][0]$_DFFE_PP_  (.D(_188_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[15][0] ),
    .QN(_019_));
 DFF_X1 \mem[15][1]$_DFFE_PP_  (.D(_189_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[15][1] ),
    .QN(_035_));
 DFF_X1 \mem[15][2]$_DFFE_PP_  (.D(_190_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[15][2] ),
    .QN(_051_));
 DFF_X1 \mem[15][3]$_DFFE_PP_  (.D(_191_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[15][3] ),
    .QN(_067_));
 DFF_X1 \mem[15][4]$_DFFE_PP_  (.D(_192_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[15][4] ),
    .QN(_083_));
 DFF_X1 \mem[15][5]$_DFFE_PP_  (.D(_193_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[15][5] ),
    .QN(_099_));
 DFF_X1 \mem[15][6]$_DFFE_PP_  (.D(_194_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[15][6] ),
    .QN(_115_));
 DFF_X1 \mem[15][7]$_DFFE_PP_  (.D(_195_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[15][7] ),
    .QN(_131_));
 DFF_X1 \mem[1][0]$_DFFE_PP_  (.D(_196_),
    .CK(clknet_4_15_0_clk),
    .Q(\mem[1][0] ),
    .QN(_005_));
 DFF_X1 \mem[1][1]$_DFFE_PP_  (.D(_197_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[1][1] ),
    .QN(_021_));
 DFF_X1 \mem[1][2]$_DFFE_PP_  (.D(_198_),
    .CK(clknet_4_15_0_clk),
    .Q(\mem[1][2] ),
    .QN(_037_));
 DFF_X1 \mem[1][3]$_DFFE_PP_  (.D(_199_),
    .CK(clknet_4_13_0_clk),
    .Q(\mem[1][3] ),
    .QN(_053_));
 DFF_X1 \mem[1][4]$_DFFE_PP_  (.D(_200_),
    .CK(clknet_4_13_0_clk),
    .Q(\mem[1][4] ),
    .QN(_069_));
 DFF_X1 \mem[1][5]$_DFFE_PP_  (.D(_201_),
    .CK(clknet_4_7_0_clk),
    .Q(\mem[1][5] ),
    .QN(_085_));
 DFF_X1 \mem[1][6]$_DFFE_PP_  (.D(_202_),
    .CK(clknet_4_5_0_clk),
    .Q(\mem[1][6] ),
    .QN(_101_));
 DFF_X1 \mem[1][7]$_DFFE_PP_  (.D(_203_),
    .CK(clknet_4_7_0_clk),
    .Q(\mem[1][7] ),
    .QN(_117_));
 DFF_X1 \mem[2][0]$_DFFE_PP_  (.D(_204_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[2][0] ),
    .QN(_006_));
 DFF_X1 \mem[2][1]$_DFFE_PP_  (.D(_205_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[2][1] ),
    .QN(_022_));
 DFF_X1 \mem[2][2]$_DFFE_PP_  (.D(_206_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[2][2] ),
    .QN(_038_));
 DFF_X1 \mem[2][3]$_DFFE_PP_  (.D(_207_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[2][3] ),
    .QN(_054_));
 DFF_X1 \mem[2][4]$_DFFE_PP_  (.D(_208_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[2][4] ),
    .QN(_070_));
 DFF_X1 \mem[2][5]$_DFFE_PP_  (.D(_209_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[2][5] ),
    .QN(_086_));
 DFF_X1 \mem[2][6]$_DFFE_PP_  (.D(_210_),
    .CK(clknet_4_0_0_clk),
    .Q(\mem[2][6] ),
    .QN(_102_));
 DFF_X1 \mem[2][7]$_DFFE_PP_  (.D(_211_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[2][7] ),
    .QN(_118_));
 DFF_X1 \mem[3][0]$_DFFE_PP_  (.D(_212_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[3][0] ),
    .QN(_007_));
 DFF_X1 \mem[3][1]$_DFFE_PP_  (.D(_213_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[3][1] ),
    .QN(_023_));
 DFF_X1 \mem[3][2]$_DFFE_PP_  (.D(_214_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[3][2] ),
    .QN(_039_));
 DFF_X1 \mem[3][3]$_DFFE_PP_  (.D(_215_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[3][3] ),
    .QN(_055_));
 DFF_X1 \mem[3][4]$_DFFE_PP_  (.D(_216_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[3][4] ),
    .QN(_071_));
 DFF_X1 \mem[3][5]$_DFFE_PP_  (.D(_217_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[3][5] ),
    .QN(_087_));
 DFF_X1 \mem[3][6]$_DFFE_PP_  (.D(_218_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[3][6] ),
    .QN(_103_));
 DFF_X1 \mem[3][7]$_DFFE_PP_  (.D(_219_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[3][7] ),
    .QN(_119_));
 DFF_X1 \mem[4][0]$_DFFE_PP_  (.D(_220_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[4][0] ),
    .QN(_008_));
 DFF_X1 \mem[4][1]$_DFFE_PP_  (.D(_221_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[4][1] ),
    .QN(_024_));
 DFF_X1 \mem[4][2]$_DFFE_PP_  (.D(_222_),
    .CK(clknet_4_13_0_clk),
    .Q(\mem[4][2] ),
    .QN(_040_));
 DFF_X1 \mem[4][3]$_DFFE_PP_  (.D(_223_),
    .CK(clknet_4_13_0_clk),
    .Q(\mem[4][3] ),
    .QN(_056_));
 DFF_X1 \mem[4][4]$_DFFE_PP_  (.D(_224_),
    .CK(clknet_4_13_0_clk),
    .Q(\mem[4][4] ),
    .QN(_072_));
 DFF_X1 \mem[4][5]$_DFFE_PP_  (.D(_225_),
    .CK(clknet_4_7_0_clk),
    .Q(\mem[4][5] ),
    .QN(_088_));
 DFF_X1 \mem[4][6]$_DFFE_PP_  (.D(_226_),
    .CK(clknet_4_5_0_clk),
    .Q(\mem[4][6] ),
    .QN(_104_));
 DFF_X1 \mem[4][7]$_DFFE_PP_  (.D(_227_),
    .CK(clknet_4_7_0_clk),
    .Q(\mem[4][7] ),
    .QN(_120_));
 DFF_X1 \mem[5][0]$_DFFE_PP_  (.D(_228_),
    .CK(clknet_4_15_0_clk),
    .Q(\mem[5][0] ),
    .QN(_009_));
 DFF_X1 \mem[5][1]$_DFFE_PP_  (.D(_229_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[5][1] ),
    .QN(_025_));
 DFF_X1 \mem[5][2]$_DFFE_PP_  (.D(_230_),
    .CK(clknet_4_15_0_clk),
    .Q(\mem[5][2] ),
    .QN(_041_));
 DFF_X1 \mem[5][3]$_DFFE_PP_  (.D(_231_),
    .CK(clknet_4_13_0_clk),
    .Q(\mem[5][3] ),
    .QN(_057_));
 DFF_X1 \mem[5][4]$_DFFE_PP_  (.D(_232_),
    .CK(clknet_4_13_0_clk),
    .Q(\mem[5][4] ),
    .QN(_073_));
 DFF_X1 \mem[5][5]$_DFFE_PP_  (.D(_233_),
    .CK(clknet_4_7_0_clk),
    .Q(\mem[5][5] ),
    .QN(_089_));
 DFF_X1 \mem[5][6]$_DFFE_PP_  (.D(_234_),
    .CK(clknet_4_7_0_clk),
    .Q(\mem[5][6] ),
    .QN(_105_));
 DFF_X1 \mem[5][7]$_DFFE_PP_  (.D(_235_),
    .CK(clknet_4_7_0_clk),
    .Q(\mem[5][7] ),
    .QN(_121_));
 DFF_X1 \mem[6][0]$_DFFE_PP_  (.D(_236_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[6][0] ),
    .QN(_010_));
 DFF_X1 \mem[6][1]$_DFFE_PP_  (.D(_237_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[6][1] ),
    .QN(_026_));
 DFF_X1 \mem[6][2]$_DFFE_PP_  (.D(_238_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[6][2] ),
    .QN(_042_));
 DFF_X1 \mem[6][3]$_DFFE_PP_  (.D(_239_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[6][3] ),
    .QN(_058_));
 DFF_X1 \mem[6][4]$_DFFE_PP_  (.D(_240_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[6][4] ),
    .QN(_074_));
 DFF_X1 \mem[6][5]$_DFFE_PP_  (.D(_241_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[6][5] ),
    .QN(_090_));
 DFF_X1 \mem[6][6]$_DFFE_PP_  (.D(_242_),
    .CK(clknet_4_1_0_clk),
    .Q(\mem[6][6] ),
    .QN(_106_));
 DFF_X1 \mem[6][7]$_DFFE_PP_  (.D(_243_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[6][7] ),
    .QN(_122_));
 DFF_X1 \mem[7][0]$_DFFE_PP_  (.D(_244_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[7][0] ),
    .QN(_011_));
 DFF_X1 \mem[7][1]$_DFFE_PP_  (.D(_245_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[7][1] ),
    .QN(_027_));
 DFF_X1 \mem[7][2]$_DFFE_PP_  (.D(_246_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[7][2] ),
    .QN(_043_));
 DFF_X1 \mem[7][3]$_DFFE_PP_  (.D(_247_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[7][3] ),
    .QN(_059_));
 DFF_X1 \mem[7][4]$_DFFE_PP_  (.D(_248_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[7][4] ),
    .QN(_075_));
 DFF_X1 \mem[7][5]$_DFFE_PP_  (.D(_249_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[7][5] ),
    .QN(_091_));
 DFF_X1 \mem[7][6]$_DFFE_PP_  (.D(_250_),
    .CK(clknet_4_1_0_clk),
    .Q(\mem[7][6] ),
    .QN(_107_));
 DFF_X1 \mem[7][7]$_DFFE_PP_  (.D(_251_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[7][7] ),
    .QN(_123_));
 DFF_X1 \mem[8][0]$_DFFE_PP_  (.D(_252_),
    .CK(clknet_4_15_0_clk),
    .Q(\mem[8][0] ),
    .QN(_012_));
 DFF_X1 \mem[8][1]$_DFFE_PP_  (.D(_253_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[8][1] ),
    .QN(_028_));
 DFF_X1 \mem[8][2]$_DFFE_PP_  (.D(_254_),
    .CK(clknet_4_15_0_clk),
    .Q(\mem[8][2] ),
    .QN(_044_));
 DFF_X1 \mem[8][3]$_DFFE_PP_  (.D(_255_),
    .CK(clknet_4_13_0_clk),
    .Q(\mem[8][3] ),
    .QN(_060_));
 DFF_X1 \mem[8][4]$_DFFE_PP_  (.D(_256_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[8][4] ),
    .QN(_076_));
 DFF_X1 \mem[8][5]$_DFFE_PP_  (.D(_257_),
    .CK(clknet_4_6_0_clk),
    .Q(\mem[8][5] ),
    .QN(_092_));
 DFF_X1 \mem[8][6]$_DFFE_PP_  (.D(_258_),
    .CK(clknet_4_5_0_clk),
    .Q(\mem[8][6] ),
    .QN(_108_));
 DFF_X1 \mem[8][7]$_DFFE_PP_  (.D(_259_),
    .CK(clknet_4_6_0_clk),
    .Q(\mem[8][7] ),
    .QN(_124_));
 DFF_X1 \mem[9][0]$_DFFE_PP_  (.D(_260_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[9][0] ),
    .QN(_013_));
 DFF_X1 \mem[9][1]$_DFFE_PP_  (.D(_261_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[9][1] ),
    .QN(_029_));
 DFF_X1 \mem[9][2]$_DFFE_PP_  (.D(_262_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[9][2] ),
    .QN(_045_));
 DFF_X1 \mem[9][3]$_DFFE_PP_  (.D(_263_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[9][3] ),
    .QN(_061_));
 DFF_X1 \mem[9][4]$_DFFE_PP_  (.D(_264_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[9][4] ),
    .QN(_077_));
 DFF_X1 \mem[9][5]$_DFFE_PP_  (.D(_265_),
    .CK(clknet_4_6_0_clk),
    .Q(\mem[9][5] ),
    .QN(_093_));
 DFF_X1 \mem[9][6]$_DFFE_PP_  (.D(_266_),
    .CK(clknet_4_5_0_clk),
    .Q(\mem[9][6] ),
    .QN(_109_));
 DFF_X1 \mem[9][7]$_DFFE_PP_  (.D(_267_),
    .CK(clknet_4_6_0_clk),
    .Q(\mem[9][7] ),
    .QN(_125_));
 DFF_X2 \rd_ptr[0]$_SDFFE_PN0P_  (.D(_268_),
    .CK(clknet_4_4_0_clk),
    .Q(\rd_ptr[0] ),
    .QN(_134_));
 DFF_X1 \rd_ptr[1]$_SDFFE_PN0P_  (.D(_137_),
    .CK(clknet_4_1_0_clk),
    .Q(\rd_ptr[1] ),
    .QN(_536_));
 DFF_X1 \rd_ptr[2]$_SDFFE_PN0P_  (.D(_138_),
    .CK(clknet_4_4_0_clk),
    .Q(\rd_ptr[2] ),
    .QN(_544_));
 DFF_X1 \rd_ptr[3]$_SDFFE_PN0P_  (.D(_139_),
    .CK(clknet_4_1_0_clk),
    .Q(\rd_ptr[3] ),
    .QN(_539_));
 DFF_X1 \rd_ptr[4]$_SDFFE_PN0P_  (.D(_269_),
    .CK(clknet_4_1_0_clk),
    .Q(\rd_ptr[4] ),
    .QN(_531_));
 DFF_X2 \wr_ptr[0]$_SDFFE_PN0P_  (.D(_270_),
    .CK(clknet_4_0_0_clk),
    .Q(\wr_ptr[0] ),
    .QN(_132_));
 DFF_X2 \wr_ptr[1]$_SDFFE_PN0P_  (.D(_271_),
    .CK(clknet_4_1_0_clk),
    .Q(\wr_ptr[1] ),
    .QN(_548_));
 DFF_X2 \wr_ptr[2]$_SDFFE_PN0P_  (.D(_272_),
    .CK(clknet_4_0_0_clk),
    .Q(\wr_ptr[2] ),
    .QN(_530_));
 DFF_X2 \wr_ptr[3]$_SDFFE_PN0P_  (.D(_273_),
    .CK(clknet_4_0_0_clk),
    .Q(\wr_ptr[3] ),
    .QN(_529_));
 DFF_X1 \wr_ptr[4]$_SDFFE_PN0P_  (.D(_274_),
    .CK(clknet_4_0_0_clk),
    .Q(\wr_ptr[4] ),
    .QN(_528_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Right_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Right_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Right_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Right_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Right_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Right_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Right_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Right_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Right_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Right_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Right_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Right_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Right_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Right_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Right_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Right_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Right_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Right_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Right_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Right_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Right_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Right_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Right_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Right_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Right_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Right_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Right_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Right_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Right_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Right_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Right_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Right_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Right_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Right_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Right_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Right_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Right_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Right_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_Right_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_Right_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_Right_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_Right_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_Right_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_Right_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_Right_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_Right_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_Right_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_Right_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_Right_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_Right_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_Right_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_Right_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_Right_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_Right_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_Right_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_Right_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_Right_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_Right_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_Right_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_Right_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_Right_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_Right_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_Right_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_Right_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_Right_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_Right_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_Right_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_Right_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_Right_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_Right_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_Right_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_Right_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_Right_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_Right_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_Right_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_Right_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Right_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Right_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Right_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Right_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Right_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Right_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Right_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Right_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Right_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Right_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Right_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Right_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Right_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Right_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Right_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Right_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_224_Right_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_225_Right_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_226_Right_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_227_Right_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_228_Right_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_229_Right_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_230_Right_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_231_Right_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_232_Right_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_233_Right_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_234_Right_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_235_Right_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_236_Right_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_237_Right_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_238_Right_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_239_Right_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_240_Right_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_241_Right_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_242_Right_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_243_Right_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_244_Right_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_245_Right_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_246_Right_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_247_Right_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_248_Right_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_249_Right_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_250_Right_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_251_Right_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_252_Right_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_253_Right_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_254_Right_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_255_Right_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_256_Right_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_257_Right_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_258_Right_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_259_Right_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_260_Right_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_261_Right_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_262_Right_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_263_Right_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_264_Right_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_265_Right_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_266_Right_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_267_Right_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_268_Right_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_269_Right_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_270_Right_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_271_Right_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_272_Right_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_273_Right_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_274_Right_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_275_Right_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_276_Right_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_277_Right_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_278_Right_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_279_Right_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_280_Right_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_281_Right_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_282_Right_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_283_Right_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_284_Right_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_285_Right_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_286_Right_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_287_Right_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_288_Right_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_289_Right_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_290_Right_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_291_Right_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_292_Right_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_293_Right_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_294_Right_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_295_Right_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_296_Right_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_297_Right_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_298_Right_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_299_Right_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_300_Right_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_301_Right_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_302_Right_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_303_Right_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_304_Right_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_305_Right_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_306_Right_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_307_Right_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_308_Right_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_309_Right_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_310_Right_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_311_Right_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_312_Right_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_313_Right_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_314_Right_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_315_Right_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_316_Right_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_317_Right_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_318_Right_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_319_Right_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_320_Right_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_321_Right_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_322_Right_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_323_Right_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_324_Right_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_325_Right_325 ();
 TAPCELL_X1 PHY_EDGE_ROW_326_Right_326 ();
 TAPCELL_X1 PHY_EDGE_ROW_327_Right_327 ();
 TAPCELL_X1 PHY_EDGE_ROW_328_Right_328 ();
 TAPCELL_X1 PHY_EDGE_ROW_329_Right_329 ();
 TAPCELL_X1 PHY_EDGE_ROW_330_Right_330 ();
 TAPCELL_X1 PHY_EDGE_ROW_331_Right_331 ();
 TAPCELL_X1 PHY_EDGE_ROW_332_Right_332 ();
 TAPCELL_X1 PHY_EDGE_ROW_333_Right_333 ();
 TAPCELL_X1 PHY_EDGE_ROW_334_Right_334 ();
 TAPCELL_X1 PHY_EDGE_ROW_335_Right_335 ();
 TAPCELL_X1 PHY_EDGE_ROW_336_Right_336 ();
 TAPCELL_X1 PHY_EDGE_ROW_337_Right_337 ();
 TAPCELL_X1 PHY_EDGE_ROW_338_Right_338 ();
 TAPCELL_X1 PHY_EDGE_ROW_339_Right_339 ();
 TAPCELL_X1 PHY_EDGE_ROW_340_Right_340 ();
 TAPCELL_X1 PHY_EDGE_ROW_341_Right_341 ();
 TAPCELL_X1 PHY_EDGE_ROW_342_Right_342 ();
 TAPCELL_X1 PHY_EDGE_ROW_343_Right_343 ();
 TAPCELL_X1 PHY_EDGE_ROW_344_Right_344 ();
 TAPCELL_X1 PHY_EDGE_ROW_345_Right_345 ();
 TAPCELL_X1 PHY_EDGE_ROW_346_Right_346 ();
 TAPCELL_X1 PHY_EDGE_ROW_347_Right_347 ();
 TAPCELL_X1 PHY_EDGE_ROW_348_Right_348 ();
 TAPCELL_X1 PHY_EDGE_ROW_349_Right_349 ();
 TAPCELL_X1 PHY_EDGE_ROW_350_Right_350 ();
 TAPCELL_X1 PHY_EDGE_ROW_351_Right_351 ();
 TAPCELL_X1 PHY_EDGE_ROW_352_Right_352 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_353 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_354 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_355 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_356 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_357 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_358 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_359 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_360 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_361 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_362 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_363 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_364 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_365 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_366 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_367 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_368 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_369 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_370 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_371 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_372 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_373 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_374 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_375 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_376 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_377 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_378 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_379 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_380 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_381 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_382 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_383 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_384 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_385 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_386 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_387 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_388 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_389 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_390 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_391 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_392 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_393 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_394 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_395 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_396 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_397 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_398 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_399 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_400 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_401 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_402 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_403 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_404 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_405 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_406 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_407 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_408 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_409 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_410 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_411 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_412 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_413 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_414 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_415 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_416 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_417 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_418 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_419 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_420 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_421 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_422 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Left_423 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Left_424 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Left_425 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Left_426 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Left_427 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Left_428 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Left_429 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Left_430 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Left_431 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_432 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_433 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_434 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_435 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_436 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_437 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_438 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_439 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_440 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Left_441 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Left_442 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Left_443 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Left_444 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Left_445 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Left_446 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Left_447 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Left_448 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Left_449 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Left_450 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Left_451 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Left_452 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Left_453 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Left_454 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Left_455 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Left_456 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Left_457 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Left_458 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Left_459 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Left_460 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Left_461 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Left_462 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Left_463 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Left_464 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Left_465 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Left_466 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Left_467 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Left_468 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Left_469 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Left_470 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Left_471 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Left_472 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Left_473 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Left_474 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Left_475 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Left_476 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Left_477 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Left_478 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Left_479 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Left_480 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Left_481 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Left_482 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Left_483 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Left_484 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Left_485 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Left_486 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Left_487 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Left_488 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Left_489 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Left_490 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Left_491 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Left_492 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Left_493 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Left_494 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Left_495 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Left_496 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Left_497 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Left_498 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Left_499 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Left_500 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Left_501 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Left_502 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Left_503 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Left_504 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Left_505 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Left_506 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Left_507 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Left_508 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Left_509 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Left_510 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Left_511 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Left_512 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Left_513 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Left_514 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Left_515 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Left_516 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Left_517 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Left_518 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Left_519 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Left_520 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Left_521 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Left_522 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_Left_523 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_Left_524 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_Left_525 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_Left_526 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_Left_527 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_Left_528 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_Left_529 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_Left_530 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_Left_531 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_Left_532 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_Left_533 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_Left_534 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_Left_535 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_Left_536 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_Left_537 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_Left_538 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_Left_539 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_Left_540 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_Left_541 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_Left_542 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_Left_543 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_Left_544 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_Left_545 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_Left_546 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_Left_547 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_Left_548 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_Left_549 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_Left_550 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_Left_551 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_Left_552 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_Left_553 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_Left_554 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_Left_555 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_Left_556 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_Left_557 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_Left_558 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_Left_559 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_Left_560 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Left_561 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Left_562 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Left_563 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Left_564 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Left_565 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Left_566 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Left_567 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Left_568 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Left_569 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Left_570 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Left_571 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Left_572 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Left_573 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Left_574 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Left_575 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Left_576 ();
 TAPCELL_X1 PHY_EDGE_ROW_224_Left_577 ();
 TAPCELL_X1 PHY_EDGE_ROW_225_Left_578 ();
 TAPCELL_X1 PHY_EDGE_ROW_226_Left_579 ();
 TAPCELL_X1 PHY_EDGE_ROW_227_Left_580 ();
 TAPCELL_X1 PHY_EDGE_ROW_228_Left_581 ();
 TAPCELL_X1 PHY_EDGE_ROW_229_Left_582 ();
 TAPCELL_X1 PHY_EDGE_ROW_230_Left_583 ();
 TAPCELL_X1 PHY_EDGE_ROW_231_Left_584 ();
 TAPCELL_X1 PHY_EDGE_ROW_232_Left_585 ();
 TAPCELL_X1 PHY_EDGE_ROW_233_Left_586 ();
 TAPCELL_X1 PHY_EDGE_ROW_234_Left_587 ();
 TAPCELL_X1 PHY_EDGE_ROW_235_Left_588 ();
 TAPCELL_X1 PHY_EDGE_ROW_236_Left_589 ();
 TAPCELL_X1 PHY_EDGE_ROW_237_Left_590 ();
 TAPCELL_X1 PHY_EDGE_ROW_238_Left_591 ();
 TAPCELL_X1 PHY_EDGE_ROW_239_Left_592 ();
 TAPCELL_X1 PHY_EDGE_ROW_240_Left_593 ();
 TAPCELL_X1 PHY_EDGE_ROW_241_Left_594 ();
 TAPCELL_X1 PHY_EDGE_ROW_242_Left_595 ();
 TAPCELL_X1 PHY_EDGE_ROW_243_Left_596 ();
 TAPCELL_X1 PHY_EDGE_ROW_244_Left_597 ();
 TAPCELL_X1 PHY_EDGE_ROW_245_Left_598 ();
 TAPCELL_X1 PHY_EDGE_ROW_246_Left_599 ();
 TAPCELL_X1 PHY_EDGE_ROW_247_Left_600 ();
 TAPCELL_X1 PHY_EDGE_ROW_248_Left_601 ();
 TAPCELL_X1 PHY_EDGE_ROW_249_Left_602 ();
 TAPCELL_X1 PHY_EDGE_ROW_250_Left_603 ();
 TAPCELL_X1 PHY_EDGE_ROW_251_Left_604 ();
 TAPCELL_X1 PHY_EDGE_ROW_252_Left_605 ();
 TAPCELL_X1 PHY_EDGE_ROW_253_Left_606 ();
 TAPCELL_X1 PHY_EDGE_ROW_254_Left_607 ();
 TAPCELL_X1 PHY_EDGE_ROW_255_Left_608 ();
 TAPCELL_X1 PHY_EDGE_ROW_256_Left_609 ();
 TAPCELL_X1 PHY_EDGE_ROW_257_Left_610 ();
 TAPCELL_X1 PHY_EDGE_ROW_258_Left_611 ();
 TAPCELL_X1 PHY_EDGE_ROW_259_Left_612 ();
 TAPCELL_X1 PHY_EDGE_ROW_260_Left_613 ();
 TAPCELL_X1 PHY_EDGE_ROW_261_Left_614 ();
 TAPCELL_X1 PHY_EDGE_ROW_262_Left_615 ();
 TAPCELL_X1 PHY_EDGE_ROW_263_Left_616 ();
 TAPCELL_X1 PHY_EDGE_ROW_264_Left_617 ();
 TAPCELL_X1 PHY_EDGE_ROW_265_Left_618 ();
 TAPCELL_X1 PHY_EDGE_ROW_266_Left_619 ();
 TAPCELL_X1 PHY_EDGE_ROW_267_Left_620 ();
 TAPCELL_X1 PHY_EDGE_ROW_268_Left_621 ();
 TAPCELL_X1 PHY_EDGE_ROW_269_Left_622 ();
 TAPCELL_X1 PHY_EDGE_ROW_270_Left_623 ();
 TAPCELL_X1 PHY_EDGE_ROW_271_Left_624 ();
 TAPCELL_X1 PHY_EDGE_ROW_272_Left_625 ();
 TAPCELL_X1 PHY_EDGE_ROW_273_Left_626 ();
 TAPCELL_X1 PHY_EDGE_ROW_274_Left_627 ();
 TAPCELL_X1 PHY_EDGE_ROW_275_Left_628 ();
 TAPCELL_X1 PHY_EDGE_ROW_276_Left_629 ();
 TAPCELL_X1 PHY_EDGE_ROW_277_Left_630 ();
 TAPCELL_X1 PHY_EDGE_ROW_278_Left_631 ();
 TAPCELL_X1 PHY_EDGE_ROW_279_Left_632 ();
 TAPCELL_X1 PHY_EDGE_ROW_280_Left_633 ();
 TAPCELL_X1 PHY_EDGE_ROW_281_Left_634 ();
 TAPCELL_X1 PHY_EDGE_ROW_282_Left_635 ();
 TAPCELL_X1 PHY_EDGE_ROW_283_Left_636 ();
 TAPCELL_X1 PHY_EDGE_ROW_284_Left_637 ();
 TAPCELL_X1 PHY_EDGE_ROW_285_Left_638 ();
 TAPCELL_X1 PHY_EDGE_ROW_286_Left_639 ();
 TAPCELL_X1 PHY_EDGE_ROW_287_Left_640 ();
 TAPCELL_X1 PHY_EDGE_ROW_288_Left_641 ();
 TAPCELL_X1 PHY_EDGE_ROW_289_Left_642 ();
 TAPCELL_X1 PHY_EDGE_ROW_290_Left_643 ();
 TAPCELL_X1 PHY_EDGE_ROW_291_Left_644 ();
 TAPCELL_X1 PHY_EDGE_ROW_292_Left_645 ();
 TAPCELL_X1 PHY_EDGE_ROW_293_Left_646 ();
 TAPCELL_X1 PHY_EDGE_ROW_294_Left_647 ();
 TAPCELL_X1 PHY_EDGE_ROW_295_Left_648 ();
 TAPCELL_X1 PHY_EDGE_ROW_296_Left_649 ();
 TAPCELL_X1 PHY_EDGE_ROW_297_Left_650 ();
 TAPCELL_X1 PHY_EDGE_ROW_298_Left_651 ();
 TAPCELL_X1 PHY_EDGE_ROW_299_Left_652 ();
 TAPCELL_X1 PHY_EDGE_ROW_300_Left_653 ();
 TAPCELL_X1 PHY_EDGE_ROW_301_Left_654 ();
 TAPCELL_X1 PHY_EDGE_ROW_302_Left_655 ();
 TAPCELL_X1 PHY_EDGE_ROW_303_Left_656 ();
 TAPCELL_X1 PHY_EDGE_ROW_304_Left_657 ();
 TAPCELL_X1 PHY_EDGE_ROW_305_Left_658 ();
 TAPCELL_X1 PHY_EDGE_ROW_306_Left_659 ();
 TAPCELL_X1 PHY_EDGE_ROW_307_Left_660 ();
 TAPCELL_X1 PHY_EDGE_ROW_308_Left_661 ();
 TAPCELL_X1 PHY_EDGE_ROW_309_Left_662 ();
 TAPCELL_X1 PHY_EDGE_ROW_310_Left_663 ();
 TAPCELL_X1 PHY_EDGE_ROW_311_Left_664 ();
 TAPCELL_X1 PHY_EDGE_ROW_312_Left_665 ();
 TAPCELL_X1 PHY_EDGE_ROW_313_Left_666 ();
 TAPCELL_X1 PHY_EDGE_ROW_314_Left_667 ();
 TAPCELL_X1 PHY_EDGE_ROW_315_Left_668 ();
 TAPCELL_X1 PHY_EDGE_ROW_316_Left_669 ();
 TAPCELL_X1 PHY_EDGE_ROW_317_Left_670 ();
 TAPCELL_X1 PHY_EDGE_ROW_318_Left_671 ();
 TAPCELL_X1 PHY_EDGE_ROW_319_Left_672 ();
 TAPCELL_X1 PHY_EDGE_ROW_320_Left_673 ();
 TAPCELL_X1 PHY_EDGE_ROW_321_Left_674 ();
 TAPCELL_X1 PHY_EDGE_ROW_322_Left_675 ();
 TAPCELL_X1 PHY_EDGE_ROW_323_Left_676 ();
 TAPCELL_X1 PHY_EDGE_ROW_324_Left_677 ();
 TAPCELL_X1 PHY_EDGE_ROW_325_Left_678 ();
 TAPCELL_X1 PHY_EDGE_ROW_326_Left_679 ();
 TAPCELL_X1 PHY_EDGE_ROW_327_Left_680 ();
 TAPCELL_X1 PHY_EDGE_ROW_328_Left_681 ();
 TAPCELL_X1 PHY_EDGE_ROW_329_Left_682 ();
 TAPCELL_X1 PHY_EDGE_ROW_330_Left_683 ();
 TAPCELL_X1 PHY_EDGE_ROW_331_Left_684 ();
 TAPCELL_X1 PHY_EDGE_ROW_332_Left_685 ();
 TAPCELL_X1 PHY_EDGE_ROW_333_Left_686 ();
 TAPCELL_X1 PHY_EDGE_ROW_334_Left_687 ();
 TAPCELL_X1 PHY_EDGE_ROW_335_Left_688 ();
 TAPCELL_X1 PHY_EDGE_ROW_336_Left_689 ();
 TAPCELL_X1 PHY_EDGE_ROW_337_Left_690 ();
 TAPCELL_X1 PHY_EDGE_ROW_338_Left_691 ();
 TAPCELL_X1 PHY_EDGE_ROW_339_Left_692 ();
 TAPCELL_X1 PHY_EDGE_ROW_340_Left_693 ();
 TAPCELL_X1 PHY_EDGE_ROW_341_Left_694 ();
 TAPCELL_X1 PHY_EDGE_ROW_342_Left_695 ();
 TAPCELL_X1 PHY_EDGE_ROW_343_Left_696 ();
 TAPCELL_X1 PHY_EDGE_ROW_344_Left_697 ();
 TAPCELL_X1 PHY_EDGE_ROW_345_Left_698 ();
 TAPCELL_X1 PHY_EDGE_ROW_346_Left_699 ();
 TAPCELL_X1 PHY_EDGE_ROW_347_Left_700 ();
 TAPCELL_X1 PHY_EDGE_ROW_348_Left_701 ();
 TAPCELL_X1 PHY_EDGE_ROW_349_Left_702 ();
 TAPCELL_X1 PHY_EDGE_ROW_350_Left_703 ();
 TAPCELL_X1 PHY_EDGE_ROW_351_Left_704 ();
 TAPCELL_X1 PHY_EDGE_ROW_352_Left_705 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_706 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_707 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_708 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_709 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_710 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_711 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_712 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_713 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_714 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_715 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_716 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_717 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_718 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_719 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_720 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_721 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_722 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_723 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_724 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_725 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_726 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_727 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_728 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_729 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_730 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_731 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_732 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_733 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_734 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_735 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_736 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_737 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_738 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_739 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_740 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_741 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_742 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_743 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_744 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_745 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_746 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_747 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_748 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_749 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_750 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_751 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_752 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_753 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_754 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_755 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_756 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_757 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_758 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_759 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_760 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_761 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_762 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_763 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_764 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_765 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_766 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_767 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_768 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_769 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_770 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_771 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_772 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_773 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_774 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_775 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_776 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_777 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_778 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_779 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_780 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_781 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_782 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_783 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_784 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_785 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_786 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_787 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_788 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_789 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_41_790 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_41_791 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_792 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_793 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_43_794 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_43_795 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_796 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_797 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_45_798 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_45_799 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_800 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_801 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_47_802 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_47_803 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_804 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_805 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_49_806 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_49_807 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_808 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_809 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_810 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_811 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_812 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_813 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_53_814 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_53_815 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_816 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_817 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_55_818 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_55_819 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_820 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_821 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_57_822 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_57_823 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_824 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_825 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_59_826 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_59_827 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_828 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_829 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_61_830 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_61_831 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_832 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_833 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_63_834 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_63_835 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_836 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_837 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_65_838 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_65_839 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_840 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_841 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_67_842 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_67_843 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_844 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_845 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_846 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_847 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_848 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_849 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_71_850 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_71_851 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_852 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_853 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_73_854 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_73_855 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_856 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_857 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_75_858 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_75_859 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_860 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_861 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_77_862 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_77_863 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_864 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_865 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_79_866 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_79_867 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_868 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_869 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_81_870 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_81_871 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_872 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_873 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_83_874 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_83_875 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_876 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_877 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_85_878 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_85_879 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_880 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_881 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_87_882 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_87_883 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_884 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_885 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_89_886 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_89_887 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_888 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_889 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_91_890 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_91_891 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_892 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_893 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_93_894 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_93_895 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_896 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_897 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_95_898 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_95_899 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_900 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_901 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_97_902 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_97_903 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_904 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_905 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_99_906 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_99_907 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_908 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_909 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_101_910 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_101_911 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_912 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_913 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_103_914 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_103_915 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_916 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_917 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_105_918 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_105_919 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_920 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_921 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_107_922 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_107_923 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_924 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_925 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_109_926 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_109_927 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_928 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_929 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_111_930 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_111_931 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_932 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_933 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_113_934 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_113_935 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_936 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_937 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_115_938 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_115_939 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_940 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_941 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_117_942 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_117_943 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_944 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_945 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_119_946 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_119_947 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_948 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_949 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_121_950 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_121_951 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_952 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_953 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_123_954 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_123_955 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_956 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_957 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_125_958 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_125_959 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_960 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_961 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_127_962 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_127_963 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_964 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_965 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_129_966 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_129_967 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_968 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_969 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_131_970 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_131_971 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_972 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_973 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_133_974 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_133_975 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_976 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_977 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_135_978 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_135_979 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_980 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_981 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_137_982 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_137_983 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_984 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_985 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_139_986 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_139_987 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_988 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_989 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_141_990 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_141_991 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_992 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_993 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_143_994 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_143_995 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_996 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_997 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_145_998 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_145_999 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_1000 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_1001 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_147_1002 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_147_1003 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_1004 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_1005 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_149_1006 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_149_1007 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_1008 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_1009 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_151_1010 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_151_1011 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_1012 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_1013 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_153_1014 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_153_1015 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_1016 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_1017 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_155_1018 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_155_1019 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_156_1020 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_156_1021 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_157_1022 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_157_1023 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_158_1024 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_158_1025 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_159_1026 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_159_1027 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_160_1028 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_160_1029 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_161_1030 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_161_1031 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_162_1032 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_162_1033 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_163_1034 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_163_1035 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_164_1036 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_164_1037 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_165_1038 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_165_1039 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_166_1040 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_166_1041 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_167_1042 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_167_1043 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_168_1044 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_168_1045 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_169_1046 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_169_1047 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_170_1048 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_170_1049 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_171_1050 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_171_1051 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_172_1052 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_172_1053 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_173_1054 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_173_1055 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_174_1056 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_174_1057 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_175_1058 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_175_1059 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_176_1060 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_176_1061 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_177_1062 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_177_1063 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_178_1064 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_178_1065 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_179_1066 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_179_1067 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_180_1068 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_180_1069 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_181_1070 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_181_1071 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_182_1072 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_182_1073 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_183_1074 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_183_1075 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_184_1076 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_184_1077 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_185_1078 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_185_1079 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_186_1080 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_186_1081 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_187_1082 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_187_1083 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_188_1084 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_188_1085 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_189_1086 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_189_1087 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_190_1088 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_190_1089 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_191_1090 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_191_1091 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_192_1092 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_192_1093 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_193_1094 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_193_1095 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_194_1096 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_194_1097 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_195_1098 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_195_1099 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_196_1100 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_196_1101 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_197_1102 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_197_1103 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_198_1104 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_198_1105 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_199_1106 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_199_1107 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_200_1108 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_200_1109 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_201_1110 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_201_1111 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_202_1112 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_202_1113 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_203_1114 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_203_1115 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_204_1116 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_204_1117 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_205_1118 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_205_1119 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_206_1120 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_206_1121 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_207_1122 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_207_1123 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_1124 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_1125 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_209_1126 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_209_1127 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_210_1128 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_210_1129 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_211_1130 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_211_1131 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_212_1132 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_212_1133 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_213_1134 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_213_1135 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_214_1136 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_214_1137 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_215_1138 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_215_1139 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_216_1140 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_216_1141 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_217_1142 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_217_1143 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_218_1144 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_218_1145 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_219_1146 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_219_1147 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_220_1148 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_220_1149 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_221_1150 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_221_1151 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_222_1152 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_222_1153 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_223_1154 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_223_1155 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_224_1156 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_224_1157 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_225_1158 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_225_1159 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_226_1160 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_226_1161 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_227_1162 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_227_1163 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_228_1164 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_228_1165 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_229_1166 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_229_1167 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_230_1168 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_230_1169 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_231_1170 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_231_1171 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_232_1172 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_232_1173 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_233_1174 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_233_1175 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_234_1176 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_234_1177 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_235_1178 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_235_1179 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_236_1180 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_236_1181 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_237_1182 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_237_1183 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_238_1184 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_238_1185 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_239_1186 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_239_1187 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_240_1188 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_240_1189 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_241_1190 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_241_1191 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_242_1192 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_242_1193 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_243_1194 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_243_1195 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_244_1196 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_244_1197 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_245_1198 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_245_1199 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_246_1200 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_246_1201 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_247_1202 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_247_1203 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_248_1204 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_248_1205 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_249_1206 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_249_1207 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_250_1208 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_250_1209 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_251_1210 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_251_1211 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_252_1212 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_252_1213 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_253_1214 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_253_1215 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_254_1216 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_254_1217 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_255_1218 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_255_1219 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_256_1220 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_256_1221 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_257_1222 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_257_1223 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_258_1224 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_258_1225 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_259_1226 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_259_1227 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_260_1228 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_260_1229 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_261_1230 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_261_1231 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_262_1232 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_262_1233 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_263_1234 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_263_1235 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_264_1236 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_264_1237 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_265_1238 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_265_1239 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_266_1240 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_266_1241 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_267_1242 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_267_1243 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_268_1244 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_268_1245 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_269_1246 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_269_1247 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_270_1248 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_270_1249 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_271_1250 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_271_1251 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_272_1252 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_272_1253 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_273_1254 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_273_1255 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_274_1256 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_274_1257 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_275_1258 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_275_1259 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_276_1260 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_276_1261 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_277_1262 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_277_1263 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_278_1264 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_278_1265 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_279_1266 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_279_1267 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_280_1268 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_280_1269 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_281_1270 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_281_1271 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_282_1272 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_282_1273 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_283_1274 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_283_1275 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_284_1276 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_284_1277 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_285_1278 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_285_1279 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_286_1280 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_286_1281 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_287_1282 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_287_1283 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_288_1284 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_288_1285 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_289_1286 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_289_1287 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_290_1288 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_290_1289 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_291_1290 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_291_1291 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_292_1292 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_292_1293 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_293_1294 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_293_1295 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_294_1296 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_294_1297 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_295_1298 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_295_1299 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_296_1300 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_296_1301 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_297_1302 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_297_1303 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_298_1304 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_298_1305 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_299_1306 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_299_1307 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_300_1308 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_300_1309 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_301_1310 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_301_1311 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_302_1312 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_302_1313 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_303_1314 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_303_1315 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_304_1316 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_304_1317 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_305_1318 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_305_1319 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_306_1320 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_306_1321 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_307_1322 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_307_1323 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_308_1324 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_308_1325 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_309_1326 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_309_1327 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_310_1328 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_310_1329 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_311_1330 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_311_1331 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_312_1332 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_312_1333 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_313_1334 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_313_1335 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_314_1336 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_314_1337 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_315_1338 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_315_1339 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_316_1340 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_316_1341 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_317_1342 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_317_1343 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_318_1344 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_318_1345 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_319_1346 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_319_1347 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_320_1348 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_320_1349 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_321_1350 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_321_1351 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_322_1352 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_322_1353 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_323_1354 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_323_1355 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_324_1356 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_324_1357 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_325_1358 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_325_1359 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_326_1360 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_326_1361 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_327_1362 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_327_1363 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_328_1364 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_328_1365 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_329_1366 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_329_1367 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_330_1368 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_330_1369 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_331_1370 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_331_1371 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_332_1372 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_332_1373 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_333_1374 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_333_1375 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_334_1376 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_334_1377 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_335_1378 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_335_1379 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_336_1380 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_336_1381 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_337_1382 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_337_1383 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_338_1384 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_338_1385 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_339_1386 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_339_1387 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_340_1388 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_340_1389 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_341_1390 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_341_1391 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_342_1392 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_342_1393 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_343_1394 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_343_1395 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_344_1396 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_344_1397 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_345_1398 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_345_1399 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_346_1400 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_346_1401 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_347_1402 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_347_1403 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_348_1404 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_348_1405 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_349_1406 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_349_1407 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_350_1408 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_350_1409 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_351_1410 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_351_1411 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_352_1412 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_352_1413 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_352_1414 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_352_1415 ();
 BUF_X4 input1 (.A(rd_en),
    .Z(net1));
 BUF_X4 input2 (.A(rst_n),
    .Z(net2));
 BUF_X1 output3 (.A(net3),
    .Z(almost_empty));
 BUF_X1 output4 (.A(net4),
    .Z(almost_full));
 BUF_X1 output5 (.A(net5),
    .Z(data_count[0]));
 BUF_X1 output6 (.A(net6),
    .Z(data_count[1]));
 BUF_X1 output7 (.A(net7),
    .Z(data_count[2]));
 BUF_X1 output8 (.A(net8),
    .Z(data_count[3]));
 BUF_X1 output9 (.A(net9),
    .Z(data_count[4]));
 BUF_X1 output10 (.A(net10),
    .Z(empty));
 BUF_X1 output11 (.A(net11),
    .Z(full));
 BUF_X1 output12 (.A(net12),
    .Z(rd_data[0]));
 BUF_X1 output13 (.A(net13),
    .Z(rd_data[1]));
 BUF_X1 output14 (.A(net14),
    .Z(rd_data[2]));
 BUF_X1 output15 (.A(net15),
    .Z(rd_data[3]));
 BUF_X1 output16 (.A(net16),
    .Z(rd_data[4]));
 BUF_X1 output17 (.A(net17),
    .Z(rd_data[5]));
 BUF_X1 output18 (.A(net18),
    .Z(rd_data[6]));
 BUF_X1 output19 (.A(net19),
    .Z(rd_data[7]));
 BUF_X1 output20 (.A(net20),
    .Z(valid));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 CLKBUF_X3 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 CLKBUF_X3 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 CLKBUF_X3 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 CLKBUF_X3 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 CLKBUF_X3 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 CLKBUF_X3 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 CLKBUF_X3 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 CLKBUF_X3 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 CLKBUF_X3 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 CLKBUF_X3 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 CLKBUF_X3 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 CLKBUF_X3 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 CLKBUF_X3 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 CLKBUF_X3 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 CLKBUF_X3 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 INV_X4 clkload0 (.A(clknet_4_0_0_clk));
 INV_X4 clkload1 (.A(clknet_4_1_0_clk));
 INV_X2 clkload2 (.A(clknet_4_2_0_clk));
 INV_X2 clkload3 (.A(clknet_4_3_0_clk));
 INV_X4 clkload4 (.A(clknet_4_4_0_clk));
 INV_X2 clkload5 (.A(clknet_4_5_0_clk));
 INV_X2 clkload6 (.A(clknet_4_6_0_clk));
 INV_X1 clkload7 (.A(clknet_4_7_0_clk));
 INV_X2 clkload8 (.A(clknet_4_9_0_clk));
 INV_X2 clkload9 (.A(clknet_4_12_0_clk));
 CLKBUF_X1 clkload10 (.A(clknet_4_14_0_clk));
 INV_X2 clkload11 (.A(clknet_4_15_0_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_193 ();
 FILLCELL_X32 FILLER_0_225 ();
 FILLCELL_X32 FILLER_0_257 ();
 FILLCELL_X32 FILLER_0_289 ();
 FILLCELL_X32 FILLER_0_321 ();
 FILLCELL_X32 FILLER_0_353 ();
 FILLCELL_X32 FILLER_0_385 ();
 FILLCELL_X32 FILLER_0_417 ();
 FILLCELL_X32 FILLER_0_449 ();
 FILLCELL_X32 FILLER_0_481 ();
 FILLCELL_X32 FILLER_0_513 ();
 FILLCELL_X32 FILLER_0_545 ();
 FILLCELL_X32 FILLER_0_577 ();
 FILLCELL_X16 FILLER_0_609 ();
 FILLCELL_X4 FILLER_0_625 ();
 FILLCELL_X2 FILLER_0_629 ();
 FILLCELL_X32 FILLER_0_632 ();
 FILLCELL_X32 FILLER_0_664 ();
 FILLCELL_X32 FILLER_0_696 ();
 FILLCELL_X32 FILLER_0_728 ();
 FILLCELL_X32 FILLER_0_760 ();
 FILLCELL_X32 FILLER_0_792 ();
 FILLCELL_X32 FILLER_0_824 ();
 FILLCELL_X32 FILLER_0_856 ();
 FILLCELL_X32 FILLER_0_888 ();
 FILLCELL_X32 FILLER_0_920 ();
 FILLCELL_X32 FILLER_0_952 ();
 FILLCELL_X32 FILLER_0_984 ();
 FILLCELL_X32 FILLER_0_1016 ();
 FILLCELL_X32 FILLER_0_1048 ();
 FILLCELL_X32 FILLER_0_1080 ();
 FILLCELL_X32 FILLER_0_1112 ();
 FILLCELL_X32 FILLER_0_1144 ();
 FILLCELL_X32 FILLER_0_1176 ();
 FILLCELL_X32 FILLER_0_1208 ();
 FILLCELL_X16 FILLER_0_1240 ();
 FILLCELL_X4 FILLER_0_1256 ();
 FILLCELL_X2 FILLER_0_1260 ();
 FILLCELL_X32 FILLER_0_1263 ();
 FILLCELL_X32 FILLER_0_1295 ();
 FILLCELL_X32 FILLER_0_1327 ();
 FILLCELL_X32 FILLER_0_1359 ();
 FILLCELL_X32 FILLER_0_1391 ();
 FILLCELL_X32 FILLER_0_1423 ();
 FILLCELL_X32 FILLER_0_1455 ();
 FILLCELL_X32 FILLER_0_1487 ();
 FILLCELL_X32 FILLER_0_1519 ();
 FILLCELL_X32 FILLER_0_1551 ();
 FILLCELL_X32 FILLER_0_1583 ();
 FILLCELL_X32 FILLER_0_1615 ();
 FILLCELL_X32 FILLER_0_1647 ();
 FILLCELL_X32 FILLER_0_1679 ();
 FILLCELL_X32 FILLER_0_1711 ();
 FILLCELL_X32 FILLER_0_1743 ();
 FILLCELL_X32 FILLER_0_1775 ();
 FILLCELL_X32 FILLER_0_1807 ();
 FILLCELL_X32 FILLER_0_1839 ();
 FILLCELL_X16 FILLER_0_1871 ();
 FILLCELL_X4 FILLER_0_1887 ();
 FILLCELL_X2 FILLER_0_1891 ();
 FILLCELL_X32 FILLER_0_1894 ();
 FILLCELL_X32 FILLER_0_1926 ();
 FILLCELL_X32 FILLER_0_1958 ();
 FILLCELL_X32 FILLER_0_1990 ();
 FILLCELL_X32 FILLER_0_2022 ();
 FILLCELL_X32 FILLER_0_2054 ();
 FILLCELL_X32 FILLER_0_2086 ();
 FILLCELL_X32 FILLER_0_2118 ();
 FILLCELL_X32 FILLER_0_2150 ();
 FILLCELL_X32 FILLER_0_2182 ();
 FILLCELL_X32 FILLER_0_2214 ();
 FILLCELL_X32 FILLER_0_2246 ();
 FILLCELL_X32 FILLER_0_2278 ();
 FILLCELL_X32 FILLER_0_2310 ();
 FILLCELL_X32 FILLER_0_2342 ();
 FILLCELL_X32 FILLER_0_2374 ();
 FILLCELL_X32 FILLER_0_2406 ();
 FILLCELL_X32 FILLER_0_2438 ();
 FILLCELL_X32 FILLER_0_2470 ();
 FILLCELL_X16 FILLER_0_2502 ();
 FILLCELL_X4 FILLER_0_2518 ();
 FILLCELL_X2 FILLER_0_2522 ();
 FILLCELL_X32 FILLER_0_2525 ();
 FILLCELL_X32 FILLER_0_2557 ();
 FILLCELL_X8 FILLER_0_2589 ();
 FILLCELL_X4 FILLER_0_2597 ();
 FILLCELL_X1 FILLER_0_2601 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X32 FILLER_1_289 ();
 FILLCELL_X32 FILLER_1_321 ();
 FILLCELL_X32 FILLER_1_353 ();
 FILLCELL_X32 FILLER_1_385 ();
 FILLCELL_X32 FILLER_1_417 ();
 FILLCELL_X32 FILLER_1_449 ();
 FILLCELL_X32 FILLER_1_481 ();
 FILLCELL_X32 FILLER_1_513 ();
 FILLCELL_X32 FILLER_1_545 ();
 FILLCELL_X32 FILLER_1_577 ();
 FILLCELL_X32 FILLER_1_609 ();
 FILLCELL_X32 FILLER_1_641 ();
 FILLCELL_X32 FILLER_1_673 ();
 FILLCELL_X32 FILLER_1_705 ();
 FILLCELL_X32 FILLER_1_737 ();
 FILLCELL_X32 FILLER_1_769 ();
 FILLCELL_X32 FILLER_1_801 ();
 FILLCELL_X32 FILLER_1_833 ();
 FILLCELL_X32 FILLER_1_865 ();
 FILLCELL_X32 FILLER_1_897 ();
 FILLCELL_X32 FILLER_1_929 ();
 FILLCELL_X32 FILLER_1_961 ();
 FILLCELL_X32 FILLER_1_993 ();
 FILLCELL_X32 FILLER_1_1025 ();
 FILLCELL_X32 FILLER_1_1057 ();
 FILLCELL_X32 FILLER_1_1089 ();
 FILLCELL_X32 FILLER_1_1121 ();
 FILLCELL_X32 FILLER_1_1153 ();
 FILLCELL_X32 FILLER_1_1185 ();
 FILLCELL_X32 FILLER_1_1217 ();
 FILLCELL_X8 FILLER_1_1249 ();
 FILLCELL_X4 FILLER_1_1257 ();
 FILLCELL_X2 FILLER_1_1261 ();
 FILLCELL_X32 FILLER_1_1264 ();
 FILLCELL_X32 FILLER_1_1296 ();
 FILLCELL_X32 FILLER_1_1328 ();
 FILLCELL_X32 FILLER_1_1360 ();
 FILLCELL_X32 FILLER_1_1392 ();
 FILLCELL_X32 FILLER_1_1424 ();
 FILLCELL_X32 FILLER_1_1456 ();
 FILLCELL_X32 FILLER_1_1488 ();
 FILLCELL_X32 FILLER_1_1520 ();
 FILLCELL_X32 FILLER_1_1552 ();
 FILLCELL_X32 FILLER_1_1584 ();
 FILLCELL_X32 FILLER_1_1616 ();
 FILLCELL_X32 FILLER_1_1648 ();
 FILLCELL_X32 FILLER_1_1680 ();
 FILLCELL_X32 FILLER_1_1712 ();
 FILLCELL_X32 FILLER_1_1744 ();
 FILLCELL_X32 FILLER_1_1776 ();
 FILLCELL_X32 FILLER_1_1808 ();
 FILLCELL_X32 FILLER_1_1840 ();
 FILLCELL_X32 FILLER_1_1872 ();
 FILLCELL_X32 FILLER_1_1904 ();
 FILLCELL_X32 FILLER_1_1936 ();
 FILLCELL_X32 FILLER_1_1968 ();
 FILLCELL_X32 FILLER_1_2000 ();
 FILLCELL_X32 FILLER_1_2032 ();
 FILLCELL_X32 FILLER_1_2064 ();
 FILLCELL_X32 FILLER_1_2096 ();
 FILLCELL_X32 FILLER_1_2128 ();
 FILLCELL_X32 FILLER_1_2160 ();
 FILLCELL_X32 FILLER_1_2192 ();
 FILLCELL_X32 FILLER_1_2224 ();
 FILLCELL_X32 FILLER_1_2256 ();
 FILLCELL_X32 FILLER_1_2288 ();
 FILLCELL_X32 FILLER_1_2320 ();
 FILLCELL_X32 FILLER_1_2352 ();
 FILLCELL_X32 FILLER_1_2384 ();
 FILLCELL_X32 FILLER_1_2416 ();
 FILLCELL_X32 FILLER_1_2448 ();
 FILLCELL_X32 FILLER_1_2480 ();
 FILLCELL_X8 FILLER_1_2512 ();
 FILLCELL_X4 FILLER_1_2520 ();
 FILLCELL_X2 FILLER_1_2524 ();
 FILLCELL_X32 FILLER_1_2527 ();
 FILLCELL_X32 FILLER_1_2559 ();
 FILLCELL_X8 FILLER_1_2591 ();
 FILLCELL_X2 FILLER_1_2599 ();
 FILLCELL_X1 FILLER_1_2601 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X32 FILLER_2_321 ();
 FILLCELL_X32 FILLER_2_353 ();
 FILLCELL_X32 FILLER_2_385 ();
 FILLCELL_X32 FILLER_2_417 ();
 FILLCELL_X32 FILLER_2_449 ();
 FILLCELL_X32 FILLER_2_481 ();
 FILLCELL_X32 FILLER_2_513 ();
 FILLCELL_X32 FILLER_2_545 ();
 FILLCELL_X32 FILLER_2_577 ();
 FILLCELL_X16 FILLER_2_609 ();
 FILLCELL_X4 FILLER_2_625 ();
 FILLCELL_X2 FILLER_2_629 ();
 FILLCELL_X32 FILLER_2_632 ();
 FILLCELL_X32 FILLER_2_664 ();
 FILLCELL_X32 FILLER_2_696 ();
 FILLCELL_X32 FILLER_2_728 ();
 FILLCELL_X32 FILLER_2_760 ();
 FILLCELL_X32 FILLER_2_792 ();
 FILLCELL_X32 FILLER_2_824 ();
 FILLCELL_X32 FILLER_2_856 ();
 FILLCELL_X32 FILLER_2_888 ();
 FILLCELL_X32 FILLER_2_920 ();
 FILLCELL_X32 FILLER_2_952 ();
 FILLCELL_X32 FILLER_2_984 ();
 FILLCELL_X32 FILLER_2_1016 ();
 FILLCELL_X32 FILLER_2_1048 ();
 FILLCELL_X32 FILLER_2_1080 ();
 FILLCELL_X32 FILLER_2_1112 ();
 FILLCELL_X32 FILLER_2_1144 ();
 FILLCELL_X32 FILLER_2_1176 ();
 FILLCELL_X32 FILLER_2_1208 ();
 FILLCELL_X32 FILLER_2_1240 ();
 FILLCELL_X32 FILLER_2_1272 ();
 FILLCELL_X32 FILLER_2_1304 ();
 FILLCELL_X32 FILLER_2_1336 ();
 FILLCELL_X32 FILLER_2_1368 ();
 FILLCELL_X32 FILLER_2_1400 ();
 FILLCELL_X32 FILLER_2_1432 ();
 FILLCELL_X32 FILLER_2_1464 ();
 FILLCELL_X32 FILLER_2_1496 ();
 FILLCELL_X32 FILLER_2_1528 ();
 FILLCELL_X32 FILLER_2_1560 ();
 FILLCELL_X32 FILLER_2_1592 ();
 FILLCELL_X32 FILLER_2_1624 ();
 FILLCELL_X32 FILLER_2_1656 ();
 FILLCELL_X32 FILLER_2_1688 ();
 FILLCELL_X32 FILLER_2_1720 ();
 FILLCELL_X32 FILLER_2_1752 ();
 FILLCELL_X32 FILLER_2_1784 ();
 FILLCELL_X32 FILLER_2_1816 ();
 FILLCELL_X32 FILLER_2_1848 ();
 FILLCELL_X8 FILLER_2_1880 ();
 FILLCELL_X4 FILLER_2_1888 ();
 FILLCELL_X2 FILLER_2_1892 ();
 FILLCELL_X32 FILLER_2_1895 ();
 FILLCELL_X32 FILLER_2_1927 ();
 FILLCELL_X32 FILLER_2_1959 ();
 FILLCELL_X32 FILLER_2_1991 ();
 FILLCELL_X32 FILLER_2_2023 ();
 FILLCELL_X32 FILLER_2_2055 ();
 FILLCELL_X32 FILLER_2_2087 ();
 FILLCELL_X32 FILLER_2_2119 ();
 FILLCELL_X32 FILLER_2_2151 ();
 FILLCELL_X32 FILLER_2_2183 ();
 FILLCELL_X32 FILLER_2_2215 ();
 FILLCELL_X32 FILLER_2_2247 ();
 FILLCELL_X32 FILLER_2_2279 ();
 FILLCELL_X32 FILLER_2_2311 ();
 FILLCELL_X32 FILLER_2_2343 ();
 FILLCELL_X32 FILLER_2_2375 ();
 FILLCELL_X32 FILLER_2_2407 ();
 FILLCELL_X32 FILLER_2_2439 ();
 FILLCELL_X32 FILLER_2_2471 ();
 FILLCELL_X32 FILLER_2_2503 ();
 FILLCELL_X32 FILLER_2_2535 ();
 FILLCELL_X32 FILLER_2_2567 ();
 FILLCELL_X2 FILLER_2_2599 ();
 FILLCELL_X1 FILLER_2_2601 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X32 FILLER_3_321 ();
 FILLCELL_X32 FILLER_3_353 ();
 FILLCELL_X32 FILLER_3_385 ();
 FILLCELL_X32 FILLER_3_417 ();
 FILLCELL_X32 FILLER_3_449 ();
 FILLCELL_X32 FILLER_3_481 ();
 FILLCELL_X32 FILLER_3_513 ();
 FILLCELL_X32 FILLER_3_545 ();
 FILLCELL_X32 FILLER_3_577 ();
 FILLCELL_X32 FILLER_3_609 ();
 FILLCELL_X32 FILLER_3_641 ();
 FILLCELL_X32 FILLER_3_673 ();
 FILLCELL_X32 FILLER_3_705 ();
 FILLCELL_X32 FILLER_3_737 ();
 FILLCELL_X32 FILLER_3_769 ();
 FILLCELL_X32 FILLER_3_801 ();
 FILLCELL_X32 FILLER_3_833 ();
 FILLCELL_X32 FILLER_3_865 ();
 FILLCELL_X32 FILLER_3_897 ();
 FILLCELL_X32 FILLER_3_929 ();
 FILLCELL_X32 FILLER_3_961 ();
 FILLCELL_X32 FILLER_3_993 ();
 FILLCELL_X32 FILLER_3_1025 ();
 FILLCELL_X32 FILLER_3_1057 ();
 FILLCELL_X32 FILLER_3_1089 ();
 FILLCELL_X32 FILLER_3_1121 ();
 FILLCELL_X32 FILLER_3_1153 ();
 FILLCELL_X32 FILLER_3_1185 ();
 FILLCELL_X32 FILLER_3_1217 ();
 FILLCELL_X8 FILLER_3_1249 ();
 FILLCELL_X4 FILLER_3_1257 ();
 FILLCELL_X2 FILLER_3_1261 ();
 FILLCELL_X32 FILLER_3_1264 ();
 FILLCELL_X32 FILLER_3_1296 ();
 FILLCELL_X32 FILLER_3_1328 ();
 FILLCELL_X32 FILLER_3_1360 ();
 FILLCELL_X32 FILLER_3_1392 ();
 FILLCELL_X32 FILLER_3_1424 ();
 FILLCELL_X32 FILLER_3_1456 ();
 FILLCELL_X32 FILLER_3_1488 ();
 FILLCELL_X32 FILLER_3_1520 ();
 FILLCELL_X32 FILLER_3_1552 ();
 FILLCELL_X32 FILLER_3_1584 ();
 FILLCELL_X32 FILLER_3_1616 ();
 FILLCELL_X32 FILLER_3_1648 ();
 FILLCELL_X32 FILLER_3_1680 ();
 FILLCELL_X32 FILLER_3_1712 ();
 FILLCELL_X32 FILLER_3_1744 ();
 FILLCELL_X32 FILLER_3_1776 ();
 FILLCELL_X32 FILLER_3_1808 ();
 FILLCELL_X32 FILLER_3_1840 ();
 FILLCELL_X32 FILLER_3_1872 ();
 FILLCELL_X32 FILLER_3_1904 ();
 FILLCELL_X32 FILLER_3_1936 ();
 FILLCELL_X32 FILLER_3_1968 ();
 FILLCELL_X32 FILLER_3_2000 ();
 FILLCELL_X32 FILLER_3_2032 ();
 FILLCELL_X32 FILLER_3_2064 ();
 FILLCELL_X32 FILLER_3_2096 ();
 FILLCELL_X32 FILLER_3_2128 ();
 FILLCELL_X32 FILLER_3_2160 ();
 FILLCELL_X32 FILLER_3_2192 ();
 FILLCELL_X32 FILLER_3_2224 ();
 FILLCELL_X32 FILLER_3_2256 ();
 FILLCELL_X32 FILLER_3_2288 ();
 FILLCELL_X32 FILLER_3_2320 ();
 FILLCELL_X32 FILLER_3_2352 ();
 FILLCELL_X32 FILLER_3_2384 ();
 FILLCELL_X32 FILLER_3_2416 ();
 FILLCELL_X32 FILLER_3_2448 ();
 FILLCELL_X32 FILLER_3_2480 ();
 FILLCELL_X8 FILLER_3_2512 ();
 FILLCELL_X4 FILLER_3_2520 ();
 FILLCELL_X2 FILLER_3_2524 ();
 FILLCELL_X32 FILLER_3_2527 ();
 FILLCELL_X32 FILLER_3_2559 ();
 FILLCELL_X8 FILLER_3_2591 ();
 FILLCELL_X2 FILLER_3_2599 ();
 FILLCELL_X1 FILLER_3_2601 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X32 FILLER_4_321 ();
 FILLCELL_X32 FILLER_4_353 ();
 FILLCELL_X32 FILLER_4_385 ();
 FILLCELL_X32 FILLER_4_417 ();
 FILLCELL_X32 FILLER_4_449 ();
 FILLCELL_X32 FILLER_4_481 ();
 FILLCELL_X32 FILLER_4_513 ();
 FILLCELL_X32 FILLER_4_545 ();
 FILLCELL_X32 FILLER_4_577 ();
 FILLCELL_X16 FILLER_4_609 ();
 FILLCELL_X4 FILLER_4_625 ();
 FILLCELL_X2 FILLER_4_629 ();
 FILLCELL_X32 FILLER_4_632 ();
 FILLCELL_X32 FILLER_4_664 ();
 FILLCELL_X32 FILLER_4_696 ();
 FILLCELL_X32 FILLER_4_728 ();
 FILLCELL_X32 FILLER_4_760 ();
 FILLCELL_X32 FILLER_4_792 ();
 FILLCELL_X32 FILLER_4_824 ();
 FILLCELL_X32 FILLER_4_856 ();
 FILLCELL_X32 FILLER_4_888 ();
 FILLCELL_X32 FILLER_4_920 ();
 FILLCELL_X32 FILLER_4_952 ();
 FILLCELL_X32 FILLER_4_984 ();
 FILLCELL_X32 FILLER_4_1016 ();
 FILLCELL_X32 FILLER_4_1048 ();
 FILLCELL_X32 FILLER_4_1080 ();
 FILLCELL_X32 FILLER_4_1112 ();
 FILLCELL_X32 FILLER_4_1144 ();
 FILLCELL_X32 FILLER_4_1176 ();
 FILLCELL_X32 FILLER_4_1208 ();
 FILLCELL_X32 FILLER_4_1240 ();
 FILLCELL_X32 FILLER_4_1272 ();
 FILLCELL_X32 FILLER_4_1304 ();
 FILLCELL_X32 FILLER_4_1336 ();
 FILLCELL_X32 FILLER_4_1368 ();
 FILLCELL_X32 FILLER_4_1400 ();
 FILLCELL_X32 FILLER_4_1432 ();
 FILLCELL_X32 FILLER_4_1464 ();
 FILLCELL_X32 FILLER_4_1496 ();
 FILLCELL_X32 FILLER_4_1528 ();
 FILLCELL_X32 FILLER_4_1560 ();
 FILLCELL_X32 FILLER_4_1592 ();
 FILLCELL_X32 FILLER_4_1624 ();
 FILLCELL_X32 FILLER_4_1656 ();
 FILLCELL_X32 FILLER_4_1688 ();
 FILLCELL_X32 FILLER_4_1720 ();
 FILLCELL_X32 FILLER_4_1752 ();
 FILLCELL_X32 FILLER_4_1784 ();
 FILLCELL_X32 FILLER_4_1816 ();
 FILLCELL_X32 FILLER_4_1848 ();
 FILLCELL_X8 FILLER_4_1880 ();
 FILLCELL_X4 FILLER_4_1888 ();
 FILLCELL_X2 FILLER_4_1892 ();
 FILLCELL_X32 FILLER_4_1895 ();
 FILLCELL_X32 FILLER_4_1927 ();
 FILLCELL_X32 FILLER_4_1959 ();
 FILLCELL_X32 FILLER_4_1991 ();
 FILLCELL_X32 FILLER_4_2023 ();
 FILLCELL_X32 FILLER_4_2055 ();
 FILLCELL_X32 FILLER_4_2087 ();
 FILLCELL_X32 FILLER_4_2119 ();
 FILLCELL_X32 FILLER_4_2151 ();
 FILLCELL_X32 FILLER_4_2183 ();
 FILLCELL_X32 FILLER_4_2215 ();
 FILLCELL_X32 FILLER_4_2247 ();
 FILLCELL_X32 FILLER_4_2279 ();
 FILLCELL_X32 FILLER_4_2311 ();
 FILLCELL_X32 FILLER_4_2343 ();
 FILLCELL_X32 FILLER_4_2375 ();
 FILLCELL_X32 FILLER_4_2407 ();
 FILLCELL_X32 FILLER_4_2439 ();
 FILLCELL_X32 FILLER_4_2471 ();
 FILLCELL_X32 FILLER_4_2503 ();
 FILLCELL_X32 FILLER_4_2535 ();
 FILLCELL_X32 FILLER_4_2567 ();
 FILLCELL_X2 FILLER_4_2599 ();
 FILLCELL_X1 FILLER_4_2601 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X32 FILLER_5_321 ();
 FILLCELL_X32 FILLER_5_353 ();
 FILLCELL_X32 FILLER_5_385 ();
 FILLCELL_X32 FILLER_5_417 ();
 FILLCELL_X32 FILLER_5_449 ();
 FILLCELL_X32 FILLER_5_481 ();
 FILLCELL_X32 FILLER_5_513 ();
 FILLCELL_X32 FILLER_5_545 ();
 FILLCELL_X32 FILLER_5_577 ();
 FILLCELL_X32 FILLER_5_609 ();
 FILLCELL_X32 FILLER_5_641 ();
 FILLCELL_X32 FILLER_5_673 ();
 FILLCELL_X32 FILLER_5_705 ();
 FILLCELL_X32 FILLER_5_737 ();
 FILLCELL_X32 FILLER_5_769 ();
 FILLCELL_X32 FILLER_5_801 ();
 FILLCELL_X32 FILLER_5_833 ();
 FILLCELL_X32 FILLER_5_865 ();
 FILLCELL_X32 FILLER_5_897 ();
 FILLCELL_X32 FILLER_5_929 ();
 FILLCELL_X32 FILLER_5_961 ();
 FILLCELL_X32 FILLER_5_993 ();
 FILLCELL_X32 FILLER_5_1025 ();
 FILLCELL_X32 FILLER_5_1057 ();
 FILLCELL_X32 FILLER_5_1089 ();
 FILLCELL_X32 FILLER_5_1121 ();
 FILLCELL_X32 FILLER_5_1153 ();
 FILLCELL_X32 FILLER_5_1185 ();
 FILLCELL_X32 FILLER_5_1217 ();
 FILLCELL_X8 FILLER_5_1249 ();
 FILLCELL_X4 FILLER_5_1257 ();
 FILLCELL_X2 FILLER_5_1261 ();
 FILLCELL_X32 FILLER_5_1264 ();
 FILLCELL_X32 FILLER_5_1296 ();
 FILLCELL_X32 FILLER_5_1328 ();
 FILLCELL_X32 FILLER_5_1360 ();
 FILLCELL_X32 FILLER_5_1392 ();
 FILLCELL_X32 FILLER_5_1424 ();
 FILLCELL_X32 FILLER_5_1456 ();
 FILLCELL_X32 FILLER_5_1488 ();
 FILLCELL_X32 FILLER_5_1520 ();
 FILLCELL_X32 FILLER_5_1552 ();
 FILLCELL_X32 FILLER_5_1584 ();
 FILLCELL_X32 FILLER_5_1616 ();
 FILLCELL_X32 FILLER_5_1648 ();
 FILLCELL_X32 FILLER_5_1680 ();
 FILLCELL_X32 FILLER_5_1712 ();
 FILLCELL_X32 FILLER_5_1744 ();
 FILLCELL_X32 FILLER_5_1776 ();
 FILLCELL_X32 FILLER_5_1808 ();
 FILLCELL_X32 FILLER_5_1840 ();
 FILLCELL_X32 FILLER_5_1872 ();
 FILLCELL_X32 FILLER_5_1904 ();
 FILLCELL_X32 FILLER_5_1936 ();
 FILLCELL_X32 FILLER_5_1968 ();
 FILLCELL_X32 FILLER_5_2000 ();
 FILLCELL_X32 FILLER_5_2032 ();
 FILLCELL_X32 FILLER_5_2064 ();
 FILLCELL_X32 FILLER_5_2096 ();
 FILLCELL_X32 FILLER_5_2128 ();
 FILLCELL_X32 FILLER_5_2160 ();
 FILLCELL_X32 FILLER_5_2192 ();
 FILLCELL_X32 FILLER_5_2224 ();
 FILLCELL_X32 FILLER_5_2256 ();
 FILLCELL_X32 FILLER_5_2288 ();
 FILLCELL_X32 FILLER_5_2320 ();
 FILLCELL_X32 FILLER_5_2352 ();
 FILLCELL_X32 FILLER_5_2384 ();
 FILLCELL_X32 FILLER_5_2416 ();
 FILLCELL_X32 FILLER_5_2448 ();
 FILLCELL_X32 FILLER_5_2480 ();
 FILLCELL_X8 FILLER_5_2512 ();
 FILLCELL_X4 FILLER_5_2520 ();
 FILLCELL_X2 FILLER_5_2524 ();
 FILLCELL_X32 FILLER_5_2527 ();
 FILLCELL_X32 FILLER_5_2559 ();
 FILLCELL_X8 FILLER_5_2591 ();
 FILLCELL_X2 FILLER_5_2599 ();
 FILLCELL_X1 FILLER_5_2601 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X32 FILLER_6_257 ();
 FILLCELL_X32 FILLER_6_289 ();
 FILLCELL_X32 FILLER_6_321 ();
 FILLCELL_X32 FILLER_6_353 ();
 FILLCELL_X32 FILLER_6_385 ();
 FILLCELL_X32 FILLER_6_417 ();
 FILLCELL_X32 FILLER_6_449 ();
 FILLCELL_X32 FILLER_6_481 ();
 FILLCELL_X32 FILLER_6_513 ();
 FILLCELL_X32 FILLER_6_545 ();
 FILLCELL_X32 FILLER_6_577 ();
 FILLCELL_X16 FILLER_6_609 ();
 FILLCELL_X4 FILLER_6_625 ();
 FILLCELL_X2 FILLER_6_629 ();
 FILLCELL_X32 FILLER_6_632 ();
 FILLCELL_X32 FILLER_6_664 ();
 FILLCELL_X32 FILLER_6_696 ();
 FILLCELL_X32 FILLER_6_728 ();
 FILLCELL_X32 FILLER_6_760 ();
 FILLCELL_X32 FILLER_6_792 ();
 FILLCELL_X32 FILLER_6_824 ();
 FILLCELL_X32 FILLER_6_856 ();
 FILLCELL_X32 FILLER_6_888 ();
 FILLCELL_X32 FILLER_6_920 ();
 FILLCELL_X32 FILLER_6_952 ();
 FILLCELL_X32 FILLER_6_984 ();
 FILLCELL_X32 FILLER_6_1016 ();
 FILLCELL_X32 FILLER_6_1048 ();
 FILLCELL_X32 FILLER_6_1080 ();
 FILLCELL_X32 FILLER_6_1112 ();
 FILLCELL_X32 FILLER_6_1144 ();
 FILLCELL_X32 FILLER_6_1176 ();
 FILLCELL_X32 FILLER_6_1208 ();
 FILLCELL_X32 FILLER_6_1240 ();
 FILLCELL_X32 FILLER_6_1272 ();
 FILLCELL_X32 FILLER_6_1304 ();
 FILLCELL_X32 FILLER_6_1336 ();
 FILLCELL_X32 FILLER_6_1368 ();
 FILLCELL_X32 FILLER_6_1400 ();
 FILLCELL_X32 FILLER_6_1432 ();
 FILLCELL_X32 FILLER_6_1464 ();
 FILLCELL_X32 FILLER_6_1496 ();
 FILLCELL_X32 FILLER_6_1528 ();
 FILLCELL_X32 FILLER_6_1560 ();
 FILLCELL_X32 FILLER_6_1592 ();
 FILLCELL_X32 FILLER_6_1624 ();
 FILLCELL_X32 FILLER_6_1656 ();
 FILLCELL_X32 FILLER_6_1688 ();
 FILLCELL_X32 FILLER_6_1720 ();
 FILLCELL_X32 FILLER_6_1752 ();
 FILLCELL_X32 FILLER_6_1784 ();
 FILLCELL_X32 FILLER_6_1816 ();
 FILLCELL_X32 FILLER_6_1848 ();
 FILLCELL_X8 FILLER_6_1880 ();
 FILLCELL_X4 FILLER_6_1888 ();
 FILLCELL_X2 FILLER_6_1892 ();
 FILLCELL_X32 FILLER_6_1895 ();
 FILLCELL_X32 FILLER_6_1927 ();
 FILLCELL_X32 FILLER_6_1959 ();
 FILLCELL_X32 FILLER_6_1991 ();
 FILLCELL_X32 FILLER_6_2023 ();
 FILLCELL_X32 FILLER_6_2055 ();
 FILLCELL_X32 FILLER_6_2087 ();
 FILLCELL_X32 FILLER_6_2119 ();
 FILLCELL_X32 FILLER_6_2151 ();
 FILLCELL_X32 FILLER_6_2183 ();
 FILLCELL_X32 FILLER_6_2215 ();
 FILLCELL_X32 FILLER_6_2247 ();
 FILLCELL_X32 FILLER_6_2279 ();
 FILLCELL_X32 FILLER_6_2311 ();
 FILLCELL_X32 FILLER_6_2343 ();
 FILLCELL_X32 FILLER_6_2375 ();
 FILLCELL_X32 FILLER_6_2407 ();
 FILLCELL_X32 FILLER_6_2439 ();
 FILLCELL_X32 FILLER_6_2471 ();
 FILLCELL_X32 FILLER_6_2503 ();
 FILLCELL_X32 FILLER_6_2535 ();
 FILLCELL_X32 FILLER_6_2567 ();
 FILLCELL_X2 FILLER_6_2599 ();
 FILLCELL_X1 FILLER_6_2601 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X32 FILLER_7_257 ();
 FILLCELL_X32 FILLER_7_289 ();
 FILLCELL_X32 FILLER_7_321 ();
 FILLCELL_X32 FILLER_7_353 ();
 FILLCELL_X32 FILLER_7_385 ();
 FILLCELL_X32 FILLER_7_417 ();
 FILLCELL_X32 FILLER_7_449 ();
 FILLCELL_X32 FILLER_7_481 ();
 FILLCELL_X32 FILLER_7_513 ();
 FILLCELL_X32 FILLER_7_545 ();
 FILLCELL_X32 FILLER_7_577 ();
 FILLCELL_X32 FILLER_7_609 ();
 FILLCELL_X32 FILLER_7_641 ();
 FILLCELL_X32 FILLER_7_673 ();
 FILLCELL_X32 FILLER_7_705 ();
 FILLCELL_X32 FILLER_7_737 ();
 FILLCELL_X32 FILLER_7_769 ();
 FILLCELL_X32 FILLER_7_801 ();
 FILLCELL_X32 FILLER_7_833 ();
 FILLCELL_X32 FILLER_7_865 ();
 FILLCELL_X32 FILLER_7_897 ();
 FILLCELL_X32 FILLER_7_929 ();
 FILLCELL_X32 FILLER_7_961 ();
 FILLCELL_X32 FILLER_7_993 ();
 FILLCELL_X32 FILLER_7_1025 ();
 FILLCELL_X32 FILLER_7_1057 ();
 FILLCELL_X32 FILLER_7_1089 ();
 FILLCELL_X32 FILLER_7_1121 ();
 FILLCELL_X32 FILLER_7_1153 ();
 FILLCELL_X32 FILLER_7_1185 ();
 FILLCELL_X32 FILLER_7_1217 ();
 FILLCELL_X8 FILLER_7_1249 ();
 FILLCELL_X4 FILLER_7_1257 ();
 FILLCELL_X2 FILLER_7_1261 ();
 FILLCELL_X32 FILLER_7_1264 ();
 FILLCELL_X32 FILLER_7_1296 ();
 FILLCELL_X32 FILLER_7_1328 ();
 FILLCELL_X32 FILLER_7_1360 ();
 FILLCELL_X32 FILLER_7_1392 ();
 FILLCELL_X32 FILLER_7_1424 ();
 FILLCELL_X32 FILLER_7_1456 ();
 FILLCELL_X32 FILLER_7_1488 ();
 FILLCELL_X32 FILLER_7_1520 ();
 FILLCELL_X32 FILLER_7_1552 ();
 FILLCELL_X32 FILLER_7_1584 ();
 FILLCELL_X32 FILLER_7_1616 ();
 FILLCELL_X32 FILLER_7_1648 ();
 FILLCELL_X32 FILLER_7_1680 ();
 FILLCELL_X32 FILLER_7_1712 ();
 FILLCELL_X32 FILLER_7_1744 ();
 FILLCELL_X32 FILLER_7_1776 ();
 FILLCELL_X32 FILLER_7_1808 ();
 FILLCELL_X32 FILLER_7_1840 ();
 FILLCELL_X32 FILLER_7_1872 ();
 FILLCELL_X32 FILLER_7_1904 ();
 FILLCELL_X32 FILLER_7_1936 ();
 FILLCELL_X32 FILLER_7_1968 ();
 FILLCELL_X32 FILLER_7_2000 ();
 FILLCELL_X32 FILLER_7_2032 ();
 FILLCELL_X32 FILLER_7_2064 ();
 FILLCELL_X32 FILLER_7_2096 ();
 FILLCELL_X32 FILLER_7_2128 ();
 FILLCELL_X32 FILLER_7_2160 ();
 FILLCELL_X32 FILLER_7_2192 ();
 FILLCELL_X32 FILLER_7_2224 ();
 FILLCELL_X32 FILLER_7_2256 ();
 FILLCELL_X32 FILLER_7_2288 ();
 FILLCELL_X32 FILLER_7_2320 ();
 FILLCELL_X32 FILLER_7_2352 ();
 FILLCELL_X32 FILLER_7_2384 ();
 FILLCELL_X32 FILLER_7_2416 ();
 FILLCELL_X32 FILLER_7_2448 ();
 FILLCELL_X32 FILLER_7_2480 ();
 FILLCELL_X8 FILLER_7_2512 ();
 FILLCELL_X4 FILLER_7_2520 ();
 FILLCELL_X2 FILLER_7_2524 ();
 FILLCELL_X32 FILLER_7_2527 ();
 FILLCELL_X32 FILLER_7_2559 ();
 FILLCELL_X8 FILLER_7_2591 ();
 FILLCELL_X2 FILLER_7_2599 ();
 FILLCELL_X1 FILLER_7_2601 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_257 ();
 FILLCELL_X32 FILLER_8_289 ();
 FILLCELL_X32 FILLER_8_321 ();
 FILLCELL_X32 FILLER_8_353 ();
 FILLCELL_X32 FILLER_8_385 ();
 FILLCELL_X32 FILLER_8_417 ();
 FILLCELL_X32 FILLER_8_449 ();
 FILLCELL_X32 FILLER_8_481 ();
 FILLCELL_X32 FILLER_8_513 ();
 FILLCELL_X32 FILLER_8_545 ();
 FILLCELL_X32 FILLER_8_577 ();
 FILLCELL_X16 FILLER_8_609 ();
 FILLCELL_X4 FILLER_8_625 ();
 FILLCELL_X2 FILLER_8_629 ();
 FILLCELL_X32 FILLER_8_632 ();
 FILLCELL_X32 FILLER_8_664 ();
 FILLCELL_X32 FILLER_8_696 ();
 FILLCELL_X32 FILLER_8_728 ();
 FILLCELL_X32 FILLER_8_760 ();
 FILLCELL_X32 FILLER_8_792 ();
 FILLCELL_X32 FILLER_8_824 ();
 FILLCELL_X32 FILLER_8_856 ();
 FILLCELL_X32 FILLER_8_888 ();
 FILLCELL_X32 FILLER_8_920 ();
 FILLCELL_X32 FILLER_8_952 ();
 FILLCELL_X32 FILLER_8_984 ();
 FILLCELL_X32 FILLER_8_1016 ();
 FILLCELL_X32 FILLER_8_1048 ();
 FILLCELL_X32 FILLER_8_1080 ();
 FILLCELL_X32 FILLER_8_1112 ();
 FILLCELL_X32 FILLER_8_1144 ();
 FILLCELL_X32 FILLER_8_1176 ();
 FILLCELL_X32 FILLER_8_1208 ();
 FILLCELL_X32 FILLER_8_1240 ();
 FILLCELL_X32 FILLER_8_1272 ();
 FILLCELL_X32 FILLER_8_1304 ();
 FILLCELL_X32 FILLER_8_1336 ();
 FILLCELL_X32 FILLER_8_1368 ();
 FILLCELL_X32 FILLER_8_1400 ();
 FILLCELL_X32 FILLER_8_1432 ();
 FILLCELL_X32 FILLER_8_1464 ();
 FILLCELL_X32 FILLER_8_1496 ();
 FILLCELL_X32 FILLER_8_1528 ();
 FILLCELL_X32 FILLER_8_1560 ();
 FILLCELL_X32 FILLER_8_1592 ();
 FILLCELL_X32 FILLER_8_1624 ();
 FILLCELL_X32 FILLER_8_1656 ();
 FILLCELL_X32 FILLER_8_1688 ();
 FILLCELL_X32 FILLER_8_1720 ();
 FILLCELL_X32 FILLER_8_1752 ();
 FILLCELL_X32 FILLER_8_1784 ();
 FILLCELL_X32 FILLER_8_1816 ();
 FILLCELL_X32 FILLER_8_1848 ();
 FILLCELL_X8 FILLER_8_1880 ();
 FILLCELL_X4 FILLER_8_1888 ();
 FILLCELL_X2 FILLER_8_1892 ();
 FILLCELL_X32 FILLER_8_1895 ();
 FILLCELL_X32 FILLER_8_1927 ();
 FILLCELL_X32 FILLER_8_1959 ();
 FILLCELL_X32 FILLER_8_1991 ();
 FILLCELL_X32 FILLER_8_2023 ();
 FILLCELL_X32 FILLER_8_2055 ();
 FILLCELL_X32 FILLER_8_2087 ();
 FILLCELL_X32 FILLER_8_2119 ();
 FILLCELL_X32 FILLER_8_2151 ();
 FILLCELL_X32 FILLER_8_2183 ();
 FILLCELL_X32 FILLER_8_2215 ();
 FILLCELL_X32 FILLER_8_2247 ();
 FILLCELL_X32 FILLER_8_2279 ();
 FILLCELL_X32 FILLER_8_2311 ();
 FILLCELL_X32 FILLER_8_2343 ();
 FILLCELL_X32 FILLER_8_2375 ();
 FILLCELL_X32 FILLER_8_2407 ();
 FILLCELL_X32 FILLER_8_2439 ();
 FILLCELL_X32 FILLER_8_2471 ();
 FILLCELL_X32 FILLER_8_2503 ();
 FILLCELL_X32 FILLER_8_2535 ();
 FILLCELL_X32 FILLER_8_2567 ();
 FILLCELL_X2 FILLER_8_2599 ();
 FILLCELL_X1 FILLER_8_2601 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X32 FILLER_9_289 ();
 FILLCELL_X32 FILLER_9_321 ();
 FILLCELL_X32 FILLER_9_353 ();
 FILLCELL_X32 FILLER_9_385 ();
 FILLCELL_X32 FILLER_9_417 ();
 FILLCELL_X32 FILLER_9_449 ();
 FILLCELL_X32 FILLER_9_481 ();
 FILLCELL_X32 FILLER_9_513 ();
 FILLCELL_X32 FILLER_9_545 ();
 FILLCELL_X32 FILLER_9_577 ();
 FILLCELL_X32 FILLER_9_609 ();
 FILLCELL_X32 FILLER_9_641 ();
 FILLCELL_X32 FILLER_9_673 ();
 FILLCELL_X32 FILLER_9_705 ();
 FILLCELL_X32 FILLER_9_737 ();
 FILLCELL_X32 FILLER_9_769 ();
 FILLCELL_X32 FILLER_9_801 ();
 FILLCELL_X32 FILLER_9_833 ();
 FILLCELL_X32 FILLER_9_865 ();
 FILLCELL_X32 FILLER_9_897 ();
 FILLCELL_X32 FILLER_9_929 ();
 FILLCELL_X32 FILLER_9_961 ();
 FILLCELL_X32 FILLER_9_993 ();
 FILLCELL_X32 FILLER_9_1025 ();
 FILLCELL_X32 FILLER_9_1057 ();
 FILLCELL_X32 FILLER_9_1089 ();
 FILLCELL_X32 FILLER_9_1121 ();
 FILLCELL_X32 FILLER_9_1153 ();
 FILLCELL_X32 FILLER_9_1185 ();
 FILLCELL_X32 FILLER_9_1217 ();
 FILLCELL_X8 FILLER_9_1249 ();
 FILLCELL_X4 FILLER_9_1257 ();
 FILLCELL_X2 FILLER_9_1261 ();
 FILLCELL_X32 FILLER_9_1264 ();
 FILLCELL_X32 FILLER_9_1296 ();
 FILLCELL_X32 FILLER_9_1328 ();
 FILLCELL_X32 FILLER_9_1360 ();
 FILLCELL_X32 FILLER_9_1392 ();
 FILLCELL_X32 FILLER_9_1424 ();
 FILLCELL_X32 FILLER_9_1456 ();
 FILLCELL_X32 FILLER_9_1488 ();
 FILLCELL_X32 FILLER_9_1520 ();
 FILLCELL_X32 FILLER_9_1552 ();
 FILLCELL_X32 FILLER_9_1584 ();
 FILLCELL_X32 FILLER_9_1616 ();
 FILLCELL_X32 FILLER_9_1648 ();
 FILLCELL_X32 FILLER_9_1680 ();
 FILLCELL_X32 FILLER_9_1712 ();
 FILLCELL_X32 FILLER_9_1744 ();
 FILLCELL_X32 FILLER_9_1776 ();
 FILLCELL_X32 FILLER_9_1808 ();
 FILLCELL_X32 FILLER_9_1840 ();
 FILLCELL_X32 FILLER_9_1872 ();
 FILLCELL_X32 FILLER_9_1904 ();
 FILLCELL_X32 FILLER_9_1936 ();
 FILLCELL_X32 FILLER_9_1968 ();
 FILLCELL_X32 FILLER_9_2000 ();
 FILLCELL_X32 FILLER_9_2032 ();
 FILLCELL_X32 FILLER_9_2064 ();
 FILLCELL_X32 FILLER_9_2096 ();
 FILLCELL_X32 FILLER_9_2128 ();
 FILLCELL_X32 FILLER_9_2160 ();
 FILLCELL_X32 FILLER_9_2192 ();
 FILLCELL_X32 FILLER_9_2224 ();
 FILLCELL_X32 FILLER_9_2256 ();
 FILLCELL_X32 FILLER_9_2288 ();
 FILLCELL_X32 FILLER_9_2320 ();
 FILLCELL_X32 FILLER_9_2352 ();
 FILLCELL_X32 FILLER_9_2384 ();
 FILLCELL_X32 FILLER_9_2416 ();
 FILLCELL_X32 FILLER_9_2448 ();
 FILLCELL_X32 FILLER_9_2480 ();
 FILLCELL_X8 FILLER_9_2512 ();
 FILLCELL_X4 FILLER_9_2520 ();
 FILLCELL_X2 FILLER_9_2524 ();
 FILLCELL_X32 FILLER_9_2527 ();
 FILLCELL_X32 FILLER_9_2559 ();
 FILLCELL_X8 FILLER_9_2591 ();
 FILLCELL_X2 FILLER_9_2599 ();
 FILLCELL_X1 FILLER_9_2601 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X32 FILLER_10_289 ();
 FILLCELL_X32 FILLER_10_321 ();
 FILLCELL_X32 FILLER_10_353 ();
 FILLCELL_X32 FILLER_10_385 ();
 FILLCELL_X32 FILLER_10_417 ();
 FILLCELL_X32 FILLER_10_449 ();
 FILLCELL_X32 FILLER_10_481 ();
 FILLCELL_X32 FILLER_10_513 ();
 FILLCELL_X32 FILLER_10_545 ();
 FILLCELL_X32 FILLER_10_577 ();
 FILLCELL_X16 FILLER_10_609 ();
 FILLCELL_X4 FILLER_10_625 ();
 FILLCELL_X2 FILLER_10_629 ();
 FILLCELL_X32 FILLER_10_632 ();
 FILLCELL_X32 FILLER_10_664 ();
 FILLCELL_X32 FILLER_10_696 ();
 FILLCELL_X32 FILLER_10_728 ();
 FILLCELL_X32 FILLER_10_760 ();
 FILLCELL_X32 FILLER_10_792 ();
 FILLCELL_X32 FILLER_10_824 ();
 FILLCELL_X32 FILLER_10_856 ();
 FILLCELL_X32 FILLER_10_888 ();
 FILLCELL_X32 FILLER_10_920 ();
 FILLCELL_X32 FILLER_10_952 ();
 FILLCELL_X32 FILLER_10_984 ();
 FILLCELL_X32 FILLER_10_1016 ();
 FILLCELL_X32 FILLER_10_1048 ();
 FILLCELL_X32 FILLER_10_1080 ();
 FILLCELL_X32 FILLER_10_1112 ();
 FILLCELL_X32 FILLER_10_1144 ();
 FILLCELL_X32 FILLER_10_1176 ();
 FILLCELL_X32 FILLER_10_1208 ();
 FILLCELL_X32 FILLER_10_1240 ();
 FILLCELL_X32 FILLER_10_1272 ();
 FILLCELL_X32 FILLER_10_1304 ();
 FILLCELL_X32 FILLER_10_1336 ();
 FILLCELL_X32 FILLER_10_1368 ();
 FILLCELL_X32 FILLER_10_1400 ();
 FILLCELL_X32 FILLER_10_1432 ();
 FILLCELL_X32 FILLER_10_1464 ();
 FILLCELL_X32 FILLER_10_1496 ();
 FILLCELL_X32 FILLER_10_1528 ();
 FILLCELL_X32 FILLER_10_1560 ();
 FILLCELL_X32 FILLER_10_1592 ();
 FILLCELL_X32 FILLER_10_1624 ();
 FILLCELL_X32 FILLER_10_1656 ();
 FILLCELL_X32 FILLER_10_1688 ();
 FILLCELL_X32 FILLER_10_1720 ();
 FILLCELL_X32 FILLER_10_1752 ();
 FILLCELL_X32 FILLER_10_1784 ();
 FILLCELL_X32 FILLER_10_1816 ();
 FILLCELL_X32 FILLER_10_1848 ();
 FILLCELL_X8 FILLER_10_1880 ();
 FILLCELL_X4 FILLER_10_1888 ();
 FILLCELL_X2 FILLER_10_1892 ();
 FILLCELL_X32 FILLER_10_1895 ();
 FILLCELL_X32 FILLER_10_1927 ();
 FILLCELL_X32 FILLER_10_1959 ();
 FILLCELL_X32 FILLER_10_1991 ();
 FILLCELL_X32 FILLER_10_2023 ();
 FILLCELL_X32 FILLER_10_2055 ();
 FILLCELL_X32 FILLER_10_2087 ();
 FILLCELL_X32 FILLER_10_2119 ();
 FILLCELL_X32 FILLER_10_2151 ();
 FILLCELL_X32 FILLER_10_2183 ();
 FILLCELL_X32 FILLER_10_2215 ();
 FILLCELL_X32 FILLER_10_2247 ();
 FILLCELL_X32 FILLER_10_2279 ();
 FILLCELL_X32 FILLER_10_2311 ();
 FILLCELL_X32 FILLER_10_2343 ();
 FILLCELL_X32 FILLER_10_2375 ();
 FILLCELL_X32 FILLER_10_2407 ();
 FILLCELL_X32 FILLER_10_2439 ();
 FILLCELL_X32 FILLER_10_2471 ();
 FILLCELL_X32 FILLER_10_2503 ();
 FILLCELL_X32 FILLER_10_2535 ();
 FILLCELL_X32 FILLER_10_2567 ();
 FILLCELL_X2 FILLER_10_2599 ();
 FILLCELL_X1 FILLER_10_2601 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X32 FILLER_11_289 ();
 FILLCELL_X32 FILLER_11_321 ();
 FILLCELL_X32 FILLER_11_353 ();
 FILLCELL_X32 FILLER_11_385 ();
 FILLCELL_X32 FILLER_11_417 ();
 FILLCELL_X32 FILLER_11_449 ();
 FILLCELL_X32 FILLER_11_481 ();
 FILLCELL_X32 FILLER_11_513 ();
 FILLCELL_X32 FILLER_11_545 ();
 FILLCELL_X32 FILLER_11_577 ();
 FILLCELL_X32 FILLER_11_609 ();
 FILLCELL_X32 FILLER_11_641 ();
 FILLCELL_X32 FILLER_11_673 ();
 FILLCELL_X32 FILLER_11_705 ();
 FILLCELL_X32 FILLER_11_737 ();
 FILLCELL_X32 FILLER_11_769 ();
 FILLCELL_X32 FILLER_11_801 ();
 FILLCELL_X32 FILLER_11_833 ();
 FILLCELL_X32 FILLER_11_865 ();
 FILLCELL_X32 FILLER_11_897 ();
 FILLCELL_X32 FILLER_11_929 ();
 FILLCELL_X32 FILLER_11_961 ();
 FILLCELL_X32 FILLER_11_993 ();
 FILLCELL_X32 FILLER_11_1025 ();
 FILLCELL_X32 FILLER_11_1057 ();
 FILLCELL_X32 FILLER_11_1089 ();
 FILLCELL_X32 FILLER_11_1121 ();
 FILLCELL_X32 FILLER_11_1153 ();
 FILLCELL_X32 FILLER_11_1185 ();
 FILLCELL_X32 FILLER_11_1217 ();
 FILLCELL_X8 FILLER_11_1249 ();
 FILLCELL_X4 FILLER_11_1257 ();
 FILLCELL_X2 FILLER_11_1261 ();
 FILLCELL_X32 FILLER_11_1264 ();
 FILLCELL_X32 FILLER_11_1296 ();
 FILLCELL_X32 FILLER_11_1328 ();
 FILLCELL_X32 FILLER_11_1360 ();
 FILLCELL_X32 FILLER_11_1392 ();
 FILLCELL_X32 FILLER_11_1424 ();
 FILLCELL_X32 FILLER_11_1456 ();
 FILLCELL_X32 FILLER_11_1488 ();
 FILLCELL_X32 FILLER_11_1520 ();
 FILLCELL_X32 FILLER_11_1552 ();
 FILLCELL_X32 FILLER_11_1584 ();
 FILLCELL_X32 FILLER_11_1616 ();
 FILLCELL_X32 FILLER_11_1648 ();
 FILLCELL_X32 FILLER_11_1680 ();
 FILLCELL_X32 FILLER_11_1712 ();
 FILLCELL_X32 FILLER_11_1744 ();
 FILLCELL_X32 FILLER_11_1776 ();
 FILLCELL_X32 FILLER_11_1808 ();
 FILLCELL_X32 FILLER_11_1840 ();
 FILLCELL_X32 FILLER_11_1872 ();
 FILLCELL_X32 FILLER_11_1904 ();
 FILLCELL_X32 FILLER_11_1936 ();
 FILLCELL_X32 FILLER_11_1968 ();
 FILLCELL_X32 FILLER_11_2000 ();
 FILLCELL_X32 FILLER_11_2032 ();
 FILLCELL_X32 FILLER_11_2064 ();
 FILLCELL_X32 FILLER_11_2096 ();
 FILLCELL_X32 FILLER_11_2128 ();
 FILLCELL_X32 FILLER_11_2160 ();
 FILLCELL_X32 FILLER_11_2192 ();
 FILLCELL_X32 FILLER_11_2224 ();
 FILLCELL_X32 FILLER_11_2256 ();
 FILLCELL_X32 FILLER_11_2288 ();
 FILLCELL_X32 FILLER_11_2320 ();
 FILLCELL_X32 FILLER_11_2352 ();
 FILLCELL_X32 FILLER_11_2384 ();
 FILLCELL_X32 FILLER_11_2416 ();
 FILLCELL_X32 FILLER_11_2448 ();
 FILLCELL_X32 FILLER_11_2480 ();
 FILLCELL_X8 FILLER_11_2512 ();
 FILLCELL_X4 FILLER_11_2520 ();
 FILLCELL_X2 FILLER_11_2524 ();
 FILLCELL_X32 FILLER_11_2527 ();
 FILLCELL_X32 FILLER_11_2559 ();
 FILLCELL_X8 FILLER_11_2591 ();
 FILLCELL_X2 FILLER_11_2599 ();
 FILLCELL_X1 FILLER_11_2601 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X32 FILLER_12_257 ();
 FILLCELL_X32 FILLER_12_289 ();
 FILLCELL_X32 FILLER_12_321 ();
 FILLCELL_X32 FILLER_12_353 ();
 FILLCELL_X32 FILLER_12_385 ();
 FILLCELL_X32 FILLER_12_417 ();
 FILLCELL_X32 FILLER_12_449 ();
 FILLCELL_X32 FILLER_12_481 ();
 FILLCELL_X32 FILLER_12_513 ();
 FILLCELL_X32 FILLER_12_545 ();
 FILLCELL_X32 FILLER_12_577 ();
 FILLCELL_X16 FILLER_12_609 ();
 FILLCELL_X4 FILLER_12_625 ();
 FILLCELL_X2 FILLER_12_629 ();
 FILLCELL_X32 FILLER_12_632 ();
 FILLCELL_X32 FILLER_12_664 ();
 FILLCELL_X32 FILLER_12_696 ();
 FILLCELL_X32 FILLER_12_728 ();
 FILLCELL_X32 FILLER_12_760 ();
 FILLCELL_X32 FILLER_12_792 ();
 FILLCELL_X32 FILLER_12_824 ();
 FILLCELL_X32 FILLER_12_856 ();
 FILLCELL_X32 FILLER_12_888 ();
 FILLCELL_X32 FILLER_12_920 ();
 FILLCELL_X32 FILLER_12_952 ();
 FILLCELL_X32 FILLER_12_984 ();
 FILLCELL_X32 FILLER_12_1016 ();
 FILLCELL_X32 FILLER_12_1048 ();
 FILLCELL_X32 FILLER_12_1080 ();
 FILLCELL_X32 FILLER_12_1112 ();
 FILLCELL_X32 FILLER_12_1144 ();
 FILLCELL_X32 FILLER_12_1176 ();
 FILLCELL_X32 FILLER_12_1208 ();
 FILLCELL_X32 FILLER_12_1240 ();
 FILLCELL_X32 FILLER_12_1272 ();
 FILLCELL_X32 FILLER_12_1304 ();
 FILLCELL_X32 FILLER_12_1336 ();
 FILLCELL_X32 FILLER_12_1368 ();
 FILLCELL_X32 FILLER_12_1400 ();
 FILLCELL_X32 FILLER_12_1432 ();
 FILLCELL_X32 FILLER_12_1464 ();
 FILLCELL_X32 FILLER_12_1496 ();
 FILLCELL_X32 FILLER_12_1528 ();
 FILLCELL_X32 FILLER_12_1560 ();
 FILLCELL_X32 FILLER_12_1592 ();
 FILLCELL_X32 FILLER_12_1624 ();
 FILLCELL_X32 FILLER_12_1656 ();
 FILLCELL_X32 FILLER_12_1688 ();
 FILLCELL_X32 FILLER_12_1720 ();
 FILLCELL_X32 FILLER_12_1752 ();
 FILLCELL_X32 FILLER_12_1784 ();
 FILLCELL_X32 FILLER_12_1816 ();
 FILLCELL_X32 FILLER_12_1848 ();
 FILLCELL_X8 FILLER_12_1880 ();
 FILLCELL_X4 FILLER_12_1888 ();
 FILLCELL_X2 FILLER_12_1892 ();
 FILLCELL_X32 FILLER_12_1895 ();
 FILLCELL_X32 FILLER_12_1927 ();
 FILLCELL_X32 FILLER_12_1959 ();
 FILLCELL_X32 FILLER_12_1991 ();
 FILLCELL_X32 FILLER_12_2023 ();
 FILLCELL_X32 FILLER_12_2055 ();
 FILLCELL_X32 FILLER_12_2087 ();
 FILLCELL_X32 FILLER_12_2119 ();
 FILLCELL_X32 FILLER_12_2151 ();
 FILLCELL_X32 FILLER_12_2183 ();
 FILLCELL_X32 FILLER_12_2215 ();
 FILLCELL_X32 FILLER_12_2247 ();
 FILLCELL_X32 FILLER_12_2279 ();
 FILLCELL_X32 FILLER_12_2311 ();
 FILLCELL_X32 FILLER_12_2343 ();
 FILLCELL_X32 FILLER_12_2375 ();
 FILLCELL_X32 FILLER_12_2407 ();
 FILLCELL_X32 FILLER_12_2439 ();
 FILLCELL_X32 FILLER_12_2471 ();
 FILLCELL_X32 FILLER_12_2503 ();
 FILLCELL_X32 FILLER_12_2535 ();
 FILLCELL_X32 FILLER_12_2567 ();
 FILLCELL_X2 FILLER_12_2599 ();
 FILLCELL_X1 FILLER_12_2601 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X32 FILLER_13_257 ();
 FILLCELL_X32 FILLER_13_289 ();
 FILLCELL_X32 FILLER_13_321 ();
 FILLCELL_X32 FILLER_13_353 ();
 FILLCELL_X32 FILLER_13_385 ();
 FILLCELL_X32 FILLER_13_417 ();
 FILLCELL_X32 FILLER_13_449 ();
 FILLCELL_X32 FILLER_13_481 ();
 FILLCELL_X32 FILLER_13_513 ();
 FILLCELL_X32 FILLER_13_545 ();
 FILLCELL_X32 FILLER_13_577 ();
 FILLCELL_X32 FILLER_13_609 ();
 FILLCELL_X32 FILLER_13_641 ();
 FILLCELL_X32 FILLER_13_673 ();
 FILLCELL_X32 FILLER_13_705 ();
 FILLCELL_X32 FILLER_13_737 ();
 FILLCELL_X32 FILLER_13_769 ();
 FILLCELL_X32 FILLER_13_801 ();
 FILLCELL_X32 FILLER_13_833 ();
 FILLCELL_X32 FILLER_13_865 ();
 FILLCELL_X32 FILLER_13_897 ();
 FILLCELL_X32 FILLER_13_929 ();
 FILLCELL_X32 FILLER_13_961 ();
 FILLCELL_X32 FILLER_13_993 ();
 FILLCELL_X32 FILLER_13_1025 ();
 FILLCELL_X32 FILLER_13_1057 ();
 FILLCELL_X32 FILLER_13_1089 ();
 FILLCELL_X32 FILLER_13_1121 ();
 FILLCELL_X32 FILLER_13_1153 ();
 FILLCELL_X32 FILLER_13_1185 ();
 FILLCELL_X32 FILLER_13_1217 ();
 FILLCELL_X8 FILLER_13_1249 ();
 FILLCELL_X4 FILLER_13_1257 ();
 FILLCELL_X2 FILLER_13_1261 ();
 FILLCELL_X32 FILLER_13_1264 ();
 FILLCELL_X32 FILLER_13_1296 ();
 FILLCELL_X32 FILLER_13_1328 ();
 FILLCELL_X32 FILLER_13_1360 ();
 FILLCELL_X32 FILLER_13_1392 ();
 FILLCELL_X32 FILLER_13_1424 ();
 FILLCELL_X32 FILLER_13_1456 ();
 FILLCELL_X32 FILLER_13_1488 ();
 FILLCELL_X32 FILLER_13_1520 ();
 FILLCELL_X32 FILLER_13_1552 ();
 FILLCELL_X32 FILLER_13_1584 ();
 FILLCELL_X32 FILLER_13_1616 ();
 FILLCELL_X32 FILLER_13_1648 ();
 FILLCELL_X32 FILLER_13_1680 ();
 FILLCELL_X32 FILLER_13_1712 ();
 FILLCELL_X32 FILLER_13_1744 ();
 FILLCELL_X32 FILLER_13_1776 ();
 FILLCELL_X32 FILLER_13_1808 ();
 FILLCELL_X32 FILLER_13_1840 ();
 FILLCELL_X32 FILLER_13_1872 ();
 FILLCELL_X32 FILLER_13_1904 ();
 FILLCELL_X32 FILLER_13_1936 ();
 FILLCELL_X32 FILLER_13_1968 ();
 FILLCELL_X32 FILLER_13_2000 ();
 FILLCELL_X32 FILLER_13_2032 ();
 FILLCELL_X32 FILLER_13_2064 ();
 FILLCELL_X32 FILLER_13_2096 ();
 FILLCELL_X32 FILLER_13_2128 ();
 FILLCELL_X32 FILLER_13_2160 ();
 FILLCELL_X32 FILLER_13_2192 ();
 FILLCELL_X32 FILLER_13_2224 ();
 FILLCELL_X32 FILLER_13_2256 ();
 FILLCELL_X32 FILLER_13_2288 ();
 FILLCELL_X32 FILLER_13_2320 ();
 FILLCELL_X32 FILLER_13_2352 ();
 FILLCELL_X32 FILLER_13_2384 ();
 FILLCELL_X32 FILLER_13_2416 ();
 FILLCELL_X32 FILLER_13_2448 ();
 FILLCELL_X32 FILLER_13_2480 ();
 FILLCELL_X8 FILLER_13_2512 ();
 FILLCELL_X4 FILLER_13_2520 ();
 FILLCELL_X2 FILLER_13_2524 ();
 FILLCELL_X32 FILLER_13_2527 ();
 FILLCELL_X32 FILLER_13_2559 ();
 FILLCELL_X8 FILLER_13_2591 ();
 FILLCELL_X2 FILLER_13_2599 ();
 FILLCELL_X1 FILLER_13_2601 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X32 FILLER_14_193 ();
 FILLCELL_X32 FILLER_14_225 ();
 FILLCELL_X32 FILLER_14_257 ();
 FILLCELL_X32 FILLER_14_289 ();
 FILLCELL_X32 FILLER_14_321 ();
 FILLCELL_X32 FILLER_14_353 ();
 FILLCELL_X32 FILLER_14_385 ();
 FILLCELL_X32 FILLER_14_417 ();
 FILLCELL_X32 FILLER_14_449 ();
 FILLCELL_X32 FILLER_14_481 ();
 FILLCELL_X32 FILLER_14_513 ();
 FILLCELL_X32 FILLER_14_545 ();
 FILLCELL_X32 FILLER_14_577 ();
 FILLCELL_X16 FILLER_14_609 ();
 FILLCELL_X4 FILLER_14_625 ();
 FILLCELL_X2 FILLER_14_629 ();
 FILLCELL_X32 FILLER_14_632 ();
 FILLCELL_X32 FILLER_14_664 ();
 FILLCELL_X32 FILLER_14_696 ();
 FILLCELL_X32 FILLER_14_728 ();
 FILLCELL_X32 FILLER_14_760 ();
 FILLCELL_X32 FILLER_14_792 ();
 FILLCELL_X32 FILLER_14_824 ();
 FILLCELL_X32 FILLER_14_856 ();
 FILLCELL_X32 FILLER_14_888 ();
 FILLCELL_X32 FILLER_14_920 ();
 FILLCELL_X32 FILLER_14_952 ();
 FILLCELL_X32 FILLER_14_984 ();
 FILLCELL_X32 FILLER_14_1016 ();
 FILLCELL_X32 FILLER_14_1048 ();
 FILLCELL_X32 FILLER_14_1080 ();
 FILLCELL_X32 FILLER_14_1112 ();
 FILLCELL_X32 FILLER_14_1144 ();
 FILLCELL_X32 FILLER_14_1176 ();
 FILLCELL_X32 FILLER_14_1208 ();
 FILLCELL_X32 FILLER_14_1240 ();
 FILLCELL_X32 FILLER_14_1272 ();
 FILLCELL_X32 FILLER_14_1304 ();
 FILLCELL_X32 FILLER_14_1336 ();
 FILLCELL_X32 FILLER_14_1368 ();
 FILLCELL_X32 FILLER_14_1400 ();
 FILLCELL_X32 FILLER_14_1432 ();
 FILLCELL_X32 FILLER_14_1464 ();
 FILLCELL_X32 FILLER_14_1496 ();
 FILLCELL_X32 FILLER_14_1528 ();
 FILLCELL_X32 FILLER_14_1560 ();
 FILLCELL_X32 FILLER_14_1592 ();
 FILLCELL_X32 FILLER_14_1624 ();
 FILLCELL_X32 FILLER_14_1656 ();
 FILLCELL_X32 FILLER_14_1688 ();
 FILLCELL_X32 FILLER_14_1720 ();
 FILLCELL_X32 FILLER_14_1752 ();
 FILLCELL_X32 FILLER_14_1784 ();
 FILLCELL_X32 FILLER_14_1816 ();
 FILLCELL_X32 FILLER_14_1848 ();
 FILLCELL_X8 FILLER_14_1880 ();
 FILLCELL_X4 FILLER_14_1888 ();
 FILLCELL_X2 FILLER_14_1892 ();
 FILLCELL_X32 FILLER_14_1895 ();
 FILLCELL_X32 FILLER_14_1927 ();
 FILLCELL_X32 FILLER_14_1959 ();
 FILLCELL_X32 FILLER_14_1991 ();
 FILLCELL_X32 FILLER_14_2023 ();
 FILLCELL_X32 FILLER_14_2055 ();
 FILLCELL_X32 FILLER_14_2087 ();
 FILLCELL_X32 FILLER_14_2119 ();
 FILLCELL_X32 FILLER_14_2151 ();
 FILLCELL_X32 FILLER_14_2183 ();
 FILLCELL_X32 FILLER_14_2215 ();
 FILLCELL_X32 FILLER_14_2247 ();
 FILLCELL_X32 FILLER_14_2279 ();
 FILLCELL_X32 FILLER_14_2311 ();
 FILLCELL_X32 FILLER_14_2343 ();
 FILLCELL_X32 FILLER_14_2375 ();
 FILLCELL_X32 FILLER_14_2407 ();
 FILLCELL_X32 FILLER_14_2439 ();
 FILLCELL_X32 FILLER_14_2471 ();
 FILLCELL_X32 FILLER_14_2503 ();
 FILLCELL_X32 FILLER_14_2535 ();
 FILLCELL_X32 FILLER_14_2567 ();
 FILLCELL_X2 FILLER_14_2599 ();
 FILLCELL_X1 FILLER_14_2601 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_15_161 ();
 FILLCELL_X32 FILLER_15_193 ();
 FILLCELL_X32 FILLER_15_225 ();
 FILLCELL_X32 FILLER_15_257 ();
 FILLCELL_X32 FILLER_15_289 ();
 FILLCELL_X32 FILLER_15_321 ();
 FILLCELL_X32 FILLER_15_353 ();
 FILLCELL_X32 FILLER_15_385 ();
 FILLCELL_X32 FILLER_15_417 ();
 FILLCELL_X32 FILLER_15_449 ();
 FILLCELL_X32 FILLER_15_481 ();
 FILLCELL_X32 FILLER_15_513 ();
 FILLCELL_X32 FILLER_15_545 ();
 FILLCELL_X32 FILLER_15_577 ();
 FILLCELL_X32 FILLER_15_609 ();
 FILLCELL_X32 FILLER_15_641 ();
 FILLCELL_X32 FILLER_15_673 ();
 FILLCELL_X32 FILLER_15_705 ();
 FILLCELL_X32 FILLER_15_737 ();
 FILLCELL_X32 FILLER_15_769 ();
 FILLCELL_X32 FILLER_15_801 ();
 FILLCELL_X32 FILLER_15_833 ();
 FILLCELL_X32 FILLER_15_865 ();
 FILLCELL_X32 FILLER_15_897 ();
 FILLCELL_X32 FILLER_15_929 ();
 FILLCELL_X32 FILLER_15_961 ();
 FILLCELL_X32 FILLER_15_993 ();
 FILLCELL_X32 FILLER_15_1025 ();
 FILLCELL_X32 FILLER_15_1057 ();
 FILLCELL_X32 FILLER_15_1089 ();
 FILLCELL_X32 FILLER_15_1121 ();
 FILLCELL_X32 FILLER_15_1153 ();
 FILLCELL_X32 FILLER_15_1185 ();
 FILLCELL_X32 FILLER_15_1217 ();
 FILLCELL_X8 FILLER_15_1249 ();
 FILLCELL_X4 FILLER_15_1257 ();
 FILLCELL_X2 FILLER_15_1261 ();
 FILLCELL_X32 FILLER_15_1264 ();
 FILLCELL_X32 FILLER_15_1296 ();
 FILLCELL_X32 FILLER_15_1328 ();
 FILLCELL_X32 FILLER_15_1360 ();
 FILLCELL_X32 FILLER_15_1392 ();
 FILLCELL_X32 FILLER_15_1424 ();
 FILLCELL_X32 FILLER_15_1456 ();
 FILLCELL_X32 FILLER_15_1488 ();
 FILLCELL_X32 FILLER_15_1520 ();
 FILLCELL_X32 FILLER_15_1552 ();
 FILLCELL_X32 FILLER_15_1584 ();
 FILLCELL_X32 FILLER_15_1616 ();
 FILLCELL_X32 FILLER_15_1648 ();
 FILLCELL_X32 FILLER_15_1680 ();
 FILLCELL_X32 FILLER_15_1712 ();
 FILLCELL_X32 FILLER_15_1744 ();
 FILLCELL_X32 FILLER_15_1776 ();
 FILLCELL_X32 FILLER_15_1808 ();
 FILLCELL_X32 FILLER_15_1840 ();
 FILLCELL_X32 FILLER_15_1872 ();
 FILLCELL_X32 FILLER_15_1904 ();
 FILLCELL_X32 FILLER_15_1936 ();
 FILLCELL_X32 FILLER_15_1968 ();
 FILLCELL_X32 FILLER_15_2000 ();
 FILLCELL_X32 FILLER_15_2032 ();
 FILLCELL_X32 FILLER_15_2064 ();
 FILLCELL_X32 FILLER_15_2096 ();
 FILLCELL_X32 FILLER_15_2128 ();
 FILLCELL_X32 FILLER_15_2160 ();
 FILLCELL_X32 FILLER_15_2192 ();
 FILLCELL_X32 FILLER_15_2224 ();
 FILLCELL_X32 FILLER_15_2256 ();
 FILLCELL_X32 FILLER_15_2288 ();
 FILLCELL_X32 FILLER_15_2320 ();
 FILLCELL_X32 FILLER_15_2352 ();
 FILLCELL_X32 FILLER_15_2384 ();
 FILLCELL_X32 FILLER_15_2416 ();
 FILLCELL_X32 FILLER_15_2448 ();
 FILLCELL_X32 FILLER_15_2480 ();
 FILLCELL_X8 FILLER_15_2512 ();
 FILLCELL_X4 FILLER_15_2520 ();
 FILLCELL_X2 FILLER_15_2524 ();
 FILLCELL_X32 FILLER_15_2527 ();
 FILLCELL_X32 FILLER_15_2559 ();
 FILLCELL_X8 FILLER_15_2591 ();
 FILLCELL_X2 FILLER_15_2599 ();
 FILLCELL_X1 FILLER_15_2601 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X32 FILLER_16_193 ();
 FILLCELL_X32 FILLER_16_225 ();
 FILLCELL_X32 FILLER_16_257 ();
 FILLCELL_X32 FILLER_16_289 ();
 FILLCELL_X32 FILLER_16_321 ();
 FILLCELL_X32 FILLER_16_353 ();
 FILLCELL_X32 FILLER_16_385 ();
 FILLCELL_X32 FILLER_16_417 ();
 FILLCELL_X32 FILLER_16_449 ();
 FILLCELL_X32 FILLER_16_481 ();
 FILLCELL_X32 FILLER_16_513 ();
 FILLCELL_X32 FILLER_16_545 ();
 FILLCELL_X32 FILLER_16_577 ();
 FILLCELL_X16 FILLER_16_609 ();
 FILLCELL_X4 FILLER_16_625 ();
 FILLCELL_X2 FILLER_16_629 ();
 FILLCELL_X32 FILLER_16_632 ();
 FILLCELL_X32 FILLER_16_664 ();
 FILLCELL_X32 FILLER_16_696 ();
 FILLCELL_X32 FILLER_16_728 ();
 FILLCELL_X32 FILLER_16_760 ();
 FILLCELL_X32 FILLER_16_792 ();
 FILLCELL_X32 FILLER_16_824 ();
 FILLCELL_X32 FILLER_16_856 ();
 FILLCELL_X32 FILLER_16_888 ();
 FILLCELL_X32 FILLER_16_920 ();
 FILLCELL_X32 FILLER_16_952 ();
 FILLCELL_X32 FILLER_16_984 ();
 FILLCELL_X32 FILLER_16_1016 ();
 FILLCELL_X32 FILLER_16_1048 ();
 FILLCELL_X32 FILLER_16_1080 ();
 FILLCELL_X32 FILLER_16_1112 ();
 FILLCELL_X32 FILLER_16_1144 ();
 FILLCELL_X32 FILLER_16_1176 ();
 FILLCELL_X32 FILLER_16_1208 ();
 FILLCELL_X32 FILLER_16_1240 ();
 FILLCELL_X32 FILLER_16_1272 ();
 FILLCELL_X32 FILLER_16_1304 ();
 FILLCELL_X32 FILLER_16_1336 ();
 FILLCELL_X32 FILLER_16_1368 ();
 FILLCELL_X32 FILLER_16_1400 ();
 FILLCELL_X32 FILLER_16_1432 ();
 FILLCELL_X32 FILLER_16_1464 ();
 FILLCELL_X32 FILLER_16_1496 ();
 FILLCELL_X32 FILLER_16_1528 ();
 FILLCELL_X32 FILLER_16_1560 ();
 FILLCELL_X32 FILLER_16_1592 ();
 FILLCELL_X32 FILLER_16_1624 ();
 FILLCELL_X32 FILLER_16_1656 ();
 FILLCELL_X32 FILLER_16_1688 ();
 FILLCELL_X32 FILLER_16_1720 ();
 FILLCELL_X32 FILLER_16_1752 ();
 FILLCELL_X32 FILLER_16_1784 ();
 FILLCELL_X32 FILLER_16_1816 ();
 FILLCELL_X32 FILLER_16_1848 ();
 FILLCELL_X8 FILLER_16_1880 ();
 FILLCELL_X4 FILLER_16_1888 ();
 FILLCELL_X2 FILLER_16_1892 ();
 FILLCELL_X32 FILLER_16_1895 ();
 FILLCELL_X32 FILLER_16_1927 ();
 FILLCELL_X32 FILLER_16_1959 ();
 FILLCELL_X32 FILLER_16_1991 ();
 FILLCELL_X32 FILLER_16_2023 ();
 FILLCELL_X32 FILLER_16_2055 ();
 FILLCELL_X32 FILLER_16_2087 ();
 FILLCELL_X32 FILLER_16_2119 ();
 FILLCELL_X32 FILLER_16_2151 ();
 FILLCELL_X32 FILLER_16_2183 ();
 FILLCELL_X32 FILLER_16_2215 ();
 FILLCELL_X32 FILLER_16_2247 ();
 FILLCELL_X32 FILLER_16_2279 ();
 FILLCELL_X32 FILLER_16_2311 ();
 FILLCELL_X32 FILLER_16_2343 ();
 FILLCELL_X32 FILLER_16_2375 ();
 FILLCELL_X32 FILLER_16_2407 ();
 FILLCELL_X32 FILLER_16_2439 ();
 FILLCELL_X32 FILLER_16_2471 ();
 FILLCELL_X32 FILLER_16_2503 ();
 FILLCELL_X32 FILLER_16_2535 ();
 FILLCELL_X32 FILLER_16_2567 ();
 FILLCELL_X2 FILLER_16_2599 ();
 FILLCELL_X1 FILLER_16_2601 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X32 FILLER_17_193 ();
 FILLCELL_X32 FILLER_17_225 ();
 FILLCELL_X32 FILLER_17_257 ();
 FILLCELL_X32 FILLER_17_289 ();
 FILLCELL_X32 FILLER_17_321 ();
 FILLCELL_X32 FILLER_17_353 ();
 FILLCELL_X32 FILLER_17_385 ();
 FILLCELL_X32 FILLER_17_417 ();
 FILLCELL_X32 FILLER_17_449 ();
 FILLCELL_X32 FILLER_17_481 ();
 FILLCELL_X32 FILLER_17_513 ();
 FILLCELL_X32 FILLER_17_545 ();
 FILLCELL_X32 FILLER_17_577 ();
 FILLCELL_X32 FILLER_17_609 ();
 FILLCELL_X32 FILLER_17_641 ();
 FILLCELL_X32 FILLER_17_673 ();
 FILLCELL_X32 FILLER_17_705 ();
 FILLCELL_X32 FILLER_17_737 ();
 FILLCELL_X32 FILLER_17_769 ();
 FILLCELL_X32 FILLER_17_801 ();
 FILLCELL_X32 FILLER_17_833 ();
 FILLCELL_X32 FILLER_17_865 ();
 FILLCELL_X32 FILLER_17_897 ();
 FILLCELL_X32 FILLER_17_929 ();
 FILLCELL_X32 FILLER_17_961 ();
 FILLCELL_X32 FILLER_17_993 ();
 FILLCELL_X32 FILLER_17_1025 ();
 FILLCELL_X32 FILLER_17_1057 ();
 FILLCELL_X32 FILLER_17_1089 ();
 FILLCELL_X32 FILLER_17_1121 ();
 FILLCELL_X32 FILLER_17_1153 ();
 FILLCELL_X32 FILLER_17_1185 ();
 FILLCELL_X32 FILLER_17_1217 ();
 FILLCELL_X8 FILLER_17_1249 ();
 FILLCELL_X4 FILLER_17_1257 ();
 FILLCELL_X2 FILLER_17_1261 ();
 FILLCELL_X32 FILLER_17_1264 ();
 FILLCELL_X32 FILLER_17_1296 ();
 FILLCELL_X32 FILLER_17_1328 ();
 FILLCELL_X32 FILLER_17_1360 ();
 FILLCELL_X32 FILLER_17_1392 ();
 FILLCELL_X32 FILLER_17_1424 ();
 FILLCELL_X32 FILLER_17_1456 ();
 FILLCELL_X32 FILLER_17_1488 ();
 FILLCELL_X32 FILLER_17_1520 ();
 FILLCELL_X32 FILLER_17_1552 ();
 FILLCELL_X32 FILLER_17_1584 ();
 FILLCELL_X32 FILLER_17_1616 ();
 FILLCELL_X32 FILLER_17_1648 ();
 FILLCELL_X32 FILLER_17_1680 ();
 FILLCELL_X32 FILLER_17_1712 ();
 FILLCELL_X32 FILLER_17_1744 ();
 FILLCELL_X32 FILLER_17_1776 ();
 FILLCELL_X32 FILLER_17_1808 ();
 FILLCELL_X32 FILLER_17_1840 ();
 FILLCELL_X32 FILLER_17_1872 ();
 FILLCELL_X32 FILLER_17_1904 ();
 FILLCELL_X32 FILLER_17_1936 ();
 FILLCELL_X32 FILLER_17_1968 ();
 FILLCELL_X32 FILLER_17_2000 ();
 FILLCELL_X32 FILLER_17_2032 ();
 FILLCELL_X32 FILLER_17_2064 ();
 FILLCELL_X32 FILLER_17_2096 ();
 FILLCELL_X32 FILLER_17_2128 ();
 FILLCELL_X32 FILLER_17_2160 ();
 FILLCELL_X32 FILLER_17_2192 ();
 FILLCELL_X32 FILLER_17_2224 ();
 FILLCELL_X32 FILLER_17_2256 ();
 FILLCELL_X32 FILLER_17_2288 ();
 FILLCELL_X32 FILLER_17_2320 ();
 FILLCELL_X32 FILLER_17_2352 ();
 FILLCELL_X32 FILLER_17_2384 ();
 FILLCELL_X32 FILLER_17_2416 ();
 FILLCELL_X32 FILLER_17_2448 ();
 FILLCELL_X32 FILLER_17_2480 ();
 FILLCELL_X8 FILLER_17_2512 ();
 FILLCELL_X4 FILLER_17_2520 ();
 FILLCELL_X2 FILLER_17_2524 ();
 FILLCELL_X32 FILLER_17_2527 ();
 FILLCELL_X32 FILLER_17_2559 ();
 FILLCELL_X8 FILLER_17_2591 ();
 FILLCELL_X2 FILLER_17_2599 ();
 FILLCELL_X1 FILLER_17_2601 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X32 FILLER_18_193 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X32 FILLER_18_257 ();
 FILLCELL_X32 FILLER_18_289 ();
 FILLCELL_X32 FILLER_18_321 ();
 FILLCELL_X32 FILLER_18_353 ();
 FILLCELL_X32 FILLER_18_385 ();
 FILLCELL_X32 FILLER_18_417 ();
 FILLCELL_X32 FILLER_18_449 ();
 FILLCELL_X32 FILLER_18_481 ();
 FILLCELL_X32 FILLER_18_513 ();
 FILLCELL_X32 FILLER_18_545 ();
 FILLCELL_X32 FILLER_18_577 ();
 FILLCELL_X16 FILLER_18_609 ();
 FILLCELL_X4 FILLER_18_625 ();
 FILLCELL_X2 FILLER_18_629 ();
 FILLCELL_X32 FILLER_18_632 ();
 FILLCELL_X32 FILLER_18_664 ();
 FILLCELL_X32 FILLER_18_696 ();
 FILLCELL_X32 FILLER_18_728 ();
 FILLCELL_X32 FILLER_18_760 ();
 FILLCELL_X32 FILLER_18_792 ();
 FILLCELL_X32 FILLER_18_824 ();
 FILLCELL_X32 FILLER_18_856 ();
 FILLCELL_X32 FILLER_18_888 ();
 FILLCELL_X32 FILLER_18_920 ();
 FILLCELL_X32 FILLER_18_952 ();
 FILLCELL_X32 FILLER_18_984 ();
 FILLCELL_X32 FILLER_18_1016 ();
 FILLCELL_X32 FILLER_18_1048 ();
 FILLCELL_X32 FILLER_18_1080 ();
 FILLCELL_X32 FILLER_18_1112 ();
 FILLCELL_X32 FILLER_18_1144 ();
 FILLCELL_X32 FILLER_18_1176 ();
 FILLCELL_X32 FILLER_18_1208 ();
 FILLCELL_X32 FILLER_18_1240 ();
 FILLCELL_X32 FILLER_18_1272 ();
 FILLCELL_X32 FILLER_18_1304 ();
 FILLCELL_X32 FILLER_18_1336 ();
 FILLCELL_X32 FILLER_18_1368 ();
 FILLCELL_X32 FILLER_18_1400 ();
 FILLCELL_X32 FILLER_18_1432 ();
 FILLCELL_X32 FILLER_18_1464 ();
 FILLCELL_X32 FILLER_18_1496 ();
 FILLCELL_X32 FILLER_18_1528 ();
 FILLCELL_X32 FILLER_18_1560 ();
 FILLCELL_X32 FILLER_18_1592 ();
 FILLCELL_X32 FILLER_18_1624 ();
 FILLCELL_X32 FILLER_18_1656 ();
 FILLCELL_X32 FILLER_18_1688 ();
 FILLCELL_X32 FILLER_18_1720 ();
 FILLCELL_X32 FILLER_18_1752 ();
 FILLCELL_X32 FILLER_18_1784 ();
 FILLCELL_X32 FILLER_18_1816 ();
 FILLCELL_X32 FILLER_18_1848 ();
 FILLCELL_X8 FILLER_18_1880 ();
 FILLCELL_X4 FILLER_18_1888 ();
 FILLCELL_X2 FILLER_18_1892 ();
 FILLCELL_X32 FILLER_18_1895 ();
 FILLCELL_X32 FILLER_18_1927 ();
 FILLCELL_X32 FILLER_18_1959 ();
 FILLCELL_X32 FILLER_18_1991 ();
 FILLCELL_X32 FILLER_18_2023 ();
 FILLCELL_X32 FILLER_18_2055 ();
 FILLCELL_X32 FILLER_18_2087 ();
 FILLCELL_X32 FILLER_18_2119 ();
 FILLCELL_X32 FILLER_18_2151 ();
 FILLCELL_X32 FILLER_18_2183 ();
 FILLCELL_X32 FILLER_18_2215 ();
 FILLCELL_X32 FILLER_18_2247 ();
 FILLCELL_X32 FILLER_18_2279 ();
 FILLCELL_X32 FILLER_18_2311 ();
 FILLCELL_X32 FILLER_18_2343 ();
 FILLCELL_X32 FILLER_18_2375 ();
 FILLCELL_X32 FILLER_18_2407 ();
 FILLCELL_X32 FILLER_18_2439 ();
 FILLCELL_X32 FILLER_18_2471 ();
 FILLCELL_X32 FILLER_18_2503 ();
 FILLCELL_X32 FILLER_18_2535 ();
 FILLCELL_X32 FILLER_18_2567 ();
 FILLCELL_X2 FILLER_18_2599 ();
 FILLCELL_X1 FILLER_18_2601 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X32 FILLER_19_193 ();
 FILLCELL_X32 FILLER_19_225 ();
 FILLCELL_X32 FILLER_19_257 ();
 FILLCELL_X32 FILLER_19_289 ();
 FILLCELL_X32 FILLER_19_321 ();
 FILLCELL_X32 FILLER_19_353 ();
 FILLCELL_X32 FILLER_19_385 ();
 FILLCELL_X32 FILLER_19_417 ();
 FILLCELL_X32 FILLER_19_449 ();
 FILLCELL_X32 FILLER_19_481 ();
 FILLCELL_X32 FILLER_19_513 ();
 FILLCELL_X32 FILLER_19_545 ();
 FILLCELL_X32 FILLER_19_577 ();
 FILLCELL_X32 FILLER_19_609 ();
 FILLCELL_X32 FILLER_19_641 ();
 FILLCELL_X32 FILLER_19_673 ();
 FILLCELL_X32 FILLER_19_705 ();
 FILLCELL_X32 FILLER_19_737 ();
 FILLCELL_X32 FILLER_19_769 ();
 FILLCELL_X32 FILLER_19_801 ();
 FILLCELL_X32 FILLER_19_833 ();
 FILLCELL_X32 FILLER_19_865 ();
 FILLCELL_X32 FILLER_19_897 ();
 FILLCELL_X32 FILLER_19_929 ();
 FILLCELL_X32 FILLER_19_961 ();
 FILLCELL_X32 FILLER_19_993 ();
 FILLCELL_X32 FILLER_19_1025 ();
 FILLCELL_X32 FILLER_19_1057 ();
 FILLCELL_X32 FILLER_19_1089 ();
 FILLCELL_X32 FILLER_19_1121 ();
 FILLCELL_X32 FILLER_19_1153 ();
 FILLCELL_X32 FILLER_19_1185 ();
 FILLCELL_X32 FILLER_19_1217 ();
 FILLCELL_X8 FILLER_19_1249 ();
 FILLCELL_X4 FILLER_19_1257 ();
 FILLCELL_X2 FILLER_19_1261 ();
 FILLCELL_X32 FILLER_19_1264 ();
 FILLCELL_X32 FILLER_19_1296 ();
 FILLCELL_X32 FILLER_19_1328 ();
 FILLCELL_X32 FILLER_19_1360 ();
 FILLCELL_X32 FILLER_19_1392 ();
 FILLCELL_X32 FILLER_19_1424 ();
 FILLCELL_X32 FILLER_19_1456 ();
 FILLCELL_X32 FILLER_19_1488 ();
 FILLCELL_X32 FILLER_19_1520 ();
 FILLCELL_X32 FILLER_19_1552 ();
 FILLCELL_X32 FILLER_19_1584 ();
 FILLCELL_X32 FILLER_19_1616 ();
 FILLCELL_X32 FILLER_19_1648 ();
 FILLCELL_X32 FILLER_19_1680 ();
 FILLCELL_X32 FILLER_19_1712 ();
 FILLCELL_X32 FILLER_19_1744 ();
 FILLCELL_X32 FILLER_19_1776 ();
 FILLCELL_X32 FILLER_19_1808 ();
 FILLCELL_X32 FILLER_19_1840 ();
 FILLCELL_X32 FILLER_19_1872 ();
 FILLCELL_X32 FILLER_19_1904 ();
 FILLCELL_X32 FILLER_19_1936 ();
 FILLCELL_X32 FILLER_19_1968 ();
 FILLCELL_X32 FILLER_19_2000 ();
 FILLCELL_X32 FILLER_19_2032 ();
 FILLCELL_X32 FILLER_19_2064 ();
 FILLCELL_X32 FILLER_19_2096 ();
 FILLCELL_X32 FILLER_19_2128 ();
 FILLCELL_X32 FILLER_19_2160 ();
 FILLCELL_X32 FILLER_19_2192 ();
 FILLCELL_X32 FILLER_19_2224 ();
 FILLCELL_X32 FILLER_19_2256 ();
 FILLCELL_X32 FILLER_19_2288 ();
 FILLCELL_X32 FILLER_19_2320 ();
 FILLCELL_X32 FILLER_19_2352 ();
 FILLCELL_X32 FILLER_19_2384 ();
 FILLCELL_X32 FILLER_19_2416 ();
 FILLCELL_X32 FILLER_19_2448 ();
 FILLCELL_X32 FILLER_19_2480 ();
 FILLCELL_X8 FILLER_19_2512 ();
 FILLCELL_X4 FILLER_19_2520 ();
 FILLCELL_X2 FILLER_19_2524 ();
 FILLCELL_X32 FILLER_19_2527 ();
 FILLCELL_X32 FILLER_19_2559 ();
 FILLCELL_X8 FILLER_19_2591 ();
 FILLCELL_X2 FILLER_19_2599 ();
 FILLCELL_X1 FILLER_19_2601 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X32 FILLER_20_193 ();
 FILLCELL_X32 FILLER_20_225 ();
 FILLCELL_X32 FILLER_20_257 ();
 FILLCELL_X32 FILLER_20_289 ();
 FILLCELL_X32 FILLER_20_321 ();
 FILLCELL_X32 FILLER_20_353 ();
 FILLCELL_X32 FILLER_20_385 ();
 FILLCELL_X32 FILLER_20_417 ();
 FILLCELL_X32 FILLER_20_449 ();
 FILLCELL_X32 FILLER_20_481 ();
 FILLCELL_X32 FILLER_20_513 ();
 FILLCELL_X32 FILLER_20_545 ();
 FILLCELL_X32 FILLER_20_577 ();
 FILLCELL_X16 FILLER_20_609 ();
 FILLCELL_X4 FILLER_20_625 ();
 FILLCELL_X2 FILLER_20_629 ();
 FILLCELL_X32 FILLER_20_632 ();
 FILLCELL_X32 FILLER_20_664 ();
 FILLCELL_X32 FILLER_20_696 ();
 FILLCELL_X32 FILLER_20_728 ();
 FILLCELL_X32 FILLER_20_760 ();
 FILLCELL_X32 FILLER_20_792 ();
 FILLCELL_X32 FILLER_20_824 ();
 FILLCELL_X32 FILLER_20_856 ();
 FILLCELL_X32 FILLER_20_888 ();
 FILLCELL_X32 FILLER_20_920 ();
 FILLCELL_X32 FILLER_20_952 ();
 FILLCELL_X32 FILLER_20_984 ();
 FILLCELL_X32 FILLER_20_1016 ();
 FILLCELL_X32 FILLER_20_1048 ();
 FILLCELL_X32 FILLER_20_1080 ();
 FILLCELL_X32 FILLER_20_1112 ();
 FILLCELL_X32 FILLER_20_1144 ();
 FILLCELL_X32 FILLER_20_1176 ();
 FILLCELL_X32 FILLER_20_1208 ();
 FILLCELL_X32 FILLER_20_1240 ();
 FILLCELL_X32 FILLER_20_1272 ();
 FILLCELL_X32 FILLER_20_1304 ();
 FILLCELL_X32 FILLER_20_1336 ();
 FILLCELL_X32 FILLER_20_1368 ();
 FILLCELL_X32 FILLER_20_1400 ();
 FILLCELL_X32 FILLER_20_1432 ();
 FILLCELL_X32 FILLER_20_1464 ();
 FILLCELL_X32 FILLER_20_1496 ();
 FILLCELL_X32 FILLER_20_1528 ();
 FILLCELL_X32 FILLER_20_1560 ();
 FILLCELL_X32 FILLER_20_1592 ();
 FILLCELL_X32 FILLER_20_1624 ();
 FILLCELL_X32 FILLER_20_1656 ();
 FILLCELL_X32 FILLER_20_1688 ();
 FILLCELL_X32 FILLER_20_1720 ();
 FILLCELL_X32 FILLER_20_1752 ();
 FILLCELL_X32 FILLER_20_1784 ();
 FILLCELL_X32 FILLER_20_1816 ();
 FILLCELL_X32 FILLER_20_1848 ();
 FILLCELL_X8 FILLER_20_1880 ();
 FILLCELL_X4 FILLER_20_1888 ();
 FILLCELL_X2 FILLER_20_1892 ();
 FILLCELL_X32 FILLER_20_1895 ();
 FILLCELL_X32 FILLER_20_1927 ();
 FILLCELL_X32 FILLER_20_1959 ();
 FILLCELL_X32 FILLER_20_1991 ();
 FILLCELL_X32 FILLER_20_2023 ();
 FILLCELL_X32 FILLER_20_2055 ();
 FILLCELL_X32 FILLER_20_2087 ();
 FILLCELL_X32 FILLER_20_2119 ();
 FILLCELL_X32 FILLER_20_2151 ();
 FILLCELL_X32 FILLER_20_2183 ();
 FILLCELL_X32 FILLER_20_2215 ();
 FILLCELL_X32 FILLER_20_2247 ();
 FILLCELL_X32 FILLER_20_2279 ();
 FILLCELL_X32 FILLER_20_2311 ();
 FILLCELL_X32 FILLER_20_2343 ();
 FILLCELL_X32 FILLER_20_2375 ();
 FILLCELL_X32 FILLER_20_2407 ();
 FILLCELL_X32 FILLER_20_2439 ();
 FILLCELL_X32 FILLER_20_2471 ();
 FILLCELL_X32 FILLER_20_2503 ();
 FILLCELL_X32 FILLER_20_2535 ();
 FILLCELL_X32 FILLER_20_2567 ();
 FILLCELL_X2 FILLER_20_2599 ();
 FILLCELL_X1 FILLER_20_2601 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X32 FILLER_21_193 ();
 FILLCELL_X32 FILLER_21_225 ();
 FILLCELL_X32 FILLER_21_257 ();
 FILLCELL_X32 FILLER_21_289 ();
 FILLCELL_X32 FILLER_21_321 ();
 FILLCELL_X32 FILLER_21_353 ();
 FILLCELL_X32 FILLER_21_385 ();
 FILLCELL_X32 FILLER_21_417 ();
 FILLCELL_X32 FILLER_21_449 ();
 FILLCELL_X32 FILLER_21_481 ();
 FILLCELL_X32 FILLER_21_513 ();
 FILLCELL_X32 FILLER_21_545 ();
 FILLCELL_X32 FILLER_21_577 ();
 FILLCELL_X32 FILLER_21_609 ();
 FILLCELL_X32 FILLER_21_641 ();
 FILLCELL_X32 FILLER_21_673 ();
 FILLCELL_X32 FILLER_21_705 ();
 FILLCELL_X32 FILLER_21_737 ();
 FILLCELL_X32 FILLER_21_769 ();
 FILLCELL_X32 FILLER_21_801 ();
 FILLCELL_X32 FILLER_21_833 ();
 FILLCELL_X32 FILLER_21_865 ();
 FILLCELL_X32 FILLER_21_897 ();
 FILLCELL_X32 FILLER_21_929 ();
 FILLCELL_X32 FILLER_21_961 ();
 FILLCELL_X32 FILLER_21_993 ();
 FILLCELL_X32 FILLER_21_1025 ();
 FILLCELL_X32 FILLER_21_1057 ();
 FILLCELL_X32 FILLER_21_1089 ();
 FILLCELL_X32 FILLER_21_1121 ();
 FILLCELL_X32 FILLER_21_1153 ();
 FILLCELL_X32 FILLER_21_1185 ();
 FILLCELL_X32 FILLER_21_1217 ();
 FILLCELL_X8 FILLER_21_1249 ();
 FILLCELL_X4 FILLER_21_1257 ();
 FILLCELL_X2 FILLER_21_1261 ();
 FILLCELL_X32 FILLER_21_1264 ();
 FILLCELL_X32 FILLER_21_1296 ();
 FILLCELL_X32 FILLER_21_1328 ();
 FILLCELL_X32 FILLER_21_1360 ();
 FILLCELL_X32 FILLER_21_1392 ();
 FILLCELL_X32 FILLER_21_1424 ();
 FILLCELL_X32 FILLER_21_1456 ();
 FILLCELL_X32 FILLER_21_1488 ();
 FILLCELL_X32 FILLER_21_1520 ();
 FILLCELL_X32 FILLER_21_1552 ();
 FILLCELL_X32 FILLER_21_1584 ();
 FILLCELL_X32 FILLER_21_1616 ();
 FILLCELL_X32 FILLER_21_1648 ();
 FILLCELL_X32 FILLER_21_1680 ();
 FILLCELL_X32 FILLER_21_1712 ();
 FILLCELL_X32 FILLER_21_1744 ();
 FILLCELL_X32 FILLER_21_1776 ();
 FILLCELL_X32 FILLER_21_1808 ();
 FILLCELL_X32 FILLER_21_1840 ();
 FILLCELL_X32 FILLER_21_1872 ();
 FILLCELL_X32 FILLER_21_1904 ();
 FILLCELL_X32 FILLER_21_1936 ();
 FILLCELL_X32 FILLER_21_1968 ();
 FILLCELL_X32 FILLER_21_2000 ();
 FILLCELL_X32 FILLER_21_2032 ();
 FILLCELL_X32 FILLER_21_2064 ();
 FILLCELL_X32 FILLER_21_2096 ();
 FILLCELL_X32 FILLER_21_2128 ();
 FILLCELL_X32 FILLER_21_2160 ();
 FILLCELL_X32 FILLER_21_2192 ();
 FILLCELL_X32 FILLER_21_2224 ();
 FILLCELL_X32 FILLER_21_2256 ();
 FILLCELL_X32 FILLER_21_2288 ();
 FILLCELL_X32 FILLER_21_2320 ();
 FILLCELL_X32 FILLER_21_2352 ();
 FILLCELL_X32 FILLER_21_2384 ();
 FILLCELL_X32 FILLER_21_2416 ();
 FILLCELL_X32 FILLER_21_2448 ();
 FILLCELL_X32 FILLER_21_2480 ();
 FILLCELL_X8 FILLER_21_2512 ();
 FILLCELL_X4 FILLER_21_2520 ();
 FILLCELL_X2 FILLER_21_2524 ();
 FILLCELL_X32 FILLER_21_2527 ();
 FILLCELL_X32 FILLER_21_2559 ();
 FILLCELL_X8 FILLER_21_2591 ();
 FILLCELL_X2 FILLER_21_2599 ();
 FILLCELL_X1 FILLER_21_2601 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X32 FILLER_22_193 ();
 FILLCELL_X32 FILLER_22_225 ();
 FILLCELL_X32 FILLER_22_257 ();
 FILLCELL_X32 FILLER_22_289 ();
 FILLCELL_X32 FILLER_22_321 ();
 FILLCELL_X32 FILLER_22_353 ();
 FILLCELL_X32 FILLER_22_385 ();
 FILLCELL_X32 FILLER_22_417 ();
 FILLCELL_X32 FILLER_22_449 ();
 FILLCELL_X32 FILLER_22_481 ();
 FILLCELL_X32 FILLER_22_513 ();
 FILLCELL_X32 FILLER_22_545 ();
 FILLCELL_X32 FILLER_22_577 ();
 FILLCELL_X16 FILLER_22_609 ();
 FILLCELL_X4 FILLER_22_625 ();
 FILLCELL_X2 FILLER_22_629 ();
 FILLCELL_X32 FILLER_22_632 ();
 FILLCELL_X32 FILLER_22_664 ();
 FILLCELL_X32 FILLER_22_696 ();
 FILLCELL_X32 FILLER_22_728 ();
 FILLCELL_X32 FILLER_22_760 ();
 FILLCELL_X32 FILLER_22_792 ();
 FILLCELL_X32 FILLER_22_824 ();
 FILLCELL_X32 FILLER_22_856 ();
 FILLCELL_X32 FILLER_22_888 ();
 FILLCELL_X32 FILLER_22_920 ();
 FILLCELL_X32 FILLER_22_952 ();
 FILLCELL_X32 FILLER_22_984 ();
 FILLCELL_X32 FILLER_22_1016 ();
 FILLCELL_X32 FILLER_22_1048 ();
 FILLCELL_X32 FILLER_22_1080 ();
 FILLCELL_X32 FILLER_22_1112 ();
 FILLCELL_X32 FILLER_22_1144 ();
 FILLCELL_X32 FILLER_22_1176 ();
 FILLCELL_X32 FILLER_22_1208 ();
 FILLCELL_X32 FILLER_22_1240 ();
 FILLCELL_X32 FILLER_22_1272 ();
 FILLCELL_X32 FILLER_22_1304 ();
 FILLCELL_X32 FILLER_22_1336 ();
 FILLCELL_X32 FILLER_22_1368 ();
 FILLCELL_X32 FILLER_22_1400 ();
 FILLCELL_X32 FILLER_22_1432 ();
 FILLCELL_X32 FILLER_22_1464 ();
 FILLCELL_X32 FILLER_22_1496 ();
 FILLCELL_X32 FILLER_22_1528 ();
 FILLCELL_X32 FILLER_22_1560 ();
 FILLCELL_X32 FILLER_22_1592 ();
 FILLCELL_X32 FILLER_22_1624 ();
 FILLCELL_X32 FILLER_22_1656 ();
 FILLCELL_X32 FILLER_22_1688 ();
 FILLCELL_X32 FILLER_22_1720 ();
 FILLCELL_X32 FILLER_22_1752 ();
 FILLCELL_X32 FILLER_22_1784 ();
 FILLCELL_X32 FILLER_22_1816 ();
 FILLCELL_X32 FILLER_22_1848 ();
 FILLCELL_X8 FILLER_22_1880 ();
 FILLCELL_X4 FILLER_22_1888 ();
 FILLCELL_X2 FILLER_22_1892 ();
 FILLCELL_X32 FILLER_22_1895 ();
 FILLCELL_X32 FILLER_22_1927 ();
 FILLCELL_X32 FILLER_22_1959 ();
 FILLCELL_X32 FILLER_22_1991 ();
 FILLCELL_X32 FILLER_22_2023 ();
 FILLCELL_X32 FILLER_22_2055 ();
 FILLCELL_X32 FILLER_22_2087 ();
 FILLCELL_X32 FILLER_22_2119 ();
 FILLCELL_X32 FILLER_22_2151 ();
 FILLCELL_X32 FILLER_22_2183 ();
 FILLCELL_X32 FILLER_22_2215 ();
 FILLCELL_X32 FILLER_22_2247 ();
 FILLCELL_X32 FILLER_22_2279 ();
 FILLCELL_X32 FILLER_22_2311 ();
 FILLCELL_X32 FILLER_22_2343 ();
 FILLCELL_X32 FILLER_22_2375 ();
 FILLCELL_X32 FILLER_22_2407 ();
 FILLCELL_X32 FILLER_22_2439 ();
 FILLCELL_X32 FILLER_22_2471 ();
 FILLCELL_X32 FILLER_22_2503 ();
 FILLCELL_X32 FILLER_22_2535 ();
 FILLCELL_X32 FILLER_22_2567 ();
 FILLCELL_X2 FILLER_22_2599 ();
 FILLCELL_X1 FILLER_22_2601 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X32 FILLER_23_225 ();
 FILLCELL_X32 FILLER_23_257 ();
 FILLCELL_X32 FILLER_23_289 ();
 FILLCELL_X32 FILLER_23_321 ();
 FILLCELL_X32 FILLER_23_353 ();
 FILLCELL_X32 FILLER_23_385 ();
 FILLCELL_X32 FILLER_23_417 ();
 FILLCELL_X32 FILLER_23_449 ();
 FILLCELL_X32 FILLER_23_481 ();
 FILLCELL_X32 FILLER_23_513 ();
 FILLCELL_X32 FILLER_23_545 ();
 FILLCELL_X32 FILLER_23_577 ();
 FILLCELL_X32 FILLER_23_609 ();
 FILLCELL_X32 FILLER_23_641 ();
 FILLCELL_X32 FILLER_23_673 ();
 FILLCELL_X32 FILLER_23_705 ();
 FILLCELL_X32 FILLER_23_737 ();
 FILLCELL_X32 FILLER_23_769 ();
 FILLCELL_X32 FILLER_23_801 ();
 FILLCELL_X32 FILLER_23_833 ();
 FILLCELL_X32 FILLER_23_865 ();
 FILLCELL_X32 FILLER_23_897 ();
 FILLCELL_X32 FILLER_23_929 ();
 FILLCELL_X32 FILLER_23_961 ();
 FILLCELL_X32 FILLER_23_993 ();
 FILLCELL_X32 FILLER_23_1025 ();
 FILLCELL_X32 FILLER_23_1057 ();
 FILLCELL_X32 FILLER_23_1089 ();
 FILLCELL_X32 FILLER_23_1121 ();
 FILLCELL_X32 FILLER_23_1153 ();
 FILLCELL_X32 FILLER_23_1185 ();
 FILLCELL_X32 FILLER_23_1217 ();
 FILLCELL_X8 FILLER_23_1249 ();
 FILLCELL_X4 FILLER_23_1257 ();
 FILLCELL_X2 FILLER_23_1261 ();
 FILLCELL_X32 FILLER_23_1264 ();
 FILLCELL_X32 FILLER_23_1296 ();
 FILLCELL_X32 FILLER_23_1328 ();
 FILLCELL_X32 FILLER_23_1360 ();
 FILLCELL_X32 FILLER_23_1392 ();
 FILLCELL_X32 FILLER_23_1424 ();
 FILLCELL_X32 FILLER_23_1456 ();
 FILLCELL_X32 FILLER_23_1488 ();
 FILLCELL_X32 FILLER_23_1520 ();
 FILLCELL_X32 FILLER_23_1552 ();
 FILLCELL_X32 FILLER_23_1584 ();
 FILLCELL_X32 FILLER_23_1616 ();
 FILLCELL_X32 FILLER_23_1648 ();
 FILLCELL_X32 FILLER_23_1680 ();
 FILLCELL_X32 FILLER_23_1712 ();
 FILLCELL_X32 FILLER_23_1744 ();
 FILLCELL_X32 FILLER_23_1776 ();
 FILLCELL_X32 FILLER_23_1808 ();
 FILLCELL_X32 FILLER_23_1840 ();
 FILLCELL_X32 FILLER_23_1872 ();
 FILLCELL_X32 FILLER_23_1904 ();
 FILLCELL_X32 FILLER_23_1936 ();
 FILLCELL_X32 FILLER_23_1968 ();
 FILLCELL_X32 FILLER_23_2000 ();
 FILLCELL_X32 FILLER_23_2032 ();
 FILLCELL_X32 FILLER_23_2064 ();
 FILLCELL_X32 FILLER_23_2096 ();
 FILLCELL_X32 FILLER_23_2128 ();
 FILLCELL_X32 FILLER_23_2160 ();
 FILLCELL_X32 FILLER_23_2192 ();
 FILLCELL_X32 FILLER_23_2224 ();
 FILLCELL_X32 FILLER_23_2256 ();
 FILLCELL_X32 FILLER_23_2288 ();
 FILLCELL_X32 FILLER_23_2320 ();
 FILLCELL_X32 FILLER_23_2352 ();
 FILLCELL_X32 FILLER_23_2384 ();
 FILLCELL_X32 FILLER_23_2416 ();
 FILLCELL_X32 FILLER_23_2448 ();
 FILLCELL_X32 FILLER_23_2480 ();
 FILLCELL_X8 FILLER_23_2512 ();
 FILLCELL_X4 FILLER_23_2520 ();
 FILLCELL_X2 FILLER_23_2524 ();
 FILLCELL_X32 FILLER_23_2527 ();
 FILLCELL_X32 FILLER_23_2559 ();
 FILLCELL_X8 FILLER_23_2591 ();
 FILLCELL_X2 FILLER_23_2599 ();
 FILLCELL_X1 FILLER_23_2601 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X32 FILLER_24_193 ();
 FILLCELL_X32 FILLER_24_225 ();
 FILLCELL_X32 FILLER_24_257 ();
 FILLCELL_X32 FILLER_24_289 ();
 FILLCELL_X32 FILLER_24_321 ();
 FILLCELL_X32 FILLER_24_353 ();
 FILLCELL_X32 FILLER_24_385 ();
 FILLCELL_X32 FILLER_24_417 ();
 FILLCELL_X32 FILLER_24_449 ();
 FILLCELL_X32 FILLER_24_481 ();
 FILLCELL_X32 FILLER_24_513 ();
 FILLCELL_X32 FILLER_24_545 ();
 FILLCELL_X32 FILLER_24_577 ();
 FILLCELL_X16 FILLER_24_609 ();
 FILLCELL_X4 FILLER_24_625 ();
 FILLCELL_X2 FILLER_24_629 ();
 FILLCELL_X32 FILLER_24_632 ();
 FILLCELL_X32 FILLER_24_664 ();
 FILLCELL_X32 FILLER_24_696 ();
 FILLCELL_X32 FILLER_24_728 ();
 FILLCELL_X32 FILLER_24_760 ();
 FILLCELL_X32 FILLER_24_792 ();
 FILLCELL_X32 FILLER_24_824 ();
 FILLCELL_X32 FILLER_24_856 ();
 FILLCELL_X32 FILLER_24_888 ();
 FILLCELL_X32 FILLER_24_920 ();
 FILLCELL_X32 FILLER_24_952 ();
 FILLCELL_X32 FILLER_24_984 ();
 FILLCELL_X32 FILLER_24_1016 ();
 FILLCELL_X32 FILLER_24_1048 ();
 FILLCELL_X32 FILLER_24_1080 ();
 FILLCELL_X32 FILLER_24_1112 ();
 FILLCELL_X32 FILLER_24_1144 ();
 FILLCELL_X32 FILLER_24_1176 ();
 FILLCELL_X32 FILLER_24_1208 ();
 FILLCELL_X32 FILLER_24_1240 ();
 FILLCELL_X32 FILLER_24_1272 ();
 FILLCELL_X32 FILLER_24_1304 ();
 FILLCELL_X32 FILLER_24_1336 ();
 FILLCELL_X32 FILLER_24_1368 ();
 FILLCELL_X32 FILLER_24_1400 ();
 FILLCELL_X32 FILLER_24_1432 ();
 FILLCELL_X32 FILLER_24_1464 ();
 FILLCELL_X32 FILLER_24_1496 ();
 FILLCELL_X32 FILLER_24_1528 ();
 FILLCELL_X32 FILLER_24_1560 ();
 FILLCELL_X32 FILLER_24_1592 ();
 FILLCELL_X32 FILLER_24_1624 ();
 FILLCELL_X32 FILLER_24_1656 ();
 FILLCELL_X32 FILLER_24_1688 ();
 FILLCELL_X32 FILLER_24_1720 ();
 FILLCELL_X32 FILLER_24_1752 ();
 FILLCELL_X32 FILLER_24_1784 ();
 FILLCELL_X32 FILLER_24_1816 ();
 FILLCELL_X32 FILLER_24_1848 ();
 FILLCELL_X8 FILLER_24_1880 ();
 FILLCELL_X4 FILLER_24_1888 ();
 FILLCELL_X2 FILLER_24_1892 ();
 FILLCELL_X32 FILLER_24_1895 ();
 FILLCELL_X32 FILLER_24_1927 ();
 FILLCELL_X32 FILLER_24_1959 ();
 FILLCELL_X32 FILLER_24_1991 ();
 FILLCELL_X32 FILLER_24_2023 ();
 FILLCELL_X32 FILLER_24_2055 ();
 FILLCELL_X32 FILLER_24_2087 ();
 FILLCELL_X32 FILLER_24_2119 ();
 FILLCELL_X32 FILLER_24_2151 ();
 FILLCELL_X32 FILLER_24_2183 ();
 FILLCELL_X32 FILLER_24_2215 ();
 FILLCELL_X32 FILLER_24_2247 ();
 FILLCELL_X32 FILLER_24_2279 ();
 FILLCELL_X32 FILLER_24_2311 ();
 FILLCELL_X32 FILLER_24_2343 ();
 FILLCELL_X32 FILLER_24_2375 ();
 FILLCELL_X32 FILLER_24_2407 ();
 FILLCELL_X32 FILLER_24_2439 ();
 FILLCELL_X32 FILLER_24_2471 ();
 FILLCELL_X32 FILLER_24_2503 ();
 FILLCELL_X32 FILLER_24_2535 ();
 FILLCELL_X32 FILLER_24_2567 ();
 FILLCELL_X2 FILLER_24_2599 ();
 FILLCELL_X1 FILLER_24_2601 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X32 FILLER_25_193 ();
 FILLCELL_X32 FILLER_25_225 ();
 FILLCELL_X32 FILLER_25_257 ();
 FILLCELL_X32 FILLER_25_289 ();
 FILLCELL_X32 FILLER_25_321 ();
 FILLCELL_X32 FILLER_25_353 ();
 FILLCELL_X32 FILLER_25_385 ();
 FILLCELL_X32 FILLER_25_417 ();
 FILLCELL_X32 FILLER_25_449 ();
 FILLCELL_X32 FILLER_25_481 ();
 FILLCELL_X32 FILLER_25_513 ();
 FILLCELL_X32 FILLER_25_545 ();
 FILLCELL_X32 FILLER_25_577 ();
 FILLCELL_X32 FILLER_25_609 ();
 FILLCELL_X32 FILLER_25_641 ();
 FILLCELL_X32 FILLER_25_673 ();
 FILLCELL_X32 FILLER_25_705 ();
 FILLCELL_X32 FILLER_25_737 ();
 FILLCELL_X32 FILLER_25_769 ();
 FILLCELL_X32 FILLER_25_801 ();
 FILLCELL_X32 FILLER_25_833 ();
 FILLCELL_X32 FILLER_25_865 ();
 FILLCELL_X32 FILLER_25_897 ();
 FILLCELL_X32 FILLER_25_929 ();
 FILLCELL_X32 FILLER_25_961 ();
 FILLCELL_X32 FILLER_25_993 ();
 FILLCELL_X32 FILLER_25_1025 ();
 FILLCELL_X32 FILLER_25_1057 ();
 FILLCELL_X32 FILLER_25_1089 ();
 FILLCELL_X32 FILLER_25_1121 ();
 FILLCELL_X32 FILLER_25_1153 ();
 FILLCELL_X32 FILLER_25_1185 ();
 FILLCELL_X32 FILLER_25_1217 ();
 FILLCELL_X8 FILLER_25_1249 ();
 FILLCELL_X4 FILLER_25_1257 ();
 FILLCELL_X2 FILLER_25_1261 ();
 FILLCELL_X32 FILLER_25_1264 ();
 FILLCELL_X32 FILLER_25_1296 ();
 FILLCELL_X32 FILLER_25_1328 ();
 FILLCELL_X32 FILLER_25_1360 ();
 FILLCELL_X32 FILLER_25_1392 ();
 FILLCELL_X32 FILLER_25_1424 ();
 FILLCELL_X32 FILLER_25_1456 ();
 FILLCELL_X32 FILLER_25_1488 ();
 FILLCELL_X32 FILLER_25_1520 ();
 FILLCELL_X32 FILLER_25_1552 ();
 FILLCELL_X32 FILLER_25_1584 ();
 FILLCELL_X32 FILLER_25_1616 ();
 FILLCELL_X32 FILLER_25_1648 ();
 FILLCELL_X32 FILLER_25_1680 ();
 FILLCELL_X32 FILLER_25_1712 ();
 FILLCELL_X32 FILLER_25_1744 ();
 FILLCELL_X32 FILLER_25_1776 ();
 FILLCELL_X32 FILLER_25_1808 ();
 FILLCELL_X32 FILLER_25_1840 ();
 FILLCELL_X32 FILLER_25_1872 ();
 FILLCELL_X32 FILLER_25_1904 ();
 FILLCELL_X32 FILLER_25_1936 ();
 FILLCELL_X32 FILLER_25_1968 ();
 FILLCELL_X32 FILLER_25_2000 ();
 FILLCELL_X32 FILLER_25_2032 ();
 FILLCELL_X32 FILLER_25_2064 ();
 FILLCELL_X32 FILLER_25_2096 ();
 FILLCELL_X32 FILLER_25_2128 ();
 FILLCELL_X32 FILLER_25_2160 ();
 FILLCELL_X32 FILLER_25_2192 ();
 FILLCELL_X32 FILLER_25_2224 ();
 FILLCELL_X32 FILLER_25_2256 ();
 FILLCELL_X32 FILLER_25_2288 ();
 FILLCELL_X32 FILLER_25_2320 ();
 FILLCELL_X32 FILLER_25_2352 ();
 FILLCELL_X32 FILLER_25_2384 ();
 FILLCELL_X32 FILLER_25_2416 ();
 FILLCELL_X32 FILLER_25_2448 ();
 FILLCELL_X32 FILLER_25_2480 ();
 FILLCELL_X8 FILLER_25_2512 ();
 FILLCELL_X4 FILLER_25_2520 ();
 FILLCELL_X2 FILLER_25_2524 ();
 FILLCELL_X32 FILLER_25_2527 ();
 FILLCELL_X32 FILLER_25_2559 ();
 FILLCELL_X8 FILLER_25_2591 ();
 FILLCELL_X2 FILLER_25_2599 ();
 FILLCELL_X1 FILLER_25_2601 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X32 FILLER_26_193 ();
 FILLCELL_X32 FILLER_26_225 ();
 FILLCELL_X32 FILLER_26_257 ();
 FILLCELL_X32 FILLER_26_289 ();
 FILLCELL_X32 FILLER_26_321 ();
 FILLCELL_X32 FILLER_26_353 ();
 FILLCELL_X32 FILLER_26_385 ();
 FILLCELL_X32 FILLER_26_417 ();
 FILLCELL_X32 FILLER_26_449 ();
 FILLCELL_X32 FILLER_26_481 ();
 FILLCELL_X32 FILLER_26_513 ();
 FILLCELL_X32 FILLER_26_545 ();
 FILLCELL_X32 FILLER_26_577 ();
 FILLCELL_X16 FILLER_26_609 ();
 FILLCELL_X4 FILLER_26_625 ();
 FILLCELL_X2 FILLER_26_629 ();
 FILLCELL_X32 FILLER_26_632 ();
 FILLCELL_X32 FILLER_26_664 ();
 FILLCELL_X32 FILLER_26_696 ();
 FILLCELL_X32 FILLER_26_728 ();
 FILLCELL_X32 FILLER_26_760 ();
 FILLCELL_X32 FILLER_26_792 ();
 FILLCELL_X32 FILLER_26_824 ();
 FILLCELL_X32 FILLER_26_856 ();
 FILLCELL_X32 FILLER_26_888 ();
 FILLCELL_X32 FILLER_26_920 ();
 FILLCELL_X32 FILLER_26_952 ();
 FILLCELL_X32 FILLER_26_984 ();
 FILLCELL_X32 FILLER_26_1016 ();
 FILLCELL_X32 FILLER_26_1048 ();
 FILLCELL_X32 FILLER_26_1080 ();
 FILLCELL_X32 FILLER_26_1112 ();
 FILLCELL_X32 FILLER_26_1144 ();
 FILLCELL_X32 FILLER_26_1176 ();
 FILLCELL_X32 FILLER_26_1208 ();
 FILLCELL_X32 FILLER_26_1240 ();
 FILLCELL_X32 FILLER_26_1272 ();
 FILLCELL_X32 FILLER_26_1304 ();
 FILLCELL_X32 FILLER_26_1336 ();
 FILLCELL_X32 FILLER_26_1368 ();
 FILLCELL_X32 FILLER_26_1400 ();
 FILLCELL_X32 FILLER_26_1432 ();
 FILLCELL_X32 FILLER_26_1464 ();
 FILLCELL_X32 FILLER_26_1496 ();
 FILLCELL_X32 FILLER_26_1528 ();
 FILLCELL_X32 FILLER_26_1560 ();
 FILLCELL_X32 FILLER_26_1592 ();
 FILLCELL_X32 FILLER_26_1624 ();
 FILLCELL_X32 FILLER_26_1656 ();
 FILLCELL_X32 FILLER_26_1688 ();
 FILLCELL_X32 FILLER_26_1720 ();
 FILLCELL_X32 FILLER_26_1752 ();
 FILLCELL_X32 FILLER_26_1784 ();
 FILLCELL_X32 FILLER_26_1816 ();
 FILLCELL_X32 FILLER_26_1848 ();
 FILLCELL_X8 FILLER_26_1880 ();
 FILLCELL_X4 FILLER_26_1888 ();
 FILLCELL_X2 FILLER_26_1892 ();
 FILLCELL_X32 FILLER_26_1895 ();
 FILLCELL_X32 FILLER_26_1927 ();
 FILLCELL_X32 FILLER_26_1959 ();
 FILLCELL_X32 FILLER_26_1991 ();
 FILLCELL_X32 FILLER_26_2023 ();
 FILLCELL_X32 FILLER_26_2055 ();
 FILLCELL_X32 FILLER_26_2087 ();
 FILLCELL_X32 FILLER_26_2119 ();
 FILLCELL_X32 FILLER_26_2151 ();
 FILLCELL_X32 FILLER_26_2183 ();
 FILLCELL_X32 FILLER_26_2215 ();
 FILLCELL_X32 FILLER_26_2247 ();
 FILLCELL_X32 FILLER_26_2279 ();
 FILLCELL_X32 FILLER_26_2311 ();
 FILLCELL_X32 FILLER_26_2343 ();
 FILLCELL_X32 FILLER_26_2375 ();
 FILLCELL_X32 FILLER_26_2407 ();
 FILLCELL_X32 FILLER_26_2439 ();
 FILLCELL_X32 FILLER_26_2471 ();
 FILLCELL_X32 FILLER_26_2503 ();
 FILLCELL_X32 FILLER_26_2535 ();
 FILLCELL_X32 FILLER_26_2567 ();
 FILLCELL_X2 FILLER_26_2599 ();
 FILLCELL_X1 FILLER_26_2601 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X32 FILLER_27_225 ();
 FILLCELL_X32 FILLER_27_257 ();
 FILLCELL_X32 FILLER_27_289 ();
 FILLCELL_X32 FILLER_27_321 ();
 FILLCELL_X32 FILLER_27_353 ();
 FILLCELL_X32 FILLER_27_385 ();
 FILLCELL_X32 FILLER_27_417 ();
 FILLCELL_X32 FILLER_27_449 ();
 FILLCELL_X32 FILLER_27_481 ();
 FILLCELL_X32 FILLER_27_513 ();
 FILLCELL_X32 FILLER_27_545 ();
 FILLCELL_X32 FILLER_27_577 ();
 FILLCELL_X32 FILLER_27_609 ();
 FILLCELL_X32 FILLER_27_641 ();
 FILLCELL_X32 FILLER_27_673 ();
 FILLCELL_X32 FILLER_27_705 ();
 FILLCELL_X32 FILLER_27_737 ();
 FILLCELL_X32 FILLER_27_769 ();
 FILLCELL_X32 FILLER_27_801 ();
 FILLCELL_X32 FILLER_27_833 ();
 FILLCELL_X32 FILLER_27_865 ();
 FILLCELL_X32 FILLER_27_897 ();
 FILLCELL_X32 FILLER_27_929 ();
 FILLCELL_X32 FILLER_27_961 ();
 FILLCELL_X32 FILLER_27_993 ();
 FILLCELL_X32 FILLER_27_1025 ();
 FILLCELL_X32 FILLER_27_1057 ();
 FILLCELL_X32 FILLER_27_1089 ();
 FILLCELL_X32 FILLER_27_1121 ();
 FILLCELL_X32 FILLER_27_1153 ();
 FILLCELL_X32 FILLER_27_1185 ();
 FILLCELL_X32 FILLER_27_1217 ();
 FILLCELL_X8 FILLER_27_1249 ();
 FILLCELL_X4 FILLER_27_1257 ();
 FILLCELL_X2 FILLER_27_1261 ();
 FILLCELL_X32 FILLER_27_1264 ();
 FILLCELL_X32 FILLER_27_1296 ();
 FILLCELL_X32 FILLER_27_1328 ();
 FILLCELL_X32 FILLER_27_1360 ();
 FILLCELL_X32 FILLER_27_1392 ();
 FILLCELL_X32 FILLER_27_1424 ();
 FILLCELL_X32 FILLER_27_1456 ();
 FILLCELL_X32 FILLER_27_1488 ();
 FILLCELL_X32 FILLER_27_1520 ();
 FILLCELL_X32 FILLER_27_1552 ();
 FILLCELL_X32 FILLER_27_1584 ();
 FILLCELL_X32 FILLER_27_1616 ();
 FILLCELL_X32 FILLER_27_1648 ();
 FILLCELL_X32 FILLER_27_1680 ();
 FILLCELL_X32 FILLER_27_1712 ();
 FILLCELL_X32 FILLER_27_1744 ();
 FILLCELL_X32 FILLER_27_1776 ();
 FILLCELL_X32 FILLER_27_1808 ();
 FILLCELL_X32 FILLER_27_1840 ();
 FILLCELL_X32 FILLER_27_1872 ();
 FILLCELL_X32 FILLER_27_1904 ();
 FILLCELL_X32 FILLER_27_1936 ();
 FILLCELL_X32 FILLER_27_1968 ();
 FILLCELL_X32 FILLER_27_2000 ();
 FILLCELL_X32 FILLER_27_2032 ();
 FILLCELL_X32 FILLER_27_2064 ();
 FILLCELL_X32 FILLER_27_2096 ();
 FILLCELL_X32 FILLER_27_2128 ();
 FILLCELL_X32 FILLER_27_2160 ();
 FILLCELL_X32 FILLER_27_2192 ();
 FILLCELL_X32 FILLER_27_2224 ();
 FILLCELL_X32 FILLER_27_2256 ();
 FILLCELL_X32 FILLER_27_2288 ();
 FILLCELL_X32 FILLER_27_2320 ();
 FILLCELL_X32 FILLER_27_2352 ();
 FILLCELL_X32 FILLER_27_2384 ();
 FILLCELL_X32 FILLER_27_2416 ();
 FILLCELL_X32 FILLER_27_2448 ();
 FILLCELL_X32 FILLER_27_2480 ();
 FILLCELL_X8 FILLER_27_2512 ();
 FILLCELL_X4 FILLER_27_2520 ();
 FILLCELL_X2 FILLER_27_2524 ();
 FILLCELL_X32 FILLER_27_2527 ();
 FILLCELL_X32 FILLER_27_2559 ();
 FILLCELL_X8 FILLER_27_2591 ();
 FILLCELL_X2 FILLER_27_2599 ();
 FILLCELL_X1 FILLER_27_2601 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X32 FILLER_28_225 ();
 FILLCELL_X32 FILLER_28_257 ();
 FILLCELL_X32 FILLER_28_289 ();
 FILLCELL_X32 FILLER_28_321 ();
 FILLCELL_X32 FILLER_28_353 ();
 FILLCELL_X32 FILLER_28_385 ();
 FILLCELL_X32 FILLER_28_417 ();
 FILLCELL_X32 FILLER_28_449 ();
 FILLCELL_X32 FILLER_28_481 ();
 FILLCELL_X32 FILLER_28_513 ();
 FILLCELL_X32 FILLER_28_545 ();
 FILLCELL_X32 FILLER_28_577 ();
 FILLCELL_X16 FILLER_28_609 ();
 FILLCELL_X4 FILLER_28_625 ();
 FILLCELL_X2 FILLER_28_629 ();
 FILLCELL_X32 FILLER_28_632 ();
 FILLCELL_X32 FILLER_28_664 ();
 FILLCELL_X32 FILLER_28_696 ();
 FILLCELL_X32 FILLER_28_728 ();
 FILLCELL_X32 FILLER_28_760 ();
 FILLCELL_X32 FILLER_28_792 ();
 FILLCELL_X32 FILLER_28_824 ();
 FILLCELL_X32 FILLER_28_856 ();
 FILLCELL_X32 FILLER_28_888 ();
 FILLCELL_X32 FILLER_28_920 ();
 FILLCELL_X32 FILLER_28_952 ();
 FILLCELL_X32 FILLER_28_984 ();
 FILLCELL_X32 FILLER_28_1016 ();
 FILLCELL_X32 FILLER_28_1048 ();
 FILLCELL_X32 FILLER_28_1080 ();
 FILLCELL_X32 FILLER_28_1112 ();
 FILLCELL_X32 FILLER_28_1144 ();
 FILLCELL_X32 FILLER_28_1176 ();
 FILLCELL_X32 FILLER_28_1208 ();
 FILLCELL_X32 FILLER_28_1240 ();
 FILLCELL_X32 FILLER_28_1272 ();
 FILLCELL_X32 FILLER_28_1304 ();
 FILLCELL_X32 FILLER_28_1336 ();
 FILLCELL_X32 FILLER_28_1368 ();
 FILLCELL_X32 FILLER_28_1400 ();
 FILLCELL_X32 FILLER_28_1432 ();
 FILLCELL_X32 FILLER_28_1464 ();
 FILLCELL_X32 FILLER_28_1496 ();
 FILLCELL_X32 FILLER_28_1528 ();
 FILLCELL_X32 FILLER_28_1560 ();
 FILLCELL_X32 FILLER_28_1592 ();
 FILLCELL_X32 FILLER_28_1624 ();
 FILLCELL_X32 FILLER_28_1656 ();
 FILLCELL_X32 FILLER_28_1688 ();
 FILLCELL_X32 FILLER_28_1720 ();
 FILLCELL_X32 FILLER_28_1752 ();
 FILLCELL_X32 FILLER_28_1784 ();
 FILLCELL_X32 FILLER_28_1816 ();
 FILLCELL_X32 FILLER_28_1848 ();
 FILLCELL_X8 FILLER_28_1880 ();
 FILLCELL_X4 FILLER_28_1888 ();
 FILLCELL_X2 FILLER_28_1892 ();
 FILLCELL_X32 FILLER_28_1895 ();
 FILLCELL_X32 FILLER_28_1927 ();
 FILLCELL_X32 FILLER_28_1959 ();
 FILLCELL_X32 FILLER_28_1991 ();
 FILLCELL_X32 FILLER_28_2023 ();
 FILLCELL_X32 FILLER_28_2055 ();
 FILLCELL_X32 FILLER_28_2087 ();
 FILLCELL_X32 FILLER_28_2119 ();
 FILLCELL_X32 FILLER_28_2151 ();
 FILLCELL_X32 FILLER_28_2183 ();
 FILLCELL_X32 FILLER_28_2215 ();
 FILLCELL_X32 FILLER_28_2247 ();
 FILLCELL_X32 FILLER_28_2279 ();
 FILLCELL_X32 FILLER_28_2311 ();
 FILLCELL_X32 FILLER_28_2343 ();
 FILLCELL_X32 FILLER_28_2375 ();
 FILLCELL_X32 FILLER_28_2407 ();
 FILLCELL_X32 FILLER_28_2439 ();
 FILLCELL_X32 FILLER_28_2471 ();
 FILLCELL_X32 FILLER_28_2503 ();
 FILLCELL_X32 FILLER_28_2535 ();
 FILLCELL_X32 FILLER_28_2567 ();
 FILLCELL_X2 FILLER_28_2599 ();
 FILLCELL_X1 FILLER_28_2601 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X32 FILLER_29_225 ();
 FILLCELL_X32 FILLER_29_257 ();
 FILLCELL_X32 FILLER_29_289 ();
 FILLCELL_X32 FILLER_29_321 ();
 FILLCELL_X32 FILLER_29_353 ();
 FILLCELL_X32 FILLER_29_385 ();
 FILLCELL_X32 FILLER_29_417 ();
 FILLCELL_X32 FILLER_29_449 ();
 FILLCELL_X32 FILLER_29_481 ();
 FILLCELL_X32 FILLER_29_513 ();
 FILLCELL_X32 FILLER_29_545 ();
 FILLCELL_X32 FILLER_29_577 ();
 FILLCELL_X32 FILLER_29_609 ();
 FILLCELL_X32 FILLER_29_641 ();
 FILLCELL_X32 FILLER_29_673 ();
 FILLCELL_X32 FILLER_29_705 ();
 FILLCELL_X32 FILLER_29_737 ();
 FILLCELL_X32 FILLER_29_769 ();
 FILLCELL_X32 FILLER_29_801 ();
 FILLCELL_X32 FILLER_29_833 ();
 FILLCELL_X32 FILLER_29_865 ();
 FILLCELL_X32 FILLER_29_897 ();
 FILLCELL_X32 FILLER_29_929 ();
 FILLCELL_X32 FILLER_29_961 ();
 FILLCELL_X32 FILLER_29_993 ();
 FILLCELL_X32 FILLER_29_1025 ();
 FILLCELL_X32 FILLER_29_1057 ();
 FILLCELL_X32 FILLER_29_1089 ();
 FILLCELL_X32 FILLER_29_1121 ();
 FILLCELL_X32 FILLER_29_1153 ();
 FILLCELL_X32 FILLER_29_1185 ();
 FILLCELL_X32 FILLER_29_1217 ();
 FILLCELL_X8 FILLER_29_1249 ();
 FILLCELL_X4 FILLER_29_1257 ();
 FILLCELL_X2 FILLER_29_1261 ();
 FILLCELL_X32 FILLER_29_1264 ();
 FILLCELL_X32 FILLER_29_1296 ();
 FILLCELL_X32 FILLER_29_1328 ();
 FILLCELL_X32 FILLER_29_1360 ();
 FILLCELL_X32 FILLER_29_1392 ();
 FILLCELL_X32 FILLER_29_1424 ();
 FILLCELL_X32 FILLER_29_1456 ();
 FILLCELL_X32 FILLER_29_1488 ();
 FILLCELL_X32 FILLER_29_1520 ();
 FILLCELL_X32 FILLER_29_1552 ();
 FILLCELL_X32 FILLER_29_1584 ();
 FILLCELL_X32 FILLER_29_1616 ();
 FILLCELL_X32 FILLER_29_1648 ();
 FILLCELL_X32 FILLER_29_1680 ();
 FILLCELL_X32 FILLER_29_1712 ();
 FILLCELL_X32 FILLER_29_1744 ();
 FILLCELL_X32 FILLER_29_1776 ();
 FILLCELL_X32 FILLER_29_1808 ();
 FILLCELL_X32 FILLER_29_1840 ();
 FILLCELL_X32 FILLER_29_1872 ();
 FILLCELL_X32 FILLER_29_1904 ();
 FILLCELL_X32 FILLER_29_1936 ();
 FILLCELL_X32 FILLER_29_1968 ();
 FILLCELL_X32 FILLER_29_2000 ();
 FILLCELL_X32 FILLER_29_2032 ();
 FILLCELL_X32 FILLER_29_2064 ();
 FILLCELL_X32 FILLER_29_2096 ();
 FILLCELL_X32 FILLER_29_2128 ();
 FILLCELL_X32 FILLER_29_2160 ();
 FILLCELL_X32 FILLER_29_2192 ();
 FILLCELL_X32 FILLER_29_2224 ();
 FILLCELL_X32 FILLER_29_2256 ();
 FILLCELL_X32 FILLER_29_2288 ();
 FILLCELL_X32 FILLER_29_2320 ();
 FILLCELL_X32 FILLER_29_2352 ();
 FILLCELL_X32 FILLER_29_2384 ();
 FILLCELL_X32 FILLER_29_2416 ();
 FILLCELL_X32 FILLER_29_2448 ();
 FILLCELL_X32 FILLER_29_2480 ();
 FILLCELL_X8 FILLER_29_2512 ();
 FILLCELL_X4 FILLER_29_2520 ();
 FILLCELL_X2 FILLER_29_2524 ();
 FILLCELL_X32 FILLER_29_2527 ();
 FILLCELL_X32 FILLER_29_2559 ();
 FILLCELL_X8 FILLER_29_2591 ();
 FILLCELL_X2 FILLER_29_2599 ();
 FILLCELL_X1 FILLER_29_2601 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X32 FILLER_30_225 ();
 FILLCELL_X32 FILLER_30_257 ();
 FILLCELL_X32 FILLER_30_289 ();
 FILLCELL_X32 FILLER_30_321 ();
 FILLCELL_X32 FILLER_30_353 ();
 FILLCELL_X32 FILLER_30_385 ();
 FILLCELL_X32 FILLER_30_417 ();
 FILLCELL_X32 FILLER_30_449 ();
 FILLCELL_X32 FILLER_30_481 ();
 FILLCELL_X32 FILLER_30_513 ();
 FILLCELL_X32 FILLER_30_545 ();
 FILLCELL_X32 FILLER_30_577 ();
 FILLCELL_X16 FILLER_30_609 ();
 FILLCELL_X4 FILLER_30_625 ();
 FILLCELL_X2 FILLER_30_629 ();
 FILLCELL_X32 FILLER_30_632 ();
 FILLCELL_X32 FILLER_30_664 ();
 FILLCELL_X32 FILLER_30_696 ();
 FILLCELL_X32 FILLER_30_728 ();
 FILLCELL_X32 FILLER_30_760 ();
 FILLCELL_X32 FILLER_30_792 ();
 FILLCELL_X32 FILLER_30_824 ();
 FILLCELL_X32 FILLER_30_856 ();
 FILLCELL_X32 FILLER_30_888 ();
 FILLCELL_X32 FILLER_30_920 ();
 FILLCELL_X32 FILLER_30_952 ();
 FILLCELL_X32 FILLER_30_984 ();
 FILLCELL_X32 FILLER_30_1016 ();
 FILLCELL_X32 FILLER_30_1048 ();
 FILLCELL_X32 FILLER_30_1080 ();
 FILLCELL_X32 FILLER_30_1112 ();
 FILLCELL_X32 FILLER_30_1144 ();
 FILLCELL_X32 FILLER_30_1176 ();
 FILLCELL_X32 FILLER_30_1208 ();
 FILLCELL_X32 FILLER_30_1240 ();
 FILLCELL_X32 FILLER_30_1272 ();
 FILLCELL_X32 FILLER_30_1304 ();
 FILLCELL_X32 FILLER_30_1336 ();
 FILLCELL_X32 FILLER_30_1368 ();
 FILLCELL_X32 FILLER_30_1400 ();
 FILLCELL_X32 FILLER_30_1432 ();
 FILLCELL_X32 FILLER_30_1464 ();
 FILLCELL_X32 FILLER_30_1496 ();
 FILLCELL_X32 FILLER_30_1528 ();
 FILLCELL_X32 FILLER_30_1560 ();
 FILLCELL_X32 FILLER_30_1592 ();
 FILLCELL_X32 FILLER_30_1624 ();
 FILLCELL_X32 FILLER_30_1656 ();
 FILLCELL_X32 FILLER_30_1688 ();
 FILLCELL_X32 FILLER_30_1720 ();
 FILLCELL_X32 FILLER_30_1752 ();
 FILLCELL_X32 FILLER_30_1784 ();
 FILLCELL_X32 FILLER_30_1816 ();
 FILLCELL_X32 FILLER_30_1848 ();
 FILLCELL_X8 FILLER_30_1880 ();
 FILLCELL_X4 FILLER_30_1888 ();
 FILLCELL_X2 FILLER_30_1892 ();
 FILLCELL_X32 FILLER_30_1895 ();
 FILLCELL_X32 FILLER_30_1927 ();
 FILLCELL_X32 FILLER_30_1959 ();
 FILLCELL_X32 FILLER_30_1991 ();
 FILLCELL_X32 FILLER_30_2023 ();
 FILLCELL_X32 FILLER_30_2055 ();
 FILLCELL_X32 FILLER_30_2087 ();
 FILLCELL_X32 FILLER_30_2119 ();
 FILLCELL_X32 FILLER_30_2151 ();
 FILLCELL_X32 FILLER_30_2183 ();
 FILLCELL_X32 FILLER_30_2215 ();
 FILLCELL_X32 FILLER_30_2247 ();
 FILLCELL_X32 FILLER_30_2279 ();
 FILLCELL_X32 FILLER_30_2311 ();
 FILLCELL_X32 FILLER_30_2343 ();
 FILLCELL_X32 FILLER_30_2375 ();
 FILLCELL_X32 FILLER_30_2407 ();
 FILLCELL_X32 FILLER_30_2439 ();
 FILLCELL_X32 FILLER_30_2471 ();
 FILLCELL_X32 FILLER_30_2503 ();
 FILLCELL_X32 FILLER_30_2535 ();
 FILLCELL_X32 FILLER_30_2567 ();
 FILLCELL_X2 FILLER_30_2599 ();
 FILLCELL_X1 FILLER_30_2601 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X32 FILLER_31_193 ();
 FILLCELL_X32 FILLER_31_225 ();
 FILLCELL_X32 FILLER_31_257 ();
 FILLCELL_X32 FILLER_31_289 ();
 FILLCELL_X32 FILLER_31_321 ();
 FILLCELL_X32 FILLER_31_353 ();
 FILLCELL_X32 FILLER_31_385 ();
 FILLCELL_X32 FILLER_31_417 ();
 FILLCELL_X32 FILLER_31_449 ();
 FILLCELL_X32 FILLER_31_481 ();
 FILLCELL_X32 FILLER_31_513 ();
 FILLCELL_X32 FILLER_31_545 ();
 FILLCELL_X32 FILLER_31_577 ();
 FILLCELL_X32 FILLER_31_609 ();
 FILLCELL_X32 FILLER_31_641 ();
 FILLCELL_X32 FILLER_31_673 ();
 FILLCELL_X32 FILLER_31_705 ();
 FILLCELL_X32 FILLER_31_737 ();
 FILLCELL_X32 FILLER_31_769 ();
 FILLCELL_X32 FILLER_31_801 ();
 FILLCELL_X32 FILLER_31_833 ();
 FILLCELL_X32 FILLER_31_865 ();
 FILLCELL_X32 FILLER_31_897 ();
 FILLCELL_X32 FILLER_31_929 ();
 FILLCELL_X32 FILLER_31_961 ();
 FILLCELL_X32 FILLER_31_993 ();
 FILLCELL_X32 FILLER_31_1025 ();
 FILLCELL_X32 FILLER_31_1057 ();
 FILLCELL_X32 FILLER_31_1089 ();
 FILLCELL_X32 FILLER_31_1121 ();
 FILLCELL_X32 FILLER_31_1153 ();
 FILLCELL_X32 FILLER_31_1185 ();
 FILLCELL_X32 FILLER_31_1217 ();
 FILLCELL_X8 FILLER_31_1249 ();
 FILLCELL_X4 FILLER_31_1257 ();
 FILLCELL_X2 FILLER_31_1261 ();
 FILLCELL_X32 FILLER_31_1264 ();
 FILLCELL_X32 FILLER_31_1296 ();
 FILLCELL_X32 FILLER_31_1328 ();
 FILLCELL_X32 FILLER_31_1360 ();
 FILLCELL_X32 FILLER_31_1392 ();
 FILLCELL_X32 FILLER_31_1424 ();
 FILLCELL_X32 FILLER_31_1456 ();
 FILLCELL_X32 FILLER_31_1488 ();
 FILLCELL_X32 FILLER_31_1520 ();
 FILLCELL_X32 FILLER_31_1552 ();
 FILLCELL_X32 FILLER_31_1584 ();
 FILLCELL_X32 FILLER_31_1616 ();
 FILLCELL_X32 FILLER_31_1648 ();
 FILLCELL_X32 FILLER_31_1680 ();
 FILLCELL_X32 FILLER_31_1712 ();
 FILLCELL_X32 FILLER_31_1744 ();
 FILLCELL_X32 FILLER_31_1776 ();
 FILLCELL_X32 FILLER_31_1808 ();
 FILLCELL_X32 FILLER_31_1840 ();
 FILLCELL_X32 FILLER_31_1872 ();
 FILLCELL_X32 FILLER_31_1904 ();
 FILLCELL_X32 FILLER_31_1936 ();
 FILLCELL_X32 FILLER_31_1968 ();
 FILLCELL_X32 FILLER_31_2000 ();
 FILLCELL_X32 FILLER_31_2032 ();
 FILLCELL_X32 FILLER_31_2064 ();
 FILLCELL_X32 FILLER_31_2096 ();
 FILLCELL_X32 FILLER_31_2128 ();
 FILLCELL_X32 FILLER_31_2160 ();
 FILLCELL_X32 FILLER_31_2192 ();
 FILLCELL_X32 FILLER_31_2224 ();
 FILLCELL_X32 FILLER_31_2256 ();
 FILLCELL_X32 FILLER_31_2288 ();
 FILLCELL_X32 FILLER_31_2320 ();
 FILLCELL_X32 FILLER_31_2352 ();
 FILLCELL_X32 FILLER_31_2384 ();
 FILLCELL_X32 FILLER_31_2416 ();
 FILLCELL_X32 FILLER_31_2448 ();
 FILLCELL_X32 FILLER_31_2480 ();
 FILLCELL_X8 FILLER_31_2512 ();
 FILLCELL_X4 FILLER_31_2520 ();
 FILLCELL_X2 FILLER_31_2524 ();
 FILLCELL_X32 FILLER_31_2527 ();
 FILLCELL_X32 FILLER_31_2559 ();
 FILLCELL_X8 FILLER_31_2591 ();
 FILLCELL_X2 FILLER_31_2599 ();
 FILLCELL_X1 FILLER_31_2601 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X32 FILLER_32_257 ();
 FILLCELL_X32 FILLER_32_289 ();
 FILLCELL_X32 FILLER_32_321 ();
 FILLCELL_X32 FILLER_32_353 ();
 FILLCELL_X32 FILLER_32_385 ();
 FILLCELL_X32 FILLER_32_417 ();
 FILLCELL_X32 FILLER_32_449 ();
 FILLCELL_X32 FILLER_32_481 ();
 FILLCELL_X32 FILLER_32_513 ();
 FILLCELL_X32 FILLER_32_545 ();
 FILLCELL_X32 FILLER_32_577 ();
 FILLCELL_X16 FILLER_32_609 ();
 FILLCELL_X4 FILLER_32_625 ();
 FILLCELL_X2 FILLER_32_629 ();
 FILLCELL_X32 FILLER_32_632 ();
 FILLCELL_X32 FILLER_32_664 ();
 FILLCELL_X32 FILLER_32_696 ();
 FILLCELL_X32 FILLER_32_728 ();
 FILLCELL_X32 FILLER_32_760 ();
 FILLCELL_X32 FILLER_32_792 ();
 FILLCELL_X32 FILLER_32_824 ();
 FILLCELL_X32 FILLER_32_856 ();
 FILLCELL_X32 FILLER_32_888 ();
 FILLCELL_X32 FILLER_32_920 ();
 FILLCELL_X32 FILLER_32_952 ();
 FILLCELL_X32 FILLER_32_984 ();
 FILLCELL_X32 FILLER_32_1016 ();
 FILLCELL_X32 FILLER_32_1048 ();
 FILLCELL_X32 FILLER_32_1080 ();
 FILLCELL_X32 FILLER_32_1112 ();
 FILLCELL_X32 FILLER_32_1144 ();
 FILLCELL_X32 FILLER_32_1176 ();
 FILLCELL_X32 FILLER_32_1208 ();
 FILLCELL_X32 FILLER_32_1240 ();
 FILLCELL_X32 FILLER_32_1272 ();
 FILLCELL_X32 FILLER_32_1304 ();
 FILLCELL_X32 FILLER_32_1336 ();
 FILLCELL_X32 FILLER_32_1368 ();
 FILLCELL_X32 FILLER_32_1400 ();
 FILLCELL_X32 FILLER_32_1432 ();
 FILLCELL_X32 FILLER_32_1464 ();
 FILLCELL_X32 FILLER_32_1496 ();
 FILLCELL_X32 FILLER_32_1528 ();
 FILLCELL_X32 FILLER_32_1560 ();
 FILLCELL_X32 FILLER_32_1592 ();
 FILLCELL_X32 FILLER_32_1624 ();
 FILLCELL_X32 FILLER_32_1656 ();
 FILLCELL_X32 FILLER_32_1688 ();
 FILLCELL_X32 FILLER_32_1720 ();
 FILLCELL_X32 FILLER_32_1752 ();
 FILLCELL_X32 FILLER_32_1784 ();
 FILLCELL_X32 FILLER_32_1816 ();
 FILLCELL_X32 FILLER_32_1848 ();
 FILLCELL_X8 FILLER_32_1880 ();
 FILLCELL_X4 FILLER_32_1888 ();
 FILLCELL_X2 FILLER_32_1892 ();
 FILLCELL_X32 FILLER_32_1895 ();
 FILLCELL_X32 FILLER_32_1927 ();
 FILLCELL_X32 FILLER_32_1959 ();
 FILLCELL_X32 FILLER_32_1991 ();
 FILLCELL_X32 FILLER_32_2023 ();
 FILLCELL_X32 FILLER_32_2055 ();
 FILLCELL_X32 FILLER_32_2087 ();
 FILLCELL_X32 FILLER_32_2119 ();
 FILLCELL_X32 FILLER_32_2151 ();
 FILLCELL_X32 FILLER_32_2183 ();
 FILLCELL_X32 FILLER_32_2215 ();
 FILLCELL_X32 FILLER_32_2247 ();
 FILLCELL_X32 FILLER_32_2279 ();
 FILLCELL_X32 FILLER_32_2311 ();
 FILLCELL_X32 FILLER_32_2343 ();
 FILLCELL_X32 FILLER_32_2375 ();
 FILLCELL_X32 FILLER_32_2407 ();
 FILLCELL_X32 FILLER_32_2439 ();
 FILLCELL_X32 FILLER_32_2471 ();
 FILLCELL_X32 FILLER_32_2503 ();
 FILLCELL_X32 FILLER_32_2535 ();
 FILLCELL_X32 FILLER_32_2567 ();
 FILLCELL_X2 FILLER_32_2599 ();
 FILLCELL_X1 FILLER_32_2601 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_225 ();
 FILLCELL_X32 FILLER_33_257 ();
 FILLCELL_X32 FILLER_33_289 ();
 FILLCELL_X32 FILLER_33_321 ();
 FILLCELL_X32 FILLER_33_353 ();
 FILLCELL_X32 FILLER_33_385 ();
 FILLCELL_X32 FILLER_33_417 ();
 FILLCELL_X32 FILLER_33_449 ();
 FILLCELL_X32 FILLER_33_481 ();
 FILLCELL_X32 FILLER_33_513 ();
 FILLCELL_X32 FILLER_33_545 ();
 FILLCELL_X32 FILLER_33_577 ();
 FILLCELL_X32 FILLER_33_609 ();
 FILLCELL_X32 FILLER_33_641 ();
 FILLCELL_X32 FILLER_33_673 ();
 FILLCELL_X32 FILLER_33_705 ();
 FILLCELL_X32 FILLER_33_737 ();
 FILLCELL_X32 FILLER_33_769 ();
 FILLCELL_X32 FILLER_33_801 ();
 FILLCELL_X32 FILLER_33_833 ();
 FILLCELL_X32 FILLER_33_865 ();
 FILLCELL_X32 FILLER_33_897 ();
 FILLCELL_X32 FILLER_33_929 ();
 FILLCELL_X32 FILLER_33_961 ();
 FILLCELL_X32 FILLER_33_993 ();
 FILLCELL_X32 FILLER_33_1025 ();
 FILLCELL_X32 FILLER_33_1057 ();
 FILLCELL_X32 FILLER_33_1089 ();
 FILLCELL_X32 FILLER_33_1121 ();
 FILLCELL_X32 FILLER_33_1153 ();
 FILLCELL_X32 FILLER_33_1185 ();
 FILLCELL_X32 FILLER_33_1217 ();
 FILLCELL_X8 FILLER_33_1249 ();
 FILLCELL_X4 FILLER_33_1257 ();
 FILLCELL_X2 FILLER_33_1261 ();
 FILLCELL_X32 FILLER_33_1264 ();
 FILLCELL_X32 FILLER_33_1296 ();
 FILLCELL_X32 FILLER_33_1328 ();
 FILLCELL_X32 FILLER_33_1360 ();
 FILLCELL_X32 FILLER_33_1392 ();
 FILLCELL_X32 FILLER_33_1424 ();
 FILLCELL_X32 FILLER_33_1456 ();
 FILLCELL_X32 FILLER_33_1488 ();
 FILLCELL_X32 FILLER_33_1520 ();
 FILLCELL_X32 FILLER_33_1552 ();
 FILLCELL_X32 FILLER_33_1584 ();
 FILLCELL_X32 FILLER_33_1616 ();
 FILLCELL_X32 FILLER_33_1648 ();
 FILLCELL_X32 FILLER_33_1680 ();
 FILLCELL_X32 FILLER_33_1712 ();
 FILLCELL_X32 FILLER_33_1744 ();
 FILLCELL_X32 FILLER_33_1776 ();
 FILLCELL_X32 FILLER_33_1808 ();
 FILLCELL_X32 FILLER_33_1840 ();
 FILLCELL_X32 FILLER_33_1872 ();
 FILLCELL_X32 FILLER_33_1904 ();
 FILLCELL_X32 FILLER_33_1936 ();
 FILLCELL_X32 FILLER_33_1968 ();
 FILLCELL_X32 FILLER_33_2000 ();
 FILLCELL_X32 FILLER_33_2032 ();
 FILLCELL_X32 FILLER_33_2064 ();
 FILLCELL_X32 FILLER_33_2096 ();
 FILLCELL_X32 FILLER_33_2128 ();
 FILLCELL_X32 FILLER_33_2160 ();
 FILLCELL_X32 FILLER_33_2192 ();
 FILLCELL_X32 FILLER_33_2224 ();
 FILLCELL_X32 FILLER_33_2256 ();
 FILLCELL_X32 FILLER_33_2288 ();
 FILLCELL_X32 FILLER_33_2320 ();
 FILLCELL_X32 FILLER_33_2352 ();
 FILLCELL_X32 FILLER_33_2384 ();
 FILLCELL_X32 FILLER_33_2416 ();
 FILLCELL_X32 FILLER_33_2448 ();
 FILLCELL_X32 FILLER_33_2480 ();
 FILLCELL_X8 FILLER_33_2512 ();
 FILLCELL_X4 FILLER_33_2520 ();
 FILLCELL_X2 FILLER_33_2524 ();
 FILLCELL_X32 FILLER_33_2527 ();
 FILLCELL_X32 FILLER_33_2559 ();
 FILLCELL_X8 FILLER_33_2591 ();
 FILLCELL_X2 FILLER_33_2599 ();
 FILLCELL_X1 FILLER_33_2601 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X32 FILLER_34_161 ();
 FILLCELL_X32 FILLER_34_193 ();
 FILLCELL_X32 FILLER_34_225 ();
 FILLCELL_X32 FILLER_34_257 ();
 FILLCELL_X32 FILLER_34_289 ();
 FILLCELL_X32 FILLER_34_321 ();
 FILLCELL_X32 FILLER_34_353 ();
 FILLCELL_X32 FILLER_34_385 ();
 FILLCELL_X32 FILLER_34_417 ();
 FILLCELL_X32 FILLER_34_449 ();
 FILLCELL_X32 FILLER_34_481 ();
 FILLCELL_X32 FILLER_34_513 ();
 FILLCELL_X32 FILLER_34_545 ();
 FILLCELL_X32 FILLER_34_577 ();
 FILLCELL_X16 FILLER_34_609 ();
 FILLCELL_X4 FILLER_34_625 ();
 FILLCELL_X2 FILLER_34_629 ();
 FILLCELL_X32 FILLER_34_632 ();
 FILLCELL_X32 FILLER_34_664 ();
 FILLCELL_X32 FILLER_34_696 ();
 FILLCELL_X32 FILLER_34_728 ();
 FILLCELL_X32 FILLER_34_760 ();
 FILLCELL_X32 FILLER_34_792 ();
 FILLCELL_X32 FILLER_34_824 ();
 FILLCELL_X32 FILLER_34_856 ();
 FILLCELL_X32 FILLER_34_888 ();
 FILLCELL_X32 FILLER_34_920 ();
 FILLCELL_X32 FILLER_34_952 ();
 FILLCELL_X32 FILLER_34_984 ();
 FILLCELL_X32 FILLER_34_1016 ();
 FILLCELL_X32 FILLER_34_1048 ();
 FILLCELL_X32 FILLER_34_1080 ();
 FILLCELL_X32 FILLER_34_1112 ();
 FILLCELL_X32 FILLER_34_1144 ();
 FILLCELL_X32 FILLER_34_1176 ();
 FILLCELL_X32 FILLER_34_1208 ();
 FILLCELL_X32 FILLER_34_1240 ();
 FILLCELL_X32 FILLER_34_1272 ();
 FILLCELL_X32 FILLER_34_1304 ();
 FILLCELL_X32 FILLER_34_1336 ();
 FILLCELL_X32 FILLER_34_1368 ();
 FILLCELL_X32 FILLER_34_1400 ();
 FILLCELL_X32 FILLER_34_1432 ();
 FILLCELL_X32 FILLER_34_1464 ();
 FILLCELL_X32 FILLER_34_1496 ();
 FILLCELL_X32 FILLER_34_1528 ();
 FILLCELL_X32 FILLER_34_1560 ();
 FILLCELL_X32 FILLER_34_1592 ();
 FILLCELL_X32 FILLER_34_1624 ();
 FILLCELL_X32 FILLER_34_1656 ();
 FILLCELL_X32 FILLER_34_1688 ();
 FILLCELL_X32 FILLER_34_1720 ();
 FILLCELL_X32 FILLER_34_1752 ();
 FILLCELL_X32 FILLER_34_1784 ();
 FILLCELL_X32 FILLER_34_1816 ();
 FILLCELL_X32 FILLER_34_1848 ();
 FILLCELL_X8 FILLER_34_1880 ();
 FILLCELL_X4 FILLER_34_1888 ();
 FILLCELL_X2 FILLER_34_1892 ();
 FILLCELL_X32 FILLER_34_1895 ();
 FILLCELL_X32 FILLER_34_1927 ();
 FILLCELL_X32 FILLER_34_1959 ();
 FILLCELL_X32 FILLER_34_1991 ();
 FILLCELL_X32 FILLER_34_2023 ();
 FILLCELL_X32 FILLER_34_2055 ();
 FILLCELL_X32 FILLER_34_2087 ();
 FILLCELL_X32 FILLER_34_2119 ();
 FILLCELL_X32 FILLER_34_2151 ();
 FILLCELL_X32 FILLER_34_2183 ();
 FILLCELL_X32 FILLER_34_2215 ();
 FILLCELL_X32 FILLER_34_2247 ();
 FILLCELL_X32 FILLER_34_2279 ();
 FILLCELL_X32 FILLER_34_2311 ();
 FILLCELL_X32 FILLER_34_2343 ();
 FILLCELL_X32 FILLER_34_2375 ();
 FILLCELL_X32 FILLER_34_2407 ();
 FILLCELL_X32 FILLER_34_2439 ();
 FILLCELL_X32 FILLER_34_2471 ();
 FILLCELL_X32 FILLER_34_2503 ();
 FILLCELL_X32 FILLER_34_2535 ();
 FILLCELL_X32 FILLER_34_2567 ();
 FILLCELL_X2 FILLER_34_2599 ();
 FILLCELL_X1 FILLER_34_2601 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X32 FILLER_35_161 ();
 FILLCELL_X32 FILLER_35_193 ();
 FILLCELL_X32 FILLER_35_225 ();
 FILLCELL_X32 FILLER_35_257 ();
 FILLCELL_X32 FILLER_35_289 ();
 FILLCELL_X32 FILLER_35_321 ();
 FILLCELL_X32 FILLER_35_353 ();
 FILLCELL_X32 FILLER_35_385 ();
 FILLCELL_X32 FILLER_35_417 ();
 FILLCELL_X32 FILLER_35_449 ();
 FILLCELL_X32 FILLER_35_481 ();
 FILLCELL_X32 FILLER_35_513 ();
 FILLCELL_X32 FILLER_35_545 ();
 FILLCELL_X32 FILLER_35_577 ();
 FILLCELL_X32 FILLER_35_609 ();
 FILLCELL_X32 FILLER_35_641 ();
 FILLCELL_X32 FILLER_35_673 ();
 FILLCELL_X32 FILLER_35_705 ();
 FILLCELL_X32 FILLER_35_737 ();
 FILLCELL_X32 FILLER_35_769 ();
 FILLCELL_X32 FILLER_35_801 ();
 FILLCELL_X32 FILLER_35_833 ();
 FILLCELL_X32 FILLER_35_865 ();
 FILLCELL_X32 FILLER_35_897 ();
 FILLCELL_X32 FILLER_35_929 ();
 FILLCELL_X32 FILLER_35_961 ();
 FILLCELL_X32 FILLER_35_993 ();
 FILLCELL_X32 FILLER_35_1025 ();
 FILLCELL_X32 FILLER_35_1057 ();
 FILLCELL_X32 FILLER_35_1089 ();
 FILLCELL_X32 FILLER_35_1121 ();
 FILLCELL_X32 FILLER_35_1153 ();
 FILLCELL_X32 FILLER_35_1185 ();
 FILLCELL_X32 FILLER_35_1217 ();
 FILLCELL_X8 FILLER_35_1249 ();
 FILLCELL_X4 FILLER_35_1257 ();
 FILLCELL_X2 FILLER_35_1261 ();
 FILLCELL_X32 FILLER_35_1264 ();
 FILLCELL_X32 FILLER_35_1296 ();
 FILLCELL_X32 FILLER_35_1328 ();
 FILLCELL_X32 FILLER_35_1360 ();
 FILLCELL_X32 FILLER_35_1392 ();
 FILLCELL_X32 FILLER_35_1424 ();
 FILLCELL_X32 FILLER_35_1456 ();
 FILLCELL_X32 FILLER_35_1488 ();
 FILLCELL_X32 FILLER_35_1520 ();
 FILLCELL_X32 FILLER_35_1552 ();
 FILLCELL_X32 FILLER_35_1584 ();
 FILLCELL_X32 FILLER_35_1616 ();
 FILLCELL_X32 FILLER_35_1648 ();
 FILLCELL_X32 FILLER_35_1680 ();
 FILLCELL_X32 FILLER_35_1712 ();
 FILLCELL_X32 FILLER_35_1744 ();
 FILLCELL_X32 FILLER_35_1776 ();
 FILLCELL_X32 FILLER_35_1808 ();
 FILLCELL_X32 FILLER_35_1840 ();
 FILLCELL_X32 FILLER_35_1872 ();
 FILLCELL_X32 FILLER_35_1904 ();
 FILLCELL_X32 FILLER_35_1936 ();
 FILLCELL_X32 FILLER_35_1968 ();
 FILLCELL_X32 FILLER_35_2000 ();
 FILLCELL_X32 FILLER_35_2032 ();
 FILLCELL_X32 FILLER_35_2064 ();
 FILLCELL_X32 FILLER_35_2096 ();
 FILLCELL_X32 FILLER_35_2128 ();
 FILLCELL_X32 FILLER_35_2160 ();
 FILLCELL_X32 FILLER_35_2192 ();
 FILLCELL_X32 FILLER_35_2224 ();
 FILLCELL_X32 FILLER_35_2256 ();
 FILLCELL_X32 FILLER_35_2288 ();
 FILLCELL_X32 FILLER_35_2320 ();
 FILLCELL_X32 FILLER_35_2352 ();
 FILLCELL_X32 FILLER_35_2384 ();
 FILLCELL_X32 FILLER_35_2416 ();
 FILLCELL_X32 FILLER_35_2448 ();
 FILLCELL_X32 FILLER_35_2480 ();
 FILLCELL_X8 FILLER_35_2512 ();
 FILLCELL_X4 FILLER_35_2520 ();
 FILLCELL_X2 FILLER_35_2524 ();
 FILLCELL_X32 FILLER_35_2527 ();
 FILLCELL_X32 FILLER_35_2559 ();
 FILLCELL_X8 FILLER_35_2591 ();
 FILLCELL_X2 FILLER_35_2599 ();
 FILLCELL_X1 FILLER_35_2601 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X32 FILLER_36_193 ();
 FILLCELL_X32 FILLER_36_225 ();
 FILLCELL_X32 FILLER_36_257 ();
 FILLCELL_X32 FILLER_36_289 ();
 FILLCELL_X32 FILLER_36_321 ();
 FILLCELL_X32 FILLER_36_353 ();
 FILLCELL_X32 FILLER_36_385 ();
 FILLCELL_X32 FILLER_36_417 ();
 FILLCELL_X32 FILLER_36_449 ();
 FILLCELL_X32 FILLER_36_481 ();
 FILLCELL_X32 FILLER_36_513 ();
 FILLCELL_X32 FILLER_36_545 ();
 FILLCELL_X32 FILLER_36_577 ();
 FILLCELL_X16 FILLER_36_609 ();
 FILLCELL_X4 FILLER_36_625 ();
 FILLCELL_X2 FILLER_36_629 ();
 FILLCELL_X32 FILLER_36_632 ();
 FILLCELL_X32 FILLER_36_664 ();
 FILLCELL_X32 FILLER_36_696 ();
 FILLCELL_X32 FILLER_36_728 ();
 FILLCELL_X32 FILLER_36_760 ();
 FILLCELL_X32 FILLER_36_792 ();
 FILLCELL_X32 FILLER_36_824 ();
 FILLCELL_X32 FILLER_36_856 ();
 FILLCELL_X32 FILLER_36_888 ();
 FILLCELL_X32 FILLER_36_920 ();
 FILLCELL_X32 FILLER_36_952 ();
 FILLCELL_X32 FILLER_36_984 ();
 FILLCELL_X32 FILLER_36_1016 ();
 FILLCELL_X32 FILLER_36_1048 ();
 FILLCELL_X32 FILLER_36_1080 ();
 FILLCELL_X32 FILLER_36_1112 ();
 FILLCELL_X32 FILLER_36_1144 ();
 FILLCELL_X32 FILLER_36_1176 ();
 FILLCELL_X32 FILLER_36_1208 ();
 FILLCELL_X32 FILLER_36_1240 ();
 FILLCELL_X32 FILLER_36_1272 ();
 FILLCELL_X32 FILLER_36_1304 ();
 FILLCELL_X32 FILLER_36_1336 ();
 FILLCELL_X32 FILLER_36_1368 ();
 FILLCELL_X32 FILLER_36_1400 ();
 FILLCELL_X32 FILLER_36_1432 ();
 FILLCELL_X32 FILLER_36_1464 ();
 FILLCELL_X32 FILLER_36_1496 ();
 FILLCELL_X32 FILLER_36_1528 ();
 FILLCELL_X32 FILLER_36_1560 ();
 FILLCELL_X32 FILLER_36_1592 ();
 FILLCELL_X32 FILLER_36_1624 ();
 FILLCELL_X32 FILLER_36_1656 ();
 FILLCELL_X32 FILLER_36_1688 ();
 FILLCELL_X32 FILLER_36_1720 ();
 FILLCELL_X32 FILLER_36_1752 ();
 FILLCELL_X32 FILLER_36_1784 ();
 FILLCELL_X32 FILLER_36_1816 ();
 FILLCELL_X32 FILLER_36_1848 ();
 FILLCELL_X8 FILLER_36_1880 ();
 FILLCELL_X4 FILLER_36_1888 ();
 FILLCELL_X2 FILLER_36_1892 ();
 FILLCELL_X32 FILLER_36_1895 ();
 FILLCELL_X32 FILLER_36_1927 ();
 FILLCELL_X32 FILLER_36_1959 ();
 FILLCELL_X32 FILLER_36_1991 ();
 FILLCELL_X32 FILLER_36_2023 ();
 FILLCELL_X32 FILLER_36_2055 ();
 FILLCELL_X32 FILLER_36_2087 ();
 FILLCELL_X32 FILLER_36_2119 ();
 FILLCELL_X32 FILLER_36_2151 ();
 FILLCELL_X32 FILLER_36_2183 ();
 FILLCELL_X32 FILLER_36_2215 ();
 FILLCELL_X32 FILLER_36_2247 ();
 FILLCELL_X32 FILLER_36_2279 ();
 FILLCELL_X32 FILLER_36_2311 ();
 FILLCELL_X32 FILLER_36_2343 ();
 FILLCELL_X32 FILLER_36_2375 ();
 FILLCELL_X32 FILLER_36_2407 ();
 FILLCELL_X32 FILLER_36_2439 ();
 FILLCELL_X32 FILLER_36_2471 ();
 FILLCELL_X32 FILLER_36_2503 ();
 FILLCELL_X32 FILLER_36_2535 ();
 FILLCELL_X32 FILLER_36_2567 ();
 FILLCELL_X2 FILLER_36_2599 ();
 FILLCELL_X1 FILLER_36_2601 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X32 FILLER_37_193 ();
 FILLCELL_X32 FILLER_37_225 ();
 FILLCELL_X32 FILLER_37_257 ();
 FILLCELL_X32 FILLER_37_289 ();
 FILLCELL_X32 FILLER_37_321 ();
 FILLCELL_X32 FILLER_37_353 ();
 FILLCELL_X32 FILLER_37_385 ();
 FILLCELL_X32 FILLER_37_417 ();
 FILLCELL_X32 FILLER_37_449 ();
 FILLCELL_X32 FILLER_37_481 ();
 FILLCELL_X32 FILLER_37_513 ();
 FILLCELL_X32 FILLER_37_545 ();
 FILLCELL_X32 FILLER_37_577 ();
 FILLCELL_X32 FILLER_37_609 ();
 FILLCELL_X32 FILLER_37_641 ();
 FILLCELL_X32 FILLER_37_673 ();
 FILLCELL_X32 FILLER_37_705 ();
 FILLCELL_X32 FILLER_37_737 ();
 FILLCELL_X32 FILLER_37_769 ();
 FILLCELL_X32 FILLER_37_801 ();
 FILLCELL_X32 FILLER_37_833 ();
 FILLCELL_X32 FILLER_37_865 ();
 FILLCELL_X32 FILLER_37_897 ();
 FILLCELL_X32 FILLER_37_929 ();
 FILLCELL_X32 FILLER_37_961 ();
 FILLCELL_X32 FILLER_37_993 ();
 FILLCELL_X32 FILLER_37_1025 ();
 FILLCELL_X32 FILLER_37_1057 ();
 FILLCELL_X32 FILLER_37_1089 ();
 FILLCELL_X32 FILLER_37_1121 ();
 FILLCELL_X32 FILLER_37_1153 ();
 FILLCELL_X32 FILLER_37_1185 ();
 FILLCELL_X32 FILLER_37_1217 ();
 FILLCELL_X8 FILLER_37_1249 ();
 FILLCELL_X4 FILLER_37_1257 ();
 FILLCELL_X2 FILLER_37_1261 ();
 FILLCELL_X32 FILLER_37_1264 ();
 FILLCELL_X32 FILLER_37_1296 ();
 FILLCELL_X32 FILLER_37_1328 ();
 FILLCELL_X32 FILLER_37_1360 ();
 FILLCELL_X32 FILLER_37_1392 ();
 FILLCELL_X32 FILLER_37_1424 ();
 FILLCELL_X32 FILLER_37_1456 ();
 FILLCELL_X32 FILLER_37_1488 ();
 FILLCELL_X32 FILLER_37_1520 ();
 FILLCELL_X32 FILLER_37_1552 ();
 FILLCELL_X32 FILLER_37_1584 ();
 FILLCELL_X32 FILLER_37_1616 ();
 FILLCELL_X32 FILLER_37_1648 ();
 FILLCELL_X32 FILLER_37_1680 ();
 FILLCELL_X32 FILLER_37_1712 ();
 FILLCELL_X32 FILLER_37_1744 ();
 FILLCELL_X32 FILLER_37_1776 ();
 FILLCELL_X32 FILLER_37_1808 ();
 FILLCELL_X32 FILLER_37_1840 ();
 FILLCELL_X32 FILLER_37_1872 ();
 FILLCELL_X32 FILLER_37_1904 ();
 FILLCELL_X32 FILLER_37_1936 ();
 FILLCELL_X32 FILLER_37_1968 ();
 FILLCELL_X32 FILLER_37_2000 ();
 FILLCELL_X32 FILLER_37_2032 ();
 FILLCELL_X32 FILLER_37_2064 ();
 FILLCELL_X32 FILLER_37_2096 ();
 FILLCELL_X32 FILLER_37_2128 ();
 FILLCELL_X32 FILLER_37_2160 ();
 FILLCELL_X32 FILLER_37_2192 ();
 FILLCELL_X32 FILLER_37_2224 ();
 FILLCELL_X32 FILLER_37_2256 ();
 FILLCELL_X32 FILLER_37_2288 ();
 FILLCELL_X32 FILLER_37_2320 ();
 FILLCELL_X32 FILLER_37_2352 ();
 FILLCELL_X32 FILLER_37_2384 ();
 FILLCELL_X32 FILLER_37_2416 ();
 FILLCELL_X32 FILLER_37_2448 ();
 FILLCELL_X32 FILLER_37_2480 ();
 FILLCELL_X8 FILLER_37_2512 ();
 FILLCELL_X4 FILLER_37_2520 ();
 FILLCELL_X2 FILLER_37_2524 ();
 FILLCELL_X32 FILLER_37_2527 ();
 FILLCELL_X32 FILLER_37_2559 ();
 FILLCELL_X8 FILLER_37_2591 ();
 FILLCELL_X2 FILLER_37_2599 ();
 FILLCELL_X1 FILLER_37_2601 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X32 FILLER_38_193 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X32 FILLER_38_257 ();
 FILLCELL_X32 FILLER_38_289 ();
 FILLCELL_X32 FILLER_38_321 ();
 FILLCELL_X32 FILLER_38_353 ();
 FILLCELL_X32 FILLER_38_385 ();
 FILLCELL_X32 FILLER_38_417 ();
 FILLCELL_X32 FILLER_38_449 ();
 FILLCELL_X32 FILLER_38_481 ();
 FILLCELL_X32 FILLER_38_513 ();
 FILLCELL_X32 FILLER_38_545 ();
 FILLCELL_X32 FILLER_38_577 ();
 FILLCELL_X16 FILLER_38_609 ();
 FILLCELL_X4 FILLER_38_625 ();
 FILLCELL_X2 FILLER_38_629 ();
 FILLCELL_X32 FILLER_38_632 ();
 FILLCELL_X32 FILLER_38_664 ();
 FILLCELL_X32 FILLER_38_696 ();
 FILLCELL_X32 FILLER_38_728 ();
 FILLCELL_X32 FILLER_38_760 ();
 FILLCELL_X32 FILLER_38_792 ();
 FILLCELL_X32 FILLER_38_824 ();
 FILLCELL_X32 FILLER_38_856 ();
 FILLCELL_X32 FILLER_38_888 ();
 FILLCELL_X32 FILLER_38_920 ();
 FILLCELL_X32 FILLER_38_952 ();
 FILLCELL_X32 FILLER_38_984 ();
 FILLCELL_X32 FILLER_38_1016 ();
 FILLCELL_X32 FILLER_38_1048 ();
 FILLCELL_X32 FILLER_38_1080 ();
 FILLCELL_X32 FILLER_38_1112 ();
 FILLCELL_X32 FILLER_38_1144 ();
 FILLCELL_X32 FILLER_38_1176 ();
 FILLCELL_X32 FILLER_38_1208 ();
 FILLCELL_X32 FILLER_38_1240 ();
 FILLCELL_X32 FILLER_38_1272 ();
 FILLCELL_X32 FILLER_38_1304 ();
 FILLCELL_X32 FILLER_38_1336 ();
 FILLCELL_X32 FILLER_38_1368 ();
 FILLCELL_X32 FILLER_38_1400 ();
 FILLCELL_X32 FILLER_38_1432 ();
 FILLCELL_X32 FILLER_38_1464 ();
 FILLCELL_X32 FILLER_38_1496 ();
 FILLCELL_X32 FILLER_38_1528 ();
 FILLCELL_X32 FILLER_38_1560 ();
 FILLCELL_X32 FILLER_38_1592 ();
 FILLCELL_X32 FILLER_38_1624 ();
 FILLCELL_X32 FILLER_38_1656 ();
 FILLCELL_X32 FILLER_38_1688 ();
 FILLCELL_X32 FILLER_38_1720 ();
 FILLCELL_X32 FILLER_38_1752 ();
 FILLCELL_X32 FILLER_38_1784 ();
 FILLCELL_X32 FILLER_38_1816 ();
 FILLCELL_X32 FILLER_38_1848 ();
 FILLCELL_X8 FILLER_38_1880 ();
 FILLCELL_X4 FILLER_38_1888 ();
 FILLCELL_X2 FILLER_38_1892 ();
 FILLCELL_X32 FILLER_38_1895 ();
 FILLCELL_X32 FILLER_38_1927 ();
 FILLCELL_X32 FILLER_38_1959 ();
 FILLCELL_X32 FILLER_38_1991 ();
 FILLCELL_X32 FILLER_38_2023 ();
 FILLCELL_X32 FILLER_38_2055 ();
 FILLCELL_X32 FILLER_38_2087 ();
 FILLCELL_X32 FILLER_38_2119 ();
 FILLCELL_X32 FILLER_38_2151 ();
 FILLCELL_X32 FILLER_38_2183 ();
 FILLCELL_X32 FILLER_38_2215 ();
 FILLCELL_X32 FILLER_38_2247 ();
 FILLCELL_X32 FILLER_38_2279 ();
 FILLCELL_X32 FILLER_38_2311 ();
 FILLCELL_X32 FILLER_38_2343 ();
 FILLCELL_X32 FILLER_38_2375 ();
 FILLCELL_X32 FILLER_38_2407 ();
 FILLCELL_X32 FILLER_38_2439 ();
 FILLCELL_X32 FILLER_38_2471 ();
 FILLCELL_X32 FILLER_38_2503 ();
 FILLCELL_X32 FILLER_38_2535 ();
 FILLCELL_X32 FILLER_38_2567 ();
 FILLCELL_X2 FILLER_38_2599 ();
 FILLCELL_X1 FILLER_38_2601 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X32 FILLER_39_193 ();
 FILLCELL_X32 FILLER_39_225 ();
 FILLCELL_X32 FILLER_39_257 ();
 FILLCELL_X32 FILLER_39_289 ();
 FILLCELL_X32 FILLER_39_321 ();
 FILLCELL_X32 FILLER_39_353 ();
 FILLCELL_X32 FILLER_39_385 ();
 FILLCELL_X32 FILLER_39_417 ();
 FILLCELL_X32 FILLER_39_449 ();
 FILLCELL_X32 FILLER_39_481 ();
 FILLCELL_X32 FILLER_39_513 ();
 FILLCELL_X32 FILLER_39_545 ();
 FILLCELL_X32 FILLER_39_577 ();
 FILLCELL_X32 FILLER_39_609 ();
 FILLCELL_X32 FILLER_39_641 ();
 FILLCELL_X32 FILLER_39_673 ();
 FILLCELL_X32 FILLER_39_705 ();
 FILLCELL_X32 FILLER_39_737 ();
 FILLCELL_X32 FILLER_39_769 ();
 FILLCELL_X32 FILLER_39_801 ();
 FILLCELL_X32 FILLER_39_833 ();
 FILLCELL_X32 FILLER_39_865 ();
 FILLCELL_X32 FILLER_39_897 ();
 FILLCELL_X32 FILLER_39_929 ();
 FILLCELL_X32 FILLER_39_961 ();
 FILLCELL_X32 FILLER_39_993 ();
 FILLCELL_X32 FILLER_39_1025 ();
 FILLCELL_X32 FILLER_39_1057 ();
 FILLCELL_X32 FILLER_39_1089 ();
 FILLCELL_X32 FILLER_39_1121 ();
 FILLCELL_X32 FILLER_39_1153 ();
 FILLCELL_X32 FILLER_39_1185 ();
 FILLCELL_X32 FILLER_39_1217 ();
 FILLCELL_X8 FILLER_39_1249 ();
 FILLCELL_X4 FILLER_39_1257 ();
 FILLCELL_X2 FILLER_39_1261 ();
 FILLCELL_X32 FILLER_39_1264 ();
 FILLCELL_X32 FILLER_39_1296 ();
 FILLCELL_X32 FILLER_39_1328 ();
 FILLCELL_X32 FILLER_39_1360 ();
 FILLCELL_X32 FILLER_39_1392 ();
 FILLCELL_X32 FILLER_39_1424 ();
 FILLCELL_X32 FILLER_39_1456 ();
 FILLCELL_X32 FILLER_39_1488 ();
 FILLCELL_X32 FILLER_39_1520 ();
 FILLCELL_X32 FILLER_39_1552 ();
 FILLCELL_X32 FILLER_39_1584 ();
 FILLCELL_X32 FILLER_39_1616 ();
 FILLCELL_X32 FILLER_39_1648 ();
 FILLCELL_X32 FILLER_39_1680 ();
 FILLCELL_X32 FILLER_39_1712 ();
 FILLCELL_X32 FILLER_39_1744 ();
 FILLCELL_X32 FILLER_39_1776 ();
 FILLCELL_X32 FILLER_39_1808 ();
 FILLCELL_X32 FILLER_39_1840 ();
 FILLCELL_X32 FILLER_39_1872 ();
 FILLCELL_X32 FILLER_39_1904 ();
 FILLCELL_X32 FILLER_39_1936 ();
 FILLCELL_X32 FILLER_39_1968 ();
 FILLCELL_X32 FILLER_39_2000 ();
 FILLCELL_X32 FILLER_39_2032 ();
 FILLCELL_X32 FILLER_39_2064 ();
 FILLCELL_X32 FILLER_39_2096 ();
 FILLCELL_X32 FILLER_39_2128 ();
 FILLCELL_X32 FILLER_39_2160 ();
 FILLCELL_X32 FILLER_39_2192 ();
 FILLCELL_X32 FILLER_39_2224 ();
 FILLCELL_X32 FILLER_39_2256 ();
 FILLCELL_X32 FILLER_39_2288 ();
 FILLCELL_X32 FILLER_39_2320 ();
 FILLCELL_X32 FILLER_39_2352 ();
 FILLCELL_X32 FILLER_39_2384 ();
 FILLCELL_X32 FILLER_39_2416 ();
 FILLCELL_X32 FILLER_39_2448 ();
 FILLCELL_X32 FILLER_39_2480 ();
 FILLCELL_X8 FILLER_39_2512 ();
 FILLCELL_X4 FILLER_39_2520 ();
 FILLCELL_X2 FILLER_39_2524 ();
 FILLCELL_X32 FILLER_39_2527 ();
 FILLCELL_X32 FILLER_39_2559 ();
 FILLCELL_X8 FILLER_39_2591 ();
 FILLCELL_X2 FILLER_39_2599 ();
 FILLCELL_X1 FILLER_39_2601 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X32 FILLER_40_193 ();
 FILLCELL_X32 FILLER_40_225 ();
 FILLCELL_X32 FILLER_40_257 ();
 FILLCELL_X32 FILLER_40_289 ();
 FILLCELL_X32 FILLER_40_321 ();
 FILLCELL_X32 FILLER_40_353 ();
 FILLCELL_X32 FILLER_40_385 ();
 FILLCELL_X32 FILLER_40_417 ();
 FILLCELL_X32 FILLER_40_449 ();
 FILLCELL_X32 FILLER_40_481 ();
 FILLCELL_X32 FILLER_40_513 ();
 FILLCELL_X32 FILLER_40_545 ();
 FILLCELL_X32 FILLER_40_577 ();
 FILLCELL_X16 FILLER_40_609 ();
 FILLCELL_X4 FILLER_40_625 ();
 FILLCELL_X2 FILLER_40_629 ();
 FILLCELL_X32 FILLER_40_632 ();
 FILLCELL_X32 FILLER_40_664 ();
 FILLCELL_X32 FILLER_40_696 ();
 FILLCELL_X32 FILLER_40_728 ();
 FILLCELL_X32 FILLER_40_760 ();
 FILLCELL_X32 FILLER_40_792 ();
 FILLCELL_X32 FILLER_40_824 ();
 FILLCELL_X32 FILLER_40_856 ();
 FILLCELL_X32 FILLER_40_888 ();
 FILLCELL_X32 FILLER_40_920 ();
 FILLCELL_X32 FILLER_40_952 ();
 FILLCELL_X32 FILLER_40_984 ();
 FILLCELL_X32 FILLER_40_1016 ();
 FILLCELL_X32 FILLER_40_1048 ();
 FILLCELL_X32 FILLER_40_1080 ();
 FILLCELL_X32 FILLER_40_1112 ();
 FILLCELL_X32 FILLER_40_1144 ();
 FILLCELL_X32 FILLER_40_1176 ();
 FILLCELL_X32 FILLER_40_1208 ();
 FILLCELL_X32 FILLER_40_1240 ();
 FILLCELL_X32 FILLER_40_1272 ();
 FILLCELL_X32 FILLER_40_1304 ();
 FILLCELL_X32 FILLER_40_1336 ();
 FILLCELL_X32 FILLER_40_1368 ();
 FILLCELL_X32 FILLER_40_1400 ();
 FILLCELL_X32 FILLER_40_1432 ();
 FILLCELL_X32 FILLER_40_1464 ();
 FILLCELL_X32 FILLER_40_1496 ();
 FILLCELL_X32 FILLER_40_1528 ();
 FILLCELL_X32 FILLER_40_1560 ();
 FILLCELL_X32 FILLER_40_1592 ();
 FILLCELL_X32 FILLER_40_1624 ();
 FILLCELL_X32 FILLER_40_1656 ();
 FILLCELL_X32 FILLER_40_1688 ();
 FILLCELL_X32 FILLER_40_1720 ();
 FILLCELL_X32 FILLER_40_1752 ();
 FILLCELL_X32 FILLER_40_1784 ();
 FILLCELL_X32 FILLER_40_1816 ();
 FILLCELL_X32 FILLER_40_1848 ();
 FILLCELL_X8 FILLER_40_1880 ();
 FILLCELL_X4 FILLER_40_1888 ();
 FILLCELL_X2 FILLER_40_1892 ();
 FILLCELL_X32 FILLER_40_1895 ();
 FILLCELL_X32 FILLER_40_1927 ();
 FILLCELL_X32 FILLER_40_1959 ();
 FILLCELL_X32 FILLER_40_1991 ();
 FILLCELL_X32 FILLER_40_2023 ();
 FILLCELL_X32 FILLER_40_2055 ();
 FILLCELL_X32 FILLER_40_2087 ();
 FILLCELL_X32 FILLER_40_2119 ();
 FILLCELL_X32 FILLER_40_2151 ();
 FILLCELL_X32 FILLER_40_2183 ();
 FILLCELL_X32 FILLER_40_2215 ();
 FILLCELL_X32 FILLER_40_2247 ();
 FILLCELL_X32 FILLER_40_2279 ();
 FILLCELL_X32 FILLER_40_2311 ();
 FILLCELL_X32 FILLER_40_2343 ();
 FILLCELL_X32 FILLER_40_2375 ();
 FILLCELL_X32 FILLER_40_2407 ();
 FILLCELL_X32 FILLER_40_2439 ();
 FILLCELL_X32 FILLER_40_2471 ();
 FILLCELL_X32 FILLER_40_2503 ();
 FILLCELL_X32 FILLER_40_2535 ();
 FILLCELL_X32 FILLER_40_2567 ();
 FILLCELL_X2 FILLER_40_2599 ();
 FILLCELL_X1 FILLER_40_2601 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X32 FILLER_41_129 ();
 FILLCELL_X32 FILLER_41_161 ();
 FILLCELL_X32 FILLER_41_193 ();
 FILLCELL_X32 FILLER_41_225 ();
 FILLCELL_X32 FILLER_41_257 ();
 FILLCELL_X32 FILLER_41_289 ();
 FILLCELL_X32 FILLER_41_321 ();
 FILLCELL_X32 FILLER_41_353 ();
 FILLCELL_X32 FILLER_41_385 ();
 FILLCELL_X32 FILLER_41_417 ();
 FILLCELL_X32 FILLER_41_449 ();
 FILLCELL_X32 FILLER_41_481 ();
 FILLCELL_X32 FILLER_41_513 ();
 FILLCELL_X32 FILLER_41_545 ();
 FILLCELL_X32 FILLER_41_577 ();
 FILLCELL_X32 FILLER_41_609 ();
 FILLCELL_X32 FILLER_41_641 ();
 FILLCELL_X32 FILLER_41_673 ();
 FILLCELL_X32 FILLER_41_705 ();
 FILLCELL_X32 FILLER_41_737 ();
 FILLCELL_X32 FILLER_41_769 ();
 FILLCELL_X32 FILLER_41_801 ();
 FILLCELL_X32 FILLER_41_833 ();
 FILLCELL_X32 FILLER_41_865 ();
 FILLCELL_X32 FILLER_41_897 ();
 FILLCELL_X32 FILLER_41_929 ();
 FILLCELL_X32 FILLER_41_961 ();
 FILLCELL_X32 FILLER_41_993 ();
 FILLCELL_X32 FILLER_41_1025 ();
 FILLCELL_X32 FILLER_41_1057 ();
 FILLCELL_X32 FILLER_41_1089 ();
 FILLCELL_X32 FILLER_41_1121 ();
 FILLCELL_X32 FILLER_41_1153 ();
 FILLCELL_X32 FILLER_41_1185 ();
 FILLCELL_X32 FILLER_41_1217 ();
 FILLCELL_X8 FILLER_41_1249 ();
 FILLCELL_X4 FILLER_41_1257 ();
 FILLCELL_X2 FILLER_41_1261 ();
 FILLCELL_X32 FILLER_41_1264 ();
 FILLCELL_X32 FILLER_41_1296 ();
 FILLCELL_X32 FILLER_41_1328 ();
 FILLCELL_X32 FILLER_41_1360 ();
 FILLCELL_X32 FILLER_41_1392 ();
 FILLCELL_X32 FILLER_41_1424 ();
 FILLCELL_X32 FILLER_41_1456 ();
 FILLCELL_X32 FILLER_41_1488 ();
 FILLCELL_X32 FILLER_41_1520 ();
 FILLCELL_X32 FILLER_41_1552 ();
 FILLCELL_X32 FILLER_41_1584 ();
 FILLCELL_X32 FILLER_41_1616 ();
 FILLCELL_X32 FILLER_41_1648 ();
 FILLCELL_X32 FILLER_41_1680 ();
 FILLCELL_X32 FILLER_41_1712 ();
 FILLCELL_X32 FILLER_41_1744 ();
 FILLCELL_X32 FILLER_41_1776 ();
 FILLCELL_X32 FILLER_41_1808 ();
 FILLCELL_X32 FILLER_41_1840 ();
 FILLCELL_X32 FILLER_41_1872 ();
 FILLCELL_X32 FILLER_41_1904 ();
 FILLCELL_X32 FILLER_41_1936 ();
 FILLCELL_X32 FILLER_41_1968 ();
 FILLCELL_X32 FILLER_41_2000 ();
 FILLCELL_X32 FILLER_41_2032 ();
 FILLCELL_X32 FILLER_41_2064 ();
 FILLCELL_X32 FILLER_41_2096 ();
 FILLCELL_X32 FILLER_41_2128 ();
 FILLCELL_X32 FILLER_41_2160 ();
 FILLCELL_X32 FILLER_41_2192 ();
 FILLCELL_X32 FILLER_41_2224 ();
 FILLCELL_X32 FILLER_41_2256 ();
 FILLCELL_X32 FILLER_41_2288 ();
 FILLCELL_X32 FILLER_41_2320 ();
 FILLCELL_X32 FILLER_41_2352 ();
 FILLCELL_X32 FILLER_41_2384 ();
 FILLCELL_X32 FILLER_41_2416 ();
 FILLCELL_X32 FILLER_41_2448 ();
 FILLCELL_X32 FILLER_41_2480 ();
 FILLCELL_X8 FILLER_41_2512 ();
 FILLCELL_X4 FILLER_41_2520 ();
 FILLCELL_X2 FILLER_41_2524 ();
 FILLCELL_X32 FILLER_41_2527 ();
 FILLCELL_X32 FILLER_41_2559 ();
 FILLCELL_X8 FILLER_41_2591 ();
 FILLCELL_X2 FILLER_41_2599 ();
 FILLCELL_X1 FILLER_41_2601 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X32 FILLER_42_129 ();
 FILLCELL_X32 FILLER_42_161 ();
 FILLCELL_X32 FILLER_42_193 ();
 FILLCELL_X32 FILLER_42_225 ();
 FILLCELL_X32 FILLER_42_257 ();
 FILLCELL_X32 FILLER_42_289 ();
 FILLCELL_X32 FILLER_42_321 ();
 FILLCELL_X32 FILLER_42_353 ();
 FILLCELL_X32 FILLER_42_385 ();
 FILLCELL_X32 FILLER_42_417 ();
 FILLCELL_X32 FILLER_42_449 ();
 FILLCELL_X32 FILLER_42_481 ();
 FILLCELL_X32 FILLER_42_513 ();
 FILLCELL_X32 FILLER_42_545 ();
 FILLCELL_X32 FILLER_42_577 ();
 FILLCELL_X16 FILLER_42_609 ();
 FILLCELL_X4 FILLER_42_625 ();
 FILLCELL_X2 FILLER_42_629 ();
 FILLCELL_X32 FILLER_42_632 ();
 FILLCELL_X32 FILLER_42_664 ();
 FILLCELL_X32 FILLER_42_696 ();
 FILLCELL_X32 FILLER_42_728 ();
 FILLCELL_X32 FILLER_42_760 ();
 FILLCELL_X32 FILLER_42_792 ();
 FILLCELL_X32 FILLER_42_824 ();
 FILLCELL_X32 FILLER_42_856 ();
 FILLCELL_X32 FILLER_42_888 ();
 FILLCELL_X32 FILLER_42_920 ();
 FILLCELL_X32 FILLER_42_952 ();
 FILLCELL_X32 FILLER_42_984 ();
 FILLCELL_X32 FILLER_42_1016 ();
 FILLCELL_X32 FILLER_42_1048 ();
 FILLCELL_X32 FILLER_42_1080 ();
 FILLCELL_X32 FILLER_42_1112 ();
 FILLCELL_X32 FILLER_42_1144 ();
 FILLCELL_X32 FILLER_42_1176 ();
 FILLCELL_X32 FILLER_42_1208 ();
 FILLCELL_X32 FILLER_42_1240 ();
 FILLCELL_X32 FILLER_42_1272 ();
 FILLCELL_X32 FILLER_42_1304 ();
 FILLCELL_X32 FILLER_42_1336 ();
 FILLCELL_X32 FILLER_42_1368 ();
 FILLCELL_X32 FILLER_42_1400 ();
 FILLCELL_X32 FILLER_42_1432 ();
 FILLCELL_X32 FILLER_42_1464 ();
 FILLCELL_X32 FILLER_42_1496 ();
 FILLCELL_X32 FILLER_42_1528 ();
 FILLCELL_X32 FILLER_42_1560 ();
 FILLCELL_X32 FILLER_42_1592 ();
 FILLCELL_X32 FILLER_42_1624 ();
 FILLCELL_X32 FILLER_42_1656 ();
 FILLCELL_X32 FILLER_42_1688 ();
 FILLCELL_X32 FILLER_42_1720 ();
 FILLCELL_X32 FILLER_42_1752 ();
 FILLCELL_X32 FILLER_42_1784 ();
 FILLCELL_X32 FILLER_42_1816 ();
 FILLCELL_X32 FILLER_42_1848 ();
 FILLCELL_X8 FILLER_42_1880 ();
 FILLCELL_X4 FILLER_42_1888 ();
 FILLCELL_X2 FILLER_42_1892 ();
 FILLCELL_X32 FILLER_42_1895 ();
 FILLCELL_X32 FILLER_42_1927 ();
 FILLCELL_X32 FILLER_42_1959 ();
 FILLCELL_X32 FILLER_42_1991 ();
 FILLCELL_X32 FILLER_42_2023 ();
 FILLCELL_X32 FILLER_42_2055 ();
 FILLCELL_X32 FILLER_42_2087 ();
 FILLCELL_X32 FILLER_42_2119 ();
 FILLCELL_X32 FILLER_42_2151 ();
 FILLCELL_X32 FILLER_42_2183 ();
 FILLCELL_X32 FILLER_42_2215 ();
 FILLCELL_X32 FILLER_42_2247 ();
 FILLCELL_X32 FILLER_42_2279 ();
 FILLCELL_X32 FILLER_42_2311 ();
 FILLCELL_X32 FILLER_42_2343 ();
 FILLCELL_X32 FILLER_42_2375 ();
 FILLCELL_X32 FILLER_42_2407 ();
 FILLCELL_X32 FILLER_42_2439 ();
 FILLCELL_X32 FILLER_42_2471 ();
 FILLCELL_X32 FILLER_42_2503 ();
 FILLCELL_X32 FILLER_42_2535 ();
 FILLCELL_X32 FILLER_42_2567 ();
 FILLCELL_X2 FILLER_42_2599 ();
 FILLCELL_X1 FILLER_42_2601 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X32 FILLER_43_97 ();
 FILLCELL_X32 FILLER_43_129 ();
 FILLCELL_X32 FILLER_43_161 ();
 FILLCELL_X32 FILLER_43_193 ();
 FILLCELL_X32 FILLER_43_225 ();
 FILLCELL_X32 FILLER_43_257 ();
 FILLCELL_X32 FILLER_43_289 ();
 FILLCELL_X32 FILLER_43_321 ();
 FILLCELL_X32 FILLER_43_353 ();
 FILLCELL_X32 FILLER_43_385 ();
 FILLCELL_X32 FILLER_43_417 ();
 FILLCELL_X32 FILLER_43_449 ();
 FILLCELL_X32 FILLER_43_481 ();
 FILLCELL_X32 FILLER_43_513 ();
 FILLCELL_X32 FILLER_43_545 ();
 FILLCELL_X32 FILLER_43_577 ();
 FILLCELL_X32 FILLER_43_609 ();
 FILLCELL_X32 FILLER_43_641 ();
 FILLCELL_X32 FILLER_43_673 ();
 FILLCELL_X32 FILLER_43_705 ();
 FILLCELL_X32 FILLER_43_737 ();
 FILLCELL_X32 FILLER_43_769 ();
 FILLCELL_X32 FILLER_43_801 ();
 FILLCELL_X32 FILLER_43_833 ();
 FILLCELL_X32 FILLER_43_865 ();
 FILLCELL_X32 FILLER_43_897 ();
 FILLCELL_X32 FILLER_43_929 ();
 FILLCELL_X32 FILLER_43_961 ();
 FILLCELL_X32 FILLER_43_993 ();
 FILLCELL_X32 FILLER_43_1025 ();
 FILLCELL_X32 FILLER_43_1057 ();
 FILLCELL_X32 FILLER_43_1089 ();
 FILLCELL_X32 FILLER_43_1121 ();
 FILLCELL_X32 FILLER_43_1153 ();
 FILLCELL_X32 FILLER_43_1185 ();
 FILLCELL_X32 FILLER_43_1217 ();
 FILLCELL_X8 FILLER_43_1249 ();
 FILLCELL_X4 FILLER_43_1257 ();
 FILLCELL_X2 FILLER_43_1261 ();
 FILLCELL_X32 FILLER_43_1264 ();
 FILLCELL_X32 FILLER_43_1296 ();
 FILLCELL_X32 FILLER_43_1328 ();
 FILLCELL_X32 FILLER_43_1360 ();
 FILLCELL_X32 FILLER_43_1392 ();
 FILLCELL_X32 FILLER_43_1424 ();
 FILLCELL_X32 FILLER_43_1456 ();
 FILLCELL_X32 FILLER_43_1488 ();
 FILLCELL_X32 FILLER_43_1520 ();
 FILLCELL_X32 FILLER_43_1552 ();
 FILLCELL_X32 FILLER_43_1584 ();
 FILLCELL_X32 FILLER_43_1616 ();
 FILLCELL_X32 FILLER_43_1648 ();
 FILLCELL_X32 FILLER_43_1680 ();
 FILLCELL_X32 FILLER_43_1712 ();
 FILLCELL_X32 FILLER_43_1744 ();
 FILLCELL_X32 FILLER_43_1776 ();
 FILLCELL_X32 FILLER_43_1808 ();
 FILLCELL_X32 FILLER_43_1840 ();
 FILLCELL_X32 FILLER_43_1872 ();
 FILLCELL_X32 FILLER_43_1904 ();
 FILLCELL_X32 FILLER_43_1936 ();
 FILLCELL_X32 FILLER_43_1968 ();
 FILLCELL_X32 FILLER_43_2000 ();
 FILLCELL_X32 FILLER_43_2032 ();
 FILLCELL_X32 FILLER_43_2064 ();
 FILLCELL_X32 FILLER_43_2096 ();
 FILLCELL_X32 FILLER_43_2128 ();
 FILLCELL_X32 FILLER_43_2160 ();
 FILLCELL_X32 FILLER_43_2192 ();
 FILLCELL_X32 FILLER_43_2224 ();
 FILLCELL_X32 FILLER_43_2256 ();
 FILLCELL_X32 FILLER_43_2288 ();
 FILLCELL_X32 FILLER_43_2320 ();
 FILLCELL_X32 FILLER_43_2352 ();
 FILLCELL_X32 FILLER_43_2384 ();
 FILLCELL_X32 FILLER_43_2416 ();
 FILLCELL_X32 FILLER_43_2448 ();
 FILLCELL_X32 FILLER_43_2480 ();
 FILLCELL_X8 FILLER_43_2512 ();
 FILLCELL_X4 FILLER_43_2520 ();
 FILLCELL_X2 FILLER_43_2524 ();
 FILLCELL_X32 FILLER_43_2527 ();
 FILLCELL_X32 FILLER_43_2559 ();
 FILLCELL_X8 FILLER_43_2591 ();
 FILLCELL_X2 FILLER_43_2599 ();
 FILLCELL_X1 FILLER_43_2601 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X32 FILLER_44_65 ();
 FILLCELL_X32 FILLER_44_97 ();
 FILLCELL_X32 FILLER_44_129 ();
 FILLCELL_X32 FILLER_44_161 ();
 FILLCELL_X32 FILLER_44_193 ();
 FILLCELL_X32 FILLER_44_225 ();
 FILLCELL_X32 FILLER_44_257 ();
 FILLCELL_X32 FILLER_44_289 ();
 FILLCELL_X32 FILLER_44_321 ();
 FILLCELL_X32 FILLER_44_353 ();
 FILLCELL_X32 FILLER_44_385 ();
 FILLCELL_X32 FILLER_44_417 ();
 FILLCELL_X32 FILLER_44_449 ();
 FILLCELL_X32 FILLER_44_481 ();
 FILLCELL_X32 FILLER_44_513 ();
 FILLCELL_X32 FILLER_44_545 ();
 FILLCELL_X32 FILLER_44_577 ();
 FILLCELL_X16 FILLER_44_609 ();
 FILLCELL_X4 FILLER_44_625 ();
 FILLCELL_X2 FILLER_44_629 ();
 FILLCELL_X32 FILLER_44_632 ();
 FILLCELL_X32 FILLER_44_664 ();
 FILLCELL_X32 FILLER_44_696 ();
 FILLCELL_X32 FILLER_44_728 ();
 FILLCELL_X32 FILLER_44_760 ();
 FILLCELL_X32 FILLER_44_792 ();
 FILLCELL_X32 FILLER_44_824 ();
 FILLCELL_X32 FILLER_44_856 ();
 FILLCELL_X32 FILLER_44_888 ();
 FILLCELL_X32 FILLER_44_920 ();
 FILLCELL_X32 FILLER_44_952 ();
 FILLCELL_X32 FILLER_44_984 ();
 FILLCELL_X32 FILLER_44_1016 ();
 FILLCELL_X32 FILLER_44_1048 ();
 FILLCELL_X32 FILLER_44_1080 ();
 FILLCELL_X32 FILLER_44_1112 ();
 FILLCELL_X32 FILLER_44_1144 ();
 FILLCELL_X32 FILLER_44_1176 ();
 FILLCELL_X32 FILLER_44_1208 ();
 FILLCELL_X32 FILLER_44_1240 ();
 FILLCELL_X32 FILLER_44_1272 ();
 FILLCELL_X32 FILLER_44_1304 ();
 FILLCELL_X32 FILLER_44_1336 ();
 FILLCELL_X32 FILLER_44_1368 ();
 FILLCELL_X32 FILLER_44_1400 ();
 FILLCELL_X32 FILLER_44_1432 ();
 FILLCELL_X32 FILLER_44_1464 ();
 FILLCELL_X32 FILLER_44_1496 ();
 FILLCELL_X32 FILLER_44_1528 ();
 FILLCELL_X32 FILLER_44_1560 ();
 FILLCELL_X32 FILLER_44_1592 ();
 FILLCELL_X32 FILLER_44_1624 ();
 FILLCELL_X32 FILLER_44_1656 ();
 FILLCELL_X32 FILLER_44_1688 ();
 FILLCELL_X32 FILLER_44_1720 ();
 FILLCELL_X32 FILLER_44_1752 ();
 FILLCELL_X32 FILLER_44_1784 ();
 FILLCELL_X32 FILLER_44_1816 ();
 FILLCELL_X32 FILLER_44_1848 ();
 FILLCELL_X8 FILLER_44_1880 ();
 FILLCELL_X4 FILLER_44_1888 ();
 FILLCELL_X2 FILLER_44_1892 ();
 FILLCELL_X32 FILLER_44_1895 ();
 FILLCELL_X32 FILLER_44_1927 ();
 FILLCELL_X32 FILLER_44_1959 ();
 FILLCELL_X32 FILLER_44_1991 ();
 FILLCELL_X32 FILLER_44_2023 ();
 FILLCELL_X32 FILLER_44_2055 ();
 FILLCELL_X32 FILLER_44_2087 ();
 FILLCELL_X32 FILLER_44_2119 ();
 FILLCELL_X32 FILLER_44_2151 ();
 FILLCELL_X32 FILLER_44_2183 ();
 FILLCELL_X32 FILLER_44_2215 ();
 FILLCELL_X32 FILLER_44_2247 ();
 FILLCELL_X32 FILLER_44_2279 ();
 FILLCELL_X32 FILLER_44_2311 ();
 FILLCELL_X32 FILLER_44_2343 ();
 FILLCELL_X32 FILLER_44_2375 ();
 FILLCELL_X32 FILLER_44_2407 ();
 FILLCELL_X32 FILLER_44_2439 ();
 FILLCELL_X32 FILLER_44_2471 ();
 FILLCELL_X32 FILLER_44_2503 ();
 FILLCELL_X32 FILLER_44_2535 ();
 FILLCELL_X32 FILLER_44_2567 ();
 FILLCELL_X2 FILLER_44_2599 ();
 FILLCELL_X1 FILLER_44_2601 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X32 FILLER_45_65 ();
 FILLCELL_X32 FILLER_45_97 ();
 FILLCELL_X32 FILLER_45_129 ();
 FILLCELL_X32 FILLER_45_161 ();
 FILLCELL_X32 FILLER_45_193 ();
 FILLCELL_X32 FILLER_45_225 ();
 FILLCELL_X32 FILLER_45_257 ();
 FILLCELL_X32 FILLER_45_289 ();
 FILLCELL_X32 FILLER_45_321 ();
 FILLCELL_X32 FILLER_45_353 ();
 FILLCELL_X32 FILLER_45_385 ();
 FILLCELL_X32 FILLER_45_417 ();
 FILLCELL_X32 FILLER_45_449 ();
 FILLCELL_X32 FILLER_45_481 ();
 FILLCELL_X32 FILLER_45_513 ();
 FILLCELL_X32 FILLER_45_545 ();
 FILLCELL_X32 FILLER_45_577 ();
 FILLCELL_X32 FILLER_45_609 ();
 FILLCELL_X32 FILLER_45_641 ();
 FILLCELL_X32 FILLER_45_673 ();
 FILLCELL_X32 FILLER_45_705 ();
 FILLCELL_X32 FILLER_45_737 ();
 FILLCELL_X32 FILLER_45_769 ();
 FILLCELL_X32 FILLER_45_801 ();
 FILLCELL_X32 FILLER_45_833 ();
 FILLCELL_X32 FILLER_45_865 ();
 FILLCELL_X32 FILLER_45_897 ();
 FILLCELL_X32 FILLER_45_929 ();
 FILLCELL_X32 FILLER_45_961 ();
 FILLCELL_X32 FILLER_45_993 ();
 FILLCELL_X32 FILLER_45_1025 ();
 FILLCELL_X32 FILLER_45_1057 ();
 FILLCELL_X32 FILLER_45_1089 ();
 FILLCELL_X32 FILLER_45_1121 ();
 FILLCELL_X32 FILLER_45_1153 ();
 FILLCELL_X32 FILLER_45_1185 ();
 FILLCELL_X32 FILLER_45_1217 ();
 FILLCELL_X8 FILLER_45_1249 ();
 FILLCELL_X4 FILLER_45_1257 ();
 FILLCELL_X2 FILLER_45_1261 ();
 FILLCELL_X32 FILLER_45_1264 ();
 FILLCELL_X32 FILLER_45_1296 ();
 FILLCELL_X32 FILLER_45_1328 ();
 FILLCELL_X32 FILLER_45_1360 ();
 FILLCELL_X32 FILLER_45_1392 ();
 FILLCELL_X32 FILLER_45_1424 ();
 FILLCELL_X32 FILLER_45_1456 ();
 FILLCELL_X32 FILLER_45_1488 ();
 FILLCELL_X32 FILLER_45_1520 ();
 FILLCELL_X32 FILLER_45_1552 ();
 FILLCELL_X32 FILLER_45_1584 ();
 FILLCELL_X32 FILLER_45_1616 ();
 FILLCELL_X32 FILLER_45_1648 ();
 FILLCELL_X32 FILLER_45_1680 ();
 FILLCELL_X32 FILLER_45_1712 ();
 FILLCELL_X32 FILLER_45_1744 ();
 FILLCELL_X32 FILLER_45_1776 ();
 FILLCELL_X32 FILLER_45_1808 ();
 FILLCELL_X32 FILLER_45_1840 ();
 FILLCELL_X32 FILLER_45_1872 ();
 FILLCELL_X32 FILLER_45_1904 ();
 FILLCELL_X32 FILLER_45_1936 ();
 FILLCELL_X32 FILLER_45_1968 ();
 FILLCELL_X32 FILLER_45_2000 ();
 FILLCELL_X32 FILLER_45_2032 ();
 FILLCELL_X32 FILLER_45_2064 ();
 FILLCELL_X32 FILLER_45_2096 ();
 FILLCELL_X32 FILLER_45_2128 ();
 FILLCELL_X32 FILLER_45_2160 ();
 FILLCELL_X32 FILLER_45_2192 ();
 FILLCELL_X32 FILLER_45_2224 ();
 FILLCELL_X32 FILLER_45_2256 ();
 FILLCELL_X32 FILLER_45_2288 ();
 FILLCELL_X32 FILLER_45_2320 ();
 FILLCELL_X32 FILLER_45_2352 ();
 FILLCELL_X32 FILLER_45_2384 ();
 FILLCELL_X32 FILLER_45_2416 ();
 FILLCELL_X32 FILLER_45_2448 ();
 FILLCELL_X32 FILLER_45_2480 ();
 FILLCELL_X8 FILLER_45_2512 ();
 FILLCELL_X4 FILLER_45_2520 ();
 FILLCELL_X2 FILLER_45_2524 ();
 FILLCELL_X32 FILLER_45_2527 ();
 FILLCELL_X32 FILLER_45_2559 ();
 FILLCELL_X8 FILLER_45_2591 ();
 FILLCELL_X2 FILLER_45_2599 ();
 FILLCELL_X1 FILLER_45_2601 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X32 FILLER_46_33 ();
 FILLCELL_X32 FILLER_46_65 ();
 FILLCELL_X32 FILLER_46_97 ();
 FILLCELL_X32 FILLER_46_129 ();
 FILLCELL_X32 FILLER_46_161 ();
 FILLCELL_X32 FILLER_46_193 ();
 FILLCELL_X32 FILLER_46_225 ();
 FILLCELL_X32 FILLER_46_257 ();
 FILLCELL_X32 FILLER_46_289 ();
 FILLCELL_X32 FILLER_46_321 ();
 FILLCELL_X32 FILLER_46_353 ();
 FILLCELL_X32 FILLER_46_385 ();
 FILLCELL_X32 FILLER_46_417 ();
 FILLCELL_X32 FILLER_46_449 ();
 FILLCELL_X32 FILLER_46_481 ();
 FILLCELL_X32 FILLER_46_513 ();
 FILLCELL_X32 FILLER_46_545 ();
 FILLCELL_X32 FILLER_46_577 ();
 FILLCELL_X16 FILLER_46_609 ();
 FILLCELL_X4 FILLER_46_625 ();
 FILLCELL_X2 FILLER_46_629 ();
 FILLCELL_X32 FILLER_46_632 ();
 FILLCELL_X32 FILLER_46_664 ();
 FILLCELL_X32 FILLER_46_696 ();
 FILLCELL_X32 FILLER_46_728 ();
 FILLCELL_X32 FILLER_46_760 ();
 FILLCELL_X32 FILLER_46_792 ();
 FILLCELL_X32 FILLER_46_824 ();
 FILLCELL_X32 FILLER_46_856 ();
 FILLCELL_X32 FILLER_46_888 ();
 FILLCELL_X32 FILLER_46_920 ();
 FILLCELL_X32 FILLER_46_952 ();
 FILLCELL_X32 FILLER_46_984 ();
 FILLCELL_X32 FILLER_46_1016 ();
 FILLCELL_X32 FILLER_46_1048 ();
 FILLCELL_X32 FILLER_46_1080 ();
 FILLCELL_X32 FILLER_46_1112 ();
 FILLCELL_X32 FILLER_46_1144 ();
 FILLCELL_X32 FILLER_46_1176 ();
 FILLCELL_X32 FILLER_46_1208 ();
 FILLCELL_X32 FILLER_46_1240 ();
 FILLCELL_X32 FILLER_46_1272 ();
 FILLCELL_X32 FILLER_46_1304 ();
 FILLCELL_X32 FILLER_46_1336 ();
 FILLCELL_X32 FILLER_46_1368 ();
 FILLCELL_X32 FILLER_46_1400 ();
 FILLCELL_X32 FILLER_46_1432 ();
 FILLCELL_X32 FILLER_46_1464 ();
 FILLCELL_X32 FILLER_46_1496 ();
 FILLCELL_X32 FILLER_46_1528 ();
 FILLCELL_X32 FILLER_46_1560 ();
 FILLCELL_X32 FILLER_46_1592 ();
 FILLCELL_X32 FILLER_46_1624 ();
 FILLCELL_X32 FILLER_46_1656 ();
 FILLCELL_X32 FILLER_46_1688 ();
 FILLCELL_X32 FILLER_46_1720 ();
 FILLCELL_X32 FILLER_46_1752 ();
 FILLCELL_X32 FILLER_46_1784 ();
 FILLCELL_X32 FILLER_46_1816 ();
 FILLCELL_X32 FILLER_46_1848 ();
 FILLCELL_X8 FILLER_46_1880 ();
 FILLCELL_X4 FILLER_46_1888 ();
 FILLCELL_X2 FILLER_46_1892 ();
 FILLCELL_X32 FILLER_46_1895 ();
 FILLCELL_X32 FILLER_46_1927 ();
 FILLCELL_X32 FILLER_46_1959 ();
 FILLCELL_X32 FILLER_46_1991 ();
 FILLCELL_X32 FILLER_46_2023 ();
 FILLCELL_X32 FILLER_46_2055 ();
 FILLCELL_X32 FILLER_46_2087 ();
 FILLCELL_X32 FILLER_46_2119 ();
 FILLCELL_X32 FILLER_46_2151 ();
 FILLCELL_X32 FILLER_46_2183 ();
 FILLCELL_X32 FILLER_46_2215 ();
 FILLCELL_X32 FILLER_46_2247 ();
 FILLCELL_X32 FILLER_46_2279 ();
 FILLCELL_X32 FILLER_46_2311 ();
 FILLCELL_X32 FILLER_46_2343 ();
 FILLCELL_X32 FILLER_46_2375 ();
 FILLCELL_X32 FILLER_46_2407 ();
 FILLCELL_X32 FILLER_46_2439 ();
 FILLCELL_X32 FILLER_46_2471 ();
 FILLCELL_X32 FILLER_46_2503 ();
 FILLCELL_X32 FILLER_46_2535 ();
 FILLCELL_X32 FILLER_46_2567 ();
 FILLCELL_X2 FILLER_46_2599 ();
 FILLCELL_X1 FILLER_46_2601 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X32 FILLER_47_33 ();
 FILLCELL_X32 FILLER_47_65 ();
 FILLCELL_X32 FILLER_47_97 ();
 FILLCELL_X32 FILLER_47_129 ();
 FILLCELL_X32 FILLER_47_161 ();
 FILLCELL_X32 FILLER_47_193 ();
 FILLCELL_X32 FILLER_47_225 ();
 FILLCELL_X32 FILLER_47_257 ();
 FILLCELL_X32 FILLER_47_289 ();
 FILLCELL_X32 FILLER_47_321 ();
 FILLCELL_X32 FILLER_47_353 ();
 FILLCELL_X32 FILLER_47_385 ();
 FILLCELL_X32 FILLER_47_417 ();
 FILLCELL_X32 FILLER_47_449 ();
 FILLCELL_X32 FILLER_47_481 ();
 FILLCELL_X32 FILLER_47_513 ();
 FILLCELL_X32 FILLER_47_545 ();
 FILLCELL_X32 FILLER_47_577 ();
 FILLCELL_X32 FILLER_47_609 ();
 FILLCELL_X32 FILLER_47_641 ();
 FILLCELL_X32 FILLER_47_673 ();
 FILLCELL_X32 FILLER_47_705 ();
 FILLCELL_X32 FILLER_47_737 ();
 FILLCELL_X32 FILLER_47_769 ();
 FILLCELL_X32 FILLER_47_801 ();
 FILLCELL_X32 FILLER_47_833 ();
 FILLCELL_X32 FILLER_47_865 ();
 FILLCELL_X32 FILLER_47_897 ();
 FILLCELL_X32 FILLER_47_929 ();
 FILLCELL_X32 FILLER_47_961 ();
 FILLCELL_X32 FILLER_47_993 ();
 FILLCELL_X32 FILLER_47_1025 ();
 FILLCELL_X32 FILLER_47_1057 ();
 FILLCELL_X32 FILLER_47_1089 ();
 FILLCELL_X32 FILLER_47_1121 ();
 FILLCELL_X32 FILLER_47_1153 ();
 FILLCELL_X32 FILLER_47_1185 ();
 FILLCELL_X32 FILLER_47_1217 ();
 FILLCELL_X8 FILLER_47_1249 ();
 FILLCELL_X4 FILLER_47_1257 ();
 FILLCELL_X2 FILLER_47_1261 ();
 FILLCELL_X32 FILLER_47_1264 ();
 FILLCELL_X32 FILLER_47_1296 ();
 FILLCELL_X32 FILLER_47_1328 ();
 FILLCELL_X32 FILLER_47_1360 ();
 FILLCELL_X32 FILLER_47_1392 ();
 FILLCELL_X32 FILLER_47_1424 ();
 FILLCELL_X32 FILLER_47_1456 ();
 FILLCELL_X32 FILLER_47_1488 ();
 FILLCELL_X32 FILLER_47_1520 ();
 FILLCELL_X32 FILLER_47_1552 ();
 FILLCELL_X32 FILLER_47_1584 ();
 FILLCELL_X32 FILLER_47_1616 ();
 FILLCELL_X32 FILLER_47_1648 ();
 FILLCELL_X32 FILLER_47_1680 ();
 FILLCELL_X32 FILLER_47_1712 ();
 FILLCELL_X32 FILLER_47_1744 ();
 FILLCELL_X32 FILLER_47_1776 ();
 FILLCELL_X32 FILLER_47_1808 ();
 FILLCELL_X32 FILLER_47_1840 ();
 FILLCELL_X32 FILLER_47_1872 ();
 FILLCELL_X32 FILLER_47_1904 ();
 FILLCELL_X32 FILLER_47_1936 ();
 FILLCELL_X32 FILLER_47_1968 ();
 FILLCELL_X32 FILLER_47_2000 ();
 FILLCELL_X32 FILLER_47_2032 ();
 FILLCELL_X32 FILLER_47_2064 ();
 FILLCELL_X32 FILLER_47_2096 ();
 FILLCELL_X32 FILLER_47_2128 ();
 FILLCELL_X32 FILLER_47_2160 ();
 FILLCELL_X32 FILLER_47_2192 ();
 FILLCELL_X32 FILLER_47_2224 ();
 FILLCELL_X32 FILLER_47_2256 ();
 FILLCELL_X32 FILLER_47_2288 ();
 FILLCELL_X32 FILLER_47_2320 ();
 FILLCELL_X32 FILLER_47_2352 ();
 FILLCELL_X32 FILLER_47_2384 ();
 FILLCELL_X32 FILLER_47_2416 ();
 FILLCELL_X32 FILLER_47_2448 ();
 FILLCELL_X32 FILLER_47_2480 ();
 FILLCELL_X8 FILLER_47_2512 ();
 FILLCELL_X4 FILLER_47_2520 ();
 FILLCELL_X2 FILLER_47_2524 ();
 FILLCELL_X32 FILLER_47_2527 ();
 FILLCELL_X32 FILLER_47_2559 ();
 FILLCELL_X8 FILLER_47_2591 ();
 FILLCELL_X2 FILLER_47_2599 ();
 FILLCELL_X1 FILLER_47_2601 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X32 FILLER_48_33 ();
 FILLCELL_X32 FILLER_48_65 ();
 FILLCELL_X32 FILLER_48_97 ();
 FILLCELL_X32 FILLER_48_129 ();
 FILLCELL_X32 FILLER_48_161 ();
 FILLCELL_X32 FILLER_48_193 ();
 FILLCELL_X32 FILLER_48_225 ();
 FILLCELL_X32 FILLER_48_257 ();
 FILLCELL_X32 FILLER_48_289 ();
 FILLCELL_X32 FILLER_48_321 ();
 FILLCELL_X32 FILLER_48_353 ();
 FILLCELL_X32 FILLER_48_385 ();
 FILLCELL_X32 FILLER_48_417 ();
 FILLCELL_X32 FILLER_48_449 ();
 FILLCELL_X32 FILLER_48_481 ();
 FILLCELL_X32 FILLER_48_513 ();
 FILLCELL_X32 FILLER_48_545 ();
 FILLCELL_X32 FILLER_48_577 ();
 FILLCELL_X16 FILLER_48_609 ();
 FILLCELL_X4 FILLER_48_625 ();
 FILLCELL_X2 FILLER_48_629 ();
 FILLCELL_X32 FILLER_48_632 ();
 FILLCELL_X32 FILLER_48_664 ();
 FILLCELL_X32 FILLER_48_696 ();
 FILLCELL_X32 FILLER_48_728 ();
 FILLCELL_X32 FILLER_48_760 ();
 FILLCELL_X32 FILLER_48_792 ();
 FILLCELL_X32 FILLER_48_824 ();
 FILLCELL_X32 FILLER_48_856 ();
 FILLCELL_X32 FILLER_48_888 ();
 FILLCELL_X32 FILLER_48_920 ();
 FILLCELL_X32 FILLER_48_952 ();
 FILLCELL_X32 FILLER_48_984 ();
 FILLCELL_X32 FILLER_48_1016 ();
 FILLCELL_X32 FILLER_48_1048 ();
 FILLCELL_X32 FILLER_48_1080 ();
 FILLCELL_X32 FILLER_48_1112 ();
 FILLCELL_X32 FILLER_48_1144 ();
 FILLCELL_X32 FILLER_48_1176 ();
 FILLCELL_X32 FILLER_48_1208 ();
 FILLCELL_X32 FILLER_48_1240 ();
 FILLCELL_X32 FILLER_48_1272 ();
 FILLCELL_X32 FILLER_48_1304 ();
 FILLCELL_X32 FILLER_48_1336 ();
 FILLCELL_X32 FILLER_48_1368 ();
 FILLCELL_X32 FILLER_48_1400 ();
 FILLCELL_X32 FILLER_48_1432 ();
 FILLCELL_X32 FILLER_48_1464 ();
 FILLCELL_X32 FILLER_48_1496 ();
 FILLCELL_X32 FILLER_48_1528 ();
 FILLCELL_X32 FILLER_48_1560 ();
 FILLCELL_X32 FILLER_48_1592 ();
 FILLCELL_X32 FILLER_48_1624 ();
 FILLCELL_X32 FILLER_48_1656 ();
 FILLCELL_X32 FILLER_48_1688 ();
 FILLCELL_X32 FILLER_48_1720 ();
 FILLCELL_X32 FILLER_48_1752 ();
 FILLCELL_X32 FILLER_48_1784 ();
 FILLCELL_X32 FILLER_48_1816 ();
 FILLCELL_X32 FILLER_48_1848 ();
 FILLCELL_X8 FILLER_48_1880 ();
 FILLCELL_X4 FILLER_48_1888 ();
 FILLCELL_X2 FILLER_48_1892 ();
 FILLCELL_X32 FILLER_48_1895 ();
 FILLCELL_X32 FILLER_48_1927 ();
 FILLCELL_X32 FILLER_48_1959 ();
 FILLCELL_X32 FILLER_48_1991 ();
 FILLCELL_X32 FILLER_48_2023 ();
 FILLCELL_X32 FILLER_48_2055 ();
 FILLCELL_X32 FILLER_48_2087 ();
 FILLCELL_X32 FILLER_48_2119 ();
 FILLCELL_X32 FILLER_48_2151 ();
 FILLCELL_X32 FILLER_48_2183 ();
 FILLCELL_X32 FILLER_48_2215 ();
 FILLCELL_X32 FILLER_48_2247 ();
 FILLCELL_X32 FILLER_48_2279 ();
 FILLCELL_X32 FILLER_48_2311 ();
 FILLCELL_X32 FILLER_48_2343 ();
 FILLCELL_X32 FILLER_48_2375 ();
 FILLCELL_X32 FILLER_48_2407 ();
 FILLCELL_X32 FILLER_48_2439 ();
 FILLCELL_X32 FILLER_48_2471 ();
 FILLCELL_X32 FILLER_48_2503 ();
 FILLCELL_X32 FILLER_48_2535 ();
 FILLCELL_X32 FILLER_48_2567 ();
 FILLCELL_X2 FILLER_48_2599 ();
 FILLCELL_X1 FILLER_48_2601 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X32 FILLER_49_33 ();
 FILLCELL_X32 FILLER_49_65 ();
 FILLCELL_X32 FILLER_49_97 ();
 FILLCELL_X32 FILLER_49_129 ();
 FILLCELL_X32 FILLER_49_161 ();
 FILLCELL_X32 FILLER_49_193 ();
 FILLCELL_X32 FILLER_49_225 ();
 FILLCELL_X32 FILLER_49_257 ();
 FILLCELL_X32 FILLER_49_289 ();
 FILLCELL_X32 FILLER_49_321 ();
 FILLCELL_X32 FILLER_49_353 ();
 FILLCELL_X32 FILLER_49_385 ();
 FILLCELL_X32 FILLER_49_417 ();
 FILLCELL_X32 FILLER_49_449 ();
 FILLCELL_X32 FILLER_49_481 ();
 FILLCELL_X32 FILLER_49_513 ();
 FILLCELL_X32 FILLER_49_545 ();
 FILLCELL_X32 FILLER_49_577 ();
 FILLCELL_X32 FILLER_49_609 ();
 FILLCELL_X32 FILLER_49_641 ();
 FILLCELL_X32 FILLER_49_673 ();
 FILLCELL_X32 FILLER_49_705 ();
 FILLCELL_X32 FILLER_49_737 ();
 FILLCELL_X32 FILLER_49_769 ();
 FILLCELL_X32 FILLER_49_801 ();
 FILLCELL_X32 FILLER_49_833 ();
 FILLCELL_X32 FILLER_49_865 ();
 FILLCELL_X32 FILLER_49_897 ();
 FILLCELL_X32 FILLER_49_929 ();
 FILLCELL_X32 FILLER_49_961 ();
 FILLCELL_X32 FILLER_49_993 ();
 FILLCELL_X32 FILLER_49_1025 ();
 FILLCELL_X32 FILLER_49_1057 ();
 FILLCELL_X32 FILLER_49_1089 ();
 FILLCELL_X32 FILLER_49_1121 ();
 FILLCELL_X32 FILLER_49_1153 ();
 FILLCELL_X32 FILLER_49_1185 ();
 FILLCELL_X32 FILLER_49_1217 ();
 FILLCELL_X8 FILLER_49_1249 ();
 FILLCELL_X4 FILLER_49_1257 ();
 FILLCELL_X2 FILLER_49_1261 ();
 FILLCELL_X32 FILLER_49_1264 ();
 FILLCELL_X32 FILLER_49_1296 ();
 FILLCELL_X32 FILLER_49_1328 ();
 FILLCELL_X32 FILLER_49_1360 ();
 FILLCELL_X32 FILLER_49_1392 ();
 FILLCELL_X32 FILLER_49_1424 ();
 FILLCELL_X32 FILLER_49_1456 ();
 FILLCELL_X32 FILLER_49_1488 ();
 FILLCELL_X32 FILLER_49_1520 ();
 FILLCELL_X32 FILLER_49_1552 ();
 FILLCELL_X32 FILLER_49_1584 ();
 FILLCELL_X32 FILLER_49_1616 ();
 FILLCELL_X32 FILLER_49_1648 ();
 FILLCELL_X32 FILLER_49_1680 ();
 FILLCELL_X32 FILLER_49_1712 ();
 FILLCELL_X32 FILLER_49_1744 ();
 FILLCELL_X32 FILLER_49_1776 ();
 FILLCELL_X32 FILLER_49_1808 ();
 FILLCELL_X32 FILLER_49_1840 ();
 FILLCELL_X32 FILLER_49_1872 ();
 FILLCELL_X32 FILLER_49_1904 ();
 FILLCELL_X32 FILLER_49_1936 ();
 FILLCELL_X32 FILLER_49_1968 ();
 FILLCELL_X32 FILLER_49_2000 ();
 FILLCELL_X32 FILLER_49_2032 ();
 FILLCELL_X32 FILLER_49_2064 ();
 FILLCELL_X32 FILLER_49_2096 ();
 FILLCELL_X32 FILLER_49_2128 ();
 FILLCELL_X32 FILLER_49_2160 ();
 FILLCELL_X32 FILLER_49_2192 ();
 FILLCELL_X32 FILLER_49_2224 ();
 FILLCELL_X32 FILLER_49_2256 ();
 FILLCELL_X32 FILLER_49_2288 ();
 FILLCELL_X32 FILLER_49_2320 ();
 FILLCELL_X32 FILLER_49_2352 ();
 FILLCELL_X32 FILLER_49_2384 ();
 FILLCELL_X32 FILLER_49_2416 ();
 FILLCELL_X32 FILLER_49_2448 ();
 FILLCELL_X32 FILLER_49_2480 ();
 FILLCELL_X8 FILLER_49_2512 ();
 FILLCELL_X4 FILLER_49_2520 ();
 FILLCELL_X2 FILLER_49_2524 ();
 FILLCELL_X32 FILLER_49_2527 ();
 FILLCELL_X32 FILLER_49_2559 ();
 FILLCELL_X8 FILLER_49_2591 ();
 FILLCELL_X2 FILLER_49_2599 ();
 FILLCELL_X1 FILLER_49_2601 ();
 FILLCELL_X32 FILLER_50_1 ();
 FILLCELL_X32 FILLER_50_33 ();
 FILLCELL_X32 FILLER_50_65 ();
 FILLCELL_X32 FILLER_50_97 ();
 FILLCELL_X32 FILLER_50_129 ();
 FILLCELL_X32 FILLER_50_161 ();
 FILLCELL_X32 FILLER_50_193 ();
 FILLCELL_X32 FILLER_50_225 ();
 FILLCELL_X32 FILLER_50_257 ();
 FILLCELL_X32 FILLER_50_289 ();
 FILLCELL_X32 FILLER_50_321 ();
 FILLCELL_X32 FILLER_50_353 ();
 FILLCELL_X32 FILLER_50_385 ();
 FILLCELL_X32 FILLER_50_417 ();
 FILLCELL_X32 FILLER_50_449 ();
 FILLCELL_X32 FILLER_50_481 ();
 FILLCELL_X32 FILLER_50_513 ();
 FILLCELL_X32 FILLER_50_545 ();
 FILLCELL_X32 FILLER_50_577 ();
 FILLCELL_X16 FILLER_50_609 ();
 FILLCELL_X4 FILLER_50_625 ();
 FILLCELL_X2 FILLER_50_629 ();
 FILLCELL_X32 FILLER_50_632 ();
 FILLCELL_X32 FILLER_50_664 ();
 FILLCELL_X32 FILLER_50_696 ();
 FILLCELL_X32 FILLER_50_728 ();
 FILLCELL_X32 FILLER_50_760 ();
 FILLCELL_X32 FILLER_50_792 ();
 FILLCELL_X32 FILLER_50_824 ();
 FILLCELL_X32 FILLER_50_856 ();
 FILLCELL_X32 FILLER_50_888 ();
 FILLCELL_X32 FILLER_50_920 ();
 FILLCELL_X32 FILLER_50_952 ();
 FILLCELL_X32 FILLER_50_984 ();
 FILLCELL_X32 FILLER_50_1016 ();
 FILLCELL_X32 FILLER_50_1048 ();
 FILLCELL_X32 FILLER_50_1080 ();
 FILLCELL_X32 FILLER_50_1112 ();
 FILLCELL_X32 FILLER_50_1144 ();
 FILLCELL_X32 FILLER_50_1176 ();
 FILLCELL_X32 FILLER_50_1208 ();
 FILLCELL_X32 FILLER_50_1240 ();
 FILLCELL_X32 FILLER_50_1272 ();
 FILLCELL_X32 FILLER_50_1304 ();
 FILLCELL_X32 FILLER_50_1336 ();
 FILLCELL_X32 FILLER_50_1368 ();
 FILLCELL_X32 FILLER_50_1400 ();
 FILLCELL_X32 FILLER_50_1432 ();
 FILLCELL_X32 FILLER_50_1464 ();
 FILLCELL_X32 FILLER_50_1496 ();
 FILLCELL_X32 FILLER_50_1528 ();
 FILLCELL_X32 FILLER_50_1560 ();
 FILLCELL_X32 FILLER_50_1592 ();
 FILLCELL_X32 FILLER_50_1624 ();
 FILLCELL_X32 FILLER_50_1656 ();
 FILLCELL_X32 FILLER_50_1688 ();
 FILLCELL_X32 FILLER_50_1720 ();
 FILLCELL_X32 FILLER_50_1752 ();
 FILLCELL_X32 FILLER_50_1784 ();
 FILLCELL_X32 FILLER_50_1816 ();
 FILLCELL_X32 FILLER_50_1848 ();
 FILLCELL_X8 FILLER_50_1880 ();
 FILLCELL_X4 FILLER_50_1888 ();
 FILLCELL_X2 FILLER_50_1892 ();
 FILLCELL_X32 FILLER_50_1895 ();
 FILLCELL_X32 FILLER_50_1927 ();
 FILLCELL_X32 FILLER_50_1959 ();
 FILLCELL_X32 FILLER_50_1991 ();
 FILLCELL_X32 FILLER_50_2023 ();
 FILLCELL_X32 FILLER_50_2055 ();
 FILLCELL_X32 FILLER_50_2087 ();
 FILLCELL_X32 FILLER_50_2119 ();
 FILLCELL_X32 FILLER_50_2151 ();
 FILLCELL_X32 FILLER_50_2183 ();
 FILLCELL_X32 FILLER_50_2215 ();
 FILLCELL_X32 FILLER_50_2247 ();
 FILLCELL_X32 FILLER_50_2279 ();
 FILLCELL_X32 FILLER_50_2311 ();
 FILLCELL_X32 FILLER_50_2343 ();
 FILLCELL_X32 FILLER_50_2375 ();
 FILLCELL_X32 FILLER_50_2407 ();
 FILLCELL_X32 FILLER_50_2439 ();
 FILLCELL_X32 FILLER_50_2471 ();
 FILLCELL_X32 FILLER_50_2503 ();
 FILLCELL_X32 FILLER_50_2535 ();
 FILLCELL_X32 FILLER_50_2567 ();
 FILLCELL_X2 FILLER_50_2599 ();
 FILLCELL_X1 FILLER_50_2601 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X32 FILLER_51_33 ();
 FILLCELL_X32 FILLER_51_65 ();
 FILLCELL_X32 FILLER_51_97 ();
 FILLCELL_X32 FILLER_51_129 ();
 FILLCELL_X32 FILLER_51_161 ();
 FILLCELL_X32 FILLER_51_193 ();
 FILLCELL_X32 FILLER_51_225 ();
 FILLCELL_X32 FILLER_51_257 ();
 FILLCELL_X32 FILLER_51_289 ();
 FILLCELL_X32 FILLER_51_321 ();
 FILLCELL_X32 FILLER_51_353 ();
 FILLCELL_X32 FILLER_51_385 ();
 FILLCELL_X32 FILLER_51_417 ();
 FILLCELL_X32 FILLER_51_449 ();
 FILLCELL_X32 FILLER_51_481 ();
 FILLCELL_X32 FILLER_51_513 ();
 FILLCELL_X32 FILLER_51_545 ();
 FILLCELL_X32 FILLER_51_577 ();
 FILLCELL_X32 FILLER_51_609 ();
 FILLCELL_X32 FILLER_51_641 ();
 FILLCELL_X32 FILLER_51_673 ();
 FILLCELL_X32 FILLER_51_705 ();
 FILLCELL_X32 FILLER_51_737 ();
 FILLCELL_X32 FILLER_51_769 ();
 FILLCELL_X32 FILLER_51_801 ();
 FILLCELL_X32 FILLER_51_833 ();
 FILLCELL_X32 FILLER_51_865 ();
 FILLCELL_X32 FILLER_51_897 ();
 FILLCELL_X32 FILLER_51_929 ();
 FILLCELL_X32 FILLER_51_961 ();
 FILLCELL_X32 FILLER_51_993 ();
 FILLCELL_X32 FILLER_51_1025 ();
 FILLCELL_X32 FILLER_51_1057 ();
 FILLCELL_X32 FILLER_51_1089 ();
 FILLCELL_X32 FILLER_51_1121 ();
 FILLCELL_X32 FILLER_51_1153 ();
 FILLCELL_X32 FILLER_51_1185 ();
 FILLCELL_X32 FILLER_51_1217 ();
 FILLCELL_X8 FILLER_51_1249 ();
 FILLCELL_X4 FILLER_51_1257 ();
 FILLCELL_X2 FILLER_51_1261 ();
 FILLCELL_X32 FILLER_51_1264 ();
 FILLCELL_X32 FILLER_51_1296 ();
 FILLCELL_X32 FILLER_51_1328 ();
 FILLCELL_X32 FILLER_51_1360 ();
 FILLCELL_X32 FILLER_51_1392 ();
 FILLCELL_X32 FILLER_51_1424 ();
 FILLCELL_X32 FILLER_51_1456 ();
 FILLCELL_X32 FILLER_51_1488 ();
 FILLCELL_X32 FILLER_51_1520 ();
 FILLCELL_X32 FILLER_51_1552 ();
 FILLCELL_X32 FILLER_51_1584 ();
 FILLCELL_X32 FILLER_51_1616 ();
 FILLCELL_X32 FILLER_51_1648 ();
 FILLCELL_X32 FILLER_51_1680 ();
 FILLCELL_X32 FILLER_51_1712 ();
 FILLCELL_X32 FILLER_51_1744 ();
 FILLCELL_X32 FILLER_51_1776 ();
 FILLCELL_X32 FILLER_51_1808 ();
 FILLCELL_X32 FILLER_51_1840 ();
 FILLCELL_X32 FILLER_51_1872 ();
 FILLCELL_X32 FILLER_51_1904 ();
 FILLCELL_X32 FILLER_51_1936 ();
 FILLCELL_X32 FILLER_51_1968 ();
 FILLCELL_X32 FILLER_51_2000 ();
 FILLCELL_X32 FILLER_51_2032 ();
 FILLCELL_X32 FILLER_51_2064 ();
 FILLCELL_X32 FILLER_51_2096 ();
 FILLCELL_X32 FILLER_51_2128 ();
 FILLCELL_X32 FILLER_51_2160 ();
 FILLCELL_X32 FILLER_51_2192 ();
 FILLCELL_X32 FILLER_51_2224 ();
 FILLCELL_X32 FILLER_51_2256 ();
 FILLCELL_X32 FILLER_51_2288 ();
 FILLCELL_X32 FILLER_51_2320 ();
 FILLCELL_X32 FILLER_51_2352 ();
 FILLCELL_X32 FILLER_51_2384 ();
 FILLCELL_X32 FILLER_51_2416 ();
 FILLCELL_X32 FILLER_51_2448 ();
 FILLCELL_X32 FILLER_51_2480 ();
 FILLCELL_X8 FILLER_51_2512 ();
 FILLCELL_X4 FILLER_51_2520 ();
 FILLCELL_X2 FILLER_51_2524 ();
 FILLCELL_X32 FILLER_51_2527 ();
 FILLCELL_X32 FILLER_51_2559 ();
 FILLCELL_X8 FILLER_51_2591 ();
 FILLCELL_X2 FILLER_51_2599 ();
 FILLCELL_X1 FILLER_51_2601 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X32 FILLER_52_33 ();
 FILLCELL_X32 FILLER_52_65 ();
 FILLCELL_X32 FILLER_52_97 ();
 FILLCELL_X32 FILLER_52_129 ();
 FILLCELL_X32 FILLER_52_161 ();
 FILLCELL_X32 FILLER_52_193 ();
 FILLCELL_X32 FILLER_52_225 ();
 FILLCELL_X32 FILLER_52_257 ();
 FILLCELL_X32 FILLER_52_289 ();
 FILLCELL_X32 FILLER_52_321 ();
 FILLCELL_X32 FILLER_52_353 ();
 FILLCELL_X32 FILLER_52_385 ();
 FILLCELL_X32 FILLER_52_417 ();
 FILLCELL_X32 FILLER_52_449 ();
 FILLCELL_X32 FILLER_52_481 ();
 FILLCELL_X32 FILLER_52_513 ();
 FILLCELL_X32 FILLER_52_545 ();
 FILLCELL_X32 FILLER_52_577 ();
 FILLCELL_X16 FILLER_52_609 ();
 FILLCELL_X4 FILLER_52_625 ();
 FILLCELL_X2 FILLER_52_629 ();
 FILLCELL_X32 FILLER_52_632 ();
 FILLCELL_X32 FILLER_52_664 ();
 FILLCELL_X32 FILLER_52_696 ();
 FILLCELL_X32 FILLER_52_728 ();
 FILLCELL_X32 FILLER_52_760 ();
 FILLCELL_X32 FILLER_52_792 ();
 FILLCELL_X32 FILLER_52_824 ();
 FILLCELL_X32 FILLER_52_856 ();
 FILLCELL_X32 FILLER_52_888 ();
 FILLCELL_X32 FILLER_52_920 ();
 FILLCELL_X32 FILLER_52_952 ();
 FILLCELL_X32 FILLER_52_984 ();
 FILLCELL_X32 FILLER_52_1016 ();
 FILLCELL_X32 FILLER_52_1048 ();
 FILLCELL_X32 FILLER_52_1080 ();
 FILLCELL_X32 FILLER_52_1112 ();
 FILLCELL_X32 FILLER_52_1144 ();
 FILLCELL_X32 FILLER_52_1176 ();
 FILLCELL_X32 FILLER_52_1208 ();
 FILLCELL_X32 FILLER_52_1240 ();
 FILLCELL_X32 FILLER_52_1272 ();
 FILLCELL_X32 FILLER_52_1304 ();
 FILLCELL_X32 FILLER_52_1336 ();
 FILLCELL_X32 FILLER_52_1368 ();
 FILLCELL_X32 FILLER_52_1400 ();
 FILLCELL_X32 FILLER_52_1432 ();
 FILLCELL_X32 FILLER_52_1464 ();
 FILLCELL_X32 FILLER_52_1496 ();
 FILLCELL_X32 FILLER_52_1528 ();
 FILLCELL_X32 FILLER_52_1560 ();
 FILLCELL_X32 FILLER_52_1592 ();
 FILLCELL_X32 FILLER_52_1624 ();
 FILLCELL_X32 FILLER_52_1656 ();
 FILLCELL_X32 FILLER_52_1688 ();
 FILLCELL_X32 FILLER_52_1720 ();
 FILLCELL_X32 FILLER_52_1752 ();
 FILLCELL_X32 FILLER_52_1784 ();
 FILLCELL_X32 FILLER_52_1816 ();
 FILLCELL_X32 FILLER_52_1848 ();
 FILLCELL_X8 FILLER_52_1880 ();
 FILLCELL_X4 FILLER_52_1888 ();
 FILLCELL_X2 FILLER_52_1892 ();
 FILLCELL_X32 FILLER_52_1895 ();
 FILLCELL_X32 FILLER_52_1927 ();
 FILLCELL_X32 FILLER_52_1959 ();
 FILLCELL_X32 FILLER_52_1991 ();
 FILLCELL_X32 FILLER_52_2023 ();
 FILLCELL_X32 FILLER_52_2055 ();
 FILLCELL_X32 FILLER_52_2087 ();
 FILLCELL_X32 FILLER_52_2119 ();
 FILLCELL_X32 FILLER_52_2151 ();
 FILLCELL_X32 FILLER_52_2183 ();
 FILLCELL_X32 FILLER_52_2215 ();
 FILLCELL_X32 FILLER_52_2247 ();
 FILLCELL_X32 FILLER_52_2279 ();
 FILLCELL_X32 FILLER_52_2311 ();
 FILLCELL_X32 FILLER_52_2343 ();
 FILLCELL_X32 FILLER_52_2375 ();
 FILLCELL_X32 FILLER_52_2407 ();
 FILLCELL_X32 FILLER_52_2439 ();
 FILLCELL_X32 FILLER_52_2471 ();
 FILLCELL_X32 FILLER_52_2503 ();
 FILLCELL_X32 FILLER_52_2535 ();
 FILLCELL_X32 FILLER_52_2567 ();
 FILLCELL_X2 FILLER_52_2599 ();
 FILLCELL_X1 FILLER_52_2601 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X32 FILLER_53_33 ();
 FILLCELL_X32 FILLER_53_65 ();
 FILLCELL_X32 FILLER_53_97 ();
 FILLCELL_X32 FILLER_53_129 ();
 FILLCELL_X32 FILLER_53_161 ();
 FILLCELL_X32 FILLER_53_193 ();
 FILLCELL_X32 FILLER_53_225 ();
 FILLCELL_X32 FILLER_53_257 ();
 FILLCELL_X32 FILLER_53_289 ();
 FILLCELL_X32 FILLER_53_321 ();
 FILLCELL_X32 FILLER_53_353 ();
 FILLCELL_X32 FILLER_53_385 ();
 FILLCELL_X32 FILLER_53_417 ();
 FILLCELL_X32 FILLER_53_449 ();
 FILLCELL_X32 FILLER_53_481 ();
 FILLCELL_X32 FILLER_53_513 ();
 FILLCELL_X32 FILLER_53_545 ();
 FILLCELL_X32 FILLER_53_577 ();
 FILLCELL_X32 FILLER_53_609 ();
 FILLCELL_X32 FILLER_53_641 ();
 FILLCELL_X32 FILLER_53_673 ();
 FILLCELL_X32 FILLER_53_705 ();
 FILLCELL_X32 FILLER_53_737 ();
 FILLCELL_X32 FILLER_53_769 ();
 FILLCELL_X32 FILLER_53_801 ();
 FILLCELL_X32 FILLER_53_833 ();
 FILLCELL_X32 FILLER_53_865 ();
 FILLCELL_X32 FILLER_53_897 ();
 FILLCELL_X32 FILLER_53_929 ();
 FILLCELL_X32 FILLER_53_961 ();
 FILLCELL_X32 FILLER_53_993 ();
 FILLCELL_X32 FILLER_53_1025 ();
 FILLCELL_X32 FILLER_53_1057 ();
 FILLCELL_X32 FILLER_53_1089 ();
 FILLCELL_X32 FILLER_53_1121 ();
 FILLCELL_X32 FILLER_53_1153 ();
 FILLCELL_X32 FILLER_53_1185 ();
 FILLCELL_X32 FILLER_53_1217 ();
 FILLCELL_X8 FILLER_53_1249 ();
 FILLCELL_X4 FILLER_53_1257 ();
 FILLCELL_X2 FILLER_53_1261 ();
 FILLCELL_X32 FILLER_53_1264 ();
 FILLCELL_X32 FILLER_53_1296 ();
 FILLCELL_X32 FILLER_53_1328 ();
 FILLCELL_X32 FILLER_53_1360 ();
 FILLCELL_X32 FILLER_53_1392 ();
 FILLCELL_X32 FILLER_53_1424 ();
 FILLCELL_X32 FILLER_53_1456 ();
 FILLCELL_X32 FILLER_53_1488 ();
 FILLCELL_X32 FILLER_53_1520 ();
 FILLCELL_X32 FILLER_53_1552 ();
 FILLCELL_X32 FILLER_53_1584 ();
 FILLCELL_X32 FILLER_53_1616 ();
 FILLCELL_X32 FILLER_53_1648 ();
 FILLCELL_X32 FILLER_53_1680 ();
 FILLCELL_X32 FILLER_53_1712 ();
 FILLCELL_X32 FILLER_53_1744 ();
 FILLCELL_X32 FILLER_53_1776 ();
 FILLCELL_X32 FILLER_53_1808 ();
 FILLCELL_X32 FILLER_53_1840 ();
 FILLCELL_X32 FILLER_53_1872 ();
 FILLCELL_X32 FILLER_53_1904 ();
 FILLCELL_X32 FILLER_53_1936 ();
 FILLCELL_X32 FILLER_53_1968 ();
 FILLCELL_X32 FILLER_53_2000 ();
 FILLCELL_X32 FILLER_53_2032 ();
 FILLCELL_X32 FILLER_53_2064 ();
 FILLCELL_X32 FILLER_53_2096 ();
 FILLCELL_X32 FILLER_53_2128 ();
 FILLCELL_X32 FILLER_53_2160 ();
 FILLCELL_X32 FILLER_53_2192 ();
 FILLCELL_X32 FILLER_53_2224 ();
 FILLCELL_X32 FILLER_53_2256 ();
 FILLCELL_X32 FILLER_53_2288 ();
 FILLCELL_X32 FILLER_53_2320 ();
 FILLCELL_X32 FILLER_53_2352 ();
 FILLCELL_X32 FILLER_53_2384 ();
 FILLCELL_X32 FILLER_53_2416 ();
 FILLCELL_X32 FILLER_53_2448 ();
 FILLCELL_X32 FILLER_53_2480 ();
 FILLCELL_X8 FILLER_53_2512 ();
 FILLCELL_X4 FILLER_53_2520 ();
 FILLCELL_X2 FILLER_53_2524 ();
 FILLCELL_X32 FILLER_53_2527 ();
 FILLCELL_X32 FILLER_53_2559 ();
 FILLCELL_X8 FILLER_53_2591 ();
 FILLCELL_X2 FILLER_53_2599 ();
 FILLCELL_X1 FILLER_53_2601 ();
 FILLCELL_X32 FILLER_54_1 ();
 FILLCELL_X32 FILLER_54_33 ();
 FILLCELL_X32 FILLER_54_65 ();
 FILLCELL_X32 FILLER_54_97 ();
 FILLCELL_X32 FILLER_54_129 ();
 FILLCELL_X32 FILLER_54_161 ();
 FILLCELL_X32 FILLER_54_193 ();
 FILLCELL_X32 FILLER_54_225 ();
 FILLCELL_X32 FILLER_54_257 ();
 FILLCELL_X32 FILLER_54_289 ();
 FILLCELL_X32 FILLER_54_321 ();
 FILLCELL_X32 FILLER_54_353 ();
 FILLCELL_X32 FILLER_54_385 ();
 FILLCELL_X32 FILLER_54_417 ();
 FILLCELL_X32 FILLER_54_449 ();
 FILLCELL_X32 FILLER_54_481 ();
 FILLCELL_X32 FILLER_54_513 ();
 FILLCELL_X32 FILLER_54_545 ();
 FILLCELL_X32 FILLER_54_577 ();
 FILLCELL_X16 FILLER_54_609 ();
 FILLCELL_X4 FILLER_54_625 ();
 FILLCELL_X2 FILLER_54_629 ();
 FILLCELL_X32 FILLER_54_632 ();
 FILLCELL_X32 FILLER_54_664 ();
 FILLCELL_X32 FILLER_54_696 ();
 FILLCELL_X32 FILLER_54_728 ();
 FILLCELL_X32 FILLER_54_760 ();
 FILLCELL_X32 FILLER_54_792 ();
 FILLCELL_X32 FILLER_54_824 ();
 FILLCELL_X32 FILLER_54_856 ();
 FILLCELL_X32 FILLER_54_888 ();
 FILLCELL_X32 FILLER_54_920 ();
 FILLCELL_X32 FILLER_54_952 ();
 FILLCELL_X32 FILLER_54_984 ();
 FILLCELL_X32 FILLER_54_1016 ();
 FILLCELL_X32 FILLER_54_1048 ();
 FILLCELL_X32 FILLER_54_1080 ();
 FILLCELL_X32 FILLER_54_1112 ();
 FILLCELL_X32 FILLER_54_1144 ();
 FILLCELL_X32 FILLER_54_1176 ();
 FILLCELL_X32 FILLER_54_1208 ();
 FILLCELL_X32 FILLER_54_1240 ();
 FILLCELL_X32 FILLER_54_1272 ();
 FILLCELL_X32 FILLER_54_1304 ();
 FILLCELL_X32 FILLER_54_1336 ();
 FILLCELL_X32 FILLER_54_1368 ();
 FILLCELL_X32 FILLER_54_1400 ();
 FILLCELL_X32 FILLER_54_1432 ();
 FILLCELL_X32 FILLER_54_1464 ();
 FILLCELL_X32 FILLER_54_1496 ();
 FILLCELL_X32 FILLER_54_1528 ();
 FILLCELL_X32 FILLER_54_1560 ();
 FILLCELL_X32 FILLER_54_1592 ();
 FILLCELL_X32 FILLER_54_1624 ();
 FILLCELL_X32 FILLER_54_1656 ();
 FILLCELL_X32 FILLER_54_1688 ();
 FILLCELL_X32 FILLER_54_1720 ();
 FILLCELL_X32 FILLER_54_1752 ();
 FILLCELL_X32 FILLER_54_1784 ();
 FILLCELL_X32 FILLER_54_1816 ();
 FILLCELL_X32 FILLER_54_1848 ();
 FILLCELL_X8 FILLER_54_1880 ();
 FILLCELL_X4 FILLER_54_1888 ();
 FILLCELL_X2 FILLER_54_1892 ();
 FILLCELL_X32 FILLER_54_1895 ();
 FILLCELL_X32 FILLER_54_1927 ();
 FILLCELL_X32 FILLER_54_1959 ();
 FILLCELL_X32 FILLER_54_1991 ();
 FILLCELL_X32 FILLER_54_2023 ();
 FILLCELL_X32 FILLER_54_2055 ();
 FILLCELL_X32 FILLER_54_2087 ();
 FILLCELL_X32 FILLER_54_2119 ();
 FILLCELL_X32 FILLER_54_2151 ();
 FILLCELL_X32 FILLER_54_2183 ();
 FILLCELL_X32 FILLER_54_2215 ();
 FILLCELL_X32 FILLER_54_2247 ();
 FILLCELL_X32 FILLER_54_2279 ();
 FILLCELL_X32 FILLER_54_2311 ();
 FILLCELL_X32 FILLER_54_2343 ();
 FILLCELL_X32 FILLER_54_2375 ();
 FILLCELL_X32 FILLER_54_2407 ();
 FILLCELL_X32 FILLER_54_2439 ();
 FILLCELL_X32 FILLER_54_2471 ();
 FILLCELL_X32 FILLER_54_2503 ();
 FILLCELL_X32 FILLER_54_2535 ();
 FILLCELL_X32 FILLER_54_2567 ();
 FILLCELL_X2 FILLER_54_2599 ();
 FILLCELL_X1 FILLER_54_2601 ();
 FILLCELL_X32 FILLER_55_1 ();
 FILLCELL_X32 FILLER_55_33 ();
 FILLCELL_X32 FILLER_55_65 ();
 FILLCELL_X32 FILLER_55_97 ();
 FILLCELL_X32 FILLER_55_129 ();
 FILLCELL_X32 FILLER_55_161 ();
 FILLCELL_X32 FILLER_55_193 ();
 FILLCELL_X32 FILLER_55_225 ();
 FILLCELL_X32 FILLER_55_257 ();
 FILLCELL_X32 FILLER_55_289 ();
 FILLCELL_X32 FILLER_55_321 ();
 FILLCELL_X32 FILLER_55_353 ();
 FILLCELL_X32 FILLER_55_385 ();
 FILLCELL_X32 FILLER_55_417 ();
 FILLCELL_X32 FILLER_55_449 ();
 FILLCELL_X32 FILLER_55_481 ();
 FILLCELL_X32 FILLER_55_513 ();
 FILLCELL_X32 FILLER_55_545 ();
 FILLCELL_X32 FILLER_55_577 ();
 FILLCELL_X32 FILLER_55_609 ();
 FILLCELL_X32 FILLER_55_641 ();
 FILLCELL_X32 FILLER_55_673 ();
 FILLCELL_X32 FILLER_55_705 ();
 FILLCELL_X32 FILLER_55_737 ();
 FILLCELL_X32 FILLER_55_769 ();
 FILLCELL_X32 FILLER_55_801 ();
 FILLCELL_X32 FILLER_55_833 ();
 FILLCELL_X32 FILLER_55_865 ();
 FILLCELL_X32 FILLER_55_897 ();
 FILLCELL_X32 FILLER_55_929 ();
 FILLCELL_X32 FILLER_55_961 ();
 FILLCELL_X32 FILLER_55_993 ();
 FILLCELL_X32 FILLER_55_1025 ();
 FILLCELL_X32 FILLER_55_1057 ();
 FILLCELL_X32 FILLER_55_1089 ();
 FILLCELL_X32 FILLER_55_1121 ();
 FILLCELL_X32 FILLER_55_1153 ();
 FILLCELL_X32 FILLER_55_1185 ();
 FILLCELL_X32 FILLER_55_1217 ();
 FILLCELL_X8 FILLER_55_1249 ();
 FILLCELL_X4 FILLER_55_1257 ();
 FILLCELL_X2 FILLER_55_1261 ();
 FILLCELL_X32 FILLER_55_1264 ();
 FILLCELL_X32 FILLER_55_1296 ();
 FILLCELL_X32 FILLER_55_1328 ();
 FILLCELL_X32 FILLER_55_1360 ();
 FILLCELL_X32 FILLER_55_1392 ();
 FILLCELL_X32 FILLER_55_1424 ();
 FILLCELL_X32 FILLER_55_1456 ();
 FILLCELL_X32 FILLER_55_1488 ();
 FILLCELL_X32 FILLER_55_1520 ();
 FILLCELL_X32 FILLER_55_1552 ();
 FILLCELL_X32 FILLER_55_1584 ();
 FILLCELL_X32 FILLER_55_1616 ();
 FILLCELL_X32 FILLER_55_1648 ();
 FILLCELL_X32 FILLER_55_1680 ();
 FILLCELL_X32 FILLER_55_1712 ();
 FILLCELL_X32 FILLER_55_1744 ();
 FILLCELL_X32 FILLER_55_1776 ();
 FILLCELL_X32 FILLER_55_1808 ();
 FILLCELL_X32 FILLER_55_1840 ();
 FILLCELL_X32 FILLER_55_1872 ();
 FILLCELL_X32 FILLER_55_1904 ();
 FILLCELL_X32 FILLER_55_1936 ();
 FILLCELL_X32 FILLER_55_1968 ();
 FILLCELL_X32 FILLER_55_2000 ();
 FILLCELL_X32 FILLER_55_2032 ();
 FILLCELL_X32 FILLER_55_2064 ();
 FILLCELL_X32 FILLER_55_2096 ();
 FILLCELL_X32 FILLER_55_2128 ();
 FILLCELL_X32 FILLER_55_2160 ();
 FILLCELL_X32 FILLER_55_2192 ();
 FILLCELL_X32 FILLER_55_2224 ();
 FILLCELL_X32 FILLER_55_2256 ();
 FILLCELL_X32 FILLER_55_2288 ();
 FILLCELL_X32 FILLER_55_2320 ();
 FILLCELL_X32 FILLER_55_2352 ();
 FILLCELL_X32 FILLER_55_2384 ();
 FILLCELL_X32 FILLER_55_2416 ();
 FILLCELL_X32 FILLER_55_2448 ();
 FILLCELL_X32 FILLER_55_2480 ();
 FILLCELL_X8 FILLER_55_2512 ();
 FILLCELL_X4 FILLER_55_2520 ();
 FILLCELL_X2 FILLER_55_2524 ();
 FILLCELL_X32 FILLER_55_2527 ();
 FILLCELL_X32 FILLER_55_2559 ();
 FILLCELL_X8 FILLER_55_2591 ();
 FILLCELL_X2 FILLER_55_2599 ();
 FILLCELL_X1 FILLER_55_2601 ();
 FILLCELL_X32 FILLER_56_1 ();
 FILLCELL_X32 FILLER_56_33 ();
 FILLCELL_X32 FILLER_56_65 ();
 FILLCELL_X32 FILLER_56_97 ();
 FILLCELL_X32 FILLER_56_129 ();
 FILLCELL_X32 FILLER_56_161 ();
 FILLCELL_X32 FILLER_56_193 ();
 FILLCELL_X32 FILLER_56_225 ();
 FILLCELL_X32 FILLER_56_257 ();
 FILLCELL_X32 FILLER_56_289 ();
 FILLCELL_X32 FILLER_56_321 ();
 FILLCELL_X32 FILLER_56_353 ();
 FILLCELL_X32 FILLER_56_385 ();
 FILLCELL_X32 FILLER_56_417 ();
 FILLCELL_X32 FILLER_56_449 ();
 FILLCELL_X32 FILLER_56_481 ();
 FILLCELL_X32 FILLER_56_513 ();
 FILLCELL_X32 FILLER_56_545 ();
 FILLCELL_X32 FILLER_56_577 ();
 FILLCELL_X16 FILLER_56_609 ();
 FILLCELL_X4 FILLER_56_625 ();
 FILLCELL_X2 FILLER_56_629 ();
 FILLCELL_X32 FILLER_56_632 ();
 FILLCELL_X32 FILLER_56_664 ();
 FILLCELL_X32 FILLER_56_696 ();
 FILLCELL_X32 FILLER_56_728 ();
 FILLCELL_X32 FILLER_56_760 ();
 FILLCELL_X32 FILLER_56_792 ();
 FILLCELL_X32 FILLER_56_824 ();
 FILLCELL_X32 FILLER_56_856 ();
 FILLCELL_X32 FILLER_56_888 ();
 FILLCELL_X32 FILLER_56_920 ();
 FILLCELL_X32 FILLER_56_952 ();
 FILLCELL_X32 FILLER_56_984 ();
 FILLCELL_X32 FILLER_56_1016 ();
 FILLCELL_X32 FILLER_56_1048 ();
 FILLCELL_X32 FILLER_56_1080 ();
 FILLCELL_X32 FILLER_56_1112 ();
 FILLCELL_X32 FILLER_56_1144 ();
 FILLCELL_X32 FILLER_56_1176 ();
 FILLCELL_X32 FILLER_56_1208 ();
 FILLCELL_X32 FILLER_56_1240 ();
 FILLCELL_X32 FILLER_56_1272 ();
 FILLCELL_X32 FILLER_56_1304 ();
 FILLCELL_X32 FILLER_56_1336 ();
 FILLCELL_X32 FILLER_56_1368 ();
 FILLCELL_X32 FILLER_56_1400 ();
 FILLCELL_X32 FILLER_56_1432 ();
 FILLCELL_X32 FILLER_56_1464 ();
 FILLCELL_X32 FILLER_56_1496 ();
 FILLCELL_X32 FILLER_56_1528 ();
 FILLCELL_X32 FILLER_56_1560 ();
 FILLCELL_X32 FILLER_56_1592 ();
 FILLCELL_X32 FILLER_56_1624 ();
 FILLCELL_X32 FILLER_56_1656 ();
 FILLCELL_X32 FILLER_56_1688 ();
 FILLCELL_X32 FILLER_56_1720 ();
 FILLCELL_X32 FILLER_56_1752 ();
 FILLCELL_X32 FILLER_56_1784 ();
 FILLCELL_X32 FILLER_56_1816 ();
 FILLCELL_X32 FILLER_56_1848 ();
 FILLCELL_X8 FILLER_56_1880 ();
 FILLCELL_X4 FILLER_56_1888 ();
 FILLCELL_X2 FILLER_56_1892 ();
 FILLCELL_X32 FILLER_56_1895 ();
 FILLCELL_X32 FILLER_56_1927 ();
 FILLCELL_X32 FILLER_56_1959 ();
 FILLCELL_X32 FILLER_56_1991 ();
 FILLCELL_X32 FILLER_56_2023 ();
 FILLCELL_X32 FILLER_56_2055 ();
 FILLCELL_X32 FILLER_56_2087 ();
 FILLCELL_X32 FILLER_56_2119 ();
 FILLCELL_X32 FILLER_56_2151 ();
 FILLCELL_X32 FILLER_56_2183 ();
 FILLCELL_X32 FILLER_56_2215 ();
 FILLCELL_X32 FILLER_56_2247 ();
 FILLCELL_X32 FILLER_56_2279 ();
 FILLCELL_X32 FILLER_56_2311 ();
 FILLCELL_X32 FILLER_56_2343 ();
 FILLCELL_X32 FILLER_56_2375 ();
 FILLCELL_X32 FILLER_56_2407 ();
 FILLCELL_X32 FILLER_56_2439 ();
 FILLCELL_X32 FILLER_56_2471 ();
 FILLCELL_X32 FILLER_56_2503 ();
 FILLCELL_X32 FILLER_56_2535 ();
 FILLCELL_X32 FILLER_56_2567 ();
 FILLCELL_X2 FILLER_56_2599 ();
 FILLCELL_X1 FILLER_56_2601 ();
 FILLCELL_X32 FILLER_57_1 ();
 FILLCELL_X32 FILLER_57_33 ();
 FILLCELL_X32 FILLER_57_65 ();
 FILLCELL_X32 FILLER_57_97 ();
 FILLCELL_X32 FILLER_57_129 ();
 FILLCELL_X32 FILLER_57_161 ();
 FILLCELL_X32 FILLER_57_193 ();
 FILLCELL_X32 FILLER_57_225 ();
 FILLCELL_X32 FILLER_57_257 ();
 FILLCELL_X32 FILLER_57_289 ();
 FILLCELL_X32 FILLER_57_321 ();
 FILLCELL_X32 FILLER_57_353 ();
 FILLCELL_X32 FILLER_57_385 ();
 FILLCELL_X32 FILLER_57_417 ();
 FILLCELL_X32 FILLER_57_449 ();
 FILLCELL_X32 FILLER_57_481 ();
 FILLCELL_X32 FILLER_57_513 ();
 FILLCELL_X32 FILLER_57_545 ();
 FILLCELL_X32 FILLER_57_577 ();
 FILLCELL_X32 FILLER_57_609 ();
 FILLCELL_X32 FILLER_57_641 ();
 FILLCELL_X32 FILLER_57_673 ();
 FILLCELL_X32 FILLER_57_705 ();
 FILLCELL_X32 FILLER_57_737 ();
 FILLCELL_X32 FILLER_57_769 ();
 FILLCELL_X32 FILLER_57_801 ();
 FILLCELL_X32 FILLER_57_833 ();
 FILLCELL_X32 FILLER_57_865 ();
 FILLCELL_X32 FILLER_57_897 ();
 FILLCELL_X32 FILLER_57_929 ();
 FILLCELL_X32 FILLER_57_961 ();
 FILLCELL_X32 FILLER_57_993 ();
 FILLCELL_X32 FILLER_57_1025 ();
 FILLCELL_X32 FILLER_57_1057 ();
 FILLCELL_X32 FILLER_57_1089 ();
 FILLCELL_X32 FILLER_57_1121 ();
 FILLCELL_X32 FILLER_57_1153 ();
 FILLCELL_X32 FILLER_57_1185 ();
 FILLCELL_X32 FILLER_57_1217 ();
 FILLCELL_X8 FILLER_57_1249 ();
 FILLCELL_X4 FILLER_57_1257 ();
 FILLCELL_X2 FILLER_57_1261 ();
 FILLCELL_X32 FILLER_57_1264 ();
 FILLCELL_X32 FILLER_57_1296 ();
 FILLCELL_X32 FILLER_57_1328 ();
 FILLCELL_X32 FILLER_57_1360 ();
 FILLCELL_X32 FILLER_57_1392 ();
 FILLCELL_X32 FILLER_57_1424 ();
 FILLCELL_X32 FILLER_57_1456 ();
 FILLCELL_X32 FILLER_57_1488 ();
 FILLCELL_X32 FILLER_57_1520 ();
 FILLCELL_X32 FILLER_57_1552 ();
 FILLCELL_X32 FILLER_57_1584 ();
 FILLCELL_X32 FILLER_57_1616 ();
 FILLCELL_X32 FILLER_57_1648 ();
 FILLCELL_X32 FILLER_57_1680 ();
 FILLCELL_X32 FILLER_57_1712 ();
 FILLCELL_X32 FILLER_57_1744 ();
 FILLCELL_X32 FILLER_57_1776 ();
 FILLCELL_X32 FILLER_57_1808 ();
 FILLCELL_X32 FILLER_57_1840 ();
 FILLCELL_X32 FILLER_57_1872 ();
 FILLCELL_X32 FILLER_57_1904 ();
 FILLCELL_X32 FILLER_57_1936 ();
 FILLCELL_X32 FILLER_57_1968 ();
 FILLCELL_X32 FILLER_57_2000 ();
 FILLCELL_X32 FILLER_57_2032 ();
 FILLCELL_X32 FILLER_57_2064 ();
 FILLCELL_X32 FILLER_57_2096 ();
 FILLCELL_X32 FILLER_57_2128 ();
 FILLCELL_X32 FILLER_57_2160 ();
 FILLCELL_X32 FILLER_57_2192 ();
 FILLCELL_X32 FILLER_57_2224 ();
 FILLCELL_X32 FILLER_57_2256 ();
 FILLCELL_X32 FILLER_57_2288 ();
 FILLCELL_X32 FILLER_57_2320 ();
 FILLCELL_X32 FILLER_57_2352 ();
 FILLCELL_X32 FILLER_57_2384 ();
 FILLCELL_X32 FILLER_57_2416 ();
 FILLCELL_X32 FILLER_57_2448 ();
 FILLCELL_X32 FILLER_57_2480 ();
 FILLCELL_X8 FILLER_57_2512 ();
 FILLCELL_X4 FILLER_57_2520 ();
 FILLCELL_X2 FILLER_57_2524 ();
 FILLCELL_X32 FILLER_57_2527 ();
 FILLCELL_X32 FILLER_57_2559 ();
 FILLCELL_X8 FILLER_57_2591 ();
 FILLCELL_X2 FILLER_57_2599 ();
 FILLCELL_X1 FILLER_57_2601 ();
 FILLCELL_X32 FILLER_58_1 ();
 FILLCELL_X32 FILLER_58_33 ();
 FILLCELL_X32 FILLER_58_65 ();
 FILLCELL_X32 FILLER_58_97 ();
 FILLCELL_X32 FILLER_58_129 ();
 FILLCELL_X32 FILLER_58_161 ();
 FILLCELL_X32 FILLER_58_193 ();
 FILLCELL_X32 FILLER_58_225 ();
 FILLCELL_X32 FILLER_58_257 ();
 FILLCELL_X32 FILLER_58_289 ();
 FILLCELL_X32 FILLER_58_321 ();
 FILLCELL_X32 FILLER_58_353 ();
 FILLCELL_X32 FILLER_58_385 ();
 FILLCELL_X32 FILLER_58_417 ();
 FILLCELL_X32 FILLER_58_449 ();
 FILLCELL_X32 FILLER_58_481 ();
 FILLCELL_X32 FILLER_58_513 ();
 FILLCELL_X32 FILLER_58_545 ();
 FILLCELL_X32 FILLER_58_577 ();
 FILLCELL_X16 FILLER_58_609 ();
 FILLCELL_X4 FILLER_58_625 ();
 FILLCELL_X2 FILLER_58_629 ();
 FILLCELL_X32 FILLER_58_632 ();
 FILLCELL_X32 FILLER_58_664 ();
 FILLCELL_X32 FILLER_58_696 ();
 FILLCELL_X32 FILLER_58_728 ();
 FILLCELL_X32 FILLER_58_760 ();
 FILLCELL_X32 FILLER_58_792 ();
 FILLCELL_X32 FILLER_58_824 ();
 FILLCELL_X32 FILLER_58_856 ();
 FILLCELL_X32 FILLER_58_888 ();
 FILLCELL_X32 FILLER_58_920 ();
 FILLCELL_X32 FILLER_58_952 ();
 FILLCELL_X32 FILLER_58_984 ();
 FILLCELL_X32 FILLER_58_1016 ();
 FILLCELL_X32 FILLER_58_1048 ();
 FILLCELL_X32 FILLER_58_1080 ();
 FILLCELL_X32 FILLER_58_1112 ();
 FILLCELL_X32 FILLER_58_1144 ();
 FILLCELL_X32 FILLER_58_1176 ();
 FILLCELL_X32 FILLER_58_1208 ();
 FILLCELL_X32 FILLER_58_1240 ();
 FILLCELL_X32 FILLER_58_1272 ();
 FILLCELL_X32 FILLER_58_1304 ();
 FILLCELL_X32 FILLER_58_1336 ();
 FILLCELL_X32 FILLER_58_1368 ();
 FILLCELL_X32 FILLER_58_1400 ();
 FILLCELL_X32 FILLER_58_1432 ();
 FILLCELL_X32 FILLER_58_1464 ();
 FILLCELL_X32 FILLER_58_1496 ();
 FILLCELL_X32 FILLER_58_1528 ();
 FILLCELL_X32 FILLER_58_1560 ();
 FILLCELL_X32 FILLER_58_1592 ();
 FILLCELL_X32 FILLER_58_1624 ();
 FILLCELL_X32 FILLER_58_1656 ();
 FILLCELL_X32 FILLER_58_1688 ();
 FILLCELL_X32 FILLER_58_1720 ();
 FILLCELL_X32 FILLER_58_1752 ();
 FILLCELL_X32 FILLER_58_1784 ();
 FILLCELL_X32 FILLER_58_1816 ();
 FILLCELL_X32 FILLER_58_1848 ();
 FILLCELL_X8 FILLER_58_1880 ();
 FILLCELL_X4 FILLER_58_1888 ();
 FILLCELL_X2 FILLER_58_1892 ();
 FILLCELL_X32 FILLER_58_1895 ();
 FILLCELL_X32 FILLER_58_1927 ();
 FILLCELL_X32 FILLER_58_1959 ();
 FILLCELL_X32 FILLER_58_1991 ();
 FILLCELL_X32 FILLER_58_2023 ();
 FILLCELL_X32 FILLER_58_2055 ();
 FILLCELL_X32 FILLER_58_2087 ();
 FILLCELL_X32 FILLER_58_2119 ();
 FILLCELL_X32 FILLER_58_2151 ();
 FILLCELL_X32 FILLER_58_2183 ();
 FILLCELL_X32 FILLER_58_2215 ();
 FILLCELL_X32 FILLER_58_2247 ();
 FILLCELL_X32 FILLER_58_2279 ();
 FILLCELL_X32 FILLER_58_2311 ();
 FILLCELL_X32 FILLER_58_2343 ();
 FILLCELL_X32 FILLER_58_2375 ();
 FILLCELL_X32 FILLER_58_2407 ();
 FILLCELL_X32 FILLER_58_2439 ();
 FILLCELL_X32 FILLER_58_2471 ();
 FILLCELL_X32 FILLER_58_2503 ();
 FILLCELL_X32 FILLER_58_2535 ();
 FILLCELL_X32 FILLER_58_2567 ();
 FILLCELL_X2 FILLER_58_2599 ();
 FILLCELL_X1 FILLER_58_2601 ();
 FILLCELL_X32 FILLER_59_1 ();
 FILLCELL_X32 FILLER_59_33 ();
 FILLCELL_X32 FILLER_59_65 ();
 FILLCELL_X32 FILLER_59_97 ();
 FILLCELL_X32 FILLER_59_129 ();
 FILLCELL_X32 FILLER_59_161 ();
 FILLCELL_X32 FILLER_59_193 ();
 FILLCELL_X32 FILLER_59_225 ();
 FILLCELL_X32 FILLER_59_257 ();
 FILLCELL_X32 FILLER_59_289 ();
 FILLCELL_X32 FILLER_59_321 ();
 FILLCELL_X32 FILLER_59_353 ();
 FILLCELL_X32 FILLER_59_385 ();
 FILLCELL_X32 FILLER_59_417 ();
 FILLCELL_X32 FILLER_59_449 ();
 FILLCELL_X32 FILLER_59_481 ();
 FILLCELL_X32 FILLER_59_513 ();
 FILLCELL_X32 FILLER_59_545 ();
 FILLCELL_X32 FILLER_59_577 ();
 FILLCELL_X32 FILLER_59_609 ();
 FILLCELL_X32 FILLER_59_641 ();
 FILLCELL_X32 FILLER_59_673 ();
 FILLCELL_X32 FILLER_59_705 ();
 FILLCELL_X32 FILLER_59_737 ();
 FILLCELL_X32 FILLER_59_769 ();
 FILLCELL_X32 FILLER_59_801 ();
 FILLCELL_X32 FILLER_59_833 ();
 FILLCELL_X32 FILLER_59_865 ();
 FILLCELL_X32 FILLER_59_897 ();
 FILLCELL_X32 FILLER_59_929 ();
 FILLCELL_X32 FILLER_59_961 ();
 FILLCELL_X32 FILLER_59_993 ();
 FILLCELL_X32 FILLER_59_1025 ();
 FILLCELL_X32 FILLER_59_1057 ();
 FILLCELL_X32 FILLER_59_1089 ();
 FILLCELL_X32 FILLER_59_1121 ();
 FILLCELL_X32 FILLER_59_1153 ();
 FILLCELL_X32 FILLER_59_1185 ();
 FILLCELL_X32 FILLER_59_1217 ();
 FILLCELL_X8 FILLER_59_1249 ();
 FILLCELL_X4 FILLER_59_1257 ();
 FILLCELL_X2 FILLER_59_1261 ();
 FILLCELL_X32 FILLER_59_1264 ();
 FILLCELL_X32 FILLER_59_1296 ();
 FILLCELL_X32 FILLER_59_1328 ();
 FILLCELL_X32 FILLER_59_1360 ();
 FILLCELL_X32 FILLER_59_1392 ();
 FILLCELL_X32 FILLER_59_1424 ();
 FILLCELL_X32 FILLER_59_1456 ();
 FILLCELL_X32 FILLER_59_1488 ();
 FILLCELL_X32 FILLER_59_1520 ();
 FILLCELL_X32 FILLER_59_1552 ();
 FILLCELL_X32 FILLER_59_1584 ();
 FILLCELL_X32 FILLER_59_1616 ();
 FILLCELL_X32 FILLER_59_1648 ();
 FILLCELL_X32 FILLER_59_1680 ();
 FILLCELL_X32 FILLER_59_1712 ();
 FILLCELL_X32 FILLER_59_1744 ();
 FILLCELL_X32 FILLER_59_1776 ();
 FILLCELL_X32 FILLER_59_1808 ();
 FILLCELL_X32 FILLER_59_1840 ();
 FILLCELL_X32 FILLER_59_1872 ();
 FILLCELL_X32 FILLER_59_1904 ();
 FILLCELL_X32 FILLER_59_1936 ();
 FILLCELL_X32 FILLER_59_1968 ();
 FILLCELL_X32 FILLER_59_2000 ();
 FILLCELL_X32 FILLER_59_2032 ();
 FILLCELL_X32 FILLER_59_2064 ();
 FILLCELL_X32 FILLER_59_2096 ();
 FILLCELL_X32 FILLER_59_2128 ();
 FILLCELL_X32 FILLER_59_2160 ();
 FILLCELL_X32 FILLER_59_2192 ();
 FILLCELL_X32 FILLER_59_2224 ();
 FILLCELL_X32 FILLER_59_2256 ();
 FILLCELL_X32 FILLER_59_2288 ();
 FILLCELL_X32 FILLER_59_2320 ();
 FILLCELL_X32 FILLER_59_2352 ();
 FILLCELL_X32 FILLER_59_2384 ();
 FILLCELL_X32 FILLER_59_2416 ();
 FILLCELL_X32 FILLER_59_2448 ();
 FILLCELL_X32 FILLER_59_2480 ();
 FILLCELL_X8 FILLER_59_2512 ();
 FILLCELL_X4 FILLER_59_2520 ();
 FILLCELL_X2 FILLER_59_2524 ();
 FILLCELL_X32 FILLER_59_2527 ();
 FILLCELL_X32 FILLER_59_2559 ();
 FILLCELL_X8 FILLER_59_2591 ();
 FILLCELL_X2 FILLER_59_2599 ();
 FILLCELL_X1 FILLER_59_2601 ();
 FILLCELL_X32 FILLER_60_1 ();
 FILLCELL_X32 FILLER_60_33 ();
 FILLCELL_X32 FILLER_60_65 ();
 FILLCELL_X32 FILLER_60_97 ();
 FILLCELL_X32 FILLER_60_129 ();
 FILLCELL_X32 FILLER_60_161 ();
 FILLCELL_X32 FILLER_60_193 ();
 FILLCELL_X32 FILLER_60_225 ();
 FILLCELL_X32 FILLER_60_257 ();
 FILLCELL_X32 FILLER_60_289 ();
 FILLCELL_X32 FILLER_60_321 ();
 FILLCELL_X32 FILLER_60_353 ();
 FILLCELL_X32 FILLER_60_385 ();
 FILLCELL_X32 FILLER_60_417 ();
 FILLCELL_X32 FILLER_60_449 ();
 FILLCELL_X32 FILLER_60_481 ();
 FILLCELL_X32 FILLER_60_513 ();
 FILLCELL_X32 FILLER_60_545 ();
 FILLCELL_X32 FILLER_60_577 ();
 FILLCELL_X16 FILLER_60_609 ();
 FILLCELL_X4 FILLER_60_625 ();
 FILLCELL_X2 FILLER_60_629 ();
 FILLCELL_X32 FILLER_60_632 ();
 FILLCELL_X32 FILLER_60_664 ();
 FILLCELL_X32 FILLER_60_696 ();
 FILLCELL_X32 FILLER_60_728 ();
 FILLCELL_X32 FILLER_60_760 ();
 FILLCELL_X32 FILLER_60_792 ();
 FILLCELL_X32 FILLER_60_824 ();
 FILLCELL_X32 FILLER_60_856 ();
 FILLCELL_X32 FILLER_60_888 ();
 FILLCELL_X32 FILLER_60_920 ();
 FILLCELL_X32 FILLER_60_952 ();
 FILLCELL_X32 FILLER_60_984 ();
 FILLCELL_X32 FILLER_60_1016 ();
 FILLCELL_X32 FILLER_60_1048 ();
 FILLCELL_X32 FILLER_60_1080 ();
 FILLCELL_X32 FILLER_60_1112 ();
 FILLCELL_X32 FILLER_60_1144 ();
 FILLCELL_X32 FILLER_60_1176 ();
 FILLCELL_X32 FILLER_60_1208 ();
 FILLCELL_X32 FILLER_60_1240 ();
 FILLCELL_X32 FILLER_60_1272 ();
 FILLCELL_X32 FILLER_60_1304 ();
 FILLCELL_X32 FILLER_60_1336 ();
 FILLCELL_X32 FILLER_60_1368 ();
 FILLCELL_X32 FILLER_60_1400 ();
 FILLCELL_X32 FILLER_60_1432 ();
 FILLCELL_X32 FILLER_60_1464 ();
 FILLCELL_X32 FILLER_60_1496 ();
 FILLCELL_X32 FILLER_60_1528 ();
 FILLCELL_X32 FILLER_60_1560 ();
 FILLCELL_X32 FILLER_60_1592 ();
 FILLCELL_X32 FILLER_60_1624 ();
 FILLCELL_X32 FILLER_60_1656 ();
 FILLCELL_X32 FILLER_60_1688 ();
 FILLCELL_X32 FILLER_60_1720 ();
 FILLCELL_X32 FILLER_60_1752 ();
 FILLCELL_X32 FILLER_60_1784 ();
 FILLCELL_X32 FILLER_60_1816 ();
 FILLCELL_X32 FILLER_60_1848 ();
 FILLCELL_X8 FILLER_60_1880 ();
 FILLCELL_X4 FILLER_60_1888 ();
 FILLCELL_X2 FILLER_60_1892 ();
 FILLCELL_X32 FILLER_60_1895 ();
 FILLCELL_X32 FILLER_60_1927 ();
 FILLCELL_X32 FILLER_60_1959 ();
 FILLCELL_X32 FILLER_60_1991 ();
 FILLCELL_X32 FILLER_60_2023 ();
 FILLCELL_X32 FILLER_60_2055 ();
 FILLCELL_X32 FILLER_60_2087 ();
 FILLCELL_X32 FILLER_60_2119 ();
 FILLCELL_X32 FILLER_60_2151 ();
 FILLCELL_X32 FILLER_60_2183 ();
 FILLCELL_X32 FILLER_60_2215 ();
 FILLCELL_X32 FILLER_60_2247 ();
 FILLCELL_X32 FILLER_60_2279 ();
 FILLCELL_X32 FILLER_60_2311 ();
 FILLCELL_X32 FILLER_60_2343 ();
 FILLCELL_X32 FILLER_60_2375 ();
 FILLCELL_X32 FILLER_60_2407 ();
 FILLCELL_X32 FILLER_60_2439 ();
 FILLCELL_X32 FILLER_60_2471 ();
 FILLCELL_X32 FILLER_60_2503 ();
 FILLCELL_X32 FILLER_60_2535 ();
 FILLCELL_X32 FILLER_60_2567 ();
 FILLCELL_X2 FILLER_60_2599 ();
 FILLCELL_X1 FILLER_60_2601 ();
 FILLCELL_X32 FILLER_61_1 ();
 FILLCELL_X32 FILLER_61_33 ();
 FILLCELL_X32 FILLER_61_65 ();
 FILLCELL_X32 FILLER_61_97 ();
 FILLCELL_X32 FILLER_61_129 ();
 FILLCELL_X32 FILLER_61_161 ();
 FILLCELL_X32 FILLER_61_193 ();
 FILLCELL_X32 FILLER_61_225 ();
 FILLCELL_X32 FILLER_61_257 ();
 FILLCELL_X32 FILLER_61_289 ();
 FILLCELL_X32 FILLER_61_321 ();
 FILLCELL_X32 FILLER_61_353 ();
 FILLCELL_X32 FILLER_61_385 ();
 FILLCELL_X32 FILLER_61_417 ();
 FILLCELL_X32 FILLER_61_449 ();
 FILLCELL_X32 FILLER_61_481 ();
 FILLCELL_X32 FILLER_61_513 ();
 FILLCELL_X32 FILLER_61_545 ();
 FILLCELL_X32 FILLER_61_577 ();
 FILLCELL_X32 FILLER_61_609 ();
 FILLCELL_X32 FILLER_61_641 ();
 FILLCELL_X32 FILLER_61_673 ();
 FILLCELL_X32 FILLER_61_705 ();
 FILLCELL_X32 FILLER_61_737 ();
 FILLCELL_X32 FILLER_61_769 ();
 FILLCELL_X32 FILLER_61_801 ();
 FILLCELL_X32 FILLER_61_833 ();
 FILLCELL_X32 FILLER_61_865 ();
 FILLCELL_X32 FILLER_61_897 ();
 FILLCELL_X32 FILLER_61_929 ();
 FILLCELL_X32 FILLER_61_961 ();
 FILLCELL_X32 FILLER_61_993 ();
 FILLCELL_X32 FILLER_61_1025 ();
 FILLCELL_X32 FILLER_61_1057 ();
 FILLCELL_X32 FILLER_61_1089 ();
 FILLCELL_X32 FILLER_61_1121 ();
 FILLCELL_X32 FILLER_61_1153 ();
 FILLCELL_X32 FILLER_61_1185 ();
 FILLCELL_X32 FILLER_61_1217 ();
 FILLCELL_X8 FILLER_61_1249 ();
 FILLCELL_X4 FILLER_61_1257 ();
 FILLCELL_X2 FILLER_61_1261 ();
 FILLCELL_X32 FILLER_61_1264 ();
 FILLCELL_X32 FILLER_61_1296 ();
 FILLCELL_X32 FILLER_61_1328 ();
 FILLCELL_X32 FILLER_61_1360 ();
 FILLCELL_X32 FILLER_61_1392 ();
 FILLCELL_X32 FILLER_61_1424 ();
 FILLCELL_X32 FILLER_61_1456 ();
 FILLCELL_X32 FILLER_61_1488 ();
 FILLCELL_X32 FILLER_61_1520 ();
 FILLCELL_X32 FILLER_61_1552 ();
 FILLCELL_X32 FILLER_61_1584 ();
 FILLCELL_X32 FILLER_61_1616 ();
 FILLCELL_X32 FILLER_61_1648 ();
 FILLCELL_X32 FILLER_61_1680 ();
 FILLCELL_X32 FILLER_61_1712 ();
 FILLCELL_X32 FILLER_61_1744 ();
 FILLCELL_X32 FILLER_61_1776 ();
 FILLCELL_X32 FILLER_61_1808 ();
 FILLCELL_X32 FILLER_61_1840 ();
 FILLCELL_X32 FILLER_61_1872 ();
 FILLCELL_X32 FILLER_61_1904 ();
 FILLCELL_X32 FILLER_61_1936 ();
 FILLCELL_X32 FILLER_61_1968 ();
 FILLCELL_X32 FILLER_61_2000 ();
 FILLCELL_X32 FILLER_61_2032 ();
 FILLCELL_X32 FILLER_61_2064 ();
 FILLCELL_X32 FILLER_61_2096 ();
 FILLCELL_X32 FILLER_61_2128 ();
 FILLCELL_X32 FILLER_61_2160 ();
 FILLCELL_X32 FILLER_61_2192 ();
 FILLCELL_X32 FILLER_61_2224 ();
 FILLCELL_X32 FILLER_61_2256 ();
 FILLCELL_X32 FILLER_61_2288 ();
 FILLCELL_X32 FILLER_61_2320 ();
 FILLCELL_X32 FILLER_61_2352 ();
 FILLCELL_X32 FILLER_61_2384 ();
 FILLCELL_X32 FILLER_61_2416 ();
 FILLCELL_X32 FILLER_61_2448 ();
 FILLCELL_X32 FILLER_61_2480 ();
 FILLCELL_X8 FILLER_61_2512 ();
 FILLCELL_X4 FILLER_61_2520 ();
 FILLCELL_X2 FILLER_61_2524 ();
 FILLCELL_X32 FILLER_61_2527 ();
 FILLCELL_X32 FILLER_61_2559 ();
 FILLCELL_X8 FILLER_61_2591 ();
 FILLCELL_X2 FILLER_61_2599 ();
 FILLCELL_X1 FILLER_61_2601 ();
 FILLCELL_X32 FILLER_62_1 ();
 FILLCELL_X32 FILLER_62_33 ();
 FILLCELL_X32 FILLER_62_65 ();
 FILLCELL_X32 FILLER_62_97 ();
 FILLCELL_X32 FILLER_62_129 ();
 FILLCELL_X32 FILLER_62_161 ();
 FILLCELL_X32 FILLER_62_193 ();
 FILLCELL_X32 FILLER_62_225 ();
 FILLCELL_X32 FILLER_62_257 ();
 FILLCELL_X32 FILLER_62_289 ();
 FILLCELL_X32 FILLER_62_321 ();
 FILLCELL_X32 FILLER_62_353 ();
 FILLCELL_X32 FILLER_62_385 ();
 FILLCELL_X32 FILLER_62_417 ();
 FILLCELL_X32 FILLER_62_449 ();
 FILLCELL_X32 FILLER_62_481 ();
 FILLCELL_X32 FILLER_62_513 ();
 FILLCELL_X32 FILLER_62_545 ();
 FILLCELL_X32 FILLER_62_577 ();
 FILLCELL_X16 FILLER_62_609 ();
 FILLCELL_X4 FILLER_62_625 ();
 FILLCELL_X2 FILLER_62_629 ();
 FILLCELL_X32 FILLER_62_632 ();
 FILLCELL_X32 FILLER_62_664 ();
 FILLCELL_X32 FILLER_62_696 ();
 FILLCELL_X32 FILLER_62_728 ();
 FILLCELL_X32 FILLER_62_760 ();
 FILLCELL_X32 FILLER_62_792 ();
 FILLCELL_X32 FILLER_62_824 ();
 FILLCELL_X32 FILLER_62_856 ();
 FILLCELL_X32 FILLER_62_888 ();
 FILLCELL_X32 FILLER_62_920 ();
 FILLCELL_X32 FILLER_62_952 ();
 FILLCELL_X32 FILLER_62_984 ();
 FILLCELL_X32 FILLER_62_1016 ();
 FILLCELL_X32 FILLER_62_1048 ();
 FILLCELL_X32 FILLER_62_1080 ();
 FILLCELL_X32 FILLER_62_1112 ();
 FILLCELL_X32 FILLER_62_1144 ();
 FILLCELL_X32 FILLER_62_1176 ();
 FILLCELL_X32 FILLER_62_1208 ();
 FILLCELL_X32 FILLER_62_1240 ();
 FILLCELL_X32 FILLER_62_1272 ();
 FILLCELL_X32 FILLER_62_1304 ();
 FILLCELL_X32 FILLER_62_1336 ();
 FILLCELL_X32 FILLER_62_1368 ();
 FILLCELL_X32 FILLER_62_1400 ();
 FILLCELL_X32 FILLER_62_1432 ();
 FILLCELL_X32 FILLER_62_1464 ();
 FILLCELL_X32 FILLER_62_1496 ();
 FILLCELL_X32 FILLER_62_1528 ();
 FILLCELL_X32 FILLER_62_1560 ();
 FILLCELL_X32 FILLER_62_1592 ();
 FILLCELL_X32 FILLER_62_1624 ();
 FILLCELL_X32 FILLER_62_1656 ();
 FILLCELL_X32 FILLER_62_1688 ();
 FILLCELL_X32 FILLER_62_1720 ();
 FILLCELL_X32 FILLER_62_1752 ();
 FILLCELL_X32 FILLER_62_1784 ();
 FILLCELL_X32 FILLER_62_1816 ();
 FILLCELL_X32 FILLER_62_1848 ();
 FILLCELL_X8 FILLER_62_1880 ();
 FILLCELL_X4 FILLER_62_1888 ();
 FILLCELL_X2 FILLER_62_1892 ();
 FILLCELL_X32 FILLER_62_1895 ();
 FILLCELL_X32 FILLER_62_1927 ();
 FILLCELL_X32 FILLER_62_1959 ();
 FILLCELL_X32 FILLER_62_1991 ();
 FILLCELL_X32 FILLER_62_2023 ();
 FILLCELL_X32 FILLER_62_2055 ();
 FILLCELL_X32 FILLER_62_2087 ();
 FILLCELL_X32 FILLER_62_2119 ();
 FILLCELL_X32 FILLER_62_2151 ();
 FILLCELL_X32 FILLER_62_2183 ();
 FILLCELL_X32 FILLER_62_2215 ();
 FILLCELL_X32 FILLER_62_2247 ();
 FILLCELL_X32 FILLER_62_2279 ();
 FILLCELL_X32 FILLER_62_2311 ();
 FILLCELL_X32 FILLER_62_2343 ();
 FILLCELL_X32 FILLER_62_2375 ();
 FILLCELL_X32 FILLER_62_2407 ();
 FILLCELL_X32 FILLER_62_2439 ();
 FILLCELL_X32 FILLER_62_2471 ();
 FILLCELL_X32 FILLER_62_2503 ();
 FILLCELL_X32 FILLER_62_2535 ();
 FILLCELL_X32 FILLER_62_2567 ();
 FILLCELL_X2 FILLER_62_2599 ();
 FILLCELL_X1 FILLER_62_2601 ();
 FILLCELL_X32 FILLER_63_1 ();
 FILLCELL_X32 FILLER_63_33 ();
 FILLCELL_X32 FILLER_63_65 ();
 FILLCELL_X32 FILLER_63_97 ();
 FILLCELL_X32 FILLER_63_129 ();
 FILLCELL_X32 FILLER_63_161 ();
 FILLCELL_X32 FILLER_63_193 ();
 FILLCELL_X32 FILLER_63_225 ();
 FILLCELL_X32 FILLER_63_257 ();
 FILLCELL_X32 FILLER_63_289 ();
 FILLCELL_X32 FILLER_63_321 ();
 FILLCELL_X32 FILLER_63_353 ();
 FILLCELL_X32 FILLER_63_385 ();
 FILLCELL_X32 FILLER_63_417 ();
 FILLCELL_X32 FILLER_63_449 ();
 FILLCELL_X32 FILLER_63_481 ();
 FILLCELL_X32 FILLER_63_513 ();
 FILLCELL_X32 FILLER_63_545 ();
 FILLCELL_X32 FILLER_63_577 ();
 FILLCELL_X32 FILLER_63_609 ();
 FILLCELL_X32 FILLER_63_641 ();
 FILLCELL_X32 FILLER_63_673 ();
 FILLCELL_X32 FILLER_63_705 ();
 FILLCELL_X32 FILLER_63_737 ();
 FILLCELL_X32 FILLER_63_769 ();
 FILLCELL_X32 FILLER_63_801 ();
 FILLCELL_X32 FILLER_63_833 ();
 FILLCELL_X32 FILLER_63_865 ();
 FILLCELL_X32 FILLER_63_897 ();
 FILLCELL_X32 FILLER_63_929 ();
 FILLCELL_X32 FILLER_63_961 ();
 FILLCELL_X32 FILLER_63_993 ();
 FILLCELL_X32 FILLER_63_1025 ();
 FILLCELL_X32 FILLER_63_1057 ();
 FILLCELL_X32 FILLER_63_1089 ();
 FILLCELL_X32 FILLER_63_1121 ();
 FILLCELL_X32 FILLER_63_1153 ();
 FILLCELL_X32 FILLER_63_1185 ();
 FILLCELL_X32 FILLER_63_1217 ();
 FILLCELL_X8 FILLER_63_1249 ();
 FILLCELL_X4 FILLER_63_1257 ();
 FILLCELL_X2 FILLER_63_1261 ();
 FILLCELL_X32 FILLER_63_1264 ();
 FILLCELL_X32 FILLER_63_1296 ();
 FILLCELL_X32 FILLER_63_1328 ();
 FILLCELL_X32 FILLER_63_1360 ();
 FILLCELL_X32 FILLER_63_1392 ();
 FILLCELL_X32 FILLER_63_1424 ();
 FILLCELL_X32 FILLER_63_1456 ();
 FILLCELL_X32 FILLER_63_1488 ();
 FILLCELL_X32 FILLER_63_1520 ();
 FILLCELL_X32 FILLER_63_1552 ();
 FILLCELL_X32 FILLER_63_1584 ();
 FILLCELL_X32 FILLER_63_1616 ();
 FILLCELL_X32 FILLER_63_1648 ();
 FILLCELL_X32 FILLER_63_1680 ();
 FILLCELL_X32 FILLER_63_1712 ();
 FILLCELL_X32 FILLER_63_1744 ();
 FILLCELL_X32 FILLER_63_1776 ();
 FILLCELL_X32 FILLER_63_1808 ();
 FILLCELL_X32 FILLER_63_1840 ();
 FILLCELL_X32 FILLER_63_1872 ();
 FILLCELL_X32 FILLER_63_1904 ();
 FILLCELL_X32 FILLER_63_1936 ();
 FILLCELL_X32 FILLER_63_1968 ();
 FILLCELL_X32 FILLER_63_2000 ();
 FILLCELL_X32 FILLER_63_2032 ();
 FILLCELL_X32 FILLER_63_2064 ();
 FILLCELL_X32 FILLER_63_2096 ();
 FILLCELL_X32 FILLER_63_2128 ();
 FILLCELL_X32 FILLER_63_2160 ();
 FILLCELL_X32 FILLER_63_2192 ();
 FILLCELL_X32 FILLER_63_2224 ();
 FILLCELL_X32 FILLER_63_2256 ();
 FILLCELL_X32 FILLER_63_2288 ();
 FILLCELL_X32 FILLER_63_2320 ();
 FILLCELL_X32 FILLER_63_2352 ();
 FILLCELL_X32 FILLER_63_2384 ();
 FILLCELL_X32 FILLER_63_2416 ();
 FILLCELL_X32 FILLER_63_2448 ();
 FILLCELL_X32 FILLER_63_2480 ();
 FILLCELL_X8 FILLER_63_2512 ();
 FILLCELL_X4 FILLER_63_2520 ();
 FILLCELL_X2 FILLER_63_2524 ();
 FILLCELL_X32 FILLER_63_2527 ();
 FILLCELL_X32 FILLER_63_2559 ();
 FILLCELL_X8 FILLER_63_2591 ();
 FILLCELL_X2 FILLER_63_2599 ();
 FILLCELL_X1 FILLER_63_2601 ();
 FILLCELL_X32 FILLER_64_1 ();
 FILLCELL_X32 FILLER_64_33 ();
 FILLCELL_X32 FILLER_64_65 ();
 FILLCELL_X32 FILLER_64_97 ();
 FILLCELL_X32 FILLER_64_129 ();
 FILLCELL_X32 FILLER_64_161 ();
 FILLCELL_X32 FILLER_64_193 ();
 FILLCELL_X32 FILLER_64_225 ();
 FILLCELL_X32 FILLER_64_257 ();
 FILLCELL_X32 FILLER_64_289 ();
 FILLCELL_X32 FILLER_64_321 ();
 FILLCELL_X32 FILLER_64_353 ();
 FILLCELL_X32 FILLER_64_385 ();
 FILLCELL_X32 FILLER_64_417 ();
 FILLCELL_X32 FILLER_64_449 ();
 FILLCELL_X32 FILLER_64_481 ();
 FILLCELL_X32 FILLER_64_513 ();
 FILLCELL_X32 FILLER_64_545 ();
 FILLCELL_X32 FILLER_64_577 ();
 FILLCELL_X16 FILLER_64_609 ();
 FILLCELL_X4 FILLER_64_625 ();
 FILLCELL_X2 FILLER_64_629 ();
 FILLCELL_X32 FILLER_64_632 ();
 FILLCELL_X32 FILLER_64_664 ();
 FILLCELL_X32 FILLER_64_696 ();
 FILLCELL_X32 FILLER_64_728 ();
 FILLCELL_X32 FILLER_64_760 ();
 FILLCELL_X32 FILLER_64_792 ();
 FILLCELL_X32 FILLER_64_824 ();
 FILLCELL_X32 FILLER_64_856 ();
 FILLCELL_X32 FILLER_64_888 ();
 FILLCELL_X32 FILLER_64_920 ();
 FILLCELL_X32 FILLER_64_952 ();
 FILLCELL_X32 FILLER_64_984 ();
 FILLCELL_X32 FILLER_64_1016 ();
 FILLCELL_X32 FILLER_64_1048 ();
 FILLCELL_X32 FILLER_64_1080 ();
 FILLCELL_X32 FILLER_64_1112 ();
 FILLCELL_X32 FILLER_64_1144 ();
 FILLCELL_X32 FILLER_64_1176 ();
 FILLCELL_X32 FILLER_64_1208 ();
 FILLCELL_X32 FILLER_64_1240 ();
 FILLCELL_X32 FILLER_64_1272 ();
 FILLCELL_X32 FILLER_64_1304 ();
 FILLCELL_X32 FILLER_64_1336 ();
 FILLCELL_X32 FILLER_64_1368 ();
 FILLCELL_X32 FILLER_64_1400 ();
 FILLCELL_X32 FILLER_64_1432 ();
 FILLCELL_X32 FILLER_64_1464 ();
 FILLCELL_X32 FILLER_64_1496 ();
 FILLCELL_X32 FILLER_64_1528 ();
 FILLCELL_X32 FILLER_64_1560 ();
 FILLCELL_X32 FILLER_64_1592 ();
 FILLCELL_X32 FILLER_64_1624 ();
 FILLCELL_X32 FILLER_64_1656 ();
 FILLCELL_X32 FILLER_64_1688 ();
 FILLCELL_X32 FILLER_64_1720 ();
 FILLCELL_X32 FILLER_64_1752 ();
 FILLCELL_X32 FILLER_64_1784 ();
 FILLCELL_X32 FILLER_64_1816 ();
 FILLCELL_X32 FILLER_64_1848 ();
 FILLCELL_X8 FILLER_64_1880 ();
 FILLCELL_X4 FILLER_64_1888 ();
 FILLCELL_X2 FILLER_64_1892 ();
 FILLCELL_X32 FILLER_64_1895 ();
 FILLCELL_X32 FILLER_64_1927 ();
 FILLCELL_X32 FILLER_64_1959 ();
 FILLCELL_X32 FILLER_64_1991 ();
 FILLCELL_X32 FILLER_64_2023 ();
 FILLCELL_X32 FILLER_64_2055 ();
 FILLCELL_X32 FILLER_64_2087 ();
 FILLCELL_X32 FILLER_64_2119 ();
 FILLCELL_X32 FILLER_64_2151 ();
 FILLCELL_X32 FILLER_64_2183 ();
 FILLCELL_X32 FILLER_64_2215 ();
 FILLCELL_X32 FILLER_64_2247 ();
 FILLCELL_X32 FILLER_64_2279 ();
 FILLCELL_X32 FILLER_64_2311 ();
 FILLCELL_X32 FILLER_64_2343 ();
 FILLCELL_X32 FILLER_64_2375 ();
 FILLCELL_X32 FILLER_64_2407 ();
 FILLCELL_X32 FILLER_64_2439 ();
 FILLCELL_X32 FILLER_64_2471 ();
 FILLCELL_X32 FILLER_64_2503 ();
 FILLCELL_X32 FILLER_64_2535 ();
 FILLCELL_X32 FILLER_64_2567 ();
 FILLCELL_X2 FILLER_64_2599 ();
 FILLCELL_X1 FILLER_64_2601 ();
 FILLCELL_X32 FILLER_65_1 ();
 FILLCELL_X32 FILLER_65_33 ();
 FILLCELL_X32 FILLER_65_65 ();
 FILLCELL_X32 FILLER_65_97 ();
 FILLCELL_X32 FILLER_65_129 ();
 FILLCELL_X32 FILLER_65_161 ();
 FILLCELL_X32 FILLER_65_193 ();
 FILLCELL_X32 FILLER_65_225 ();
 FILLCELL_X32 FILLER_65_257 ();
 FILLCELL_X32 FILLER_65_289 ();
 FILLCELL_X32 FILLER_65_321 ();
 FILLCELL_X32 FILLER_65_353 ();
 FILLCELL_X32 FILLER_65_385 ();
 FILLCELL_X32 FILLER_65_417 ();
 FILLCELL_X32 FILLER_65_449 ();
 FILLCELL_X32 FILLER_65_481 ();
 FILLCELL_X32 FILLER_65_513 ();
 FILLCELL_X32 FILLER_65_545 ();
 FILLCELL_X32 FILLER_65_577 ();
 FILLCELL_X32 FILLER_65_609 ();
 FILLCELL_X32 FILLER_65_641 ();
 FILLCELL_X32 FILLER_65_673 ();
 FILLCELL_X32 FILLER_65_705 ();
 FILLCELL_X32 FILLER_65_737 ();
 FILLCELL_X32 FILLER_65_769 ();
 FILLCELL_X32 FILLER_65_801 ();
 FILLCELL_X32 FILLER_65_833 ();
 FILLCELL_X32 FILLER_65_865 ();
 FILLCELL_X32 FILLER_65_897 ();
 FILLCELL_X32 FILLER_65_929 ();
 FILLCELL_X32 FILLER_65_961 ();
 FILLCELL_X32 FILLER_65_993 ();
 FILLCELL_X32 FILLER_65_1025 ();
 FILLCELL_X32 FILLER_65_1057 ();
 FILLCELL_X32 FILLER_65_1089 ();
 FILLCELL_X32 FILLER_65_1121 ();
 FILLCELL_X32 FILLER_65_1153 ();
 FILLCELL_X32 FILLER_65_1185 ();
 FILLCELL_X32 FILLER_65_1217 ();
 FILLCELL_X8 FILLER_65_1249 ();
 FILLCELL_X4 FILLER_65_1257 ();
 FILLCELL_X2 FILLER_65_1261 ();
 FILLCELL_X32 FILLER_65_1264 ();
 FILLCELL_X32 FILLER_65_1296 ();
 FILLCELL_X32 FILLER_65_1328 ();
 FILLCELL_X32 FILLER_65_1360 ();
 FILLCELL_X32 FILLER_65_1392 ();
 FILLCELL_X32 FILLER_65_1424 ();
 FILLCELL_X32 FILLER_65_1456 ();
 FILLCELL_X32 FILLER_65_1488 ();
 FILLCELL_X32 FILLER_65_1520 ();
 FILLCELL_X32 FILLER_65_1552 ();
 FILLCELL_X32 FILLER_65_1584 ();
 FILLCELL_X32 FILLER_65_1616 ();
 FILLCELL_X32 FILLER_65_1648 ();
 FILLCELL_X32 FILLER_65_1680 ();
 FILLCELL_X32 FILLER_65_1712 ();
 FILLCELL_X32 FILLER_65_1744 ();
 FILLCELL_X32 FILLER_65_1776 ();
 FILLCELL_X32 FILLER_65_1808 ();
 FILLCELL_X32 FILLER_65_1840 ();
 FILLCELL_X32 FILLER_65_1872 ();
 FILLCELL_X32 FILLER_65_1904 ();
 FILLCELL_X32 FILLER_65_1936 ();
 FILLCELL_X32 FILLER_65_1968 ();
 FILLCELL_X32 FILLER_65_2000 ();
 FILLCELL_X32 FILLER_65_2032 ();
 FILLCELL_X32 FILLER_65_2064 ();
 FILLCELL_X32 FILLER_65_2096 ();
 FILLCELL_X32 FILLER_65_2128 ();
 FILLCELL_X32 FILLER_65_2160 ();
 FILLCELL_X32 FILLER_65_2192 ();
 FILLCELL_X32 FILLER_65_2224 ();
 FILLCELL_X32 FILLER_65_2256 ();
 FILLCELL_X32 FILLER_65_2288 ();
 FILLCELL_X32 FILLER_65_2320 ();
 FILLCELL_X32 FILLER_65_2352 ();
 FILLCELL_X32 FILLER_65_2384 ();
 FILLCELL_X32 FILLER_65_2416 ();
 FILLCELL_X32 FILLER_65_2448 ();
 FILLCELL_X32 FILLER_65_2480 ();
 FILLCELL_X8 FILLER_65_2512 ();
 FILLCELL_X4 FILLER_65_2520 ();
 FILLCELL_X2 FILLER_65_2524 ();
 FILLCELL_X32 FILLER_65_2527 ();
 FILLCELL_X32 FILLER_65_2559 ();
 FILLCELL_X8 FILLER_65_2591 ();
 FILLCELL_X2 FILLER_65_2599 ();
 FILLCELL_X1 FILLER_65_2601 ();
 FILLCELL_X32 FILLER_66_1 ();
 FILLCELL_X32 FILLER_66_33 ();
 FILLCELL_X32 FILLER_66_65 ();
 FILLCELL_X32 FILLER_66_97 ();
 FILLCELL_X32 FILLER_66_129 ();
 FILLCELL_X32 FILLER_66_161 ();
 FILLCELL_X32 FILLER_66_193 ();
 FILLCELL_X32 FILLER_66_225 ();
 FILLCELL_X32 FILLER_66_257 ();
 FILLCELL_X32 FILLER_66_289 ();
 FILLCELL_X32 FILLER_66_321 ();
 FILLCELL_X32 FILLER_66_353 ();
 FILLCELL_X32 FILLER_66_385 ();
 FILLCELL_X32 FILLER_66_417 ();
 FILLCELL_X32 FILLER_66_449 ();
 FILLCELL_X32 FILLER_66_481 ();
 FILLCELL_X32 FILLER_66_513 ();
 FILLCELL_X32 FILLER_66_545 ();
 FILLCELL_X32 FILLER_66_577 ();
 FILLCELL_X16 FILLER_66_609 ();
 FILLCELL_X4 FILLER_66_625 ();
 FILLCELL_X2 FILLER_66_629 ();
 FILLCELL_X32 FILLER_66_632 ();
 FILLCELL_X32 FILLER_66_664 ();
 FILLCELL_X32 FILLER_66_696 ();
 FILLCELL_X32 FILLER_66_728 ();
 FILLCELL_X32 FILLER_66_760 ();
 FILLCELL_X32 FILLER_66_792 ();
 FILLCELL_X32 FILLER_66_824 ();
 FILLCELL_X32 FILLER_66_856 ();
 FILLCELL_X32 FILLER_66_888 ();
 FILLCELL_X32 FILLER_66_920 ();
 FILLCELL_X32 FILLER_66_952 ();
 FILLCELL_X32 FILLER_66_984 ();
 FILLCELL_X32 FILLER_66_1016 ();
 FILLCELL_X32 FILLER_66_1048 ();
 FILLCELL_X32 FILLER_66_1080 ();
 FILLCELL_X32 FILLER_66_1112 ();
 FILLCELL_X32 FILLER_66_1144 ();
 FILLCELL_X32 FILLER_66_1176 ();
 FILLCELL_X32 FILLER_66_1208 ();
 FILLCELL_X32 FILLER_66_1240 ();
 FILLCELL_X32 FILLER_66_1272 ();
 FILLCELL_X32 FILLER_66_1304 ();
 FILLCELL_X32 FILLER_66_1336 ();
 FILLCELL_X32 FILLER_66_1368 ();
 FILLCELL_X32 FILLER_66_1400 ();
 FILLCELL_X32 FILLER_66_1432 ();
 FILLCELL_X32 FILLER_66_1464 ();
 FILLCELL_X32 FILLER_66_1496 ();
 FILLCELL_X32 FILLER_66_1528 ();
 FILLCELL_X32 FILLER_66_1560 ();
 FILLCELL_X32 FILLER_66_1592 ();
 FILLCELL_X32 FILLER_66_1624 ();
 FILLCELL_X32 FILLER_66_1656 ();
 FILLCELL_X32 FILLER_66_1688 ();
 FILLCELL_X32 FILLER_66_1720 ();
 FILLCELL_X32 FILLER_66_1752 ();
 FILLCELL_X32 FILLER_66_1784 ();
 FILLCELL_X32 FILLER_66_1816 ();
 FILLCELL_X32 FILLER_66_1848 ();
 FILLCELL_X8 FILLER_66_1880 ();
 FILLCELL_X4 FILLER_66_1888 ();
 FILLCELL_X2 FILLER_66_1892 ();
 FILLCELL_X32 FILLER_66_1895 ();
 FILLCELL_X32 FILLER_66_1927 ();
 FILLCELL_X32 FILLER_66_1959 ();
 FILLCELL_X32 FILLER_66_1991 ();
 FILLCELL_X32 FILLER_66_2023 ();
 FILLCELL_X32 FILLER_66_2055 ();
 FILLCELL_X32 FILLER_66_2087 ();
 FILLCELL_X32 FILLER_66_2119 ();
 FILLCELL_X32 FILLER_66_2151 ();
 FILLCELL_X32 FILLER_66_2183 ();
 FILLCELL_X32 FILLER_66_2215 ();
 FILLCELL_X32 FILLER_66_2247 ();
 FILLCELL_X32 FILLER_66_2279 ();
 FILLCELL_X32 FILLER_66_2311 ();
 FILLCELL_X32 FILLER_66_2343 ();
 FILLCELL_X32 FILLER_66_2375 ();
 FILLCELL_X32 FILLER_66_2407 ();
 FILLCELL_X32 FILLER_66_2439 ();
 FILLCELL_X32 FILLER_66_2471 ();
 FILLCELL_X32 FILLER_66_2503 ();
 FILLCELL_X32 FILLER_66_2535 ();
 FILLCELL_X32 FILLER_66_2567 ();
 FILLCELL_X2 FILLER_66_2599 ();
 FILLCELL_X1 FILLER_66_2601 ();
 FILLCELL_X32 FILLER_67_1 ();
 FILLCELL_X32 FILLER_67_33 ();
 FILLCELL_X32 FILLER_67_65 ();
 FILLCELL_X32 FILLER_67_97 ();
 FILLCELL_X32 FILLER_67_129 ();
 FILLCELL_X32 FILLER_67_161 ();
 FILLCELL_X32 FILLER_67_193 ();
 FILLCELL_X32 FILLER_67_225 ();
 FILLCELL_X32 FILLER_67_257 ();
 FILLCELL_X32 FILLER_67_289 ();
 FILLCELL_X32 FILLER_67_321 ();
 FILLCELL_X32 FILLER_67_353 ();
 FILLCELL_X32 FILLER_67_385 ();
 FILLCELL_X32 FILLER_67_417 ();
 FILLCELL_X32 FILLER_67_449 ();
 FILLCELL_X32 FILLER_67_481 ();
 FILLCELL_X32 FILLER_67_513 ();
 FILLCELL_X32 FILLER_67_545 ();
 FILLCELL_X32 FILLER_67_577 ();
 FILLCELL_X32 FILLER_67_609 ();
 FILLCELL_X32 FILLER_67_641 ();
 FILLCELL_X32 FILLER_67_673 ();
 FILLCELL_X32 FILLER_67_705 ();
 FILLCELL_X32 FILLER_67_737 ();
 FILLCELL_X32 FILLER_67_769 ();
 FILLCELL_X32 FILLER_67_801 ();
 FILLCELL_X32 FILLER_67_833 ();
 FILLCELL_X32 FILLER_67_865 ();
 FILLCELL_X32 FILLER_67_897 ();
 FILLCELL_X32 FILLER_67_929 ();
 FILLCELL_X32 FILLER_67_961 ();
 FILLCELL_X32 FILLER_67_993 ();
 FILLCELL_X32 FILLER_67_1025 ();
 FILLCELL_X32 FILLER_67_1057 ();
 FILLCELL_X32 FILLER_67_1089 ();
 FILLCELL_X32 FILLER_67_1121 ();
 FILLCELL_X32 FILLER_67_1153 ();
 FILLCELL_X32 FILLER_67_1185 ();
 FILLCELL_X32 FILLER_67_1217 ();
 FILLCELL_X8 FILLER_67_1249 ();
 FILLCELL_X4 FILLER_67_1257 ();
 FILLCELL_X2 FILLER_67_1261 ();
 FILLCELL_X32 FILLER_67_1264 ();
 FILLCELL_X32 FILLER_67_1296 ();
 FILLCELL_X32 FILLER_67_1328 ();
 FILLCELL_X32 FILLER_67_1360 ();
 FILLCELL_X32 FILLER_67_1392 ();
 FILLCELL_X32 FILLER_67_1424 ();
 FILLCELL_X32 FILLER_67_1456 ();
 FILLCELL_X32 FILLER_67_1488 ();
 FILLCELL_X32 FILLER_67_1520 ();
 FILLCELL_X32 FILLER_67_1552 ();
 FILLCELL_X32 FILLER_67_1584 ();
 FILLCELL_X32 FILLER_67_1616 ();
 FILLCELL_X32 FILLER_67_1648 ();
 FILLCELL_X32 FILLER_67_1680 ();
 FILLCELL_X32 FILLER_67_1712 ();
 FILLCELL_X32 FILLER_67_1744 ();
 FILLCELL_X32 FILLER_67_1776 ();
 FILLCELL_X32 FILLER_67_1808 ();
 FILLCELL_X32 FILLER_67_1840 ();
 FILLCELL_X32 FILLER_67_1872 ();
 FILLCELL_X32 FILLER_67_1904 ();
 FILLCELL_X32 FILLER_67_1936 ();
 FILLCELL_X32 FILLER_67_1968 ();
 FILLCELL_X32 FILLER_67_2000 ();
 FILLCELL_X32 FILLER_67_2032 ();
 FILLCELL_X32 FILLER_67_2064 ();
 FILLCELL_X32 FILLER_67_2096 ();
 FILLCELL_X32 FILLER_67_2128 ();
 FILLCELL_X32 FILLER_67_2160 ();
 FILLCELL_X32 FILLER_67_2192 ();
 FILLCELL_X32 FILLER_67_2224 ();
 FILLCELL_X32 FILLER_67_2256 ();
 FILLCELL_X32 FILLER_67_2288 ();
 FILLCELL_X32 FILLER_67_2320 ();
 FILLCELL_X32 FILLER_67_2352 ();
 FILLCELL_X32 FILLER_67_2384 ();
 FILLCELL_X32 FILLER_67_2416 ();
 FILLCELL_X32 FILLER_67_2448 ();
 FILLCELL_X32 FILLER_67_2480 ();
 FILLCELL_X8 FILLER_67_2512 ();
 FILLCELL_X4 FILLER_67_2520 ();
 FILLCELL_X2 FILLER_67_2524 ();
 FILLCELL_X32 FILLER_67_2527 ();
 FILLCELL_X32 FILLER_67_2559 ();
 FILLCELL_X8 FILLER_67_2591 ();
 FILLCELL_X2 FILLER_67_2599 ();
 FILLCELL_X1 FILLER_67_2601 ();
 FILLCELL_X32 FILLER_68_1 ();
 FILLCELL_X32 FILLER_68_33 ();
 FILLCELL_X32 FILLER_68_65 ();
 FILLCELL_X32 FILLER_68_97 ();
 FILLCELL_X32 FILLER_68_129 ();
 FILLCELL_X32 FILLER_68_161 ();
 FILLCELL_X32 FILLER_68_193 ();
 FILLCELL_X32 FILLER_68_225 ();
 FILLCELL_X32 FILLER_68_257 ();
 FILLCELL_X32 FILLER_68_289 ();
 FILLCELL_X32 FILLER_68_321 ();
 FILLCELL_X32 FILLER_68_353 ();
 FILLCELL_X32 FILLER_68_385 ();
 FILLCELL_X32 FILLER_68_417 ();
 FILLCELL_X32 FILLER_68_449 ();
 FILLCELL_X32 FILLER_68_481 ();
 FILLCELL_X32 FILLER_68_513 ();
 FILLCELL_X32 FILLER_68_545 ();
 FILLCELL_X32 FILLER_68_577 ();
 FILLCELL_X16 FILLER_68_609 ();
 FILLCELL_X4 FILLER_68_625 ();
 FILLCELL_X2 FILLER_68_629 ();
 FILLCELL_X32 FILLER_68_632 ();
 FILLCELL_X32 FILLER_68_664 ();
 FILLCELL_X32 FILLER_68_696 ();
 FILLCELL_X32 FILLER_68_728 ();
 FILLCELL_X32 FILLER_68_760 ();
 FILLCELL_X32 FILLER_68_792 ();
 FILLCELL_X32 FILLER_68_824 ();
 FILLCELL_X32 FILLER_68_856 ();
 FILLCELL_X32 FILLER_68_888 ();
 FILLCELL_X32 FILLER_68_920 ();
 FILLCELL_X32 FILLER_68_952 ();
 FILLCELL_X32 FILLER_68_984 ();
 FILLCELL_X32 FILLER_68_1016 ();
 FILLCELL_X32 FILLER_68_1048 ();
 FILLCELL_X32 FILLER_68_1080 ();
 FILLCELL_X32 FILLER_68_1112 ();
 FILLCELL_X32 FILLER_68_1144 ();
 FILLCELL_X32 FILLER_68_1176 ();
 FILLCELL_X32 FILLER_68_1208 ();
 FILLCELL_X32 FILLER_68_1240 ();
 FILLCELL_X32 FILLER_68_1272 ();
 FILLCELL_X32 FILLER_68_1304 ();
 FILLCELL_X32 FILLER_68_1336 ();
 FILLCELL_X32 FILLER_68_1368 ();
 FILLCELL_X32 FILLER_68_1400 ();
 FILLCELL_X32 FILLER_68_1432 ();
 FILLCELL_X32 FILLER_68_1464 ();
 FILLCELL_X32 FILLER_68_1496 ();
 FILLCELL_X32 FILLER_68_1528 ();
 FILLCELL_X32 FILLER_68_1560 ();
 FILLCELL_X32 FILLER_68_1592 ();
 FILLCELL_X32 FILLER_68_1624 ();
 FILLCELL_X32 FILLER_68_1656 ();
 FILLCELL_X32 FILLER_68_1688 ();
 FILLCELL_X32 FILLER_68_1720 ();
 FILLCELL_X32 FILLER_68_1752 ();
 FILLCELL_X32 FILLER_68_1784 ();
 FILLCELL_X32 FILLER_68_1816 ();
 FILLCELL_X32 FILLER_68_1848 ();
 FILLCELL_X8 FILLER_68_1880 ();
 FILLCELL_X4 FILLER_68_1888 ();
 FILLCELL_X2 FILLER_68_1892 ();
 FILLCELL_X32 FILLER_68_1895 ();
 FILLCELL_X32 FILLER_68_1927 ();
 FILLCELL_X32 FILLER_68_1959 ();
 FILLCELL_X32 FILLER_68_1991 ();
 FILLCELL_X32 FILLER_68_2023 ();
 FILLCELL_X32 FILLER_68_2055 ();
 FILLCELL_X32 FILLER_68_2087 ();
 FILLCELL_X32 FILLER_68_2119 ();
 FILLCELL_X32 FILLER_68_2151 ();
 FILLCELL_X32 FILLER_68_2183 ();
 FILLCELL_X32 FILLER_68_2215 ();
 FILLCELL_X32 FILLER_68_2247 ();
 FILLCELL_X32 FILLER_68_2279 ();
 FILLCELL_X32 FILLER_68_2311 ();
 FILLCELL_X32 FILLER_68_2343 ();
 FILLCELL_X32 FILLER_68_2375 ();
 FILLCELL_X32 FILLER_68_2407 ();
 FILLCELL_X32 FILLER_68_2439 ();
 FILLCELL_X32 FILLER_68_2471 ();
 FILLCELL_X32 FILLER_68_2503 ();
 FILLCELL_X32 FILLER_68_2535 ();
 FILLCELL_X32 FILLER_68_2567 ();
 FILLCELL_X2 FILLER_68_2599 ();
 FILLCELL_X1 FILLER_68_2601 ();
 FILLCELL_X32 FILLER_69_1 ();
 FILLCELL_X32 FILLER_69_33 ();
 FILLCELL_X32 FILLER_69_65 ();
 FILLCELL_X32 FILLER_69_97 ();
 FILLCELL_X32 FILLER_69_129 ();
 FILLCELL_X32 FILLER_69_161 ();
 FILLCELL_X32 FILLER_69_193 ();
 FILLCELL_X32 FILLER_69_225 ();
 FILLCELL_X32 FILLER_69_257 ();
 FILLCELL_X32 FILLER_69_289 ();
 FILLCELL_X32 FILLER_69_321 ();
 FILLCELL_X32 FILLER_69_353 ();
 FILLCELL_X32 FILLER_69_385 ();
 FILLCELL_X32 FILLER_69_417 ();
 FILLCELL_X32 FILLER_69_449 ();
 FILLCELL_X32 FILLER_69_481 ();
 FILLCELL_X32 FILLER_69_513 ();
 FILLCELL_X32 FILLER_69_545 ();
 FILLCELL_X32 FILLER_69_577 ();
 FILLCELL_X32 FILLER_69_609 ();
 FILLCELL_X32 FILLER_69_641 ();
 FILLCELL_X32 FILLER_69_673 ();
 FILLCELL_X32 FILLER_69_705 ();
 FILLCELL_X32 FILLER_69_737 ();
 FILLCELL_X32 FILLER_69_769 ();
 FILLCELL_X32 FILLER_69_801 ();
 FILLCELL_X32 FILLER_69_833 ();
 FILLCELL_X32 FILLER_69_865 ();
 FILLCELL_X32 FILLER_69_897 ();
 FILLCELL_X32 FILLER_69_929 ();
 FILLCELL_X32 FILLER_69_961 ();
 FILLCELL_X32 FILLER_69_993 ();
 FILLCELL_X32 FILLER_69_1025 ();
 FILLCELL_X32 FILLER_69_1057 ();
 FILLCELL_X32 FILLER_69_1089 ();
 FILLCELL_X32 FILLER_69_1121 ();
 FILLCELL_X32 FILLER_69_1153 ();
 FILLCELL_X32 FILLER_69_1185 ();
 FILLCELL_X32 FILLER_69_1217 ();
 FILLCELL_X8 FILLER_69_1249 ();
 FILLCELL_X4 FILLER_69_1257 ();
 FILLCELL_X2 FILLER_69_1261 ();
 FILLCELL_X32 FILLER_69_1264 ();
 FILLCELL_X32 FILLER_69_1296 ();
 FILLCELL_X32 FILLER_69_1328 ();
 FILLCELL_X32 FILLER_69_1360 ();
 FILLCELL_X32 FILLER_69_1392 ();
 FILLCELL_X32 FILLER_69_1424 ();
 FILLCELL_X32 FILLER_69_1456 ();
 FILLCELL_X32 FILLER_69_1488 ();
 FILLCELL_X32 FILLER_69_1520 ();
 FILLCELL_X32 FILLER_69_1552 ();
 FILLCELL_X32 FILLER_69_1584 ();
 FILLCELL_X32 FILLER_69_1616 ();
 FILLCELL_X32 FILLER_69_1648 ();
 FILLCELL_X32 FILLER_69_1680 ();
 FILLCELL_X32 FILLER_69_1712 ();
 FILLCELL_X32 FILLER_69_1744 ();
 FILLCELL_X32 FILLER_69_1776 ();
 FILLCELL_X32 FILLER_69_1808 ();
 FILLCELL_X32 FILLER_69_1840 ();
 FILLCELL_X32 FILLER_69_1872 ();
 FILLCELL_X32 FILLER_69_1904 ();
 FILLCELL_X32 FILLER_69_1936 ();
 FILLCELL_X32 FILLER_69_1968 ();
 FILLCELL_X32 FILLER_69_2000 ();
 FILLCELL_X32 FILLER_69_2032 ();
 FILLCELL_X32 FILLER_69_2064 ();
 FILLCELL_X32 FILLER_69_2096 ();
 FILLCELL_X32 FILLER_69_2128 ();
 FILLCELL_X32 FILLER_69_2160 ();
 FILLCELL_X32 FILLER_69_2192 ();
 FILLCELL_X32 FILLER_69_2224 ();
 FILLCELL_X32 FILLER_69_2256 ();
 FILLCELL_X32 FILLER_69_2288 ();
 FILLCELL_X32 FILLER_69_2320 ();
 FILLCELL_X32 FILLER_69_2352 ();
 FILLCELL_X32 FILLER_69_2384 ();
 FILLCELL_X32 FILLER_69_2416 ();
 FILLCELL_X32 FILLER_69_2448 ();
 FILLCELL_X32 FILLER_69_2480 ();
 FILLCELL_X8 FILLER_69_2512 ();
 FILLCELL_X4 FILLER_69_2520 ();
 FILLCELL_X2 FILLER_69_2524 ();
 FILLCELL_X32 FILLER_69_2527 ();
 FILLCELL_X32 FILLER_69_2559 ();
 FILLCELL_X8 FILLER_69_2591 ();
 FILLCELL_X2 FILLER_69_2599 ();
 FILLCELL_X1 FILLER_69_2601 ();
 FILLCELL_X32 FILLER_70_1 ();
 FILLCELL_X32 FILLER_70_33 ();
 FILLCELL_X32 FILLER_70_65 ();
 FILLCELL_X32 FILLER_70_97 ();
 FILLCELL_X32 FILLER_70_129 ();
 FILLCELL_X32 FILLER_70_161 ();
 FILLCELL_X32 FILLER_70_193 ();
 FILLCELL_X32 FILLER_70_225 ();
 FILLCELL_X32 FILLER_70_257 ();
 FILLCELL_X32 FILLER_70_289 ();
 FILLCELL_X32 FILLER_70_321 ();
 FILLCELL_X32 FILLER_70_353 ();
 FILLCELL_X32 FILLER_70_385 ();
 FILLCELL_X32 FILLER_70_417 ();
 FILLCELL_X32 FILLER_70_449 ();
 FILLCELL_X32 FILLER_70_481 ();
 FILLCELL_X32 FILLER_70_513 ();
 FILLCELL_X32 FILLER_70_545 ();
 FILLCELL_X32 FILLER_70_577 ();
 FILLCELL_X16 FILLER_70_609 ();
 FILLCELL_X4 FILLER_70_625 ();
 FILLCELL_X2 FILLER_70_629 ();
 FILLCELL_X32 FILLER_70_632 ();
 FILLCELL_X32 FILLER_70_664 ();
 FILLCELL_X32 FILLER_70_696 ();
 FILLCELL_X32 FILLER_70_728 ();
 FILLCELL_X32 FILLER_70_760 ();
 FILLCELL_X32 FILLER_70_792 ();
 FILLCELL_X32 FILLER_70_824 ();
 FILLCELL_X32 FILLER_70_856 ();
 FILLCELL_X32 FILLER_70_888 ();
 FILLCELL_X32 FILLER_70_920 ();
 FILLCELL_X32 FILLER_70_952 ();
 FILLCELL_X32 FILLER_70_984 ();
 FILLCELL_X32 FILLER_70_1016 ();
 FILLCELL_X32 FILLER_70_1048 ();
 FILLCELL_X32 FILLER_70_1080 ();
 FILLCELL_X32 FILLER_70_1112 ();
 FILLCELL_X32 FILLER_70_1144 ();
 FILLCELL_X32 FILLER_70_1176 ();
 FILLCELL_X32 FILLER_70_1208 ();
 FILLCELL_X32 FILLER_70_1240 ();
 FILLCELL_X32 FILLER_70_1272 ();
 FILLCELL_X32 FILLER_70_1304 ();
 FILLCELL_X32 FILLER_70_1336 ();
 FILLCELL_X32 FILLER_70_1368 ();
 FILLCELL_X32 FILLER_70_1400 ();
 FILLCELL_X32 FILLER_70_1432 ();
 FILLCELL_X32 FILLER_70_1464 ();
 FILLCELL_X32 FILLER_70_1496 ();
 FILLCELL_X32 FILLER_70_1528 ();
 FILLCELL_X32 FILLER_70_1560 ();
 FILLCELL_X32 FILLER_70_1592 ();
 FILLCELL_X32 FILLER_70_1624 ();
 FILLCELL_X32 FILLER_70_1656 ();
 FILLCELL_X32 FILLER_70_1688 ();
 FILLCELL_X32 FILLER_70_1720 ();
 FILLCELL_X32 FILLER_70_1752 ();
 FILLCELL_X32 FILLER_70_1784 ();
 FILLCELL_X32 FILLER_70_1816 ();
 FILLCELL_X32 FILLER_70_1848 ();
 FILLCELL_X8 FILLER_70_1880 ();
 FILLCELL_X4 FILLER_70_1888 ();
 FILLCELL_X2 FILLER_70_1892 ();
 FILLCELL_X32 FILLER_70_1895 ();
 FILLCELL_X32 FILLER_70_1927 ();
 FILLCELL_X32 FILLER_70_1959 ();
 FILLCELL_X32 FILLER_70_1991 ();
 FILLCELL_X32 FILLER_70_2023 ();
 FILLCELL_X32 FILLER_70_2055 ();
 FILLCELL_X32 FILLER_70_2087 ();
 FILLCELL_X32 FILLER_70_2119 ();
 FILLCELL_X32 FILLER_70_2151 ();
 FILLCELL_X32 FILLER_70_2183 ();
 FILLCELL_X32 FILLER_70_2215 ();
 FILLCELL_X32 FILLER_70_2247 ();
 FILLCELL_X32 FILLER_70_2279 ();
 FILLCELL_X32 FILLER_70_2311 ();
 FILLCELL_X32 FILLER_70_2343 ();
 FILLCELL_X32 FILLER_70_2375 ();
 FILLCELL_X32 FILLER_70_2407 ();
 FILLCELL_X32 FILLER_70_2439 ();
 FILLCELL_X32 FILLER_70_2471 ();
 FILLCELL_X32 FILLER_70_2503 ();
 FILLCELL_X32 FILLER_70_2535 ();
 FILLCELL_X32 FILLER_70_2567 ();
 FILLCELL_X2 FILLER_70_2599 ();
 FILLCELL_X1 FILLER_70_2601 ();
 FILLCELL_X32 FILLER_71_1 ();
 FILLCELL_X32 FILLER_71_33 ();
 FILLCELL_X32 FILLER_71_65 ();
 FILLCELL_X32 FILLER_71_97 ();
 FILLCELL_X32 FILLER_71_129 ();
 FILLCELL_X32 FILLER_71_161 ();
 FILLCELL_X32 FILLER_71_193 ();
 FILLCELL_X32 FILLER_71_225 ();
 FILLCELL_X32 FILLER_71_257 ();
 FILLCELL_X32 FILLER_71_289 ();
 FILLCELL_X32 FILLER_71_321 ();
 FILLCELL_X32 FILLER_71_353 ();
 FILLCELL_X32 FILLER_71_385 ();
 FILLCELL_X32 FILLER_71_417 ();
 FILLCELL_X32 FILLER_71_449 ();
 FILLCELL_X32 FILLER_71_481 ();
 FILLCELL_X32 FILLER_71_513 ();
 FILLCELL_X32 FILLER_71_545 ();
 FILLCELL_X32 FILLER_71_577 ();
 FILLCELL_X32 FILLER_71_609 ();
 FILLCELL_X32 FILLER_71_641 ();
 FILLCELL_X32 FILLER_71_673 ();
 FILLCELL_X32 FILLER_71_705 ();
 FILLCELL_X32 FILLER_71_737 ();
 FILLCELL_X32 FILLER_71_769 ();
 FILLCELL_X32 FILLER_71_801 ();
 FILLCELL_X32 FILLER_71_833 ();
 FILLCELL_X32 FILLER_71_865 ();
 FILLCELL_X32 FILLER_71_897 ();
 FILLCELL_X32 FILLER_71_929 ();
 FILLCELL_X32 FILLER_71_961 ();
 FILLCELL_X32 FILLER_71_993 ();
 FILLCELL_X32 FILLER_71_1025 ();
 FILLCELL_X32 FILLER_71_1057 ();
 FILLCELL_X32 FILLER_71_1089 ();
 FILLCELL_X32 FILLER_71_1121 ();
 FILLCELL_X32 FILLER_71_1153 ();
 FILLCELL_X32 FILLER_71_1185 ();
 FILLCELL_X32 FILLER_71_1217 ();
 FILLCELL_X8 FILLER_71_1249 ();
 FILLCELL_X4 FILLER_71_1257 ();
 FILLCELL_X2 FILLER_71_1261 ();
 FILLCELL_X32 FILLER_71_1264 ();
 FILLCELL_X32 FILLER_71_1296 ();
 FILLCELL_X32 FILLER_71_1328 ();
 FILLCELL_X32 FILLER_71_1360 ();
 FILLCELL_X32 FILLER_71_1392 ();
 FILLCELL_X32 FILLER_71_1424 ();
 FILLCELL_X32 FILLER_71_1456 ();
 FILLCELL_X32 FILLER_71_1488 ();
 FILLCELL_X32 FILLER_71_1520 ();
 FILLCELL_X32 FILLER_71_1552 ();
 FILLCELL_X32 FILLER_71_1584 ();
 FILLCELL_X32 FILLER_71_1616 ();
 FILLCELL_X32 FILLER_71_1648 ();
 FILLCELL_X32 FILLER_71_1680 ();
 FILLCELL_X32 FILLER_71_1712 ();
 FILLCELL_X32 FILLER_71_1744 ();
 FILLCELL_X32 FILLER_71_1776 ();
 FILLCELL_X32 FILLER_71_1808 ();
 FILLCELL_X32 FILLER_71_1840 ();
 FILLCELL_X32 FILLER_71_1872 ();
 FILLCELL_X32 FILLER_71_1904 ();
 FILLCELL_X32 FILLER_71_1936 ();
 FILLCELL_X32 FILLER_71_1968 ();
 FILLCELL_X32 FILLER_71_2000 ();
 FILLCELL_X32 FILLER_71_2032 ();
 FILLCELL_X32 FILLER_71_2064 ();
 FILLCELL_X32 FILLER_71_2096 ();
 FILLCELL_X32 FILLER_71_2128 ();
 FILLCELL_X32 FILLER_71_2160 ();
 FILLCELL_X32 FILLER_71_2192 ();
 FILLCELL_X32 FILLER_71_2224 ();
 FILLCELL_X32 FILLER_71_2256 ();
 FILLCELL_X32 FILLER_71_2288 ();
 FILLCELL_X32 FILLER_71_2320 ();
 FILLCELL_X32 FILLER_71_2352 ();
 FILLCELL_X32 FILLER_71_2384 ();
 FILLCELL_X32 FILLER_71_2416 ();
 FILLCELL_X32 FILLER_71_2448 ();
 FILLCELL_X32 FILLER_71_2480 ();
 FILLCELL_X8 FILLER_71_2512 ();
 FILLCELL_X4 FILLER_71_2520 ();
 FILLCELL_X2 FILLER_71_2524 ();
 FILLCELL_X32 FILLER_71_2527 ();
 FILLCELL_X32 FILLER_71_2559 ();
 FILLCELL_X8 FILLER_71_2591 ();
 FILLCELL_X2 FILLER_71_2599 ();
 FILLCELL_X1 FILLER_71_2601 ();
 FILLCELL_X32 FILLER_72_1 ();
 FILLCELL_X32 FILLER_72_33 ();
 FILLCELL_X32 FILLER_72_65 ();
 FILLCELL_X32 FILLER_72_97 ();
 FILLCELL_X32 FILLER_72_129 ();
 FILLCELL_X32 FILLER_72_161 ();
 FILLCELL_X32 FILLER_72_193 ();
 FILLCELL_X32 FILLER_72_225 ();
 FILLCELL_X32 FILLER_72_257 ();
 FILLCELL_X32 FILLER_72_289 ();
 FILLCELL_X32 FILLER_72_321 ();
 FILLCELL_X32 FILLER_72_353 ();
 FILLCELL_X32 FILLER_72_385 ();
 FILLCELL_X32 FILLER_72_417 ();
 FILLCELL_X32 FILLER_72_449 ();
 FILLCELL_X32 FILLER_72_481 ();
 FILLCELL_X32 FILLER_72_513 ();
 FILLCELL_X32 FILLER_72_545 ();
 FILLCELL_X32 FILLER_72_577 ();
 FILLCELL_X16 FILLER_72_609 ();
 FILLCELL_X4 FILLER_72_625 ();
 FILLCELL_X2 FILLER_72_629 ();
 FILLCELL_X32 FILLER_72_632 ();
 FILLCELL_X32 FILLER_72_664 ();
 FILLCELL_X32 FILLER_72_696 ();
 FILLCELL_X32 FILLER_72_728 ();
 FILLCELL_X32 FILLER_72_760 ();
 FILLCELL_X32 FILLER_72_792 ();
 FILLCELL_X32 FILLER_72_824 ();
 FILLCELL_X32 FILLER_72_856 ();
 FILLCELL_X32 FILLER_72_888 ();
 FILLCELL_X32 FILLER_72_920 ();
 FILLCELL_X32 FILLER_72_952 ();
 FILLCELL_X32 FILLER_72_984 ();
 FILLCELL_X32 FILLER_72_1016 ();
 FILLCELL_X32 FILLER_72_1048 ();
 FILLCELL_X32 FILLER_72_1080 ();
 FILLCELL_X32 FILLER_72_1112 ();
 FILLCELL_X32 FILLER_72_1144 ();
 FILLCELL_X32 FILLER_72_1176 ();
 FILLCELL_X32 FILLER_72_1208 ();
 FILLCELL_X32 FILLER_72_1240 ();
 FILLCELL_X32 FILLER_72_1272 ();
 FILLCELL_X32 FILLER_72_1304 ();
 FILLCELL_X32 FILLER_72_1336 ();
 FILLCELL_X32 FILLER_72_1368 ();
 FILLCELL_X32 FILLER_72_1400 ();
 FILLCELL_X32 FILLER_72_1432 ();
 FILLCELL_X32 FILLER_72_1464 ();
 FILLCELL_X32 FILLER_72_1496 ();
 FILLCELL_X32 FILLER_72_1528 ();
 FILLCELL_X32 FILLER_72_1560 ();
 FILLCELL_X32 FILLER_72_1592 ();
 FILLCELL_X32 FILLER_72_1624 ();
 FILLCELL_X32 FILLER_72_1656 ();
 FILLCELL_X32 FILLER_72_1688 ();
 FILLCELL_X32 FILLER_72_1720 ();
 FILLCELL_X32 FILLER_72_1752 ();
 FILLCELL_X32 FILLER_72_1784 ();
 FILLCELL_X32 FILLER_72_1816 ();
 FILLCELL_X32 FILLER_72_1848 ();
 FILLCELL_X8 FILLER_72_1880 ();
 FILLCELL_X4 FILLER_72_1888 ();
 FILLCELL_X2 FILLER_72_1892 ();
 FILLCELL_X32 FILLER_72_1895 ();
 FILLCELL_X32 FILLER_72_1927 ();
 FILLCELL_X32 FILLER_72_1959 ();
 FILLCELL_X32 FILLER_72_1991 ();
 FILLCELL_X32 FILLER_72_2023 ();
 FILLCELL_X32 FILLER_72_2055 ();
 FILLCELL_X32 FILLER_72_2087 ();
 FILLCELL_X32 FILLER_72_2119 ();
 FILLCELL_X32 FILLER_72_2151 ();
 FILLCELL_X32 FILLER_72_2183 ();
 FILLCELL_X32 FILLER_72_2215 ();
 FILLCELL_X32 FILLER_72_2247 ();
 FILLCELL_X32 FILLER_72_2279 ();
 FILLCELL_X32 FILLER_72_2311 ();
 FILLCELL_X32 FILLER_72_2343 ();
 FILLCELL_X32 FILLER_72_2375 ();
 FILLCELL_X32 FILLER_72_2407 ();
 FILLCELL_X32 FILLER_72_2439 ();
 FILLCELL_X32 FILLER_72_2471 ();
 FILLCELL_X32 FILLER_72_2503 ();
 FILLCELL_X32 FILLER_72_2535 ();
 FILLCELL_X32 FILLER_72_2567 ();
 FILLCELL_X2 FILLER_72_2599 ();
 FILLCELL_X1 FILLER_72_2601 ();
 FILLCELL_X32 FILLER_73_1 ();
 FILLCELL_X32 FILLER_73_33 ();
 FILLCELL_X32 FILLER_73_65 ();
 FILLCELL_X32 FILLER_73_97 ();
 FILLCELL_X32 FILLER_73_129 ();
 FILLCELL_X32 FILLER_73_161 ();
 FILLCELL_X32 FILLER_73_193 ();
 FILLCELL_X32 FILLER_73_225 ();
 FILLCELL_X32 FILLER_73_257 ();
 FILLCELL_X32 FILLER_73_289 ();
 FILLCELL_X32 FILLER_73_321 ();
 FILLCELL_X32 FILLER_73_353 ();
 FILLCELL_X32 FILLER_73_385 ();
 FILLCELL_X32 FILLER_73_417 ();
 FILLCELL_X32 FILLER_73_449 ();
 FILLCELL_X32 FILLER_73_481 ();
 FILLCELL_X32 FILLER_73_513 ();
 FILLCELL_X32 FILLER_73_545 ();
 FILLCELL_X32 FILLER_73_577 ();
 FILLCELL_X32 FILLER_73_609 ();
 FILLCELL_X32 FILLER_73_641 ();
 FILLCELL_X32 FILLER_73_673 ();
 FILLCELL_X32 FILLER_73_705 ();
 FILLCELL_X32 FILLER_73_737 ();
 FILLCELL_X32 FILLER_73_769 ();
 FILLCELL_X32 FILLER_73_801 ();
 FILLCELL_X32 FILLER_73_833 ();
 FILLCELL_X32 FILLER_73_865 ();
 FILLCELL_X32 FILLER_73_897 ();
 FILLCELL_X32 FILLER_73_929 ();
 FILLCELL_X32 FILLER_73_961 ();
 FILLCELL_X32 FILLER_73_993 ();
 FILLCELL_X32 FILLER_73_1025 ();
 FILLCELL_X32 FILLER_73_1057 ();
 FILLCELL_X32 FILLER_73_1089 ();
 FILLCELL_X32 FILLER_73_1121 ();
 FILLCELL_X32 FILLER_73_1153 ();
 FILLCELL_X32 FILLER_73_1185 ();
 FILLCELL_X32 FILLER_73_1217 ();
 FILLCELL_X8 FILLER_73_1249 ();
 FILLCELL_X4 FILLER_73_1257 ();
 FILLCELL_X2 FILLER_73_1261 ();
 FILLCELL_X32 FILLER_73_1264 ();
 FILLCELL_X32 FILLER_73_1296 ();
 FILLCELL_X32 FILLER_73_1328 ();
 FILLCELL_X32 FILLER_73_1360 ();
 FILLCELL_X32 FILLER_73_1392 ();
 FILLCELL_X32 FILLER_73_1424 ();
 FILLCELL_X32 FILLER_73_1456 ();
 FILLCELL_X32 FILLER_73_1488 ();
 FILLCELL_X32 FILLER_73_1520 ();
 FILLCELL_X32 FILLER_73_1552 ();
 FILLCELL_X32 FILLER_73_1584 ();
 FILLCELL_X32 FILLER_73_1616 ();
 FILLCELL_X32 FILLER_73_1648 ();
 FILLCELL_X32 FILLER_73_1680 ();
 FILLCELL_X32 FILLER_73_1712 ();
 FILLCELL_X32 FILLER_73_1744 ();
 FILLCELL_X32 FILLER_73_1776 ();
 FILLCELL_X32 FILLER_73_1808 ();
 FILLCELL_X32 FILLER_73_1840 ();
 FILLCELL_X32 FILLER_73_1872 ();
 FILLCELL_X32 FILLER_73_1904 ();
 FILLCELL_X32 FILLER_73_1936 ();
 FILLCELL_X32 FILLER_73_1968 ();
 FILLCELL_X32 FILLER_73_2000 ();
 FILLCELL_X32 FILLER_73_2032 ();
 FILLCELL_X32 FILLER_73_2064 ();
 FILLCELL_X32 FILLER_73_2096 ();
 FILLCELL_X32 FILLER_73_2128 ();
 FILLCELL_X32 FILLER_73_2160 ();
 FILLCELL_X32 FILLER_73_2192 ();
 FILLCELL_X32 FILLER_73_2224 ();
 FILLCELL_X32 FILLER_73_2256 ();
 FILLCELL_X32 FILLER_73_2288 ();
 FILLCELL_X32 FILLER_73_2320 ();
 FILLCELL_X32 FILLER_73_2352 ();
 FILLCELL_X32 FILLER_73_2384 ();
 FILLCELL_X32 FILLER_73_2416 ();
 FILLCELL_X32 FILLER_73_2448 ();
 FILLCELL_X32 FILLER_73_2480 ();
 FILLCELL_X8 FILLER_73_2512 ();
 FILLCELL_X4 FILLER_73_2520 ();
 FILLCELL_X2 FILLER_73_2524 ();
 FILLCELL_X32 FILLER_73_2527 ();
 FILLCELL_X32 FILLER_73_2559 ();
 FILLCELL_X8 FILLER_73_2591 ();
 FILLCELL_X2 FILLER_73_2599 ();
 FILLCELL_X1 FILLER_73_2601 ();
 FILLCELL_X32 FILLER_74_1 ();
 FILLCELL_X32 FILLER_74_33 ();
 FILLCELL_X32 FILLER_74_65 ();
 FILLCELL_X32 FILLER_74_97 ();
 FILLCELL_X32 FILLER_74_129 ();
 FILLCELL_X32 FILLER_74_161 ();
 FILLCELL_X32 FILLER_74_193 ();
 FILLCELL_X32 FILLER_74_225 ();
 FILLCELL_X32 FILLER_74_257 ();
 FILLCELL_X32 FILLER_74_289 ();
 FILLCELL_X32 FILLER_74_321 ();
 FILLCELL_X32 FILLER_74_353 ();
 FILLCELL_X32 FILLER_74_385 ();
 FILLCELL_X32 FILLER_74_417 ();
 FILLCELL_X32 FILLER_74_449 ();
 FILLCELL_X32 FILLER_74_481 ();
 FILLCELL_X32 FILLER_74_513 ();
 FILLCELL_X32 FILLER_74_545 ();
 FILLCELL_X32 FILLER_74_577 ();
 FILLCELL_X16 FILLER_74_609 ();
 FILLCELL_X4 FILLER_74_625 ();
 FILLCELL_X2 FILLER_74_629 ();
 FILLCELL_X32 FILLER_74_632 ();
 FILLCELL_X32 FILLER_74_664 ();
 FILLCELL_X32 FILLER_74_696 ();
 FILLCELL_X32 FILLER_74_728 ();
 FILLCELL_X32 FILLER_74_760 ();
 FILLCELL_X32 FILLER_74_792 ();
 FILLCELL_X32 FILLER_74_824 ();
 FILLCELL_X32 FILLER_74_856 ();
 FILLCELL_X32 FILLER_74_888 ();
 FILLCELL_X32 FILLER_74_920 ();
 FILLCELL_X32 FILLER_74_952 ();
 FILLCELL_X32 FILLER_74_984 ();
 FILLCELL_X32 FILLER_74_1016 ();
 FILLCELL_X32 FILLER_74_1048 ();
 FILLCELL_X32 FILLER_74_1080 ();
 FILLCELL_X32 FILLER_74_1112 ();
 FILLCELL_X32 FILLER_74_1144 ();
 FILLCELL_X32 FILLER_74_1176 ();
 FILLCELL_X32 FILLER_74_1208 ();
 FILLCELL_X32 FILLER_74_1240 ();
 FILLCELL_X32 FILLER_74_1272 ();
 FILLCELL_X32 FILLER_74_1304 ();
 FILLCELL_X32 FILLER_74_1336 ();
 FILLCELL_X32 FILLER_74_1368 ();
 FILLCELL_X32 FILLER_74_1400 ();
 FILLCELL_X32 FILLER_74_1432 ();
 FILLCELL_X32 FILLER_74_1464 ();
 FILLCELL_X32 FILLER_74_1496 ();
 FILLCELL_X32 FILLER_74_1528 ();
 FILLCELL_X32 FILLER_74_1560 ();
 FILLCELL_X32 FILLER_74_1592 ();
 FILLCELL_X32 FILLER_74_1624 ();
 FILLCELL_X32 FILLER_74_1656 ();
 FILLCELL_X32 FILLER_74_1688 ();
 FILLCELL_X32 FILLER_74_1720 ();
 FILLCELL_X32 FILLER_74_1752 ();
 FILLCELL_X32 FILLER_74_1784 ();
 FILLCELL_X32 FILLER_74_1816 ();
 FILLCELL_X32 FILLER_74_1848 ();
 FILLCELL_X8 FILLER_74_1880 ();
 FILLCELL_X4 FILLER_74_1888 ();
 FILLCELL_X2 FILLER_74_1892 ();
 FILLCELL_X32 FILLER_74_1895 ();
 FILLCELL_X32 FILLER_74_1927 ();
 FILLCELL_X32 FILLER_74_1959 ();
 FILLCELL_X32 FILLER_74_1991 ();
 FILLCELL_X32 FILLER_74_2023 ();
 FILLCELL_X32 FILLER_74_2055 ();
 FILLCELL_X32 FILLER_74_2087 ();
 FILLCELL_X32 FILLER_74_2119 ();
 FILLCELL_X32 FILLER_74_2151 ();
 FILLCELL_X32 FILLER_74_2183 ();
 FILLCELL_X32 FILLER_74_2215 ();
 FILLCELL_X32 FILLER_74_2247 ();
 FILLCELL_X32 FILLER_74_2279 ();
 FILLCELL_X32 FILLER_74_2311 ();
 FILLCELL_X32 FILLER_74_2343 ();
 FILLCELL_X32 FILLER_74_2375 ();
 FILLCELL_X32 FILLER_74_2407 ();
 FILLCELL_X32 FILLER_74_2439 ();
 FILLCELL_X32 FILLER_74_2471 ();
 FILLCELL_X32 FILLER_74_2503 ();
 FILLCELL_X32 FILLER_74_2535 ();
 FILLCELL_X32 FILLER_74_2567 ();
 FILLCELL_X2 FILLER_74_2599 ();
 FILLCELL_X1 FILLER_74_2601 ();
 FILLCELL_X32 FILLER_75_1 ();
 FILLCELL_X32 FILLER_75_33 ();
 FILLCELL_X32 FILLER_75_65 ();
 FILLCELL_X32 FILLER_75_97 ();
 FILLCELL_X32 FILLER_75_129 ();
 FILLCELL_X32 FILLER_75_161 ();
 FILLCELL_X32 FILLER_75_193 ();
 FILLCELL_X32 FILLER_75_225 ();
 FILLCELL_X32 FILLER_75_257 ();
 FILLCELL_X32 FILLER_75_289 ();
 FILLCELL_X32 FILLER_75_321 ();
 FILLCELL_X32 FILLER_75_353 ();
 FILLCELL_X32 FILLER_75_385 ();
 FILLCELL_X32 FILLER_75_417 ();
 FILLCELL_X32 FILLER_75_449 ();
 FILLCELL_X32 FILLER_75_481 ();
 FILLCELL_X32 FILLER_75_513 ();
 FILLCELL_X32 FILLER_75_545 ();
 FILLCELL_X32 FILLER_75_577 ();
 FILLCELL_X32 FILLER_75_609 ();
 FILLCELL_X32 FILLER_75_641 ();
 FILLCELL_X32 FILLER_75_673 ();
 FILLCELL_X32 FILLER_75_705 ();
 FILLCELL_X32 FILLER_75_737 ();
 FILLCELL_X32 FILLER_75_769 ();
 FILLCELL_X32 FILLER_75_801 ();
 FILLCELL_X32 FILLER_75_833 ();
 FILLCELL_X32 FILLER_75_865 ();
 FILLCELL_X32 FILLER_75_897 ();
 FILLCELL_X32 FILLER_75_929 ();
 FILLCELL_X32 FILLER_75_961 ();
 FILLCELL_X32 FILLER_75_993 ();
 FILLCELL_X32 FILLER_75_1025 ();
 FILLCELL_X32 FILLER_75_1057 ();
 FILLCELL_X32 FILLER_75_1089 ();
 FILLCELL_X32 FILLER_75_1121 ();
 FILLCELL_X32 FILLER_75_1153 ();
 FILLCELL_X32 FILLER_75_1185 ();
 FILLCELL_X32 FILLER_75_1217 ();
 FILLCELL_X8 FILLER_75_1249 ();
 FILLCELL_X4 FILLER_75_1257 ();
 FILLCELL_X2 FILLER_75_1261 ();
 FILLCELL_X32 FILLER_75_1264 ();
 FILLCELL_X32 FILLER_75_1296 ();
 FILLCELL_X32 FILLER_75_1328 ();
 FILLCELL_X32 FILLER_75_1360 ();
 FILLCELL_X32 FILLER_75_1392 ();
 FILLCELL_X32 FILLER_75_1424 ();
 FILLCELL_X32 FILLER_75_1456 ();
 FILLCELL_X32 FILLER_75_1488 ();
 FILLCELL_X32 FILLER_75_1520 ();
 FILLCELL_X32 FILLER_75_1552 ();
 FILLCELL_X32 FILLER_75_1584 ();
 FILLCELL_X32 FILLER_75_1616 ();
 FILLCELL_X32 FILLER_75_1648 ();
 FILLCELL_X32 FILLER_75_1680 ();
 FILLCELL_X32 FILLER_75_1712 ();
 FILLCELL_X32 FILLER_75_1744 ();
 FILLCELL_X32 FILLER_75_1776 ();
 FILLCELL_X32 FILLER_75_1808 ();
 FILLCELL_X32 FILLER_75_1840 ();
 FILLCELL_X32 FILLER_75_1872 ();
 FILLCELL_X32 FILLER_75_1904 ();
 FILLCELL_X32 FILLER_75_1936 ();
 FILLCELL_X32 FILLER_75_1968 ();
 FILLCELL_X32 FILLER_75_2000 ();
 FILLCELL_X32 FILLER_75_2032 ();
 FILLCELL_X32 FILLER_75_2064 ();
 FILLCELL_X32 FILLER_75_2096 ();
 FILLCELL_X32 FILLER_75_2128 ();
 FILLCELL_X32 FILLER_75_2160 ();
 FILLCELL_X32 FILLER_75_2192 ();
 FILLCELL_X32 FILLER_75_2224 ();
 FILLCELL_X32 FILLER_75_2256 ();
 FILLCELL_X32 FILLER_75_2288 ();
 FILLCELL_X32 FILLER_75_2320 ();
 FILLCELL_X32 FILLER_75_2352 ();
 FILLCELL_X32 FILLER_75_2384 ();
 FILLCELL_X32 FILLER_75_2416 ();
 FILLCELL_X32 FILLER_75_2448 ();
 FILLCELL_X32 FILLER_75_2480 ();
 FILLCELL_X8 FILLER_75_2512 ();
 FILLCELL_X4 FILLER_75_2520 ();
 FILLCELL_X2 FILLER_75_2524 ();
 FILLCELL_X32 FILLER_75_2527 ();
 FILLCELL_X32 FILLER_75_2559 ();
 FILLCELL_X8 FILLER_75_2591 ();
 FILLCELL_X2 FILLER_75_2599 ();
 FILLCELL_X1 FILLER_75_2601 ();
 FILLCELL_X32 FILLER_76_1 ();
 FILLCELL_X32 FILLER_76_33 ();
 FILLCELL_X32 FILLER_76_65 ();
 FILLCELL_X32 FILLER_76_97 ();
 FILLCELL_X32 FILLER_76_129 ();
 FILLCELL_X32 FILLER_76_161 ();
 FILLCELL_X32 FILLER_76_193 ();
 FILLCELL_X32 FILLER_76_225 ();
 FILLCELL_X32 FILLER_76_257 ();
 FILLCELL_X32 FILLER_76_289 ();
 FILLCELL_X32 FILLER_76_321 ();
 FILLCELL_X32 FILLER_76_353 ();
 FILLCELL_X32 FILLER_76_385 ();
 FILLCELL_X32 FILLER_76_417 ();
 FILLCELL_X32 FILLER_76_449 ();
 FILLCELL_X32 FILLER_76_481 ();
 FILLCELL_X32 FILLER_76_513 ();
 FILLCELL_X32 FILLER_76_545 ();
 FILLCELL_X32 FILLER_76_577 ();
 FILLCELL_X16 FILLER_76_609 ();
 FILLCELL_X4 FILLER_76_625 ();
 FILLCELL_X2 FILLER_76_629 ();
 FILLCELL_X32 FILLER_76_632 ();
 FILLCELL_X32 FILLER_76_664 ();
 FILLCELL_X32 FILLER_76_696 ();
 FILLCELL_X32 FILLER_76_728 ();
 FILLCELL_X32 FILLER_76_760 ();
 FILLCELL_X32 FILLER_76_792 ();
 FILLCELL_X32 FILLER_76_824 ();
 FILLCELL_X32 FILLER_76_856 ();
 FILLCELL_X32 FILLER_76_888 ();
 FILLCELL_X32 FILLER_76_920 ();
 FILLCELL_X32 FILLER_76_952 ();
 FILLCELL_X32 FILLER_76_984 ();
 FILLCELL_X32 FILLER_76_1016 ();
 FILLCELL_X32 FILLER_76_1048 ();
 FILLCELL_X32 FILLER_76_1080 ();
 FILLCELL_X32 FILLER_76_1112 ();
 FILLCELL_X32 FILLER_76_1144 ();
 FILLCELL_X32 FILLER_76_1176 ();
 FILLCELL_X32 FILLER_76_1208 ();
 FILLCELL_X32 FILLER_76_1240 ();
 FILLCELL_X32 FILLER_76_1272 ();
 FILLCELL_X32 FILLER_76_1304 ();
 FILLCELL_X32 FILLER_76_1336 ();
 FILLCELL_X32 FILLER_76_1368 ();
 FILLCELL_X32 FILLER_76_1400 ();
 FILLCELL_X32 FILLER_76_1432 ();
 FILLCELL_X32 FILLER_76_1464 ();
 FILLCELL_X32 FILLER_76_1496 ();
 FILLCELL_X32 FILLER_76_1528 ();
 FILLCELL_X32 FILLER_76_1560 ();
 FILLCELL_X32 FILLER_76_1592 ();
 FILLCELL_X32 FILLER_76_1624 ();
 FILLCELL_X32 FILLER_76_1656 ();
 FILLCELL_X32 FILLER_76_1688 ();
 FILLCELL_X32 FILLER_76_1720 ();
 FILLCELL_X32 FILLER_76_1752 ();
 FILLCELL_X32 FILLER_76_1784 ();
 FILLCELL_X32 FILLER_76_1816 ();
 FILLCELL_X32 FILLER_76_1848 ();
 FILLCELL_X8 FILLER_76_1880 ();
 FILLCELL_X4 FILLER_76_1888 ();
 FILLCELL_X2 FILLER_76_1892 ();
 FILLCELL_X32 FILLER_76_1895 ();
 FILLCELL_X32 FILLER_76_1927 ();
 FILLCELL_X32 FILLER_76_1959 ();
 FILLCELL_X32 FILLER_76_1991 ();
 FILLCELL_X32 FILLER_76_2023 ();
 FILLCELL_X32 FILLER_76_2055 ();
 FILLCELL_X32 FILLER_76_2087 ();
 FILLCELL_X32 FILLER_76_2119 ();
 FILLCELL_X32 FILLER_76_2151 ();
 FILLCELL_X32 FILLER_76_2183 ();
 FILLCELL_X32 FILLER_76_2215 ();
 FILLCELL_X32 FILLER_76_2247 ();
 FILLCELL_X32 FILLER_76_2279 ();
 FILLCELL_X32 FILLER_76_2311 ();
 FILLCELL_X32 FILLER_76_2343 ();
 FILLCELL_X32 FILLER_76_2375 ();
 FILLCELL_X32 FILLER_76_2407 ();
 FILLCELL_X32 FILLER_76_2439 ();
 FILLCELL_X32 FILLER_76_2471 ();
 FILLCELL_X32 FILLER_76_2503 ();
 FILLCELL_X32 FILLER_76_2535 ();
 FILLCELL_X32 FILLER_76_2567 ();
 FILLCELL_X2 FILLER_76_2599 ();
 FILLCELL_X1 FILLER_76_2601 ();
 FILLCELL_X32 FILLER_77_1 ();
 FILLCELL_X32 FILLER_77_33 ();
 FILLCELL_X32 FILLER_77_65 ();
 FILLCELL_X32 FILLER_77_97 ();
 FILLCELL_X32 FILLER_77_129 ();
 FILLCELL_X32 FILLER_77_161 ();
 FILLCELL_X32 FILLER_77_193 ();
 FILLCELL_X32 FILLER_77_225 ();
 FILLCELL_X32 FILLER_77_257 ();
 FILLCELL_X32 FILLER_77_289 ();
 FILLCELL_X32 FILLER_77_321 ();
 FILLCELL_X32 FILLER_77_353 ();
 FILLCELL_X32 FILLER_77_385 ();
 FILLCELL_X32 FILLER_77_417 ();
 FILLCELL_X32 FILLER_77_449 ();
 FILLCELL_X32 FILLER_77_481 ();
 FILLCELL_X32 FILLER_77_513 ();
 FILLCELL_X32 FILLER_77_545 ();
 FILLCELL_X32 FILLER_77_577 ();
 FILLCELL_X32 FILLER_77_609 ();
 FILLCELL_X32 FILLER_77_641 ();
 FILLCELL_X32 FILLER_77_673 ();
 FILLCELL_X32 FILLER_77_705 ();
 FILLCELL_X32 FILLER_77_737 ();
 FILLCELL_X32 FILLER_77_769 ();
 FILLCELL_X32 FILLER_77_801 ();
 FILLCELL_X32 FILLER_77_833 ();
 FILLCELL_X32 FILLER_77_865 ();
 FILLCELL_X32 FILLER_77_897 ();
 FILLCELL_X32 FILLER_77_929 ();
 FILLCELL_X32 FILLER_77_961 ();
 FILLCELL_X32 FILLER_77_993 ();
 FILLCELL_X32 FILLER_77_1025 ();
 FILLCELL_X32 FILLER_77_1057 ();
 FILLCELL_X32 FILLER_77_1089 ();
 FILLCELL_X32 FILLER_77_1121 ();
 FILLCELL_X32 FILLER_77_1153 ();
 FILLCELL_X32 FILLER_77_1185 ();
 FILLCELL_X32 FILLER_77_1217 ();
 FILLCELL_X8 FILLER_77_1249 ();
 FILLCELL_X4 FILLER_77_1257 ();
 FILLCELL_X2 FILLER_77_1261 ();
 FILLCELL_X32 FILLER_77_1264 ();
 FILLCELL_X32 FILLER_77_1296 ();
 FILLCELL_X32 FILLER_77_1328 ();
 FILLCELL_X32 FILLER_77_1360 ();
 FILLCELL_X32 FILLER_77_1392 ();
 FILLCELL_X32 FILLER_77_1424 ();
 FILLCELL_X32 FILLER_77_1456 ();
 FILLCELL_X32 FILLER_77_1488 ();
 FILLCELL_X32 FILLER_77_1520 ();
 FILLCELL_X32 FILLER_77_1552 ();
 FILLCELL_X32 FILLER_77_1584 ();
 FILLCELL_X32 FILLER_77_1616 ();
 FILLCELL_X32 FILLER_77_1648 ();
 FILLCELL_X32 FILLER_77_1680 ();
 FILLCELL_X32 FILLER_77_1712 ();
 FILLCELL_X32 FILLER_77_1744 ();
 FILLCELL_X32 FILLER_77_1776 ();
 FILLCELL_X32 FILLER_77_1808 ();
 FILLCELL_X32 FILLER_77_1840 ();
 FILLCELL_X32 FILLER_77_1872 ();
 FILLCELL_X32 FILLER_77_1904 ();
 FILLCELL_X32 FILLER_77_1936 ();
 FILLCELL_X32 FILLER_77_1968 ();
 FILLCELL_X32 FILLER_77_2000 ();
 FILLCELL_X32 FILLER_77_2032 ();
 FILLCELL_X32 FILLER_77_2064 ();
 FILLCELL_X32 FILLER_77_2096 ();
 FILLCELL_X32 FILLER_77_2128 ();
 FILLCELL_X32 FILLER_77_2160 ();
 FILLCELL_X32 FILLER_77_2192 ();
 FILLCELL_X32 FILLER_77_2224 ();
 FILLCELL_X32 FILLER_77_2256 ();
 FILLCELL_X32 FILLER_77_2288 ();
 FILLCELL_X32 FILLER_77_2320 ();
 FILLCELL_X32 FILLER_77_2352 ();
 FILLCELL_X32 FILLER_77_2384 ();
 FILLCELL_X32 FILLER_77_2416 ();
 FILLCELL_X32 FILLER_77_2448 ();
 FILLCELL_X32 FILLER_77_2480 ();
 FILLCELL_X8 FILLER_77_2512 ();
 FILLCELL_X4 FILLER_77_2520 ();
 FILLCELL_X2 FILLER_77_2524 ();
 FILLCELL_X32 FILLER_77_2527 ();
 FILLCELL_X32 FILLER_77_2559 ();
 FILLCELL_X8 FILLER_77_2591 ();
 FILLCELL_X2 FILLER_77_2599 ();
 FILLCELL_X1 FILLER_77_2601 ();
 FILLCELL_X32 FILLER_78_1 ();
 FILLCELL_X32 FILLER_78_33 ();
 FILLCELL_X32 FILLER_78_65 ();
 FILLCELL_X32 FILLER_78_97 ();
 FILLCELL_X32 FILLER_78_129 ();
 FILLCELL_X32 FILLER_78_161 ();
 FILLCELL_X32 FILLER_78_193 ();
 FILLCELL_X32 FILLER_78_225 ();
 FILLCELL_X32 FILLER_78_257 ();
 FILLCELL_X32 FILLER_78_289 ();
 FILLCELL_X32 FILLER_78_321 ();
 FILLCELL_X32 FILLER_78_353 ();
 FILLCELL_X32 FILLER_78_385 ();
 FILLCELL_X32 FILLER_78_417 ();
 FILLCELL_X32 FILLER_78_449 ();
 FILLCELL_X32 FILLER_78_481 ();
 FILLCELL_X32 FILLER_78_513 ();
 FILLCELL_X32 FILLER_78_545 ();
 FILLCELL_X32 FILLER_78_577 ();
 FILLCELL_X16 FILLER_78_609 ();
 FILLCELL_X4 FILLER_78_625 ();
 FILLCELL_X2 FILLER_78_629 ();
 FILLCELL_X32 FILLER_78_632 ();
 FILLCELL_X32 FILLER_78_664 ();
 FILLCELL_X32 FILLER_78_696 ();
 FILLCELL_X32 FILLER_78_728 ();
 FILLCELL_X32 FILLER_78_760 ();
 FILLCELL_X32 FILLER_78_792 ();
 FILLCELL_X32 FILLER_78_824 ();
 FILLCELL_X32 FILLER_78_856 ();
 FILLCELL_X32 FILLER_78_888 ();
 FILLCELL_X32 FILLER_78_920 ();
 FILLCELL_X32 FILLER_78_952 ();
 FILLCELL_X32 FILLER_78_984 ();
 FILLCELL_X32 FILLER_78_1016 ();
 FILLCELL_X32 FILLER_78_1048 ();
 FILLCELL_X32 FILLER_78_1080 ();
 FILLCELL_X32 FILLER_78_1112 ();
 FILLCELL_X32 FILLER_78_1144 ();
 FILLCELL_X32 FILLER_78_1176 ();
 FILLCELL_X32 FILLER_78_1208 ();
 FILLCELL_X32 FILLER_78_1240 ();
 FILLCELL_X32 FILLER_78_1272 ();
 FILLCELL_X32 FILLER_78_1304 ();
 FILLCELL_X32 FILLER_78_1336 ();
 FILLCELL_X32 FILLER_78_1368 ();
 FILLCELL_X32 FILLER_78_1400 ();
 FILLCELL_X32 FILLER_78_1432 ();
 FILLCELL_X32 FILLER_78_1464 ();
 FILLCELL_X32 FILLER_78_1496 ();
 FILLCELL_X32 FILLER_78_1528 ();
 FILLCELL_X32 FILLER_78_1560 ();
 FILLCELL_X32 FILLER_78_1592 ();
 FILLCELL_X32 FILLER_78_1624 ();
 FILLCELL_X32 FILLER_78_1656 ();
 FILLCELL_X32 FILLER_78_1688 ();
 FILLCELL_X32 FILLER_78_1720 ();
 FILLCELL_X32 FILLER_78_1752 ();
 FILLCELL_X32 FILLER_78_1784 ();
 FILLCELL_X32 FILLER_78_1816 ();
 FILLCELL_X32 FILLER_78_1848 ();
 FILLCELL_X8 FILLER_78_1880 ();
 FILLCELL_X4 FILLER_78_1888 ();
 FILLCELL_X2 FILLER_78_1892 ();
 FILLCELL_X32 FILLER_78_1895 ();
 FILLCELL_X32 FILLER_78_1927 ();
 FILLCELL_X32 FILLER_78_1959 ();
 FILLCELL_X32 FILLER_78_1991 ();
 FILLCELL_X32 FILLER_78_2023 ();
 FILLCELL_X32 FILLER_78_2055 ();
 FILLCELL_X32 FILLER_78_2087 ();
 FILLCELL_X32 FILLER_78_2119 ();
 FILLCELL_X32 FILLER_78_2151 ();
 FILLCELL_X32 FILLER_78_2183 ();
 FILLCELL_X32 FILLER_78_2215 ();
 FILLCELL_X32 FILLER_78_2247 ();
 FILLCELL_X32 FILLER_78_2279 ();
 FILLCELL_X32 FILLER_78_2311 ();
 FILLCELL_X32 FILLER_78_2343 ();
 FILLCELL_X32 FILLER_78_2375 ();
 FILLCELL_X32 FILLER_78_2407 ();
 FILLCELL_X32 FILLER_78_2439 ();
 FILLCELL_X32 FILLER_78_2471 ();
 FILLCELL_X32 FILLER_78_2503 ();
 FILLCELL_X32 FILLER_78_2535 ();
 FILLCELL_X32 FILLER_78_2567 ();
 FILLCELL_X2 FILLER_78_2599 ();
 FILLCELL_X1 FILLER_78_2601 ();
 FILLCELL_X32 FILLER_79_1 ();
 FILLCELL_X32 FILLER_79_33 ();
 FILLCELL_X32 FILLER_79_65 ();
 FILLCELL_X32 FILLER_79_97 ();
 FILLCELL_X32 FILLER_79_129 ();
 FILLCELL_X32 FILLER_79_161 ();
 FILLCELL_X32 FILLER_79_193 ();
 FILLCELL_X32 FILLER_79_225 ();
 FILLCELL_X32 FILLER_79_257 ();
 FILLCELL_X32 FILLER_79_289 ();
 FILLCELL_X32 FILLER_79_321 ();
 FILLCELL_X32 FILLER_79_353 ();
 FILLCELL_X32 FILLER_79_385 ();
 FILLCELL_X32 FILLER_79_417 ();
 FILLCELL_X32 FILLER_79_449 ();
 FILLCELL_X32 FILLER_79_481 ();
 FILLCELL_X32 FILLER_79_513 ();
 FILLCELL_X32 FILLER_79_545 ();
 FILLCELL_X32 FILLER_79_577 ();
 FILLCELL_X32 FILLER_79_609 ();
 FILLCELL_X32 FILLER_79_641 ();
 FILLCELL_X32 FILLER_79_673 ();
 FILLCELL_X32 FILLER_79_705 ();
 FILLCELL_X32 FILLER_79_737 ();
 FILLCELL_X32 FILLER_79_769 ();
 FILLCELL_X32 FILLER_79_801 ();
 FILLCELL_X32 FILLER_79_833 ();
 FILLCELL_X32 FILLER_79_865 ();
 FILLCELL_X32 FILLER_79_897 ();
 FILLCELL_X32 FILLER_79_929 ();
 FILLCELL_X32 FILLER_79_961 ();
 FILLCELL_X32 FILLER_79_993 ();
 FILLCELL_X32 FILLER_79_1025 ();
 FILLCELL_X32 FILLER_79_1057 ();
 FILLCELL_X32 FILLER_79_1089 ();
 FILLCELL_X32 FILLER_79_1121 ();
 FILLCELL_X32 FILLER_79_1153 ();
 FILLCELL_X32 FILLER_79_1185 ();
 FILLCELL_X32 FILLER_79_1217 ();
 FILLCELL_X8 FILLER_79_1249 ();
 FILLCELL_X4 FILLER_79_1257 ();
 FILLCELL_X2 FILLER_79_1261 ();
 FILLCELL_X32 FILLER_79_1264 ();
 FILLCELL_X32 FILLER_79_1296 ();
 FILLCELL_X32 FILLER_79_1328 ();
 FILLCELL_X32 FILLER_79_1360 ();
 FILLCELL_X32 FILLER_79_1392 ();
 FILLCELL_X32 FILLER_79_1424 ();
 FILLCELL_X32 FILLER_79_1456 ();
 FILLCELL_X32 FILLER_79_1488 ();
 FILLCELL_X32 FILLER_79_1520 ();
 FILLCELL_X32 FILLER_79_1552 ();
 FILLCELL_X32 FILLER_79_1584 ();
 FILLCELL_X32 FILLER_79_1616 ();
 FILLCELL_X32 FILLER_79_1648 ();
 FILLCELL_X32 FILLER_79_1680 ();
 FILLCELL_X32 FILLER_79_1712 ();
 FILLCELL_X32 FILLER_79_1744 ();
 FILLCELL_X32 FILLER_79_1776 ();
 FILLCELL_X32 FILLER_79_1808 ();
 FILLCELL_X32 FILLER_79_1840 ();
 FILLCELL_X32 FILLER_79_1872 ();
 FILLCELL_X32 FILLER_79_1904 ();
 FILLCELL_X32 FILLER_79_1936 ();
 FILLCELL_X32 FILLER_79_1968 ();
 FILLCELL_X32 FILLER_79_2000 ();
 FILLCELL_X32 FILLER_79_2032 ();
 FILLCELL_X32 FILLER_79_2064 ();
 FILLCELL_X32 FILLER_79_2096 ();
 FILLCELL_X32 FILLER_79_2128 ();
 FILLCELL_X32 FILLER_79_2160 ();
 FILLCELL_X32 FILLER_79_2192 ();
 FILLCELL_X32 FILLER_79_2224 ();
 FILLCELL_X32 FILLER_79_2256 ();
 FILLCELL_X32 FILLER_79_2288 ();
 FILLCELL_X32 FILLER_79_2320 ();
 FILLCELL_X32 FILLER_79_2352 ();
 FILLCELL_X32 FILLER_79_2384 ();
 FILLCELL_X32 FILLER_79_2416 ();
 FILLCELL_X32 FILLER_79_2448 ();
 FILLCELL_X32 FILLER_79_2480 ();
 FILLCELL_X8 FILLER_79_2512 ();
 FILLCELL_X4 FILLER_79_2520 ();
 FILLCELL_X2 FILLER_79_2524 ();
 FILLCELL_X32 FILLER_79_2527 ();
 FILLCELL_X32 FILLER_79_2559 ();
 FILLCELL_X8 FILLER_79_2591 ();
 FILLCELL_X2 FILLER_79_2599 ();
 FILLCELL_X1 FILLER_79_2601 ();
 FILLCELL_X32 FILLER_80_1 ();
 FILLCELL_X32 FILLER_80_33 ();
 FILLCELL_X32 FILLER_80_65 ();
 FILLCELL_X32 FILLER_80_97 ();
 FILLCELL_X32 FILLER_80_129 ();
 FILLCELL_X32 FILLER_80_161 ();
 FILLCELL_X32 FILLER_80_193 ();
 FILLCELL_X32 FILLER_80_225 ();
 FILLCELL_X32 FILLER_80_257 ();
 FILLCELL_X32 FILLER_80_289 ();
 FILLCELL_X32 FILLER_80_321 ();
 FILLCELL_X32 FILLER_80_353 ();
 FILLCELL_X32 FILLER_80_385 ();
 FILLCELL_X32 FILLER_80_417 ();
 FILLCELL_X32 FILLER_80_449 ();
 FILLCELL_X32 FILLER_80_481 ();
 FILLCELL_X32 FILLER_80_513 ();
 FILLCELL_X32 FILLER_80_545 ();
 FILLCELL_X32 FILLER_80_577 ();
 FILLCELL_X16 FILLER_80_609 ();
 FILLCELL_X4 FILLER_80_625 ();
 FILLCELL_X2 FILLER_80_629 ();
 FILLCELL_X32 FILLER_80_632 ();
 FILLCELL_X32 FILLER_80_664 ();
 FILLCELL_X32 FILLER_80_696 ();
 FILLCELL_X32 FILLER_80_728 ();
 FILLCELL_X32 FILLER_80_760 ();
 FILLCELL_X32 FILLER_80_792 ();
 FILLCELL_X32 FILLER_80_824 ();
 FILLCELL_X32 FILLER_80_856 ();
 FILLCELL_X32 FILLER_80_888 ();
 FILLCELL_X32 FILLER_80_920 ();
 FILLCELL_X32 FILLER_80_952 ();
 FILLCELL_X32 FILLER_80_984 ();
 FILLCELL_X32 FILLER_80_1016 ();
 FILLCELL_X32 FILLER_80_1048 ();
 FILLCELL_X32 FILLER_80_1080 ();
 FILLCELL_X32 FILLER_80_1112 ();
 FILLCELL_X32 FILLER_80_1144 ();
 FILLCELL_X32 FILLER_80_1176 ();
 FILLCELL_X32 FILLER_80_1208 ();
 FILLCELL_X32 FILLER_80_1240 ();
 FILLCELL_X32 FILLER_80_1272 ();
 FILLCELL_X32 FILLER_80_1304 ();
 FILLCELL_X32 FILLER_80_1336 ();
 FILLCELL_X32 FILLER_80_1368 ();
 FILLCELL_X32 FILLER_80_1400 ();
 FILLCELL_X32 FILLER_80_1432 ();
 FILLCELL_X32 FILLER_80_1464 ();
 FILLCELL_X32 FILLER_80_1496 ();
 FILLCELL_X32 FILLER_80_1528 ();
 FILLCELL_X32 FILLER_80_1560 ();
 FILLCELL_X32 FILLER_80_1592 ();
 FILLCELL_X32 FILLER_80_1624 ();
 FILLCELL_X32 FILLER_80_1656 ();
 FILLCELL_X32 FILLER_80_1688 ();
 FILLCELL_X32 FILLER_80_1720 ();
 FILLCELL_X32 FILLER_80_1752 ();
 FILLCELL_X32 FILLER_80_1784 ();
 FILLCELL_X32 FILLER_80_1816 ();
 FILLCELL_X32 FILLER_80_1848 ();
 FILLCELL_X8 FILLER_80_1880 ();
 FILLCELL_X4 FILLER_80_1888 ();
 FILLCELL_X2 FILLER_80_1892 ();
 FILLCELL_X32 FILLER_80_1895 ();
 FILLCELL_X32 FILLER_80_1927 ();
 FILLCELL_X32 FILLER_80_1959 ();
 FILLCELL_X32 FILLER_80_1991 ();
 FILLCELL_X32 FILLER_80_2023 ();
 FILLCELL_X32 FILLER_80_2055 ();
 FILLCELL_X32 FILLER_80_2087 ();
 FILLCELL_X32 FILLER_80_2119 ();
 FILLCELL_X32 FILLER_80_2151 ();
 FILLCELL_X32 FILLER_80_2183 ();
 FILLCELL_X32 FILLER_80_2215 ();
 FILLCELL_X32 FILLER_80_2247 ();
 FILLCELL_X32 FILLER_80_2279 ();
 FILLCELL_X32 FILLER_80_2311 ();
 FILLCELL_X32 FILLER_80_2343 ();
 FILLCELL_X32 FILLER_80_2375 ();
 FILLCELL_X32 FILLER_80_2407 ();
 FILLCELL_X32 FILLER_80_2439 ();
 FILLCELL_X32 FILLER_80_2471 ();
 FILLCELL_X32 FILLER_80_2503 ();
 FILLCELL_X32 FILLER_80_2535 ();
 FILLCELL_X32 FILLER_80_2567 ();
 FILLCELL_X2 FILLER_80_2599 ();
 FILLCELL_X1 FILLER_80_2601 ();
 FILLCELL_X32 FILLER_81_1 ();
 FILLCELL_X32 FILLER_81_33 ();
 FILLCELL_X32 FILLER_81_65 ();
 FILLCELL_X32 FILLER_81_97 ();
 FILLCELL_X32 FILLER_81_129 ();
 FILLCELL_X32 FILLER_81_161 ();
 FILLCELL_X32 FILLER_81_193 ();
 FILLCELL_X32 FILLER_81_225 ();
 FILLCELL_X32 FILLER_81_257 ();
 FILLCELL_X32 FILLER_81_289 ();
 FILLCELL_X32 FILLER_81_321 ();
 FILLCELL_X32 FILLER_81_353 ();
 FILLCELL_X32 FILLER_81_385 ();
 FILLCELL_X32 FILLER_81_417 ();
 FILLCELL_X32 FILLER_81_449 ();
 FILLCELL_X32 FILLER_81_481 ();
 FILLCELL_X32 FILLER_81_513 ();
 FILLCELL_X32 FILLER_81_545 ();
 FILLCELL_X32 FILLER_81_577 ();
 FILLCELL_X32 FILLER_81_609 ();
 FILLCELL_X32 FILLER_81_641 ();
 FILLCELL_X32 FILLER_81_673 ();
 FILLCELL_X32 FILLER_81_705 ();
 FILLCELL_X32 FILLER_81_737 ();
 FILLCELL_X32 FILLER_81_769 ();
 FILLCELL_X32 FILLER_81_801 ();
 FILLCELL_X32 FILLER_81_833 ();
 FILLCELL_X32 FILLER_81_865 ();
 FILLCELL_X32 FILLER_81_897 ();
 FILLCELL_X32 FILLER_81_929 ();
 FILLCELL_X32 FILLER_81_961 ();
 FILLCELL_X32 FILLER_81_993 ();
 FILLCELL_X32 FILLER_81_1025 ();
 FILLCELL_X32 FILLER_81_1057 ();
 FILLCELL_X32 FILLER_81_1089 ();
 FILLCELL_X32 FILLER_81_1121 ();
 FILLCELL_X32 FILLER_81_1153 ();
 FILLCELL_X32 FILLER_81_1185 ();
 FILLCELL_X32 FILLER_81_1217 ();
 FILLCELL_X8 FILLER_81_1249 ();
 FILLCELL_X4 FILLER_81_1257 ();
 FILLCELL_X2 FILLER_81_1261 ();
 FILLCELL_X32 FILLER_81_1264 ();
 FILLCELL_X32 FILLER_81_1296 ();
 FILLCELL_X32 FILLER_81_1328 ();
 FILLCELL_X32 FILLER_81_1360 ();
 FILLCELL_X32 FILLER_81_1392 ();
 FILLCELL_X32 FILLER_81_1424 ();
 FILLCELL_X32 FILLER_81_1456 ();
 FILLCELL_X32 FILLER_81_1488 ();
 FILLCELL_X32 FILLER_81_1520 ();
 FILLCELL_X32 FILLER_81_1552 ();
 FILLCELL_X32 FILLER_81_1584 ();
 FILLCELL_X32 FILLER_81_1616 ();
 FILLCELL_X32 FILLER_81_1648 ();
 FILLCELL_X32 FILLER_81_1680 ();
 FILLCELL_X32 FILLER_81_1712 ();
 FILLCELL_X32 FILLER_81_1744 ();
 FILLCELL_X32 FILLER_81_1776 ();
 FILLCELL_X32 FILLER_81_1808 ();
 FILLCELL_X32 FILLER_81_1840 ();
 FILLCELL_X32 FILLER_81_1872 ();
 FILLCELL_X32 FILLER_81_1904 ();
 FILLCELL_X32 FILLER_81_1936 ();
 FILLCELL_X32 FILLER_81_1968 ();
 FILLCELL_X32 FILLER_81_2000 ();
 FILLCELL_X32 FILLER_81_2032 ();
 FILLCELL_X32 FILLER_81_2064 ();
 FILLCELL_X32 FILLER_81_2096 ();
 FILLCELL_X32 FILLER_81_2128 ();
 FILLCELL_X32 FILLER_81_2160 ();
 FILLCELL_X32 FILLER_81_2192 ();
 FILLCELL_X32 FILLER_81_2224 ();
 FILLCELL_X32 FILLER_81_2256 ();
 FILLCELL_X32 FILLER_81_2288 ();
 FILLCELL_X32 FILLER_81_2320 ();
 FILLCELL_X32 FILLER_81_2352 ();
 FILLCELL_X32 FILLER_81_2384 ();
 FILLCELL_X32 FILLER_81_2416 ();
 FILLCELL_X32 FILLER_81_2448 ();
 FILLCELL_X32 FILLER_81_2480 ();
 FILLCELL_X8 FILLER_81_2512 ();
 FILLCELL_X4 FILLER_81_2520 ();
 FILLCELL_X2 FILLER_81_2524 ();
 FILLCELL_X32 FILLER_81_2527 ();
 FILLCELL_X32 FILLER_81_2559 ();
 FILLCELL_X8 FILLER_81_2591 ();
 FILLCELL_X2 FILLER_81_2599 ();
 FILLCELL_X1 FILLER_81_2601 ();
 FILLCELL_X32 FILLER_82_1 ();
 FILLCELL_X32 FILLER_82_33 ();
 FILLCELL_X32 FILLER_82_65 ();
 FILLCELL_X32 FILLER_82_97 ();
 FILLCELL_X32 FILLER_82_129 ();
 FILLCELL_X32 FILLER_82_161 ();
 FILLCELL_X32 FILLER_82_193 ();
 FILLCELL_X32 FILLER_82_225 ();
 FILLCELL_X32 FILLER_82_257 ();
 FILLCELL_X32 FILLER_82_289 ();
 FILLCELL_X32 FILLER_82_321 ();
 FILLCELL_X32 FILLER_82_353 ();
 FILLCELL_X32 FILLER_82_385 ();
 FILLCELL_X32 FILLER_82_417 ();
 FILLCELL_X32 FILLER_82_449 ();
 FILLCELL_X32 FILLER_82_481 ();
 FILLCELL_X32 FILLER_82_513 ();
 FILLCELL_X32 FILLER_82_545 ();
 FILLCELL_X32 FILLER_82_577 ();
 FILLCELL_X16 FILLER_82_609 ();
 FILLCELL_X4 FILLER_82_625 ();
 FILLCELL_X2 FILLER_82_629 ();
 FILLCELL_X32 FILLER_82_632 ();
 FILLCELL_X32 FILLER_82_664 ();
 FILLCELL_X32 FILLER_82_696 ();
 FILLCELL_X32 FILLER_82_728 ();
 FILLCELL_X32 FILLER_82_760 ();
 FILLCELL_X32 FILLER_82_792 ();
 FILLCELL_X32 FILLER_82_824 ();
 FILLCELL_X32 FILLER_82_856 ();
 FILLCELL_X32 FILLER_82_888 ();
 FILLCELL_X32 FILLER_82_920 ();
 FILLCELL_X32 FILLER_82_952 ();
 FILLCELL_X32 FILLER_82_984 ();
 FILLCELL_X32 FILLER_82_1016 ();
 FILLCELL_X32 FILLER_82_1048 ();
 FILLCELL_X32 FILLER_82_1080 ();
 FILLCELL_X32 FILLER_82_1112 ();
 FILLCELL_X32 FILLER_82_1144 ();
 FILLCELL_X32 FILLER_82_1176 ();
 FILLCELL_X32 FILLER_82_1208 ();
 FILLCELL_X32 FILLER_82_1240 ();
 FILLCELL_X32 FILLER_82_1272 ();
 FILLCELL_X32 FILLER_82_1304 ();
 FILLCELL_X32 FILLER_82_1336 ();
 FILLCELL_X32 FILLER_82_1368 ();
 FILLCELL_X32 FILLER_82_1400 ();
 FILLCELL_X32 FILLER_82_1432 ();
 FILLCELL_X32 FILLER_82_1464 ();
 FILLCELL_X32 FILLER_82_1496 ();
 FILLCELL_X32 FILLER_82_1528 ();
 FILLCELL_X32 FILLER_82_1560 ();
 FILLCELL_X32 FILLER_82_1592 ();
 FILLCELL_X32 FILLER_82_1624 ();
 FILLCELL_X32 FILLER_82_1656 ();
 FILLCELL_X32 FILLER_82_1688 ();
 FILLCELL_X32 FILLER_82_1720 ();
 FILLCELL_X32 FILLER_82_1752 ();
 FILLCELL_X32 FILLER_82_1784 ();
 FILLCELL_X32 FILLER_82_1816 ();
 FILLCELL_X32 FILLER_82_1848 ();
 FILLCELL_X8 FILLER_82_1880 ();
 FILLCELL_X4 FILLER_82_1888 ();
 FILLCELL_X2 FILLER_82_1892 ();
 FILLCELL_X32 FILLER_82_1895 ();
 FILLCELL_X32 FILLER_82_1927 ();
 FILLCELL_X32 FILLER_82_1959 ();
 FILLCELL_X32 FILLER_82_1991 ();
 FILLCELL_X32 FILLER_82_2023 ();
 FILLCELL_X32 FILLER_82_2055 ();
 FILLCELL_X32 FILLER_82_2087 ();
 FILLCELL_X32 FILLER_82_2119 ();
 FILLCELL_X32 FILLER_82_2151 ();
 FILLCELL_X32 FILLER_82_2183 ();
 FILLCELL_X32 FILLER_82_2215 ();
 FILLCELL_X32 FILLER_82_2247 ();
 FILLCELL_X32 FILLER_82_2279 ();
 FILLCELL_X32 FILLER_82_2311 ();
 FILLCELL_X32 FILLER_82_2343 ();
 FILLCELL_X32 FILLER_82_2375 ();
 FILLCELL_X32 FILLER_82_2407 ();
 FILLCELL_X32 FILLER_82_2439 ();
 FILLCELL_X32 FILLER_82_2471 ();
 FILLCELL_X32 FILLER_82_2503 ();
 FILLCELL_X32 FILLER_82_2535 ();
 FILLCELL_X32 FILLER_82_2567 ();
 FILLCELL_X2 FILLER_82_2599 ();
 FILLCELL_X1 FILLER_82_2601 ();
 FILLCELL_X32 FILLER_83_1 ();
 FILLCELL_X32 FILLER_83_33 ();
 FILLCELL_X32 FILLER_83_65 ();
 FILLCELL_X32 FILLER_83_97 ();
 FILLCELL_X32 FILLER_83_129 ();
 FILLCELL_X32 FILLER_83_161 ();
 FILLCELL_X32 FILLER_83_193 ();
 FILLCELL_X32 FILLER_83_225 ();
 FILLCELL_X32 FILLER_83_257 ();
 FILLCELL_X32 FILLER_83_289 ();
 FILLCELL_X32 FILLER_83_321 ();
 FILLCELL_X32 FILLER_83_353 ();
 FILLCELL_X32 FILLER_83_385 ();
 FILLCELL_X32 FILLER_83_417 ();
 FILLCELL_X32 FILLER_83_449 ();
 FILLCELL_X32 FILLER_83_481 ();
 FILLCELL_X32 FILLER_83_513 ();
 FILLCELL_X32 FILLER_83_545 ();
 FILLCELL_X32 FILLER_83_577 ();
 FILLCELL_X32 FILLER_83_609 ();
 FILLCELL_X32 FILLER_83_641 ();
 FILLCELL_X32 FILLER_83_673 ();
 FILLCELL_X32 FILLER_83_705 ();
 FILLCELL_X32 FILLER_83_737 ();
 FILLCELL_X32 FILLER_83_769 ();
 FILLCELL_X32 FILLER_83_801 ();
 FILLCELL_X32 FILLER_83_833 ();
 FILLCELL_X32 FILLER_83_865 ();
 FILLCELL_X32 FILLER_83_897 ();
 FILLCELL_X32 FILLER_83_929 ();
 FILLCELL_X32 FILLER_83_961 ();
 FILLCELL_X32 FILLER_83_993 ();
 FILLCELL_X32 FILLER_83_1025 ();
 FILLCELL_X32 FILLER_83_1057 ();
 FILLCELL_X32 FILLER_83_1089 ();
 FILLCELL_X32 FILLER_83_1121 ();
 FILLCELL_X32 FILLER_83_1153 ();
 FILLCELL_X32 FILLER_83_1185 ();
 FILLCELL_X32 FILLER_83_1217 ();
 FILLCELL_X8 FILLER_83_1249 ();
 FILLCELL_X4 FILLER_83_1257 ();
 FILLCELL_X2 FILLER_83_1261 ();
 FILLCELL_X32 FILLER_83_1264 ();
 FILLCELL_X32 FILLER_83_1296 ();
 FILLCELL_X32 FILLER_83_1328 ();
 FILLCELL_X32 FILLER_83_1360 ();
 FILLCELL_X32 FILLER_83_1392 ();
 FILLCELL_X32 FILLER_83_1424 ();
 FILLCELL_X32 FILLER_83_1456 ();
 FILLCELL_X32 FILLER_83_1488 ();
 FILLCELL_X32 FILLER_83_1520 ();
 FILLCELL_X32 FILLER_83_1552 ();
 FILLCELL_X32 FILLER_83_1584 ();
 FILLCELL_X32 FILLER_83_1616 ();
 FILLCELL_X32 FILLER_83_1648 ();
 FILLCELL_X32 FILLER_83_1680 ();
 FILLCELL_X32 FILLER_83_1712 ();
 FILLCELL_X32 FILLER_83_1744 ();
 FILLCELL_X32 FILLER_83_1776 ();
 FILLCELL_X32 FILLER_83_1808 ();
 FILLCELL_X32 FILLER_83_1840 ();
 FILLCELL_X32 FILLER_83_1872 ();
 FILLCELL_X32 FILLER_83_1904 ();
 FILLCELL_X32 FILLER_83_1936 ();
 FILLCELL_X32 FILLER_83_1968 ();
 FILLCELL_X32 FILLER_83_2000 ();
 FILLCELL_X32 FILLER_83_2032 ();
 FILLCELL_X32 FILLER_83_2064 ();
 FILLCELL_X32 FILLER_83_2096 ();
 FILLCELL_X32 FILLER_83_2128 ();
 FILLCELL_X32 FILLER_83_2160 ();
 FILLCELL_X32 FILLER_83_2192 ();
 FILLCELL_X32 FILLER_83_2224 ();
 FILLCELL_X32 FILLER_83_2256 ();
 FILLCELL_X32 FILLER_83_2288 ();
 FILLCELL_X32 FILLER_83_2320 ();
 FILLCELL_X32 FILLER_83_2352 ();
 FILLCELL_X32 FILLER_83_2384 ();
 FILLCELL_X32 FILLER_83_2416 ();
 FILLCELL_X32 FILLER_83_2448 ();
 FILLCELL_X32 FILLER_83_2480 ();
 FILLCELL_X8 FILLER_83_2512 ();
 FILLCELL_X4 FILLER_83_2520 ();
 FILLCELL_X2 FILLER_83_2524 ();
 FILLCELL_X32 FILLER_83_2527 ();
 FILLCELL_X32 FILLER_83_2559 ();
 FILLCELL_X8 FILLER_83_2591 ();
 FILLCELL_X2 FILLER_83_2599 ();
 FILLCELL_X1 FILLER_83_2601 ();
 FILLCELL_X32 FILLER_84_1 ();
 FILLCELL_X32 FILLER_84_33 ();
 FILLCELL_X32 FILLER_84_65 ();
 FILLCELL_X32 FILLER_84_97 ();
 FILLCELL_X32 FILLER_84_129 ();
 FILLCELL_X32 FILLER_84_161 ();
 FILLCELL_X32 FILLER_84_193 ();
 FILLCELL_X32 FILLER_84_225 ();
 FILLCELL_X32 FILLER_84_257 ();
 FILLCELL_X32 FILLER_84_289 ();
 FILLCELL_X32 FILLER_84_321 ();
 FILLCELL_X32 FILLER_84_353 ();
 FILLCELL_X32 FILLER_84_385 ();
 FILLCELL_X32 FILLER_84_417 ();
 FILLCELL_X32 FILLER_84_449 ();
 FILLCELL_X32 FILLER_84_481 ();
 FILLCELL_X32 FILLER_84_513 ();
 FILLCELL_X32 FILLER_84_545 ();
 FILLCELL_X32 FILLER_84_577 ();
 FILLCELL_X16 FILLER_84_609 ();
 FILLCELL_X4 FILLER_84_625 ();
 FILLCELL_X2 FILLER_84_629 ();
 FILLCELL_X32 FILLER_84_632 ();
 FILLCELL_X32 FILLER_84_664 ();
 FILLCELL_X32 FILLER_84_696 ();
 FILLCELL_X32 FILLER_84_728 ();
 FILLCELL_X32 FILLER_84_760 ();
 FILLCELL_X32 FILLER_84_792 ();
 FILLCELL_X32 FILLER_84_824 ();
 FILLCELL_X32 FILLER_84_856 ();
 FILLCELL_X32 FILLER_84_888 ();
 FILLCELL_X32 FILLER_84_920 ();
 FILLCELL_X32 FILLER_84_952 ();
 FILLCELL_X32 FILLER_84_984 ();
 FILLCELL_X32 FILLER_84_1016 ();
 FILLCELL_X32 FILLER_84_1048 ();
 FILLCELL_X32 FILLER_84_1080 ();
 FILLCELL_X32 FILLER_84_1112 ();
 FILLCELL_X32 FILLER_84_1144 ();
 FILLCELL_X32 FILLER_84_1176 ();
 FILLCELL_X32 FILLER_84_1208 ();
 FILLCELL_X32 FILLER_84_1240 ();
 FILLCELL_X32 FILLER_84_1272 ();
 FILLCELL_X32 FILLER_84_1304 ();
 FILLCELL_X32 FILLER_84_1336 ();
 FILLCELL_X32 FILLER_84_1368 ();
 FILLCELL_X32 FILLER_84_1400 ();
 FILLCELL_X32 FILLER_84_1432 ();
 FILLCELL_X32 FILLER_84_1464 ();
 FILLCELL_X32 FILLER_84_1496 ();
 FILLCELL_X32 FILLER_84_1528 ();
 FILLCELL_X32 FILLER_84_1560 ();
 FILLCELL_X32 FILLER_84_1592 ();
 FILLCELL_X32 FILLER_84_1624 ();
 FILLCELL_X32 FILLER_84_1656 ();
 FILLCELL_X32 FILLER_84_1688 ();
 FILLCELL_X32 FILLER_84_1720 ();
 FILLCELL_X32 FILLER_84_1752 ();
 FILLCELL_X32 FILLER_84_1784 ();
 FILLCELL_X32 FILLER_84_1816 ();
 FILLCELL_X32 FILLER_84_1848 ();
 FILLCELL_X8 FILLER_84_1880 ();
 FILLCELL_X4 FILLER_84_1888 ();
 FILLCELL_X2 FILLER_84_1892 ();
 FILLCELL_X32 FILLER_84_1895 ();
 FILLCELL_X32 FILLER_84_1927 ();
 FILLCELL_X32 FILLER_84_1959 ();
 FILLCELL_X32 FILLER_84_1991 ();
 FILLCELL_X32 FILLER_84_2023 ();
 FILLCELL_X32 FILLER_84_2055 ();
 FILLCELL_X32 FILLER_84_2087 ();
 FILLCELL_X32 FILLER_84_2119 ();
 FILLCELL_X32 FILLER_84_2151 ();
 FILLCELL_X32 FILLER_84_2183 ();
 FILLCELL_X32 FILLER_84_2215 ();
 FILLCELL_X32 FILLER_84_2247 ();
 FILLCELL_X32 FILLER_84_2279 ();
 FILLCELL_X32 FILLER_84_2311 ();
 FILLCELL_X32 FILLER_84_2343 ();
 FILLCELL_X32 FILLER_84_2375 ();
 FILLCELL_X32 FILLER_84_2407 ();
 FILLCELL_X32 FILLER_84_2439 ();
 FILLCELL_X32 FILLER_84_2471 ();
 FILLCELL_X32 FILLER_84_2503 ();
 FILLCELL_X32 FILLER_84_2535 ();
 FILLCELL_X32 FILLER_84_2567 ();
 FILLCELL_X2 FILLER_84_2599 ();
 FILLCELL_X1 FILLER_84_2601 ();
 FILLCELL_X32 FILLER_85_1 ();
 FILLCELL_X32 FILLER_85_33 ();
 FILLCELL_X32 FILLER_85_65 ();
 FILLCELL_X32 FILLER_85_97 ();
 FILLCELL_X32 FILLER_85_129 ();
 FILLCELL_X32 FILLER_85_161 ();
 FILLCELL_X32 FILLER_85_193 ();
 FILLCELL_X32 FILLER_85_225 ();
 FILLCELL_X32 FILLER_85_257 ();
 FILLCELL_X32 FILLER_85_289 ();
 FILLCELL_X32 FILLER_85_321 ();
 FILLCELL_X32 FILLER_85_353 ();
 FILLCELL_X32 FILLER_85_385 ();
 FILLCELL_X32 FILLER_85_417 ();
 FILLCELL_X32 FILLER_85_449 ();
 FILLCELL_X32 FILLER_85_481 ();
 FILLCELL_X32 FILLER_85_513 ();
 FILLCELL_X32 FILLER_85_545 ();
 FILLCELL_X32 FILLER_85_577 ();
 FILLCELL_X32 FILLER_85_609 ();
 FILLCELL_X32 FILLER_85_641 ();
 FILLCELL_X32 FILLER_85_673 ();
 FILLCELL_X32 FILLER_85_705 ();
 FILLCELL_X32 FILLER_85_737 ();
 FILLCELL_X32 FILLER_85_769 ();
 FILLCELL_X32 FILLER_85_801 ();
 FILLCELL_X32 FILLER_85_833 ();
 FILLCELL_X32 FILLER_85_865 ();
 FILLCELL_X32 FILLER_85_897 ();
 FILLCELL_X32 FILLER_85_929 ();
 FILLCELL_X32 FILLER_85_961 ();
 FILLCELL_X32 FILLER_85_993 ();
 FILLCELL_X32 FILLER_85_1025 ();
 FILLCELL_X32 FILLER_85_1057 ();
 FILLCELL_X32 FILLER_85_1089 ();
 FILLCELL_X32 FILLER_85_1121 ();
 FILLCELL_X32 FILLER_85_1153 ();
 FILLCELL_X32 FILLER_85_1185 ();
 FILLCELL_X32 FILLER_85_1217 ();
 FILLCELL_X8 FILLER_85_1249 ();
 FILLCELL_X4 FILLER_85_1257 ();
 FILLCELL_X2 FILLER_85_1261 ();
 FILLCELL_X32 FILLER_85_1264 ();
 FILLCELL_X32 FILLER_85_1296 ();
 FILLCELL_X32 FILLER_85_1328 ();
 FILLCELL_X32 FILLER_85_1360 ();
 FILLCELL_X32 FILLER_85_1392 ();
 FILLCELL_X32 FILLER_85_1424 ();
 FILLCELL_X32 FILLER_85_1456 ();
 FILLCELL_X32 FILLER_85_1488 ();
 FILLCELL_X32 FILLER_85_1520 ();
 FILLCELL_X32 FILLER_85_1552 ();
 FILLCELL_X32 FILLER_85_1584 ();
 FILLCELL_X32 FILLER_85_1616 ();
 FILLCELL_X32 FILLER_85_1648 ();
 FILLCELL_X32 FILLER_85_1680 ();
 FILLCELL_X32 FILLER_85_1712 ();
 FILLCELL_X32 FILLER_85_1744 ();
 FILLCELL_X32 FILLER_85_1776 ();
 FILLCELL_X32 FILLER_85_1808 ();
 FILLCELL_X32 FILLER_85_1840 ();
 FILLCELL_X32 FILLER_85_1872 ();
 FILLCELL_X32 FILLER_85_1904 ();
 FILLCELL_X32 FILLER_85_1936 ();
 FILLCELL_X32 FILLER_85_1968 ();
 FILLCELL_X32 FILLER_85_2000 ();
 FILLCELL_X32 FILLER_85_2032 ();
 FILLCELL_X32 FILLER_85_2064 ();
 FILLCELL_X32 FILLER_85_2096 ();
 FILLCELL_X32 FILLER_85_2128 ();
 FILLCELL_X32 FILLER_85_2160 ();
 FILLCELL_X32 FILLER_85_2192 ();
 FILLCELL_X32 FILLER_85_2224 ();
 FILLCELL_X32 FILLER_85_2256 ();
 FILLCELL_X32 FILLER_85_2288 ();
 FILLCELL_X32 FILLER_85_2320 ();
 FILLCELL_X32 FILLER_85_2352 ();
 FILLCELL_X32 FILLER_85_2384 ();
 FILLCELL_X32 FILLER_85_2416 ();
 FILLCELL_X32 FILLER_85_2448 ();
 FILLCELL_X32 FILLER_85_2480 ();
 FILLCELL_X8 FILLER_85_2512 ();
 FILLCELL_X4 FILLER_85_2520 ();
 FILLCELL_X2 FILLER_85_2524 ();
 FILLCELL_X32 FILLER_85_2527 ();
 FILLCELL_X32 FILLER_85_2559 ();
 FILLCELL_X8 FILLER_85_2591 ();
 FILLCELL_X2 FILLER_85_2599 ();
 FILLCELL_X1 FILLER_85_2601 ();
 FILLCELL_X32 FILLER_86_1 ();
 FILLCELL_X32 FILLER_86_33 ();
 FILLCELL_X32 FILLER_86_65 ();
 FILLCELL_X32 FILLER_86_97 ();
 FILLCELL_X32 FILLER_86_129 ();
 FILLCELL_X32 FILLER_86_161 ();
 FILLCELL_X32 FILLER_86_193 ();
 FILLCELL_X32 FILLER_86_225 ();
 FILLCELL_X32 FILLER_86_257 ();
 FILLCELL_X32 FILLER_86_289 ();
 FILLCELL_X32 FILLER_86_321 ();
 FILLCELL_X32 FILLER_86_353 ();
 FILLCELL_X32 FILLER_86_385 ();
 FILLCELL_X32 FILLER_86_417 ();
 FILLCELL_X32 FILLER_86_449 ();
 FILLCELL_X32 FILLER_86_481 ();
 FILLCELL_X32 FILLER_86_513 ();
 FILLCELL_X32 FILLER_86_545 ();
 FILLCELL_X32 FILLER_86_577 ();
 FILLCELL_X16 FILLER_86_609 ();
 FILLCELL_X4 FILLER_86_625 ();
 FILLCELL_X2 FILLER_86_629 ();
 FILLCELL_X32 FILLER_86_632 ();
 FILLCELL_X32 FILLER_86_664 ();
 FILLCELL_X32 FILLER_86_696 ();
 FILLCELL_X32 FILLER_86_728 ();
 FILLCELL_X32 FILLER_86_760 ();
 FILLCELL_X32 FILLER_86_792 ();
 FILLCELL_X32 FILLER_86_824 ();
 FILLCELL_X32 FILLER_86_856 ();
 FILLCELL_X32 FILLER_86_888 ();
 FILLCELL_X32 FILLER_86_920 ();
 FILLCELL_X32 FILLER_86_952 ();
 FILLCELL_X32 FILLER_86_984 ();
 FILLCELL_X32 FILLER_86_1016 ();
 FILLCELL_X32 FILLER_86_1048 ();
 FILLCELL_X32 FILLER_86_1080 ();
 FILLCELL_X32 FILLER_86_1112 ();
 FILLCELL_X32 FILLER_86_1144 ();
 FILLCELL_X32 FILLER_86_1176 ();
 FILLCELL_X32 FILLER_86_1208 ();
 FILLCELL_X32 FILLER_86_1240 ();
 FILLCELL_X32 FILLER_86_1272 ();
 FILLCELL_X32 FILLER_86_1304 ();
 FILLCELL_X32 FILLER_86_1336 ();
 FILLCELL_X32 FILLER_86_1368 ();
 FILLCELL_X32 FILLER_86_1400 ();
 FILLCELL_X32 FILLER_86_1432 ();
 FILLCELL_X32 FILLER_86_1464 ();
 FILLCELL_X32 FILLER_86_1496 ();
 FILLCELL_X32 FILLER_86_1528 ();
 FILLCELL_X32 FILLER_86_1560 ();
 FILLCELL_X32 FILLER_86_1592 ();
 FILLCELL_X32 FILLER_86_1624 ();
 FILLCELL_X32 FILLER_86_1656 ();
 FILLCELL_X32 FILLER_86_1688 ();
 FILLCELL_X32 FILLER_86_1720 ();
 FILLCELL_X32 FILLER_86_1752 ();
 FILLCELL_X32 FILLER_86_1784 ();
 FILLCELL_X32 FILLER_86_1816 ();
 FILLCELL_X32 FILLER_86_1848 ();
 FILLCELL_X8 FILLER_86_1880 ();
 FILLCELL_X4 FILLER_86_1888 ();
 FILLCELL_X2 FILLER_86_1892 ();
 FILLCELL_X32 FILLER_86_1895 ();
 FILLCELL_X32 FILLER_86_1927 ();
 FILLCELL_X32 FILLER_86_1959 ();
 FILLCELL_X32 FILLER_86_1991 ();
 FILLCELL_X32 FILLER_86_2023 ();
 FILLCELL_X32 FILLER_86_2055 ();
 FILLCELL_X32 FILLER_86_2087 ();
 FILLCELL_X32 FILLER_86_2119 ();
 FILLCELL_X32 FILLER_86_2151 ();
 FILLCELL_X32 FILLER_86_2183 ();
 FILLCELL_X32 FILLER_86_2215 ();
 FILLCELL_X32 FILLER_86_2247 ();
 FILLCELL_X32 FILLER_86_2279 ();
 FILLCELL_X32 FILLER_86_2311 ();
 FILLCELL_X32 FILLER_86_2343 ();
 FILLCELL_X32 FILLER_86_2375 ();
 FILLCELL_X32 FILLER_86_2407 ();
 FILLCELL_X32 FILLER_86_2439 ();
 FILLCELL_X32 FILLER_86_2471 ();
 FILLCELL_X32 FILLER_86_2503 ();
 FILLCELL_X32 FILLER_86_2535 ();
 FILLCELL_X32 FILLER_86_2567 ();
 FILLCELL_X2 FILLER_86_2599 ();
 FILLCELL_X1 FILLER_86_2601 ();
 FILLCELL_X32 FILLER_87_1 ();
 FILLCELL_X32 FILLER_87_33 ();
 FILLCELL_X32 FILLER_87_65 ();
 FILLCELL_X32 FILLER_87_97 ();
 FILLCELL_X32 FILLER_87_129 ();
 FILLCELL_X32 FILLER_87_161 ();
 FILLCELL_X32 FILLER_87_193 ();
 FILLCELL_X32 FILLER_87_225 ();
 FILLCELL_X32 FILLER_87_257 ();
 FILLCELL_X32 FILLER_87_289 ();
 FILLCELL_X32 FILLER_87_321 ();
 FILLCELL_X32 FILLER_87_353 ();
 FILLCELL_X32 FILLER_87_385 ();
 FILLCELL_X32 FILLER_87_417 ();
 FILLCELL_X32 FILLER_87_449 ();
 FILLCELL_X32 FILLER_87_481 ();
 FILLCELL_X32 FILLER_87_513 ();
 FILLCELL_X32 FILLER_87_545 ();
 FILLCELL_X32 FILLER_87_577 ();
 FILLCELL_X32 FILLER_87_609 ();
 FILLCELL_X32 FILLER_87_641 ();
 FILLCELL_X32 FILLER_87_673 ();
 FILLCELL_X32 FILLER_87_705 ();
 FILLCELL_X32 FILLER_87_737 ();
 FILLCELL_X32 FILLER_87_769 ();
 FILLCELL_X32 FILLER_87_801 ();
 FILLCELL_X32 FILLER_87_833 ();
 FILLCELL_X32 FILLER_87_865 ();
 FILLCELL_X32 FILLER_87_897 ();
 FILLCELL_X32 FILLER_87_929 ();
 FILLCELL_X32 FILLER_87_961 ();
 FILLCELL_X32 FILLER_87_993 ();
 FILLCELL_X32 FILLER_87_1025 ();
 FILLCELL_X32 FILLER_87_1057 ();
 FILLCELL_X32 FILLER_87_1089 ();
 FILLCELL_X32 FILLER_87_1121 ();
 FILLCELL_X32 FILLER_87_1153 ();
 FILLCELL_X32 FILLER_87_1185 ();
 FILLCELL_X32 FILLER_87_1217 ();
 FILLCELL_X8 FILLER_87_1249 ();
 FILLCELL_X4 FILLER_87_1257 ();
 FILLCELL_X2 FILLER_87_1261 ();
 FILLCELL_X32 FILLER_87_1264 ();
 FILLCELL_X32 FILLER_87_1296 ();
 FILLCELL_X32 FILLER_87_1328 ();
 FILLCELL_X32 FILLER_87_1360 ();
 FILLCELL_X32 FILLER_87_1392 ();
 FILLCELL_X32 FILLER_87_1424 ();
 FILLCELL_X32 FILLER_87_1456 ();
 FILLCELL_X32 FILLER_87_1488 ();
 FILLCELL_X32 FILLER_87_1520 ();
 FILLCELL_X32 FILLER_87_1552 ();
 FILLCELL_X32 FILLER_87_1584 ();
 FILLCELL_X32 FILLER_87_1616 ();
 FILLCELL_X32 FILLER_87_1648 ();
 FILLCELL_X32 FILLER_87_1680 ();
 FILLCELL_X32 FILLER_87_1712 ();
 FILLCELL_X32 FILLER_87_1744 ();
 FILLCELL_X32 FILLER_87_1776 ();
 FILLCELL_X32 FILLER_87_1808 ();
 FILLCELL_X32 FILLER_87_1840 ();
 FILLCELL_X32 FILLER_87_1872 ();
 FILLCELL_X32 FILLER_87_1904 ();
 FILLCELL_X32 FILLER_87_1936 ();
 FILLCELL_X32 FILLER_87_1968 ();
 FILLCELL_X32 FILLER_87_2000 ();
 FILLCELL_X32 FILLER_87_2032 ();
 FILLCELL_X32 FILLER_87_2064 ();
 FILLCELL_X32 FILLER_87_2096 ();
 FILLCELL_X32 FILLER_87_2128 ();
 FILLCELL_X32 FILLER_87_2160 ();
 FILLCELL_X32 FILLER_87_2192 ();
 FILLCELL_X32 FILLER_87_2224 ();
 FILLCELL_X32 FILLER_87_2256 ();
 FILLCELL_X32 FILLER_87_2288 ();
 FILLCELL_X32 FILLER_87_2320 ();
 FILLCELL_X32 FILLER_87_2352 ();
 FILLCELL_X32 FILLER_87_2384 ();
 FILLCELL_X32 FILLER_87_2416 ();
 FILLCELL_X32 FILLER_87_2448 ();
 FILLCELL_X32 FILLER_87_2480 ();
 FILLCELL_X8 FILLER_87_2512 ();
 FILLCELL_X4 FILLER_87_2520 ();
 FILLCELL_X2 FILLER_87_2524 ();
 FILLCELL_X32 FILLER_87_2527 ();
 FILLCELL_X32 FILLER_87_2559 ();
 FILLCELL_X8 FILLER_87_2591 ();
 FILLCELL_X2 FILLER_87_2599 ();
 FILLCELL_X1 FILLER_87_2601 ();
 FILLCELL_X32 FILLER_88_1 ();
 FILLCELL_X32 FILLER_88_33 ();
 FILLCELL_X32 FILLER_88_65 ();
 FILLCELL_X32 FILLER_88_97 ();
 FILLCELL_X32 FILLER_88_129 ();
 FILLCELL_X32 FILLER_88_161 ();
 FILLCELL_X32 FILLER_88_193 ();
 FILLCELL_X32 FILLER_88_225 ();
 FILLCELL_X32 FILLER_88_257 ();
 FILLCELL_X32 FILLER_88_289 ();
 FILLCELL_X32 FILLER_88_321 ();
 FILLCELL_X32 FILLER_88_353 ();
 FILLCELL_X32 FILLER_88_385 ();
 FILLCELL_X32 FILLER_88_417 ();
 FILLCELL_X32 FILLER_88_449 ();
 FILLCELL_X32 FILLER_88_481 ();
 FILLCELL_X32 FILLER_88_513 ();
 FILLCELL_X32 FILLER_88_545 ();
 FILLCELL_X32 FILLER_88_577 ();
 FILLCELL_X16 FILLER_88_609 ();
 FILLCELL_X4 FILLER_88_625 ();
 FILLCELL_X2 FILLER_88_629 ();
 FILLCELL_X32 FILLER_88_632 ();
 FILLCELL_X32 FILLER_88_664 ();
 FILLCELL_X32 FILLER_88_696 ();
 FILLCELL_X32 FILLER_88_728 ();
 FILLCELL_X32 FILLER_88_760 ();
 FILLCELL_X32 FILLER_88_792 ();
 FILLCELL_X32 FILLER_88_824 ();
 FILLCELL_X32 FILLER_88_856 ();
 FILLCELL_X32 FILLER_88_888 ();
 FILLCELL_X32 FILLER_88_920 ();
 FILLCELL_X32 FILLER_88_952 ();
 FILLCELL_X32 FILLER_88_984 ();
 FILLCELL_X32 FILLER_88_1016 ();
 FILLCELL_X32 FILLER_88_1048 ();
 FILLCELL_X32 FILLER_88_1080 ();
 FILLCELL_X32 FILLER_88_1112 ();
 FILLCELL_X32 FILLER_88_1144 ();
 FILLCELL_X32 FILLER_88_1176 ();
 FILLCELL_X32 FILLER_88_1208 ();
 FILLCELL_X32 FILLER_88_1240 ();
 FILLCELL_X32 FILLER_88_1272 ();
 FILLCELL_X32 FILLER_88_1304 ();
 FILLCELL_X32 FILLER_88_1336 ();
 FILLCELL_X32 FILLER_88_1368 ();
 FILLCELL_X32 FILLER_88_1400 ();
 FILLCELL_X32 FILLER_88_1432 ();
 FILLCELL_X32 FILLER_88_1464 ();
 FILLCELL_X32 FILLER_88_1496 ();
 FILLCELL_X32 FILLER_88_1528 ();
 FILLCELL_X32 FILLER_88_1560 ();
 FILLCELL_X32 FILLER_88_1592 ();
 FILLCELL_X32 FILLER_88_1624 ();
 FILLCELL_X32 FILLER_88_1656 ();
 FILLCELL_X32 FILLER_88_1688 ();
 FILLCELL_X32 FILLER_88_1720 ();
 FILLCELL_X32 FILLER_88_1752 ();
 FILLCELL_X32 FILLER_88_1784 ();
 FILLCELL_X32 FILLER_88_1816 ();
 FILLCELL_X32 FILLER_88_1848 ();
 FILLCELL_X8 FILLER_88_1880 ();
 FILLCELL_X4 FILLER_88_1888 ();
 FILLCELL_X2 FILLER_88_1892 ();
 FILLCELL_X32 FILLER_88_1895 ();
 FILLCELL_X32 FILLER_88_1927 ();
 FILLCELL_X32 FILLER_88_1959 ();
 FILLCELL_X32 FILLER_88_1991 ();
 FILLCELL_X32 FILLER_88_2023 ();
 FILLCELL_X32 FILLER_88_2055 ();
 FILLCELL_X32 FILLER_88_2087 ();
 FILLCELL_X32 FILLER_88_2119 ();
 FILLCELL_X32 FILLER_88_2151 ();
 FILLCELL_X32 FILLER_88_2183 ();
 FILLCELL_X32 FILLER_88_2215 ();
 FILLCELL_X32 FILLER_88_2247 ();
 FILLCELL_X32 FILLER_88_2279 ();
 FILLCELL_X32 FILLER_88_2311 ();
 FILLCELL_X32 FILLER_88_2343 ();
 FILLCELL_X32 FILLER_88_2375 ();
 FILLCELL_X32 FILLER_88_2407 ();
 FILLCELL_X32 FILLER_88_2439 ();
 FILLCELL_X32 FILLER_88_2471 ();
 FILLCELL_X32 FILLER_88_2503 ();
 FILLCELL_X32 FILLER_88_2535 ();
 FILLCELL_X32 FILLER_88_2567 ();
 FILLCELL_X2 FILLER_88_2599 ();
 FILLCELL_X1 FILLER_88_2601 ();
 FILLCELL_X32 FILLER_89_1 ();
 FILLCELL_X32 FILLER_89_33 ();
 FILLCELL_X32 FILLER_89_65 ();
 FILLCELL_X32 FILLER_89_97 ();
 FILLCELL_X32 FILLER_89_129 ();
 FILLCELL_X32 FILLER_89_161 ();
 FILLCELL_X32 FILLER_89_193 ();
 FILLCELL_X32 FILLER_89_225 ();
 FILLCELL_X32 FILLER_89_257 ();
 FILLCELL_X32 FILLER_89_289 ();
 FILLCELL_X32 FILLER_89_321 ();
 FILLCELL_X32 FILLER_89_353 ();
 FILLCELL_X32 FILLER_89_385 ();
 FILLCELL_X32 FILLER_89_417 ();
 FILLCELL_X32 FILLER_89_449 ();
 FILLCELL_X32 FILLER_89_481 ();
 FILLCELL_X32 FILLER_89_513 ();
 FILLCELL_X32 FILLER_89_545 ();
 FILLCELL_X32 FILLER_89_577 ();
 FILLCELL_X32 FILLER_89_609 ();
 FILLCELL_X32 FILLER_89_641 ();
 FILLCELL_X32 FILLER_89_673 ();
 FILLCELL_X32 FILLER_89_705 ();
 FILLCELL_X32 FILLER_89_737 ();
 FILLCELL_X32 FILLER_89_769 ();
 FILLCELL_X32 FILLER_89_801 ();
 FILLCELL_X32 FILLER_89_833 ();
 FILLCELL_X32 FILLER_89_865 ();
 FILLCELL_X32 FILLER_89_897 ();
 FILLCELL_X32 FILLER_89_929 ();
 FILLCELL_X32 FILLER_89_961 ();
 FILLCELL_X32 FILLER_89_993 ();
 FILLCELL_X32 FILLER_89_1025 ();
 FILLCELL_X32 FILLER_89_1057 ();
 FILLCELL_X32 FILLER_89_1089 ();
 FILLCELL_X32 FILLER_89_1121 ();
 FILLCELL_X32 FILLER_89_1153 ();
 FILLCELL_X32 FILLER_89_1185 ();
 FILLCELL_X32 FILLER_89_1217 ();
 FILLCELL_X8 FILLER_89_1249 ();
 FILLCELL_X4 FILLER_89_1257 ();
 FILLCELL_X2 FILLER_89_1261 ();
 FILLCELL_X32 FILLER_89_1264 ();
 FILLCELL_X32 FILLER_89_1296 ();
 FILLCELL_X32 FILLER_89_1328 ();
 FILLCELL_X32 FILLER_89_1360 ();
 FILLCELL_X32 FILLER_89_1392 ();
 FILLCELL_X32 FILLER_89_1424 ();
 FILLCELL_X32 FILLER_89_1456 ();
 FILLCELL_X32 FILLER_89_1488 ();
 FILLCELL_X32 FILLER_89_1520 ();
 FILLCELL_X32 FILLER_89_1552 ();
 FILLCELL_X32 FILLER_89_1584 ();
 FILLCELL_X32 FILLER_89_1616 ();
 FILLCELL_X32 FILLER_89_1648 ();
 FILLCELL_X32 FILLER_89_1680 ();
 FILLCELL_X32 FILLER_89_1712 ();
 FILLCELL_X32 FILLER_89_1744 ();
 FILLCELL_X32 FILLER_89_1776 ();
 FILLCELL_X32 FILLER_89_1808 ();
 FILLCELL_X32 FILLER_89_1840 ();
 FILLCELL_X32 FILLER_89_1872 ();
 FILLCELL_X32 FILLER_89_1904 ();
 FILLCELL_X32 FILLER_89_1936 ();
 FILLCELL_X32 FILLER_89_1968 ();
 FILLCELL_X32 FILLER_89_2000 ();
 FILLCELL_X32 FILLER_89_2032 ();
 FILLCELL_X32 FILLER_89_2064 ();
 FILLCELL_X32 FILLER_89_2096 ();
 FILLCELL_X32 FILLER_89_2128 ();
 FILLCELL_X32 FILLER_89_2160 ();
 FILLCELL_X32 FILLER_89_2192 ();
 FILLCELL_X32 FILLER_89_2224 ();
 FILLCELL_X32 FILLER_89_2256 ();
 FILLCELL_X32 FILLER_89_2288 ();
 FILLCELL_X32 FILLER_89_2320 ();
 FILLCELL_X32 FILLER_89_2352 ();
 FILLCELL_X32 FILLER_89_2384 ();
 FILLCELL_X32 FILLER_89_2416 ();
 FILLCELL_X32 FILLER_89_2448 ();
 FILLCELL_X32 FILLER_89_2480 ();
 FILLCELL_X8 FILLER_89_2512 ();
 FILLCELL_X4 FILLER_89_2520 ();
 FILLCELL_X2 FILLER_89_2524 ();
 FILLCELL_X32 FILLER_89_2527 ();
 FILLCELL_X32 FILLER_89_2559 ();
 FILLCELL_X8 FILLER_89_2591 ();
 FILLCELL_X2 FILLER_89_2599 ();
 FILLCELL_X1 FILLER_89_2601 ();
 FILLCELL_X32 FILLER_90_1 ();
 FILLCELL_X32 FILLER_90_33 ();
 FILLCELL_X32 FILLER_90_65 ();
 FILLCELL_X32 FILLER_90_97 ();
 FILLCELL_X32 FILLER_90_129 ();
 FILLCELL_X32 FILLER_90_161 ();
 FILLCELL_X32 FILLER_90_193 ();
 FILLCELL_X32 FILLER_90_225 ();
 FILLCELL_X32 FILLER_90_257 ();
 FILLCELL_X32 FILLER_90_289 ();
 FILLCELL_X32 FILLER_90_321 ();
 FILLCELL_X32 FILLER_90_353 ();
 FILLCELL_X32 FILLER_90_385 ();
 FILLCELL_X32 FILLER_90_417 ();
 FILLCELL_X32 FILLER_90_449 ();
 FILLCELL_X32 FILLER_90_481 ();
 FILLCELL_X32 FILLER_90_513 ();
 FILLCELL_X32 FILLER_90_545 ();
 FILLCELL_X32 FILLER_90_577 ();
 FILLCELL_X16 FILLER_90_609 ();
 FILLCELL_X4 FILLER_90_625 ();
 FILLCELL_X2 FILLER_90_629 ();
 FILLCELL_X32 FILLER_90_632 ();
 FILLCELL_X32 FILLER_90_664 ();
 FILLCELL_X32 FILLER_90_696 ();
 FILLCELL_X32 FILLER_90_728 ();
 FILLCELL_X32 FILLER_90_760 ();
 FILLCELL_X32 FILLER_90_792 ();
 FILLCELL_X32 FILLER_90_824 ();
 FILLCELL_X32 FILLER_90_856 ();
 FILLCELL_X32 FILLER_90_888 ();
 FILLCELL_X32 FILLER_90_920 ();
 FILLCELL_X32 FILLER_90_952 ();
 FILLCELL_X32 FILLER_90_984 ();
 FILLCELL_X32 FILLER_90_1016 ();
 FILLCELL_X32 FILLER_90_1048 ();
 FILLCELL_X32 FILLER_90_1080 ();
 FILLCELL_X32 FILLER_90_1112 ();
 FILLCELL_X32 FILLER_90_1144 ();
 FILLCELL_X32 FILLER_90_1176 ();
 FILLCELL_X32 FILLER_90_1208 ();
 FILLCELL_X32 FILLER_90_1240 ();
 FILLCELL_X32 FILLER_90_1272 ();
 FILLCELL_X32 FILLER_90_1304 ();
 FILLCELL_X32 FILLER_90_1336 ();
 FILLCELL_X32 FILLER_90_1368 ();
 FILLCELL_X32 FILLER_90_1400 ();
 FILLCELL_X32 FILLER_90_1432 ();
 FILLCELL_X32 FILLER_90_1464 ();
 FILLCELL_X32 FILLER_90_1496 ();
 FILLCELL_X32 FILLER_90_1528 ();
 FILLCELL_X32 FILLER_90_1560 ();
 FILLCELL_X32 FILLER_90_1592 ();
 FILLCELL_X32 FILLER_90_1624 ();
 FILLCELL_X32 FILLER_90_1656 ();
 FILLCELL_X32 FILLER_90_1688 ();
 FILLCELL_X32 FILLER_90_1720 ();
 FILLCELL_X32 FILLER_90_1752 ();
 FILLCELL_X32 FILLER_90_1784 ();
 FILLCELL_X32 FILLER_90_1816 ();
 FILLCELL_X32 FILLER_90_1848 ();
 FILLCELL_X8 FILLER_90_1880 ();
 FILLCELL_X4 FILLER_90_1888 ();
 FILLCELL_X2 FILLER_90_1892 ();
 FILLCELL_X32 FILLER_90_1895 ();
 FILLCELL_X32 FILLER_90_1927 ();
 FILLCELL_X32 FILLER_90_1959 ();
 FILLCELL_X32 FILLER_90_1991 ();
 FILLCELL_X32 FILLER_90_2023 ();
 FILLCELL_X32 FILLER_90_2055 ();
 FILLCELL_X32 FILLER_90_2087 ();
 FILLCELL_X32 FILLER_90_2119 ();
 FILLCELL_X32 FILLER_90_2151 ();
 FILLCELL_X32 FILLER_90_2183 ();
 FILLCELL_X32 FILLER_90_2215 ();
 FILLCELL_X32 FILLER_90_2247 ();
 FILLCELL_X32 FILLER_90_2279 ();
 FILLCELL_X32 FILLER_90_2311 ();
 FILLCELL_X32 FILLER_90_2343 ();
 FILLCELL_X32 FILLER_90_2375 ();
 FILLCELL_X32 FILLER_90_2407 ();
 FILLCELL_X32 FILLER_90_2439 ();
 FILLCELL_X32 FILLER_90_2471 ();
 FILLCELL_X32 FILLER_90_2503 ();
 FILLCELL_X32 FILLER_90_2535 ();
 FILLCELL_X32 FILLER_90_2567 ();
 FILLCELL_X2 FILLER_90_2599 ();
 FILLCELL_X1 FILLER_90_2601 ();
 FILLCELL_X32 FILLER_91_1 ();
 FILLCELL_X32 FILLER_91_33 ();
 FILLCELL_X32 FILLER_91_65 ();
 FILLCELL_X32 FILLER_91_97 ();
 FILLCELL_X32 FILLER_91_129 ();
 FILLCELL_X32 FILLER_91_161 ();
 FILLCELL_X32 FILLER_91_193 ();
 FILLCELL_X32 FILLER_91_225 ();
 FILLCELL_X32 FILLER_91_257 ();
 FILLCELL_X32 FILLER_91_289 ();
 FILLCELL_X32 FILLER_91_321 ();
 FILLCELL_X32 FILLER_91_353 ();
 FILLCELL_X32 FILLER_91_385 ();
 FILLCELL_X32 FILLER_91_417 ();
 FILLCELL_X32 FILLER_91_449 ();
 FILLCELL_X32 FILLER_91_481 ();
 FILLCELL_X32 FILLER_91_513 ();
 FILLCELL_X32 FILLER_91_545 ();
 FILLCELL_X32 FILLER_91_577 ();
 FILLCELL_X32 FILLER_91_609 ();
 FILLCELL_X32 FILLER_91_641 ();
 FILLCELL_X32 FILLER_91_673 ();
 FILLCELL_X32 FILLER_91_705 ();
 FILLCELL_X32 FILLER_91_737 ();
 FILLCELL_X32 FILLER_91_769 ();
 FILLCELL_X32 FILLER_91_801 ();
 FILLCELL_X32 FILLER_91_833 ();
 FILLCELL_X32 FILLER_91_865 ();
 FILLCELL_X32 FILLER_91_897 ();
 FILLCELL_X32 FILLER_91_929 ();
 FILLCELL_X32 FILLER_91_961 ();
 FILLCELL_X32 FILLER_91_993 ();
 FILLCELL_X32 FILLER_91_1025 ();
 FILLCELL_X32 FILLER_91_1057 ();
 FILLCELL_X32 FILLER_91_1089 ();
 FILLCELL_X32 FILLER_91_1121 ();
 FILLCELL_X32 FILLER_91_1153 ();
 FILLCELL_X32 FILLER_91_1185 ();
 FILLCELL_X32 FILLER_91_1217 ();
 FILLCELL_X8 FILLER_91_1249 ();
 FILLCELL_X4 FILLER_91_1257 ();
 FILLCELL_X2 FILLER_91_1261 ();
 FILLCELL_X32 FILLER_91_1264 ();
 FILLCELL_X32 FILLER_91_1296 ();
 FILLCELL_X32 FILLER_91_1328 ();
 FILLCELL_X32 FILLER_91_1360 ();
 FILLCELL_X32 FILLER_91_1392 ();
 FILLCELL_X32 FILLER_91_1424 ();
 FILLCELL_X32 FILLER_91_1456 ();
 FILLCELL_X32 FILLER_91_1488 ();
 FILLCELL_X32 FILLER_91_1520 ();
 FILLCELL_X32 FILLER_91_1552 ();
 FILLCELL_X32 FILLER_91_1584 ();
 FILLCELL_X32 FILLER_91_1616 ();
 FILLCELL_X32 FILLER_91_1648 ();
 FILLCELL_X32 FILLER_91_1680 ();
 FILLCELL_X32 FILLER_91_1712 ();
 FILLCELL_X32 FILLER_91_1744 ();
 FILLCELL_X32 FILLER_91_1776 ();
 FILLCELL_X32 FILLER_91_1808 ();
 FILLCELL_X32 FILLER_91_1840 ();
 FILLCELL_X32 FILLER_91_1872 ();
 FILLCELL_X32 FILLER_91_1904 ();
 FILLCELL_X32 FILLER_91_1936 ();
 FILLCELL_X32 FILLER_91_1968 ();
 FILLCELL_X32 FILLER_91_2000 ();
 FILLCELL_X32 FILLER_91_2032 ();
 FILLCELL_X32 FILLER_91_2064 ();
 FILLCELL_X32 FILLER_91_2096 ();
 FILLCELL_X32 FILLER_91_2128 ();
 FILLCELL_X32 FILLER_91_2160 ();
 FILLCELL_X32 FILLER_91_2192 ();
 FILLCELL_X32 FILLER_91_2224 ();
 FILLCELL_X32 FILLER_91_2256 ();
 FILLCELL_X32 FILLER_91_2288 ();
 FILLCELL_X32 FILLER_91_2320 ();
 FILLCELL_X32 FILLER_91_2352 ();
 FILLCELL_X32 FILLER_91_2384 ();
 FILLCELL_X32 FILLER_91_2416 ();
 FILLCELL_X32 FILLER_91_2448 ();
 FILLCELL_X32 FILLER_91_2480 ();
 FILLCELL_X8 FILLER_91_2512 ();
 FILLCELL_X4 FILLER_91_2520 ();
 FILLCELL_X2 FILLER_91_2524 ();
 FILLCELL_X32 FILLER_91_2527 ();
 FILLCELL_X32 FILLER_91_2559 ();
 FILLCELL_X8 FILLER_91_2591 ();
 FILLCELL_X2 FILLER_91_2599 ();
 FILLCELL_X1 FILLER_91_2601 ();
 FILLCELL_X32 FILLER_92_1 ();
 FILLCELL_X32 FILLER_92_33 ();
 FILLCELL_X32 FILLER_92_65 ();
 FILLCELL_X32 FILLER_92_97 ();
 FILLCELL_X32 FILLER_92_129 ();
 FILLCELL_X32 FILLER_92_161 ();
 FILLCELL_X32 FILLER_92_193 ();
 FILLCELL_X32 FILLER_92_225 ();
 FILLCELL_X32 FILLER_92_257 ();
 FILLCELL_X32 FILLER_92_289 ();
 FILLCELL_X32 FILLER_92_321 ();
 FILLCELL_X32 FILLER_92_353 ();
 FILLCELL_X32 FILLER_92_385 ();
 FILLCELL_X32 FILLER_92_417 ();
 FILLCELL_X32 FILLER_92_449 ();
 FILLCELL_X32 FILLER_92_481 ();
 FILLCELL_X32 FILLER_92_513 ();
 FILLCELL_X32 FILLER_92_545 ();
 FILLCELL_X32 FILLER_92_577 ();
 FILLCELL_X16 FILLER_92_609 ();
 FILLCELL_X4 FILLER_92_625 ();
 FILLCELL_X2 FILLER_92_629 ();
 FILLCELL_X32 FILLER_92_632 ();
 FILLCELL_X32 FILLER_92_664 ();
 FILLCELL_X32 FILLER_92_696 ();
 FILLCELL_X32 FILLER_92_728 ();
 FILLCELL_X32 FILLER_92_760 ();
 FILLCELL_X32 FILLER_92_792 ();
 FILLCELL_X32 FILLER_92_824 ();
 FILLCELL_X32 FILLER_92_856 ();
 FILLCELL_X32 FILLER_92_888 ();
 FILLCELL_X32 FILLER_92_920 ();
 FILLCELL_X32 FILLER_92_952 ();
 FILLCELL_X32 FILLER_92_984 ();
 FILLCELL_X32 FILLER_92_1016 ();
 FILLCELL_X32 FILLER_92_1048 ();
 FILLCELL_X32 FILLER_92_1080 ();
 FILLCELL_X32 FILLER_92_1112 ();
 FILLCELL_X32 FILLER_92_1144 ();
 FILLCELL_X32 FILLER_92_1176 ();
 FILLCELL_X32 FILLER_92_1208 ();
 FILLCELL_X32 FILLER_92_1240 ();
 FILLCELL_X32 FILLER_92_1272 ();
 FILLCELL_X32 FILLER_92_1304 ();
 FILLCELL_X32 FILLER_92_1336 ();
 FILLCELL_X32 FILLER_92_1368 ();
 FILLCELL_X32 FILLER_92_1400 ();
 FILLCELL_X32 FILLER_92_1432 ();
 FILLCELL_X32 FILLER_92_1464 ();
 FILLCELL_X32 FILLER_92_1496 ();
 FILLCELL_X32 FILLER_92_1528 ();
 FILLCELL_X32 FILLER_92_1560 ();
 FILLCELL_X32 FILLER_92_1592 ();
 FILLCELL_X32 FILLER_92_1624 ();
 FILLCELL_X32 FILLER_92_1656 ();
 FILLCELL_X32 FILLER_92_1688 ();
 FILLCELL_X32 FILLER_92_1720 ();
 FILLCELL_X32 FILLER_92_1752 ();
 FILLCELL_X32 FILLER_92_1784 ();
 FILLCELL_X32 FILLER_92_1816 ();
 FILLCELL_X32 FILLER_92_1848 ();
 FILLCELL_X8 FILLER_92_1880 ();
 FILLCELL_X4 FILLER_92_1888 ();
 FILLCELL_X2 FILLER_92_1892 ();
 FILLCELL_X32 FILLER_92_1895 ();
 FILLCELL_X32 FILLER_92_1927 ();
 FILLCELL_X32 FILLER_92_1959 ();
 FILLCELL_X32 FILLER_92_1991 ();
 FILLCELL_X32 FILLER_92_2023 ();
 FILLCELL_X32 FILLER_92_2055 ();
 FILLCELL_X32 FILLER_92_2087 ();
 FILLCELL_X32 FILLER_92_2119 ();
 FILLCELL_X32 FILLER_92_2151 ();
 FILLCELL_X32 FILLER_92_2183 ();
 FILLCELL_X32 FILLER_92_2215 ();
 FILLCELL_X32 FILLER_92_2247 ();
 FILLCELL_X32 FILLER_92_2279 ();
 FILLCELL_X32 FILLER_92_2311 ();
 FILLCELL_X32 FILLER_92_2343 ();
 FILLCELL_X32 FILLER_92_2375 ();
 FILLCELL_X32 FILLER_92_2407 ();
 FILLCELL_X32 FILLER_92_2439 ();
 FILLCELL_X32 FILLER_92_2471 ();
 FILLCELL_X32 FILLER_92_2503 ();
 FILLCELL_X32 FILLER_92_2535 ();
 FILLCELL_X32 FILLER_92_2567 ();
 FILLCELL_X2 FILLER_92_2599 ();
 FILLCELL_X1 FILLER_92_2601 ();
 FILLCELL_X32 FILLER_93_1 ();
 FILLCELL_X32 FILLER_93_33 ();
 FILLCELL_X32 FILLER_93_65 ();
 FILLCELL_X32 FILLER_93_97 ();
 FILLCELL_X32 FILLER_93_129 ();
 FILLCELL_X32 FILLER_93_161 ();
 FILLCELL_X32 FILLER_93_193 ();
 FILLCELL_X32 FILLER_93_225 ();
 FILLCELL_X32 FILLER_93_257 ();
 FILLCELL_X32 FILLER_93_289 ();
 FILLCELL_X32 FILLER_93_321 ();
 FILLCELL_X32 FILLER_93_353 ();
 FILLCELL_X32 FILLER_93_385 ();
 FILLCELL_X32 FILLER_93_417 ();
 FILLCELL_X32 FILLER_93_449 ();
 FILLCELL_X32 FILLER_93_481 ();
 FILLCELL_X32 FILLER_93_513 ();
 FILLCELL_X32 FILLER_93_545 ();
 FILLCELL_X32 FILLER_93_577 ();
 FILLCELL_X32 FILLER_93_609 ();
 FILLCELL_X32 FILLER_93_641 ();
 FILLCELL_X32 FILLER_93_673 ();
 FILLCELL_X32 FILLER_93_705 ();
 FILLCELL_X32 FILLER_93_737 ();
 FILLCELL_X32 FILLER_93_769 ();
 FILLCELL_X32 FILLER_93_801 ();
 FILLCELL_X32 FILLER_93_833 ();
 FILLCELL_X32 FILLER_93_865 ();
 FILLCELL_X32 FILLER_93_897 ();
 FILLCELL_X32 FILLER_93_929 ();
 FILLCELL_X32 FILLER_93_961 ();
 FILLCELL_X32 FILLER_93_993 ();
 FILLCELL_X32 FILLER_93_1025 ();
 FILLCELL_X32 FILLER_93_1057 ();
 FILLCELL_X32 FILLER_93_1089 ();
 FILLCELL_X32 FILLER_93_1121 ();
 FILLCELL_X32 FILLER_93_1153 ();
 FILLCELL_X32 FILLER_93_1185 ();
 FILLCELL_X32 FILLER_93_1217 ();
 FILLCELL_X8 FILLER_93_1249 ();
 FILLCELL_X4 FILLER_93_1257 ();
 FILLCELL_X2 FILLER_93_1261 ();
 FILLCELL_X32 FILLER_93_1264 ();
 FILLCELL_X32 FILLER_93_1296 ();
 FILLCELL_X32 FILLER_93_1328 ();
 FILLCELL_X32 FILLER_93_1360 ();
 FILLCELL_X32 FILLER_93_1392 ();
 FILLCELL_X32 FILLER_93_1424 ();
 FILLCELL_X32 FILLER_93_1456 ();
 FILLCELL_X32 FILLER_93_1488 ();
 FILLCELL_X32 FILLER_93_1520 ();
 FILLCELL_X32 FILLER_93_1552 ();
 FILLCELL_X32 FILLER_93_1584 ();
 FILLCELL_X32 FILLER_93_1616 ();
 FILLCELL_X32 FILLER_93_1648 ();
 FILLCELL_X32 FILLER_93_1680 ();
 FILLCELL_X32 FILLER_93_1712 ();
 FILLCELL_X32 FILLER_93_1744 ();
 FILLCELL_X32 FILLER_93_1776 ();
 FILLCELL_X32 FILLER_93_1808 ();
 FILLCELL_X32 FILLER_93_1840 ();
 FILLCELL_X32 FILLER_93_1872 ();
 FILLCELL_X32 FILLER_93_1904 ();
 FILLCELL_X32 FILLER_93_1936 ();
 FILLCELL_X32 FILLER_93_1968 ();
 FILLCELL_X32 FILLER_93_2000 ();
 FILLCELL_X32 FILLER_93_2032 ();
 FILLCELL_X32 FILLER_93_2064 ();
 FILLCELL_X32 FILLER_93_2096 ();
 FILLCELL_X32 FILLER_93_2128 ();
 FILLCELL_X32 FILLER_93_2160 ();
 FILLCELL_X32 FILLER_93_2192 ();
 FILLCELL_X32 FILLER_93_2224 ();
 FILLCELL_X32 FILLER_93_2256 ();
 FILLCELL_X32 FILLER_93_2288 ();
 FILLCELL_X32 FILLER_93_2320 ();
 FILLCELL_X32 FILLER_93_2352 ();
 FILLCELL_X32 FILLER_93_2384 ();
 FILLCELL_X32 FILLER_93_2416 ();
 FILLCELL_X32 FILLER_93_2448 ();
 FILLCELL_X32 FILLER_93_2480 ();
 FILLCELL_X8 FILLER_93_2512 ();
 FILLCELL_X4 FILLER_93_2520 ();
 FILLCELL_X2 FILLER_93_2524 ();
 FILLCELL_X32 FILLER_93_2527 ();
 FILLCELL_X32 FILLER_93_2559 ();
 FILLCELL_X8 FILLER_93_2591 ();
 FILLCELL_X2 FILLER_93_2599 ();
 FILLCELL_X1 FILLER_93_2601 ();
 FILLCELL_X32 FILLER_94_1 ();
 FILLCELL_X32 FILLER_94_33 ();
 FILLCELL_X32 FILLER_94_65 ();
 FILLCELL_X32 FILLER_94_97 ();
 FILLCELL_X32 FILLER_94_129 ();
 FILLCELL_X32 FILLER_94_161 ();
 FILLCELL_X32 FILLER_94_193 ();
 FILLCELL_X32 FILLER_94_225 ();
 FILLCELL_X32 FILLER_94_257 ();
 FILLCELL_X32 FILLER_94_289 ();
 FILLCELL_X32 FILLER_94_321 ();
 FILLCELL_X32 FILLER_94_353 ();
 FILLCELL_X32 FILLER_94_385 ();
 FILLCELL_X32 FILLER_94_417 ();
 FILLCELL_X32 FILLER_94_449 ();
 FILLCELL_X32 FILLER_94_481 ();
 FILLCELL_X32 FILLER_94_513 ();
 FILLCELL_X32 FILLER_94_545 ();
 FILLCELL_X32 FILLER_94_577 ();
 FILLCELL_X16 FILLER_94_609 ();
 FILLCELL_X4 FILLER_94_625 ();
 FILLCELL_X2 FILLER_94_629 ();
 FILLCELL_X32 FILLER_94_632 ();
 FILLCELL_X32 FILLER_94_664 ();
 FILLCELL_X32 FILLER_94_696 ();
 FILLCELL_X32 FILLER_94_728 ();
 FILLCELL_X32 FILLER_94_760 ();
 FILLCELL_X32 FILLER_94_792 ();
 FILLCELL_X32 FILLER_94_824 ();
 FILLCELL_X32 FILLER_94_856 ();
 FILLCELL_X32 FILLER_94_888 ();
 FILLCELL_X32 FILLER_94_920 ();
 FILLCELL_X32 FILLER_94_952 ();
 FILLCELL_X32 FILLER_94_984 ();
 FILLCELL_X32 FILLER_94_1016 ();
 FILLCELL_X32 FILLER_94_1048 ();
 FILLCELL_X32 FILLER_94_1080 ();
 FILLCELL_X32 FILLER_94_1112 ();
 FILLCELL_X32 FILLER_94_1144 ();
 FILLCELL_X32 FILLER_94_1176 ();
 FILLCELL_X32 FILLER_94_1208 ();
 FILLCELL_X32 FILLER_94_1240 ();
 FILLCELL_X32 FILLER_94_1272 ();
 FILLCELL_X32 FILLER_94_1304 ();
 FILLCELL_X32 FILLER_94_1336 ();
 FILLCELL_X32 FILLER_94_1368 ();
 FILLCELL_X32 FILLER_94_1400 ();
 FILLCELL_X32 FILLER_94_1432 ();
 FILLCELL_X32 FILLER_94_1464 ();
 FILLCELL_X32 FILLER_94_1496 ();
 FILLCELL_X32 FILLER_94_1528 ();
 FILLCELL_X32 FILLER_94_1560 ();
 FILLCELL_X32 FILLER_94_1592 ();
 FILLCELL_X32 FILLER_94_1624 ();
 FILLCELL_X32 FILLER_94_1656 ();
 FILLCELL_X32 FILLER_94_1688 ();
 FILLCELL_X32 FILLER_94_1720 ();
 FILLCELL_X32 FILLER_94_1752 ();
 FILLCELL_X32 FILLER_94_1784 ();
 FILLCELL_X32 FILLER_94_1816 ();
 FILLCELL_X32 FILLER_94_1848 ();
 FILLCELL_X8 FILLER_94_1880 ();
 FILLCELL_X4 FILLER_94_1888 ();
 FILLCELL_X2 FILLER_94_1892 ();
 FILLCELL_X32 FILLER_94_1895 ();
 FILLCELL_X32 FILLER_94_1927 ();
 FILLCELL_X32 FILLER_94_1959 ();
 FILLCELL_X32 FILLER_94_1991 ();
 FILLCELL_X32 FILLER_94_2023 ();
 FILLCELL_X32 FILLER_94_2055 ();
 FILLCELL_X32 FILLER_94_2087 ();
 FILLCELL_X32 FILLER_94_2119 ();
 FILLCELL_X32 FILLER_94_2151 ();
 FILLCELL_X32 FILLER_94_2183 ();
 FILLCELL_X32 FILLER_94_2215 ();
 FILLCELL_X32 FILLER_94_2247 ();
 FILLCELL_X32 FILLER_94_2279 ();
 FILLCELL_X32 FILLER_94_2311 ();
 FILLCELL_X32 FILLER_94_2343 ();
 FILLCELL_X32 FILLER_94_2375 ();
 FILLCELL_X32 FILLER_94_2407 ();
 FILLCELL_X32 FILLER_94_2439 ();
 FILLCELL_X32 FILLER_94_2471 ();
 FILLCELL_X32 FILLER_94_2503 ();
 FILLCELL_X32 FILLER_94_2535 ();
 FILLCELL_X32 FILLER_94_2567 ();
 FILLCELL_X2 FILLER_94_2599 ();
 FILLCELL_X1 FILLER_94_2601 ();
 FILLCELL_X32 FILLER_95_1 ();
 FILLCELL_X32 FILLER_95_33 ();
 FILLCELL_X32 FILLER_95_65 ();
 FILLCELL_X32 FILLER_95_97 ();
 FILLCELL_X32 FILLER_95_129 ();
 FILLCELL_X32 FILLER_95_161 ();
 FILLCELL_X32 FILLER_95_193 ();
 FILLCELL_X32 FILLER_95_225 ();
 FILLCELL_X32 FILLER_95_257 ();
 FILLCELL_X32 FILLER_95_289 ();
 FILLCELL_X32 FILLER_95_321 ();
 FILLCELL_X32 FILLER_95_353 ();
 FILLCELL_X32 FILLER_95_385 ();
 FILLCELL_X32 FILLER_95_417 ();
 FILLCELL_X32 FILLER_95_449 ();
 FILLCELL_X32 FILLER_95_481 ();
 FILLCELL_X32 FILLER_95_513 ();
 FILLCELL_X32 FILLER_95_545 ();
 FILLCELL_X32 FILLER_95_577 ();
 FILLCELL_X32 FILLER_95_609 ();
 FILLCELL_X32 FILLER_95_641 ();
 FILLCELL_X32 FILLER_95_673 ();
 FILLCELL_X32 FILLER_95_705 ();
 FILLCELL_X32 FILLER_95_737 ();
 FILLCELL_X32 FILLER_95_769 ();
 FILLCELL_X32 FILLER_95_801 ();
 FILLCELL_X32 FILLER_95_833 ();
 FILLCELL_X32 FILLER_95_865 ();
 FILLCELL_X32 FILLER_95_897 ();
 FILLCELL_X32 FILLER_95_929 ();
 FILLCELL_X32 FILLER_95_961 ();
 FILLCELL_X32 FILLER_95_993 ();
 FILLCELL_X32 FILLER_95_1025 ();
 FILLCELL_X32 FILLER_95_1057 ();
 FILLCELL_X32 FILLER_95_1089 ();
 FILLCELL_X32 FILLER_95_1121 ();
 FILLCELL_X32 FILLER_95_1153 ();
 FILLCELL_X32 FILLER_95_1185 ();
 FILLCELL_X32 FILLER_95_1217 ();
 FILLCELL_X8 FILLER_95_1249 ();
 FILLCELL_X4 FILLER_95_1257 ();
 FILLCELL_X2 FILLER_95_1261 ();
 FILLCELL_X32 FILLER_95_1264 ();
 FILLCELL_X32 FILLER_95_1296 ();
 FILLCELL_X32 FILLER_95_1328 ();
 FILLCELL_X32 FILLER_95_1360 ();
 FILLCELL_X32 FILLER_95_1392 ();
 FILLCELL_X32 FILLER_95_1424 ();
 FILLCELL_X32 FILLER_95_1456 ();
 FILLCELL_X32 FILLER_95_1488 ();
 FILLCELL_X32 FILLER_95_1520 ();
 FILLCELL_X32 FILLER_95_1552 ();
 FILLCELL_X32 FILLER_95_1584 ();
 FILLCELL_X32 FILLER_95_1616 ();
 FILLCELL_X32 FILLER_95_1648 ();
 FILLCELL_X32 FILLER_95_1680 ();
 FILLCELL_X32 FILLER_95_1712 ();
 FILLCELL_X32 FILLER_95_1744 ();
 FILLCELL_X32 FILLER_95_1776 ();
 FILLCELL_X32 FILLER_95_1808 ();
 FILLCELL_X32 FILLER_95_1840 ();
 FILLCELL_X32 FILLER_95_1872 ();
 FILLCELL_X32 FILLER_95_1904 ();
 FILLCELL_X32 FILLER_95_1936 ();
 FILLCELL_X32 FILLER_95_1968 ();
 FILLCELL_X32 FILLER_95_2000 ();
 FILLCELL_X32 FILLER_95_2032 ();
 FILLCELL_X32 FILLER_95_2064 ();
 FILLCELL_X32 FILLER_95_2096 ();
 FILLCELL_X32 FILLER_95_2128 ();
 FILLCELL_X32 FILLER_95_2160 ();
 FILLCELL_X32 FILLER_95_2192 ();
 FILLCELL_X32 FILLER_95_2224 ();
 FILLCELL_X32 FILLER_95_2256 ();
 FILLCELL_X32 FILLER_95_2288 ();
 FILLCELL_X32 FILLER_95_2320 ();
 FILLCELL_X32 FILLER_95_2352 ();
 FILLCELL_X32 FILLER_95_2384 ();
 FILLCELL_X32 FILLER_95_2416 ();
 FILLCELL_X32 FILLER_95_2448 ();
 FILLCELL_X32 FILLER_95_2480 ();
 FILLCELL_X8 FILLER_95_2512 ();
 FILLCELL_X4 FILLER_95_2520 ();
 FILLCELL_X2 FILLER_95_2524 ();
 FILLCELL_X32 FILLER_95_2527 ();
 FILLCELL_X32 FILLER_95_2559 ();
 FILLCELL_X8 FILLER_95_2591 ();
 FILLCELL_X2 FILLER_95_2599 ();
 FILLCELL_X1 FILLER_95_2601 ();
 FILLCELL_X32 FILLER_96_1 ();
 FILLCELL_X32 FILLER_96_33 ();
 FILLCELL_X32 FILLER_96_65 ();
 FILLCELL_X32 FILLER_96_97 ();
 FILLCELL_X32 FILLER_96_129 ();
 FILLCELL_X32 FILLER_96_161 ();
 FILLCELL_X32 FILLER_96_193 ();
 FILLCELL_X32 FILLER_96_225 ();
 FILLCELL_X32 FILLER_96_257 ();
 FILLCELL_X32 FILLER_96_289 ();
 FILLCELL_X32 FILLER_96_321 ();
 FILLCELL_X32 FILLER_96_353 ();
 FILLCELL_X32 FILLER_96_385 ();
 FILLCELL_X32 FILLER_96_417 ();
 FILLCELL_X32 FILLER_96_449 ();
 FILLCELL_X32 FILLER_96_481 ();
 FILLCELL_X32 FILLER_96_513 ();
 FILLCELL_X32 FILLER_96_545 ();
 FILLCELL_X32 FILLER_96_577 ();
 FILLCELL_X16 FILLER_96_609 ();
 FILLCELL_X4 FILLER_96_625 ();
 FILLCELL_X2 FILLER_96_629 ();
 FILLCELL_X32 FILLER_96_632 ();
 FILLCELL_X32 FILLER_96_664 ();
 FILLCELL_X32 FILLER_96_696 ();
 FILLCELL_X32 FILLER_96_728 ();
 FILLCELL_X32 FILLER_96_760 ();
 FILLCELL_X32 FILLER_96_792 ();
 FILLCELL_X32 FILLER_96_824 ();
 FILLCELL_X32 FILLER_96_856 ();
 FILLCELL_X32 FILLER_96_888 ();
 FILLCELL_X32 FILLER_96_920 ();
 FILLCELL_X32 FILLER_96_952 ();
 FILLCELL_X32 FILLER_96_984 ();
 FILLCELL_X32 FILLER_96_1016 ();
 FILLCELL_X32 FILLER_96_1048 ();
 FILLCELL_X32 FILLER_96_1080 ();
 FILLCELL_X32 FILLER_96_1112 ();
 FILLCELL_X32 FILLER_96_1144 ();
 FILLCELL_X32 FILLER_96_1176 ();
 FILLCELL_X32 FILLER_96_1208 ();
 FILLCELL_X32 FILLER_96_1240 ();
 FILLCELL_X32 FILLER_96_1272 ();
 FILLCELL_X32 FILLER_96_1304 ();
 FILLCELL_X32 FILLER_96_1336 ();
 FILLCELL_X32 FILLER_96_1368 ();
 FILLCELL_X32 FILLER_96_1400 ();
 FILLCELL_X32 FILLER_96_1432 ();
 FILLCELL_X32 FILLER_96_1464 ();
 FILLCELL_X32 FILLER_96_1496 ();
 FILLCELL_X32 FILLER_96_1528 ();
 FILLCELL_X32 FILLER_96_1560 ();
 FILLCELL_X32 FILLER_96_1592 ();
 FILLCELL_X32 FILLER_96_1624 ();
 FILLCELL_X32 FILLER_96_1656 ();
 FILLCELL_X32 FILLER_96_1688 ();
 FILLCELL_X32 FILLER_96_1720 ();
 FILLCELL_X32 FILLER_96_1752 ();
 FILLCELL_X32 FILLER_96_1784 ();
 FILLCELL_X32 FILLER_96_1816 ();
 FILLCELL_X32 FILLER_96_1848 ();
 FILLCELL_X8 FILLER_96_1880 ();
 FILLCELL_X4 FILLER_96_1888 ();
 FILLCELL_X2 FILLER_96_1892 ();
 FILLCELL_X32 FILLER_96_1895 ();
 FILLCELL_X32 FILLER_96_1927 ();
 FILLCELL_X32 FILLER_96_1959 ();
 FILLCELL_X32 FILLER_96_1991 ();
 FILLCELL_X32 FILLER_96_2023 ();
 FILLCELL_X32 FILLER_96_2055 ();
 FILLCELL_X32 FILLER_96_2087 ();
 FILLCELL_X32 FILLER_96_2119 ();
 FILLCELL_X32 FILLER_96_2151 ();
 FILLCELL_X32 FILLER_96_2183 ();
 FILLCELL_X32 FILLER_96_2215 ();
 FILLCELL_X32 FILLER_96_2247 ();
 FILLCELL_X32 FILLER_96_2279 ();
 FILLCELL_X32 FILLER_96_2311 ();
 FILLCELL_X32 FILLER_96_2343 ();
 FILLCELL_X32 FILLER_96_2375 ();
 FILLCELL_X32 FILLER_96_2407 ();
 FILLCELL_X32 FILLER_96_2439 ();
 FILLCELL_X32 FILLER_96_2471 ();
 FILLCELL_X32 FILLER_96_2503 ();
 FILLCELL_X32 FILLER_96_2535 ();
 FILLCELL_X32 FILLER_96_2567 ();
 FILLCELL_X2 FILLER_96_2599 ();
 FILLCELL_X1 FILLER_96_2601 ();
 FILLCELL_X32 FILLER_97_1 ();
 FILLCELL_X32 FILLER_97_33 ();
 FILLCELL_X32 FILLER_97_65 ();
 FILLCELL_X32 FILLER_97_97 ();
 FILLCELL_X32 FILLER_97_129 ();
 FILLCELL_X32 FILLER_97_161 ();
 FILLCELL_X32 FILLER_97_193 ();
 FILLCELL_X32 FILLER_97_225 ();
 FILLCELL_X32 FILLER_97_257 ();
 FILLCELL_X32 FILLER_97_289 ();
 FILLCELL_X32 FILLER_97_321 ();
 FILLCELL_X32 FILLER_97_353 ();
 FILLCELL_X32 FILLER_97_385 ();
 FILLCELL_X32 FILLER_97_417 ();
 FILLCELL_X32 FILLER_97_449 ();
 FILLCELL_X32 FILLER_97_481 ();
 FILLCELL_X32 FILLER_97_513 ();
 FILLCELL_X32 FILLER_97_545 ();
 FILLCELL_X32 FILLER_97_577 ();
 FILLCELL_X32 FILLER_97_609 ();
 FILLCELL_X32 FILLER_97_641 ();
 FILLCELL_X32 FILLER_97_673 ();
 FILLCELL_X32 FILLER_97_705 ();
 FILLCELL_X32 FILLER_97_737 ();
 FILLCELL_X32 FILLER_97_769 ();
 FILLCELL_X32 FILLER_97_801 ();
 FILLCELL_X32 FILLER_97_833 ();
 FILLCELL_X32 FILLER_97_865 ();
 FILLCELL_X32 FILLER_97_897 ();
 FILLCELL_X32 FILLER_97_929 ();
 FILLCELL_X32 FILLER_97_961 ();
 FILLCELL_X32 FILLER_97_993 ();
 FILLCELL_X32 FILLER_97_1025 ();
 FILLCELL_X32 FILLER_97_1057 ();
 FILLCELL_X32 FILLER_97_1089 ();
 FILLCELL_X32 FILLER_97_1121 ();
 FILLCELL_X32 FILLER_97_1153 ();
 FILLCELL_X32 FILLER_97_1185 ();
 FILLCELL_X32 FILLER_97_1217 ();
 FILLCELL_X8 FILLER_97_1249 ();
 FILLCELL_X4 FILLER_97_1257 ();
 FILLCELL_X2 FILLER_97_1261 ();
 FILLCELL_X32 FILLER_97_1264 ();
 FILLCELL_X32 FILLER_97_1296 ();
 FILLCELL_X32 FILLER_97_1328 ();
 FILLCELL_X32 FILLER_97_1360 ();
 FILLCELL_X32 FILLER_97_1392 ();
 FILLCELL_X32 FILLER_97_1424 ();
 FILLCELL_X32 FILLER_97_1456 ();
 FILLCELL_X32 FILLER_97_1488 ();
 FILLCELL_X32 FILLER_97_1520 ();
 FILLCELL_X32 FILLER_97_1552 ();
 FILLCELL_X32 FILLER_97_1584 ();
 FILLCELL_X32 FILLER_97_1616 ();
 FILLCELL_X32 FILLER_97_1648 ();
 FILLCELL_X32 FILLER_97_1680 ();
 FILLCELL_X32 FILLER_97_1712 ();
 FILLCELL_X32 FILLER_97_1744 ();
 FILLCELL_X32 FILLER_97_1776 ();
 FILLCELL_X32 FILLER_97_1808 ();
 FILLCELL_X32 FILLER_97_1840 ();
 FILLCELL_X32 FILLER_97_1872 ();
 FILLCELL_X32 FILLER_97_1904 ();
 FILLCELL_X32 FILLER_97_1936 ();
 FILLCELL_X32 FILLER_97_1968 ();
 FILLCELL_X32 FILLER_97_2000 ();
 FILLCELL_X32 FILLER_97_2032 ();
 FILLCELL_X32 FILLER_97_2064 ();
 FILLCELL_X32 FILLER_97_2096 ();
 FILLCELL_X32 FILLER_97_2128 ();
 FILLCELL_X32 FILLER_97_2160 ();
 FILLCELL_X32 FILLER_97_2192 ();
 FILLCELL_X32 FILLER_97_2224 ();
 FILLCELL_X32 FILLER_97_2256 ();
 FILLCELL_X32 FILLER_97_2288 ();
 FILLCELL_X32 FILLER_97_2320 ();
 FILLCELL_X32 FILLER_97_2352 ();
 FILLCELL_X32 FILLER_97_2384 ();
 FILLCELL_X32 FILLER_97_2416 ();
 FILLCELL_X32 FILLER_97_2448 ();
 FILLCELL_X32 FILLER_97_2480 ();
 FILLCELL_X8 FILLER_97_2512 ();
 FILLCELL_X4 FILLER_97_2520 ();
 FILLCELL_X2 FILLER_97_2524 ();
 FILLCELL_X32 FILLER_97_2527 ();
 FILLCELL_X32 FILLER_97_2559 ();
 FILLCELL_X8 FILLER_97_2591 ();
 FILLCELL_X2 FILLER_97_2599 ();
 FILLCELL_X1 FILLER_97_2601 ();
 FILLCELL_X32 FILLER_98_1 ();
 FILLCELL_X32 FILLER_98_33 ();
 FILLCELL_X32 FILLER_98_65 ();
 FILLCELL_X32 FILLER_98_97 ();
 FILLCELL_X32 FILLER_98_129 ();
 FILLCELL_X32 FILLER_98_161 ();
 FILLCELL_X32 FILLER_98_193 ();
 FILLCELL_X32 FILLER_98_225 ();
 FILLCELL_X32 FILLER_98_257 ();
 FILLCELL_X32 FILLER_98_289 ();
 FILLCELL_X32 FILLER_98_321 ();
 FILLCELL_X32 FILLER_98_353 ();
 FILLCELL_X32 FILLER_98_385 ();
 FILLCELL_X32 FILLER_98_417 ();
 FILLCELL_X32 FILLER_98_449 ();
 FILLCELL_X32 FILLER_98_481 ();
 FILLCELL_X32 FILLER_98_513 ();
 FILLCELL_X32 FILLER_98_545 ();
 FILLCELL_X32 FILLER_98_577 ();
 FILLCELL_X16 FILLER_98_609 ();
 FILLCELL_X4 FILLER_98_625 ();
 FILLCELL_X2 FILLER_98_629 ();
 FILLCELL_X32 FILLER_98_632 ();
 FILLCELL_X32 FILLER_98_664 ();
 FILLCELL_X32 FILLER_98_696 ();
 FILLCELL_X32 FILLER_98_728 ();
 FILLCELL_X32 FILLER_98_760 ();
 FILLCELL_X32 FILLER_98_792 ();
 FILLCELL_X32 FILLER_98_824 ();
 FILLCELL_X32 FILLER_98_856 ();
 FILLCELL_X32 FILLER_98_888 ();
 FILLCELL_X32 FILLER_98_920 ();
 FILLCELL_X32 FILLER_98_952 ();
 FILLCELL_X32 FILLER_98_984 ();
 FILLCELL_X32 FILLER_98_1016 ();
 FILLCELL_X32 FILLER_98_1048 ();
 FILLCELL_X32 FILLER_98_1080 ();
 FILLCELL_X32 FILLER_98_1112 ();
 FILLCELL_X32 FILLER_98_1144 ();
 FILLCELL_X32 FILLER_98_1176 ();
 FILLCELL_X32 FILLER_98_1208 ();
 FILLCELL_X32 FILLER_98_1240 ();
 FILLCELL_X32 FILLER_98_1272 ();
 FILLCELL_X32 FILLER_98_1304 ();
 FILLCELL_X32 FILLER_98_1336 ();
 FILLCELL_X32 FILLER_98_1368 ();
 FILLCELL_X32 FILLER_98_1400 ();
 FILLCELL_X32 FILLER_98_1432 ();
 FILLCELL_X32 FILLER_98_1464 ();
 FILLCELL_X32 FILLER_98_1496 ();
 FILLCELL_X32 FILLER_98_1528 ();
 FILLCELL_X32 FILLER_98_1560 ();
 FILLCELL_X32 FILLER_98_1592 ();
 FILLCELL_X32 FILLER_98_1624 ();
 FILLCELL_X32 FILLER_98_1656 ();
 FILLCELL_X32 FILLER_98_1688 ();
 FILLCELL_X32 FILLER_98_1720 ();
 FILLCELL_X32 FILLER_98_1752 ();
 FILLCELL_X32 FILLER_98_1784 ();
 FILLCELL_X32 FILLER_98_1816 ();
 FILLCELL_X32 FILLER_98_1848 ();
 FILLCELL_X8 FILLER_98_1880 ();
 FILLCELL_X4 FILLER_98_1888 ();
 FILLCELL_X2 FILLER_98_1892 ();
 FILLCELL_X32 FILLER_98_1895 ();
 FILLCELL_X32 FILLER_98_1927 ();
 FILLCELL_X32 FILLER_98_1959 ();
 FILLCELL_X32 FILLER_98_1991 ();
 FILLCELL_X32 FILLER_98_2023 ();
 FILLCELL_X32 FILLER_98_2055 ();
 FILLCELL_X32 FILLER_98_2087 ();
 FILLCELL_X32 FILLER_98_2119 ();
 FILLCELL_X32 FILLER_98_2151 ();
 FILLCELL_X32 FILLER_98_2183 ();
 FILLCELL_X32 FILLER_98_2215 ();
 FILLCELL_X32 FILLER_98_2247 ();
 FILLCELL_X32 FILLER_98_2279 ();
 FILLCELL_X32 FILLER_98_2311 ();
 FILLCELL_X32 FILLER_98_2343 ();
 FILLCELL_X32 FILLER_98_2375 ();
 FILLCELL_X32 FILLER_98_2407 ();
 FILLCELL_X32 FILLER_98_2439 ();
 FILLCELL_X32 FILLER_98_2471 ();
 FILLCELL_X32 FILLER_98_2503 ();
 FILLCELL_X32 FILLER_98_2535 ();
 FILLCELL_X32 FILLER_98_2567 ();
 FILLCELL_X2 FILLER_98_2599 ();
 FILLCELL_X1 FILLER_98_2601 ();
 FILLCELL_X32 FILLER_99_1 ();
 FILLCELL_X32 FILLER_99_33 ();
 FILLCELL_X32 FILLER_99_65 ();
 FILLCELL_X32 FILLER_99_97 ();
 FILLCELL_X32 FILLER_99_129 ();
 FILLCELL_X32 FILLER_99_161 ();
 FILLCELL_X32 FILLER_99_193 ();
 FILLCELL_X32 FILLER_99_225 ();
 FILLCELL_X32 FILLER_99_257 ();
 FILLCELL_X32 FILLER_99_289 ();
 FILLCELL_X32 FILLER_99_321 ();
 FILLCELL_X32 FILLER_99_353 ();
 FILLCELL_X32 FILLER_99_385 ();
 FILLCELL_X32 FILLER_99_417 ();
 FILLCELL_X32 FILLER_99_449 ();
 FILLCELL_X32 FILLER_99_481 ();
 FILLCELL_X32 FILLER_99_513 ();
 FILLCELL_X32 FILLER_99_545 ();
 FILLCELL_X32 FILLER_99_577 ();
 FILLCELL_X32 FILLER_99_609 ();
 FILLCELL_X32 FILLER_99_641 ();
 FILLCELL_X32 FILLER_99_673 ();
 FILLCELL_X32 FILLER_99_705 ();
 FILLCELL_X32 FILLER_99_737 ();
 FILLCELL_X32 FILLER_99_769 ();
 FILLCELL_X32 FILLER_99_801 ();
 FILLCELL_X32 FILLER_99_833 ();
 FILLCELL_X32 FILLER_99_865 ();
 FILLCELL_X32 FILLER_99_897 ();
 FILLCELL_X32 FILLER_99_929 ();
 FILLCELL_X32 FILLER_99_961 ();
 FILLCELL_X32 FILLER_99_993 ();
 FILLCELL_X32 FILLER_99_1025 ();
 FILLCELL_X32 FILLER_99_1057 ();
 FILLCELL_X32 FILLER_99_1089 ();
 FILLCELL_X32 FILLER_99_1121 ();
 FILLCELL_X32 FILLER_99_1153 ();
 FILLCELL_X32 FILLER_99_1185 ();
 FILLCELL_X32 FILLER_99_1217 ();
 FILLCELL_X8 FILLER_99_1249 ();
 FILLCELL_X4 FILLER_99_1257 ();
 FILLCELL_X2 FILLER_99_1261 ();
 FILLCELL_X32 FILLER_99_1264 ();
 FILLCELL_X32 FILLER_99_1296 ();
 FILLCELL_X32 FILLER_99_1328 ();
 FILLCELL_X32 FILLER_99_1360 ();
 FILLCELL_X32 FILLER_99_1392 ();
 FILLCELL_X32 FILLER_99_1424 ();
 FILLCELL_X32 FILLER_99_1456 ();
 FILLCELL_X32 FILLER_99_1488 ();
 FILLCELL_X32 FILLER_99_1520 ();
 FILLCELL_X32 FILLER_99_1552 ();
 FILLCELL_X32 FILLER_99_1584 ();
 FILLCELL_X32 FILLER_99_1616 ();
 FILLCELL_X32 FILLER_99_1648 ();
 FILLCELL_X32 FILLER_99_1680 ();
 FILLCELL_X32 FILLER_99_1712 ();
 FILLCELL_X32 FILLER_99_1744 ();
 FILLCELL_X32 FILLER_99_1776 ();
 FILLCELL_X32 FILLER_99_1808 ();
 FILLCELL_X32 FILLER_99_1840 ();
 FILLCELL_X32 FILLER_99_1872 ();
 FILLCELL_X32 FILLER_99_1904 ();
 FILLCELL_X32 FILLER_99_1936 ();
 FILLCELL_X32 FILLER_99_1968 ();
 FILLCELL_X32 FILLER_99_2000 ();
 FILLCELL_X32 FILLER_99_2032 ();
 FILLCELL_X32 FILLER_99_2064 ();
 FILLCELL_X32 FILLER_99_2096 ();
 FILLCELL_X32 FILLER_99_2128 ();
 FILLCELL_X32 FILLER_99_2160 ();
 FILLCELL_X32 FILLER_99_2192 ();
 FILLCELL_X32 FILLER_99_2224 ();
 FILLCELL_X32 FILLER_99_2256 ();
 FILLCELL_X32 FILLER_99_2288 ();
 FILLCELL_X32 FILLER_99_2320 ();
 FILLCELL_X32 FILLER_99_2352 ();
 FILLCELL_X32 FILLER_99_2384 ();
 FILLCELL_X32 FILLER_99_2416 ();
 FILLCELL_X32 FILLER_99_2448 ();
 FILLCELL_X32 FILLER_99_2480 ();
 FILLCELL_X8 FILLER_99_2512 ();
 FILLCELL_X4 FILLER_99_2520 ();
 FILLCELL_X2 FILLER_99_2524 ();
 FILLCELL_X32 FILLER_99_2527 ();
 FILLCELL_X32 FILLER_99_2559 ();
 FILLCELL_X8 FILLER_99_2591 ();
 FILLCELL_X2 FILLER_99_2599 ();
 FILLCELL_X1 FILLER_99_2601 ();
 FILLCELL_X32 FILLER_100_1 ();
 FILLCELL_X32 FILLER_100_33 ();
 FILLCELL_X32 FILLER_100_65 ();
 FILLCELL_X32 FILLER_100_97 ();
 FILLCELL_X32 FILLER_100_129 ();
 FILLCELL_X32 FILLER_100_161 ();
 FILLCELL_X32 FILLER_100_193 ();
 FILLCELL_X32 FILLER_100_225 ();
 FILLCELL_X32 FILLER_100_257 ();
 FILLCELL_X32 FILLER_100_289 ();
 FILLCELL_X32 FILLER_100_321 ();
 FILLCELL_X32 FILLER_100_353 ();
 FILLCELL_X32 FILLER_100_385 ();
 FILLCELL_X32 FILLER_100_417 ();
 FILLCELL_X32 FILLER_100_449 ();
 FILLCELL_X32 FILLER_100_481 ();
 FILLCELL_X32 FILLER_100_513 ();
 FILLCELL_X32 FILLER_100_545 ();
 FILLCELL_X32 FILLER_100_577 ();
 FILLCELL_X16 FILLER_100_609 ();
 FILLCELL_X4 FILLER_100_625 ();
 FILLCELL_X2 FILLER_100_629 ();
 FILLCELL_X32 FILLER_100_632 ();
 FILLCELL_X32 FILLER_100_664 ();
 FILLCELL_X32 FILLER_100_696 ();
 FILLCELL_X32 FILLER_100_728 ();
 FILLCELL_X32 FILLER_100_760 ();
 FILLCELL_X32 FILLER_100_792 ();
 FILLCELL_X32 FILLER_100_824 ();
 FILLCELL_X32 FILLER_100_856 ();
 FILLCELL_X32 FILLER_100_888 ();
 FILLCELL_X32 FILLER_100_920 ();
 FILLCELL_X32 FILLER_100_952 ();
 FILLCELL_X32 FILLER_100_984 ();
 FILLCELL_X32 FILLER_100_1016 ();
 FILLCELL_X32 FILLER_100_1048 ();
 FILLCELL_X32 FILLER_100_1080 ();
 FILLCELL_X32 FILLER_100_1112 ();
 FILLCELL_X32 FILLER_100_1144 ();
 FILLCELL_X32 FILLER_100_1176 ();
 FILLCELL_X32 FILLER_100_1208 ();
 FILLCELL_X32 FILLER_100_1240 ();
 FILLCELL_X32 FILLER_100_1272 ();
 FILLCELL_X32 FILLER_100_1304 ();
 FILLCELL_X32 FILLER_100_1336 ();
 FILLCELL_X32 FILLER_100_1368 ();
 FILLCELL_X32 FILLER_100_1400 ();
 FILLCELL_X32 FILLER_100_1432 ();
 FILLCELL_X32 FILLER_100_1464 ();
 FILLCELL_X32 FILLER_100_1496 ();
 FILLCELL_X32 FILLER_100_1528 ();
 FILLCELL_X32 FILLER_100_1560 ();
 FILLCELL_X32 FILLER_100_1592 ();
 FILLCELL_X32 FILLER_100_1624 ();
 FILLCELL_X32 FILLER_100_1656 ();
 FILLCELL_X32 FILLER_100_1688 ();
 FILLCELL_X32 FILLER_100_1720 ();
 FILLCELL_X32 FILLER_100_1752 ();
 FILLCELL_X32 FILLER_100_1784 ();
 FILLCELL_X32 FILLER_100_1816 ();
 FILLCELL_X32 FILLER_100_1848 ();
 FILLCELL_X8 FILLER_100_1880 ();
 FILLCELL_X4 FILLER_100_1888 ();
 FILLCELL_X2 FILLER_100_1892 ();
 FILLCELL_X32 FILLER_100_1895 ();
 FILLCELL_X32 FILLER_100_1927 ();
 FILLCELL_X32 FILLER_100_1959 ();
 FILLCELL_X32 FILLER_100_1991 ();
 FILLCELL_X32 FILLER_100_2023 ();
 FILLCELL_X32 FILLER_100_2055 ();
 FILLCELL_X32 FILLER_100_2087 ();
 FILLCELL_X32 FILLER_100_2119 ();
 FILLCELL_X32 FILLER_100_2151 ();
 FILLCELL_X32 FILLER_100_2183 ();
 FILLCELL_X32 FILLER_100_2215 ();
 FILLCELL_X32 FILLER_100_2247 ();
 FILLCELL_X32 FILLER_100_2279 ();
 FILLCELL_X32 FILLER_100_2311 ();
 FILLCELL_X32 FILLER_100_2343 ();
 FILLCELL_X32 FILLER_100_2375 ();
 FILLCELL_X32 FILLER_100_2407 ();
 FILLCELL_X32 FILLER_100_2439 ();
 FILLCELL_X32 FILLER_100_2471 ();
 FILLCELL_X32 FILLER_100_2503 ();
 FILLCELL_X32 FILLER_100_2535 ();
 FILLCELL_X32 FILLER_100_2567 ();
 FILLCELL_X2 FILLER_100_2599 ();
 FILLCELL_X1 FILLER_100_2601 ();
 FILLCELL_X32 FILLER_101_1 ();
 FILLCELL_X32 FILLER_101_33 ();
 FILLCELL_X32 FILLER_101_65 ();
 FILLCELL_X32 FILLER_101_97 ();
 FILLCELL_X32 FILLER_101_129 ();
 FILLCELL_X32 FILLER_101_161 ();
 FILLCELL_X32 FILLER_101_193 ();
 FILLCELL_X32 FILLER_101_225 ();
 FILLCELL_X32 FILLER_101_257 ();
 FILLCELL_X32 FILLER_101_289 ();
 FILLCELL_X32 FILLER_101_321 ();
 FILLCELL_X32 FILLER_101_353 ();
 FILLCELL_X32 FILLER_101_385 ();
 FILLCELL_X32 FILLER_101_417 ();
 FILLCELL_X32 FILLER_101_449 ();
 FILLCELL_X32 FILLER_101_481 ();
 FILLCELL_X32 FILLER_101_513 ();
 FILLCELL_X32 FILLER_101_545 ();
 FILLCELL_X32 FILLER_101_577 ();
 FILLCELL_X32 FILLER_101_609 ();
 FILLCELL_X32 FILLER_101_641 ();
 FILLCELL_X32 FILLER_101_673 ();
 FILLCELL_X32 FILLER_101_705 ();
 FILLCELL_X32 FILLER_101_737 ();
 FILLCELL_X32 FILLER_101_769 ();
 FILLCELL_X32 FILLER_101_801 ();
 FILLCELL_X32 FILLER_101_833 ();
 FILLCELL_X32 FILLER_101_865 ();
 FILLCELL_X32 FILLER_101_897 ();
 FILLCELL_X32 FILLER_101_929 ();
 FILLCELL_X32 FILLER_101_961 ();
 FILLCELL_X32 FILLER_101_993 ();
 FILLCELL_X32 FILLER_101_1025 ();
 FILLCELL_X32 FILLER_101_1057 ();
 FILLCELL_X32 FILLER_101_1089 ();
 FILLCELL_X32 FILLER_101_1121 ();
 FILLCELL_X32 FILLER_101_1153 ();
 FILLCELL_X32 FILLER_101_1185 ();
 FILLCELL_X32 FILLER_101_1217 ();
 FILLCELL_X8 FILLER_101_1249 ();
 FILLCELL_X4 FILLER_101_1257 ();
 FILLCELL_X2 FILLER_101_1261 ();
 FILLCELL_X32 FILLER_101_1264 ();
 FILLCELL_X32 FILLER_101_1296 ();
 FILLCELL_X32 FILLER_101_1328 ();
 FILLCELL_X32 FILLER_101_1360 ();
 FILLCELL_X32 FILLER_101_1392 ();
 FILLCELL_X32 FILLER_101_1424 ();
 FILLCELL_X32 FILLER_101_1456 ();
 FILLCELL_X32 FILLER_101_1488 ();
 FILLCELL_X32 FILLER_101_1520 ();
 FILLCELL_X32 FILLER_101_1552 ();
 FILLCELL_X32 FILLER_101_1584 ();
 FILLCELL_X32 FILLER_101_1616 ();
 FILLCELL_X32 FILLER_101_1648 ();
 FILLCELL_X32 FILLER_101_1680 ();
 FILLCELL_X32 FILLER_101_1712 ();
 FILLCELL_X32 FILLER_101_1744 ();
 FILLCELL_X32 FILLER_101_1776 ();
 FILLCELL_X32 FILLER_101_1808 ();
 FILLCELL_X32 FILLER_101_1840 ();
 FILLCELL_X32 FILLER_101_1872 ();
 FILLCELL_X32 FILLER_101_1904 ();
 FILLCELL_X32 FILLER_101_1936 ();
 FILLCELL_X32 FILLER_101_1968 ();
 FILLCELL_X32 FILLER_101_2000 ();
 FILLCELL_X32 FILLER_101_2032 ();
 FILLCELL_X32 FILLER_101_2064 ();
 FILLCELL_X32 FILLER_101_2096 ();
 FILLCELL_X32 FILLER_101_2128 ();
 FILLCELL_X32 FILLER_101_2160 ();
 FILLCELL_X32 FILLER_101_2192 ();
 FILLCELL_X32 FILLER_101_2224 ();
 FILLCELL_X32 FILLER_101_2256 ();
 FILLCELL_X32 FILLER_101_2288 ();
 FILLCELL_X32 FILLER_101_2320 ();
 FILLCELL_X32 FILLER_101_2352 ();
 FILLCELL_X32 FILLER_101_2384 ();
 FILLCELL_X32 FILLER_101_2416 ();
 FILLCELL_X32 FILLER_101_2448 ();
 FILLCELL_X32 FILLER_101_2480 ();
 FILLCELL_X8 FILLER_101_2512 ();
 FILLCELL_X4 FILLER_101_2520 ();
 FILLCELL_X2 FILLER_101_2524 ();
 FILLCELL_X32 FILLER_101_2527 ();
 FILLCELL_X32 FILLER_101_2559 ();
 FILLCELL_X8 FILLER_101_2591 ();
 FILLCELL_X2 FILLER_101_2599 ();
 FILLCELL_X1 FILLER_101_2601 ();
 FILLCELL_X32 FILLER_102_1 ();
 FILLCELL_X32 FILLER_102_33 ();
 FILLCELL_X32 FILLER_102_65 ();
 FILLCELL_X32 FILLER_102_97 ();
 FILLCELL_X32 FILLER_102_129 ();
 FILLCELL_X32 FILLER_102_161 ();
 FILLCELL_X32 FILLER_102_193 ();
 FILLCELL_X32 FILLER_102_225 ();
 FILLCELL_X32 FILLER_102_257 ();
 FILLCELL_X32 FILLER_102_289 ();
 FILLCELL_X32 FILLER_102_321 ();
 FILLCELL_X32 FILLER_102_353 ();
 FILLCELL_X32 FILLER_102_385 ();
 FILLCELL_X32 FILLER_102_417 ();
 FILLCELL_X32 FILLER_102_449 ();
 FILLCELL_X32 FILLER_102_481 ();
 FILLCELL_X32 FILLER_102_513 ();
 FILLCELL_X32 FILLER_102_545 ();
 FILLCELL_X32 FILLER_102_577 ();
 FILLCELL_X16 FILLER_102_609 ();
 FILLCELL_X4 FILLER_102_625 ();
 FILLCELL_X2 FILLER_102_629 ();
 FILLCELL_X32 FILLER_102_632 ();
 FILLCELL_X32 FILLER_102_664 ();
 FILLCELL_X32 FILLER_102_696 ();
 FILLCELL_X32 FILLER_102_728 ();
 FILLCELL_X32 FILLER_102_760 ();
 FILLCELL_X32 FILLER_102_792 ();
 FILLCELL_X32 FILLER_102_824 ();
 FILLCELL_X32 FILLER_102_856 ();
 FILLCELL_X32 FILLER_102_888 ();
 FILLCELL_X32 FILLER_102_920 ();
 FILLCELL_X32 FILLER_102_952 ();
 FILLCELL_X32 FILLER_102_984 ();
 FILLCELL_X32 FILLER_102_1016 ();
 FILLCELL_X32 FILLER_102_1048 ();
 FILLCELL_X32 FILLER_102_1080 ();
 FILLCELL_X32 FILLER_102_1112 ();
 FILLCELL_X32 FILLER_102_1144 ();
 FILLCELL_X32 FILLER_102_1176 ();
 FILLCELL_X32 FILLER_102_1208 ();
 FILLCELL_X32 FILLER_102_1240 ();
 FILLCELL_X32 FILLER_102_1272 ();
 FILLCELL_X32 FILLER_102_1304 ();
 FILLCELL_X32 FILLER_102_1336 ();
 FILLCELL_X32 FILLER_102_1368 ();
 FILLCELL_X32 FILLER_102_1400 ();
 FILLCELL_X32 FILLER_102_1432 ();
 FILLCELL_X32 FILLER_102_1464 ();
 FILLCELL_X32 FILLER_102_1496 ();
 FILLCELL_X32 FILLER_102_1528 ();
 FILLCELL_X32 FILLER_102_1560 ();
 FILLCELL_X32 FILLER_102_1592 ();
 FILLCELL_X32 FILLER_102_1624 ();
 FILLCELL_X32 FILLER_102_1656 ();
 FILLCELL_X32 FILLER_102_1688 ();
 FILLCELL_X32 FILLER_102_1720 ();
 FILLCELL_X32 FILLER_102_1752 ();
 FILLCELL_X32 FILLER_102_1784 ();
 FILLCELL_X32 FILLER_102_1816 ();
 FILLCELL_X32 FILLER_102_1848 ();
 FILLCELL_X8 FILLER_102_1880 ();
 FILLCELL_X4 FILLER_102_1888 ();
 FILLCELL_X2 FILLER_102_1892 ();
 FILLCELL_X32 FILLER_102_1895 ();
 FILLCELL_X32 FILLER_102_1927 ();
 FILLCELL_X32 FILLER_102_1959 ();
 FILLCELL_X32 FILLER_102_1991 ();
 FILLCELL_X32 FILLER_102_2023 ();
 FILLCELL_X32 FILLER_102_2055 ();
 FILLCELL_X32 FILLER_102_2087 ();
 FILLCELL_X32 FILLER_102_2119 ();
 FILLCELL_X32 FILLER_102_2151 ();
 FILLCELL_X32 FILLER_102_2183 ();
 FILLCELL_X32 FILLER_102_2215 ();
 FILLCELL_X32 FILLER_102_2247 ();
 FILLCELL_X32 FILLER_102_2279 ();
 FILLCELL_X32 FILLER_102_2311 ();
 FILLCELL_X32 FILLER_102_2343 ();
 FILLCELL_X32 FILLER_102_2375 ();
 FILLCELL_X32 FILLER_102_2407 ();
 FILLCELL_X32 FILLER_102_2439 ();
 FILLCELL_X32 FILLER_102_2471 ();
 FILLCELL_X32 FILLER_102_2503 ();
 FILLCELL_X32 FILLER_102_2535 ();
 FILLCELL_X32 FILLER_102_2567 ();
 FILLCELL_X2 FILLER_102_2599 ();
 FILLCELL_X1 FILLER_102_2601 ();
 FILLCELL_X32 FILLER_103_1 ();
 FILLCELL_X32 FILLER_103_33 ();
 FILLCELL_X32 FILLER_103_65 ();
 FILLCELL_X32 FILLER_103_97 ();
 FILLCELL_X32 FILLER_103_129 ();
 FILLCELL_X32 FILLER_103_161 ();
 FILLCELL_X32 FILLER_103_193 ();
 FILLCELL_X32 FILLER_103_225 ();
 FILLCELL_X32 FILLER_103_257 ();
 FILLCELL_X32 FILLER_103_289 ();
 FILLCELL_X32 FILLER_103_321 ();
 FILLCELL_X32 FILLER_103_353 ();
 FILLCELL_X32 FILLER_103_385 ();
 FILLCELL_X32 FILLER_103_417 ();
 FILLCELL_X32 FILLER_103_449 ();
 FILLCELL_X32 FILLER_103_481 ();
 FILLCELL_X32 FILLER_103_513 ();
 FILLCELL_X32 FILLER_103_545 ();
 FILLCELL_X32 FILLER_103_577 ();
 FILLCELL_X32 FILLER_103_609 ();
 FILLCELL_X32 FILLER_103_641 ();
 FILLCELL_X32 FILLER_103_673 ();
 FILLCELL_X32 FILLER_103_705 ();
 FILLCELL_X32 FILLER_103_737 ();
 FILLCELL_X32 FILLER_103_769 ();
 FILLCELL_X32 FILLER_103_801 ();
 FILLCELL_X32 FILLER_103_833 ();
 FILLCELL_X32 FILLER_103_865 ();
 FILLCELL_X32 FILLER_103_897 ();
 FILLCELL_X32 FILLER_103_929 ();
 FILLCELL_X32 FILLER_103_961 ();
 FILLCELL_X32 FILLER_103_993 ();
 FILLCELL_X32 FILLER_103_1025 ();
 FILLCELL_X32 FILLER_103_1057 ();
 FILLCELL_X32 FILLER_103_1089 ();
 FILLCELL_X32 FILLER_103_1121 ();
 FILLCELL_X32 FILLER_103_1153 ();
 FILLCELL_X32 FILLER_103_1185 ();
 FILLCELL_X32 FILLER_103_1217 ();
 FILLCELL_X8 FILLER_103_1249 ();
 FILLCELL_X4 FILLER_103_1257 ();
 FILLCELL_X2 FILLER_103_1261 ();
 FILLCELL_X32 FILLER_103_1264 ();
 FILLCELL_X32 FILLER_103_1296 ();
 FILLCELL_X32 FILLER_103_1328 ();
 FILLCELL_X32 FILLER_103_1360 ();
 FILLCELL_X32 FILLER_103_1392 ();
 FILLCELL_X32 FILLER_103_1424 ();
 FILLCELL_X32 FILLER_103_1456 ();
 FILLCELL_X32 FILLER_103_1488 ();
 FILLCELL_X32 FILLER_103_1520 ();
 FILLCELL_X32 FILLER_103_1552 ();
 FILLCELL_X32 FILLER_103_1584 ();
 FILLCELL_X32 FILLER_103_1616 ();
 FILLCELL_X32 FILLER_103_1648 ();
 FILLCELL_X32 FILLER_103_1680 ();
 FILLCELL_X32 FILLER_103_1712 ();
 FILLCELL_X32 FILLER_103_1744 ();
 FILLCELL_X32 FILLER_103_1776 ();
 FILLCELL_X32 FILLER_103_1808 ();
 FILLCELL_X32 FILLER_103_1840 ();
 FILLCELL_X32 FILLER_103_1872 ();
 FILLCELL_X32 FILLER_103_1904 ();
 FILLCELL_X32 FILLER_103_1936 ();
 FILLCELL_X32 FILLER_103_1968 ();
 FILLCELL_X32 FILLER_103_2000 ();
 FILLCELL_X32 FILLER_103_2032 ();
 FILLCELL_X32 FILLER_103_2064 ();
 FILLCELL_X32 FILLER_103_2096 ();
 FILLCELL_X32 FILLER_103_2128 ();
 FILLCELL_X32 FILLER_103_2160 ();
 FILLCELL_X32 FILLER_103_2192 ();
 FILLCELL_X32 FILLER_103_2224 ();
 FILLCELL_X32 FILLER_103_2256 ();
 FILLCELL_X32 FILLER_103_2288 ();
 FILLCELL_X32 FILLER_103_2320 ();
 FILLCELL_X32 FILLER_103_2352 ();
 FILLCELL_X32 FILLER_103_2384 ();
 FILLCELL_X32 FILLER_103_2416 ();
 FILLCELL_X32 FILLER_103_2448 ();
 FILLCELL_X32 FILLER_103_2480 ();
 FILLCELL_X8 FILLER_103_2512 ();
 FILLCELL_X4 FILLER_103_2520 ();
 FILLCELL_X2 FILLER_103_2524 ();
 FILLCELL_X32 FILLER_103_2527 ();
 FILLCELL_X32 FILLER_103_2559 ();
 FILLCELL_X8 FILLER_103_2591 ();
 FILLCELL_X2 FILLER_103_2599 ();
 FILLCELL_X1 FILLER_103_2601 ();
 FILLCELL_X32 FILLER_104_1 ();
 FILLCELL_X32 FILLER_104_33 ();
 FILLCELL_X32 FILLER_104_65 ();
 FILLCELL_X32 FILLER_104_97 ();
 FILLCELL_X32 FILLER_104_129 ();
 FILLCELL_X32 FILLER_104_161 ();
 FILLCELL_X32 FILLER_104_193 ();
 FILLCELL_X32 FILLER_104_225 ();
 FILLCELL_X32 FILLER_104_257 ();
 FILLCELL_X32 FILLER_104_289 ();
 FILLCELL_X32 FILLER_104_321 ();
 FILLCELL_X32 FILLER_104_353 ();
 FILLCELL_X32 FILLER_104_385 ();
 FILLCELL_X32 FILLER_104_417 ();
 FILLCELL_X32 FILLER_104_449 ();
 FILLCELL_X32 FILLER_104_481 ();
 FILLCELL_X32 FILLER_104_513 ();
 FILLCELL_X32 FILLER_104_545 ();
 FILLCELL_X32 FILLER_104_577 ();
 FILLCELL_X16 FILLER_104_609 ();
 FILLCELL_X4 FILLER_104_625 ();
 FILLCELL_X2 FILLER_104_629 ();
 FILLCELL_X32 FILLER_104_632 ();
 FILLCELL_X32 FILLER_104_664 ();
 FILLCELL_X32 FILLER_104_696 ();
 FILLCELL_X32 FILLER_104_728 ();
 FILLCELL_X32 FILLER_104_760 ();
 FILLCELL_X32 FILLER_104_792 ();
 FILLCELL_X32 FILLER_104_824 ();
 FILLCELL_X32 FILLER_104_856 ();
 FILLCELL_X32 FILLER_104_888 ();
 FILLCELL_X32 FILLER_104_920 ();
 FILLCELL_X32 FILLER_104_952 ();
 FILLCELL_X32 FILLER_104_984 ();
 FILLCELL_X32 FILLER_104_1016 ();
 FILLCELL_X32 FILLER_104_1048 ();
 FILLCELL_X32 FILLER_104_1080 ();
 FILLCELL_X32 FILLER_104_1112 ();
 FILLCELL_X32 FILLER_104_1144 ();
 FILLCELL_X32 FILLER_104_1176 ();
 FILLCELL_X32 FILLER_104_1208 ();
 FILLCELL_X32 FILLER_104_1240 ();
 FILLCELL_X32 FILLER_104_1272 ();
 FILLCELL_X32 FILLER_104_1304 ();
 FILLCELL_X32 FILLER_104_1336 ();
 FILLCELL_X32 FILLER_104_1368 ();
 FILLCELL_X32 FILLER_104_1400 ();
 FILLCELL_X32 FILLER_104_1432 ();
 FILLCELL_X32 FILLER_104_1464 ();
 FILLCELL_X32 FILLER_104_1496 ();
 FILLCELL_X32 FILLER_104_1528 ();
 FILLCELL_X32 FILLER_104_1560 ();
 FILLCELL_X32 FILLER_104_1592 ();
 FILLCELL_X32 FILLER_104_1624 ();
 FILLCELL_X32 FILLER_104_1656 ();
 FILLCELL_X32 FILLER_104_1688 ();
 FILLCELL_X32 FILLER_104_1720 ();
 FILLCELL_X32 FILLER_104_1752 ();
 FILLCELL_X32 FILLER_104_1784 ();
 FILLCELL_X32 FILLER_104_1816 ();
 FILLCELL_X32 FILLER_104_1848 ();
 FILLCELL_X8 FILLER_104_1880 ();
 FILLCELL_X4 FILLER_104_1888 ();
 FILLCELL_X2 FILLER_104_1892 ();
 FILLCELL_X32 FILLER_104_1895 ();
 FILLCELL_X32 FILLER_104_1927 ();
 FILLCELL_X32 FILLER_104_1959 ();
 FILLCELL_X32 FILLER_104_1991 ();
 FILLCELL_X32 FILLER_104_2023 ();
 FILLCELL_X32 FILLER_104_2055 ();
 FILLCELL_X32 FILLER_104_2087 ();
 FILLCELL_X32 FILLER_104_2119 ();
 FILLCELL_X32 FILLER_104_2151 ();
 FILLCELL_X32 FILLER_104_2183 ();
 FILLCELL_X32 FILLER_104_2215 ();
 FILLCELL_X32 FILLER_104_2247 ();
 FILLCELL_X32 FILLER_104_2279 ();
 FILLCELL_X32 FILLER_104_2311 ();
 FILLCELL_X32 FILLER_104_2343 ();
 FILLCELL_X32 FILLER_104_2375 ();
 FILLCELL_X32 FILLER_104_2407 ();
 FILLCELL_X32 FILLER_104_2439 ();
 FILLCELL_X32 FILLER_104_2471 ();
 FILLCELL_X32 FILLER_104_2503 ();
 FILLCELL_X32 FILLER_104_2535 ();
 FILLCELL_X32 FILLER_104_2567 ();
 FILLCELL_X2 FILLER_104_2599 ();
 FILLCELL_X1 FILLER_104_2601 ();
 FILLCELL_X32 FILLER_105_1 ();
 FILLCELL_X32 FILLER_105_33 ();
 FILLCELL_X32 FILLER_105_65 ();
 FILLCELL_X32 FILLER_105_97 ();
 FILLCELL_X32 FILLER_105_129 ();
 FILLCELL_X32 FILLER_105_161 ();
 FILLCELL_X32 FILLER_105_193 ();
 FILLCELL_X32 FILLER_105_225 ();
 FILLCELL_X32 FILLER_105_257 ();
 FILLCELL_X32 FILLER_105_289 ();
 FILLCELL_X32 FILLER_105_321 ();
 FILLCELL_X32 FILLER_105_353 ();
 FILLCELL_X32 FILLER_105_385 ();
 FILLCELL_X32 FILLER_105_417 ();
 FILLCELL_X32 FILLER_105_449 ();
 FILLCELL_X32 FILLER_105_481 ();
 FILLCELL_X32 FILLER_105_513 ();
 FILLCELL_X32 FILLER_105_545 ();
 FILLCELL_X32 FILLER_105_577 ();
 FILLCELL_X32 FILLER_105_609 ();
 FILLCELL_X32 FILLER_105_641 ();
 FILLCELL_X32 FILLER_105_673 ();
 FILLCELL_X32 FILLER_105_705 ();
 FILLCELL_X32 FILLER_105_737 ();
 FILLCELL_X32 FILLER_105_769 ();
 FILLCELL_X32 FILLER_105_801 ();
 FILLCELL_X32 FILLER_105_833 ();
 FILLCELL_X32 FILLER_105_865 ();
 FILLCELL_X32 FILLER_105_897 ();
 FILLCELL_X32 FILLER_105_929 ();
 FILLCELL_X32 FILLER_105_961 ();
 FILLCELL_X32 FILLER_105_993 ();
 FILLCELL_X32 FILLER_105_1025 ();
 FILLCELL_X32 FILLER_105_1057 ();
 FILLCELL_X32 FILLER_105_1089 ();
 FILLCELL_X32 FILLER_105_1121 ();
 FILLCELL_X32 FILLER_105_1153 ();
 FILLCELL_X32 FILLER_105_1185 ();
 FILLCELL_X32 FILLER_105_1217 ();
 FILLCELL_X8 FILLER_105_1249 ();
 FILLCELL_X4 FILLER_105_1257 ();
 FILLCELL_X2 FILLER_105_1261 ();
 FILLCELL_X32 FILLER_105_1264 ();
 FILLCELL_X32 FILLER_105_1296 ();
 FILLCELL_X32 FILLER_105_1328 ();
 FILLCELL_X32 FILLER_105_1360 ();
 FILLCELL_X32 FILLER_105_1392 ();
 FILLCELL_X32 FILLER_105_1424 ();
 FILLCELL_X32 FILLER_105_1456 ();
 FILLCELL_X32 FILLER_105_1488 ();
 FILLCELL_X32 FILLER_105_1520 ();
 FILLCELL_X32 FILLER_105_1552 ();
 FILLCELL_X32 FILLER_105_1584 ();
 FILLCELL_X32 FILLER_105_1616 ();
 FILLCELL_X32 FILLER_105_1648 ();
 FILLCELL_X32 FILLER_105_1680 ();
 FILLCELL_X32 FILLER_105_1712 ();
 FILLCELL_X32 FILLER_105_1744 ();
 FILLCELL_X32 FILLER_105_1776 ();
 FILLCELL_X32 FILLER_105_1808 ();
 FILLCELL_X32 FILLER_105_1840 ();
 FILLCELL_X32 FILLER_105_1872 ();
 FILLCELL_X32 FILLER_105_1904 ();
 FILLCELL_X32 FILLER_105_1936 ();
 FILLCELL_X32 FILLER_105_1968 ();
 FILLCELL_X32 FILLER_105_2000 ();
 FILLCELL_X32 FILLER_105_2032 ();
 FILLCELL_X32 FILLER_105_2064 ();
 FILLCELL_X32 FILLER_105_2096 ();
 FILLCELL_X32 FILLER_105_2128 ();
 FILLCELL_X32 FILLER_105_2160 ();
 FILLCELL_X32 FILLER_105_2192 ();
 FILLCELL_X32 FILLER_105_2224 ();
 FILLCELL_X32 FILLER_105_2256 ();
 FILLCELL_X32 FILLER_105_2288 ();
 FILLCELL_X32 FILLER_105_2320 ();
 FILLCELL_X32 FILLER_105_2352 ();
 FILLCELL_X32 FILLER_105_2384 ();
 FILLCELL_X32 FILLER_105_2416 ();
 FILLCELL_X32 FILLER_105_2448 ();
 FILLCELL_X32 FILLER_105_2480 ();
 FILLCELL_X8 FILLER_105_2512 ();
 FILLCELL_X4 FILLER_105_2520 ();
 FILLCELL_X2 FILLER_105_2524 ();
 FILLCELL_X32 FILLER_105_2527 ();
 FILLCELL_X32 FILLER_105_2559 ();
 FILLCELL_X8 FILLER_105_2591 ();
 FILLCELL_X2 FILLER_105_2599 ();
 FILLCELL_X1 FILLER_105_2601 ();
 FILLCELL_X32 FILLER_106_1 ();
 FILLCELL_X32 FILLER_106_33 ();
 FILLCELL_X32 FILLER_106_65 ();
 FILLCELL_X32 FILLER_106_97 ();
 FILLCELL_X32 FILLER_106_129 ();
 FILLCELL_X32 FILLER_106_161 ();
 FILLCELL_X32 FILLER_106_193 ();
 FILLCELL_X32 FILLER_106_225 ();
 FILLCELL_X32 FILLER_106_257 ();
 FILLCELL_X32 FILLER_106_289 ();
 FILLCELL_X32 FILLER_106_321 ();
 FILLCELL_X32 FILLER_106_353 ();
 FILLCELL_X32 FILLER_106_385 ();
 FILLCELL_X32 FILLER_106_417 ();
 FILLCELL_X32 FILLER_106_449 ();
 FILLCELL_X32 FILLER_106_481 ();
 FILLCELL_X32 FILLER_106_513 ();
 FILLCELL_X32 FILLER_106_545 ();
 FILLCELL_X32 FILLER_106_577 ();
 FILLCELL_X16 FILLER_106_609 ();
 FILLCELL_X4 FILLER_106_625 ();
 FILLCELL_X2 FILLER_106_629 ();
 FILLCELL_X32 FILLER_106_632 ();
 FILLCELL_X32 FILLER_106_664 ();
 FILLCELL_X32 FILLER_106_696 ();
 FILLCELL_X32 FILLER_106_728 ();
 FILLCELL_X32 FILLER_106_760 ();
 FILLCELL_X32 FILLER_106_792 ();
 FILLCELL_X32 FILLER_106_824 ();
 FILLCELL_X32 FILLER_106_856 ();
 FILLCELL_X32 FILLER_106_888 ();
 FILLCELL_X32 FILLER_106_920 ();
 FILLCELL_X32 FILLER_106_952 ();
 FILLCELL_X32 FILLER_106_984 ();
 FILLCELL_X32 FILLER_106_1016 ();
 FILLCELL_X32 FILLER_106_1048 ();
 FILLCELL_X32 FILLER_106_1080 ();
 FILLCELL_X32 FILLER_106_1112 ();
 FILLCELL_X32 FILLER_106_1144 ();
 FILLCELL_X32 FILLER_106_1176 ();
 FILLCELL_X32 FILLER_106_1208 ();
 FILLCELL_X32 FILLER_106_1240 ();
 FILLCELL_X32 FILLER_106_1272 ();
 FILLCELL_X32 FILLER_106_1304 ();
 FILLCELL_X32 FILLER_106_1336 ();
 FILLCELL_X32 FILLER_106_1368 ();
 FILLCELL_X32 FILLER_106_1400 ();
 FILLCELL_X32 FILLER_106_1432 ();
 FILLCELL_X32 FILLER_106_1464 ();
 FILLCELL_X32 FILLER_106_1496 ();
 FILLCELL_X32 FILLER_106_1528 ();
 FILLCELL_X32 FILLER_106_1560 ();
 FILLCELL_X32 FILLER_106_1592 ();
 FILLCELL_X32 FILLER_106_1624 ();
 FILLCELL_X32 FILLER_106_1656 ();
 FILLCELL_X32 FILLER_106_1688 ();
 FILLCELL_X32 FILLER_106_1720 ();
 FILLCELL_X32 FILLER_106_1752 ();
 FILLCELL_X32 FILLER_106_1784 ();
 FILLCELL_X32 FILLER_106_1816 ();
 FILLCELL_X32 FILLER_106_1848 ();
 FILLCELL_X8 FILLER_106_1880 ();
 FILLCELL_X4 FILLER_106_1888 ();
 FILLCELL_X2 FILLER_106_1892 ();
 FILLCELL_X32 FILLER_106_1895 ();
 FILLCELL_X32 FILLER_106_1927 ();
 FILLCELL_X32 FILLER_106_1959 ();
 FILLCELL_X32 FILLER_106_1991 ();
 FILLCELL_X32 FILLER_106_2023 ();
 FILLCELL_X32 FILLER_106_2055 ();
 FILLCELL_X32 FILLER_106_2087 ();
 FILLCELL_X32 FILLER_106_2119 ();
 FILLCELL_X32 FILLER_106_2151 ();
 FILLCELL_X32 FILLER_106_2183 ();
 FILLCELL_X32 FILLER_106_2215 ();
 FILLCELL_X32 FILLER_106_2247 ();
 FILLCELL_X32 FILLER_106_2279 ();
 FILLCELL_X32 FILLER_106_2311 ();
 FILLCELL_X32 FILLER_106_2343 ();
 FILLCELL_X32 FILLER_106_2375 ();
 FILLCELL_X32 FILLER_106_2407 ();
 FILLCELL_X32 FILLER_106_2439 ();
 FILLCELL_X32 FILLER_106_2471 ();
 FILLCELL_X32 FILLER_106_2503 ();
 FILLCELL_X32 FILLER_106_2535 ();
 FILLCELL_X32 FILLER_106_2567 ();
 FILLCELL_X2 FILLER_106_2599 ();
 FILLCELL_X1 FILLER_106_2601 ();
 FILLCELL_X32 FILLER_107_1 ();
 FILLCELL_X32 FILLER_107_33 ();
 FILLCELL_X32 FILLER_107_65 ();
 FILLCELL_X32 FILLER_107_97 ();
 FILLCELL_X32 FILLER_107_129 ();
 FILLCELL_X32 FILLER_107_161 ();
 FILLCELL_X32 FILLER_107_193 ();
 FILLCELL_X32 FILLER_107_225 ();
 FILLCELL_X32 FILLER_107_257 ();
 FILLCELL_X32 FILLER_107_289 ();
 FILLCELL_X32 FILLER_107_321 ();
 FILLCELL_X32 FILLER_107_353 ();
 FILLCELL_X32 FILLER_107_385 ();
 FILLCELL_X32 FILLER_107_417 ();
 FILLCELL_X32 FILLER_107_449 ();
 FILLCELL_X32 FILLER_107_481 ();
 FILLCELL_X32 FILLER_107_513 ();
 FILLCELL_X32 FILLER_107_545 ();
 FILLCELL_X32 FILLER_107_577 ();
 FILLCELL_X32 FILLER_107_609 ();
 FILLCELL_X32 FILLER_107_641 ();
 FILLCELL_X32 FILLER_107_673 ();
 FILLCELL_X32 FILLER_107_705 ();
 FILLCELL_X32 FILLER_107_737 ();
 FILLCELL_X32 FILLER_107_769 ();
 FILLCELL_X32 FILLER_107_801 ();
 FILLCELL_X32 FILLER_107_833 ();
 FILLCELL_X32 FILLER_107_865 ();
 FILLCELL_X32 FILLER_107_897 ();
 FILLCELL_X32 FILLER_107_929 ();
 FILLCELL_X32 FILLER_107_961 ();
 FILLCELL_X32 FILLER_107_993 ();
 FILLCELL_X32 FILLER_107_1025 ();
 FILLCELL_X32 FILLER_107_1057 ();
 FILLCELL_X32 FILLER_107_1089 ();
 FILLCELL_X32 FILLER_107_1121 ();
 FILLCELL_X32 FILLER_107_1153 ();
 FILLCELL_X32 FILLER_107_1185 ();
 FILLCELL_X32 FILLER_107_1217 ();
 FILLCELL_X8 FILLER_107_1249 ();
 FILLCELL_X4 FILLER_107_1257 ();
 FILLCELL_X2 FILLER_107_1261 ();
 FILLCELL_X32 FILLER_107_1264 ();
 FILLCELL_X32 FILLER_107_1296 ();
 FILLCELL_X32 FILLER_107_1328 ();
 FILLCELL_X32 FILLER_107_1360 ();
 FILLCELL_X32 FILLER_107_1392 ();
 FILLCELL_X32 FILLER_107_1424 ();
 FILLCELL_X32 FILLER_107_1456 ();
 FILLCELL_X32 FILLER_107_1488 ();
 FILLCELL_X32 FILLER_107_1520 ();
 FILLCELL_X32 FILLER_107_1552 ();
 FILLCELL_X32 FILLER_107_1584 ();
 FILLCELL_X32 FILLER_107_1616 ();
 FILLCELL_X32 FILLER_107_1648 ();
 FILLCELL_X32 FILLER_107_1680 ();
 FILLCELL_X32 FILLER_107_1712 ();
 FILLCELL_X32 FILLER_107_1744 ();
 FILLCELL_X32 FILLER_107_1776 ();
 FILLCELL_X32 FILLER_107_1808 ();
 FILLCELL_X32 FILLER_107_1840 ();
 FILLCELL_X32 FILLER_107_1872 ();
 FILLCELL_X32 FILLER_107_1904 ();
 FILLCELL_X32 FILLER_107_1936 ();
 FILLCELL_X32 FILLER_107_1968 ();
 FILLCELL_X32 FILLER_107_2000 ();
 FILLCELL_X32 FILLER_107_2032 ();
 FILLCELL_X32 FILLER_107_2064 ();
 FILLCELL_X32 FILLER_107_2096 ();
 FILLCELL_X32 FILLER_107_2128 ();
 FILLCELL_X32 FILLER_107_2160 ();
 FILLCELL_X32 FILLER_107_2192 ();
 FILLCELL_X32 FILLER_107_2224 ();
 FILLCELL_X32 FILLER_107_2256 ();
 FILLCELL_X32 FILLER_107_2288 ();
 FILLCELL_X32 FILLER_107_2320 ();
 FILLCELL_X32 FILLER_107_2352 ();
 FILLCELL_X32 FILLER_107_2384 ();
 FILLCELL_X32 FILLER_107_2416 ();
 FILLCELL_X32 FILLER_107_2448 ();
 FILLCELL_X32 FILLER_107_2480 ();
 FILLCELL_X8 FILLER_107_2512 ();
 FILLCELL_X4 FILLER_107_2520 ();
 FILLCELL_X2 FILLER_107_2524 ();
 FILLCELL_X32 FILLER_107_2527 ();
 FILLCELL_X32 FILLER_107_2559 ();
 FILLCELL_X8 FILLER_107_2591 ();
 FILLCELL_X2 FILLER_107_2599 ();
 FILLCELL_X1 FILLER_107_2601 ();
 FILLCELL_X32 FILLER_108_1 ();
 FILLCELL_X32 FILLER_108_33 ();
 FILLCELL_X32 FILLER_108_65 ();
 FILLCELL_X32 FILLER_108_97 ();
 FILLCELL_X32 FILLER_108_129 ();
 FILLCELL_X32 FILLER_108_161 ();
 FILLCELL_X32 FILLER_108_193 ();
 FILLCELL_X32 FILLER_108_225 ();
 FILLCELL_X32 FILLER_108_257 ();
 FILLCELL_X32 FILLER_108_289 ();
 FILLCELL_X32 FILLER_108_321 ();
 FILLCELL_X32 FILLER_108_353 ();
 FILLCELL_X32 FILLER_108_385 ();
 FILLCELL_X32 FILLER_108_417 ();
 FILLCELL_X32 FILLER_108_449 ();
 FILLCELL_X32 FILLER_108_481 ();
 FILLCELL_X32 FILLER_108_513 ();
 FILLCELL_X32 FILLER_108_545 ();
 FILLCELL_X32 FILLER_108_577 ();
 FILLCELL_X16 FILLER_108_609 ();
 FILLCELL_X4 FILLER_108_625 ();
 FILLCELL_X2 FILLER_108_629 ();
 FILLCELL_X32 FILLER_108_632 ();
 FILLCELL_X32 FILLER_108_664 ();
 FILLCELL_X32 FILLER_108_696 ();
 FILLCELL_X32 FILLER_108_728 ();
 FILLCELL_X32 FILLER_108_760 ();
 FILLCELL_X32 FILLER_108_792 ();
 FILLCELL_X32 FILLER_108_824 ();
 FILLCELL_X32 FILLER_108_856 ();
 FILLCELL_X32 FILLER_108_888 ();
 FILLCELL_X32 FILLER_108_920 ();
 FILLCELL_X32 FILLER_108_952 ();
 FILLCELL_X32 FILLER_108_984 ();
 FILLCELL_X32 FILLER_108_1016 ();
 FILLCELL_X32 FILLER_108_1048 ();
 FILLCELL_X32 FILLER_108_1080 ();
 FILLCELL_X32 FILLER_108_1112 ();
 FILLCELL_X32 FILLER_108_1144 ();
 FILLCELL_X32 FILLER_108_1176 ();
 FILLCELL_X32 FILLER_108_1208 ();
 FILLCELL_X32 FILLER_108_1240 ();
 FILLCELL_X32 FILLER_108_1272 ();
 FILLCELL_X32 FILLER_108_1304 ();
 FILLCELL_X32 FILLER_108_1336 ();
 FILLCELL_X32 FILLER_108_1368 ();
 FILLCELL_X32 FILLER_108_1400 ();
 FILLCELL_X32 FILLER_108_1432 ();
 FILLCELL_X32 FILLER_108_1464 ();
 FILLCELL_X32 FILLER_108_1496 ();
 FILLCELL_X32 FILLER_108_1528 ();
 FILLCELL_X32 FILLER_108_1560 ();
 FILLCELL_X32 FILLER_108_1592 ();
 FILLCELL_X32 FILLER_108_1624 ();
 FILLCELL_X32 FILLER_108_1656 ();
 FILLCELL_X32 FILLER_108_1688 ();
 FILLCELL_X32 FILLER_108_1720 ();
 FILLCELL_X32 FILLER_108_1752 ();
 FILLCELL_X32 FILLER_108_1784 ();
 FILLCELL_X32 FILLER_108_1816 ();
 FILLCELL_X32 FILLER_108_1848 ();
 FILLCELL_X8 FILLER_108_1880 ();
 FILLCELL_X4 FILLER_108_1888 ();
 FILLCELL_X2 FILLER_108_1892 ();
 FILLCELL_X32 FILLER_108_1895 ();
 FILLCELL_X32 FILLER_108_1927 ();
 FILLCELL_X32 FILLER_108_1959 ();
 FILLCELL_X32 FILLER_108_1991 ();
 FILLCELL_X32 FILLER_108_2023 ();
 FILLCELL_X32 FILLER_108_2055 ();
 FILLCELL_X32 FILLER_108_2087 ();
 FILLCELL_X32 FILLER_108_2119 ();
 FILLCELL_X32 FILLER_108_2151 ();
 FILLCELL_X32 FILLER_108_2183 ();
 FILLCELL_X32 FILLER_108_2215 ();
 FILLCELL_X32 FILLER_108_2247 ();
 FILLCELL_X32 FILLER_108_2279 ();
 FILLCELL_X32 FILLER_108_2311 ();
 FILLCELL_X32 FILLER_108_2343 ();
 FILLCELL_X32 FILLER_108_2375 ();
 FILLCELL_X32 FILLER_108_2407 ();
 FILLCELL_X32 FILLER_108_2439 ();
 FILLCELL_X32 FILLER_108_2471 ();
 FILLCELL_X32 FILLER_108_2503 ();
 FILLCELL_X32 FILLER_108_2535 ();
 FILLCELL_X32 FILLER_108_2567 ();
 FILLCELL_X2 FILLER_108_2599 ();
 FILLCELL_X1 FILLER_108_2601 ();
 FILLCELL_X32 FILLER_109_1 ();
 FILLCELL_X32 FILLER_109_33 ();
 FILLCELL_X32 FILLER_109_65 ();
 FILLCELL_X32 FILLER_109_97 ();
 FILLCELL_X32 FILLER_109_129 ();
 FILLCELL_X32 FILLER_109_161 ();
 FILLCELL_X32 FILLER_109_193 ();
 FILLCELL_X32 FILLER_109_225 ();
 FILLCELL_X32 FILLER_109_257 ();
 FILLCELL_X32 FILLER_109_289 ();
 FILLCELL_X32 FILLER_109_321 ();
 FILLCELL_X32 FILLER_109_353 ();
 FILLCELL_X32 FILLER_109_385 ();
 FILLCELL_X32 FILLER_109_417 ();
 FILLCELL_X32 FILLER_109_449 ();
 FILLCELL_X32 FILLER_109_481 ();
 FILLCELL_X32 FILLER_109_513 ();
 FILLCELL_X32 FILLER_109_545 ();
 FILLCELL_X32 FILLER_109_577 ();
 FILLCELL_X32 FILLER_109_609 ();
 FILLCELL_X32 FILLER_109_641 ();
 FILLCELL_X32 FILLER_109_673 ();
 FILLCELL_X32 FILLER_109_705 ();
 FILLCELL_X32 FILLER_109_737 ();
 FILLCELL_X32 FILLER_109_769 ();
 FILLCELL_X32 FILLER_109_801 ();
 FILLCELL_X32 FILLER_109_833 ();
 FILLCELL_X32 FILLER_109_865 ();
 FILLCELL_X32 FILLER_109_897 ();
 FILLCELL_X32 FILLER_109_929 ();
 FILLCELL_X32 FILLER_109_961 ();
 FILLCELL_X32 FILLER_109_993 ();
 FILLCELL_X32 FILLER_109_1025 ();
 FILLCELL_X32 FILLER_109_1057 ();
 FILLCELL_X32 FILLER_109_1089 ();
 FILLCELL_X32 FILLER_109_1121 ();
 FILLCELL_X32 FILLER_109_1153 ();
 FILLCELL_X32 FILLER_109_1185 ();
 FILLCELL_X32 FILLER_109_1217 ();
 FILLCELL_X8 FILLER_109_1249 ();
 FILLCELL_X4 FILLER_109_1257 ();
 FILLCELL_X2 FILLER_109_1261 ();
 FILLCELL_X32 FILLER_109_1264 ();
 FILLCELL_X32 FILLER_109_1296 ();
 FILLCELL_X32 FILLER_109_1328 ();
 FILLCELL_X32 FILLER_109_1360 ();
 FILLCELL_X32 FILLER_109_1392 ();
 FILLCELL_X32 FILLER_109_1424 ();
 FILLCELL_X32 FILLER_109_1456 ();
 FILLCELL_X32 FILLER_109_1488 ();
 FILLCELL_X32 FILLER_109_1520 ();
 FILLCELL_X32 FILLER_109_1552 ();
 FILLCELL_X32 FILLER_109_1584 ();
 FILLCELL_X32 FILLER_109_1616 ();
 FILLCELL_X32 FILLER_109_1648 ();
 FILLCELL_X32 FILLER_109_1680 ();
 FILLCELL_X32 FILLER_109_1712 ();
 FILLCELL_X32 FILLER_109_1744 ();
 FILLCELL_X32 FILLER_109_1776 ();
 FILLCELL_X32 FILLER_109_1808 ();
 FILLCELL_X32 FILLER_109_1840 ();
 FILLCELL_X32 FILLER_109_1872 ();
 FILLCELL_X32 FILLER_109_1904 ();
 FILLCELL_X32 FILLER_109_1936 ();
 FILLCELL_X32 FILLER_109_1968 ();
 FILLCELL_X32 FILLER_109_2000 ();
 FILLCELL_X32 FILLER_109_2032 ();
 FILLCELL_X32 FILLER_109_2064 ();
 FILLCELL_X32 FILLER_109_2096 ();
 FILLCELL_X32 FILLER_109_2128 ();
 FILLCELL_X32 FILLER_109_2160 ();
 FILLCELL_X32 FILLER_109_2192 ();
 FILLCELL_X32 FILLER_109_2224 ();
 FILLCELL_X32 FILLER_109_2256 ();
 FILLCELL_X32 FILLER_109_2288 ();
 FILLCELL_X32 FILLER_109_2320 ();
 FILLCELL_X32 FILLER_109_2352 ();
 FILLCELL_X32 FILLER_109_2384 ();
 FILLCELL_X32 FILLER_109_2416 ();
 FILLCELL_X32 FILLER_109_2448 ();
 FILLCELL_X32 FILLER_109_2480 ();
 FILLCELL_X8 FILLER_109_2512 ();
 FILLCELL_X4 FILLER_109_2520 ();
 FILLCELL_X2 FILLER_109_2524 ();
 FILLCELL_X32 FILLER_109_2527 ();
 FILLCELL_X32 FILLER_109_2559 ();
 FILLCELL_X8 FILLER_109_2591 ();
 FILLCELL_X2 FILLER_109_2599 ();
 FILLCELL_X1 FILLER_109_2601 ();
 FILLCELL_X32 FILLER_110_1 ();
 FILLCELL_X32 FILLER_110_33 ();
 FILLCELL_X32 FILLER_110_65 ();
 FILLCELL_X32 FILLER_110_97 ();
 FILLCELL_X32 FILLER_110_129 ();
 FILLCELL_X32 FILLER_110_161 ();
 FILLCELL_X32 FILLER_110_193 ();
 FILLCELL_X32 FILLER_110_225 ();
 FILLCELL_X32 FILLER_110_257 ();
 FILLCELL_X32 FILLER_110_289 ();
 FILLCELL_X32 FILLER_110_321 ();
 FILLCELL_X32 FILLER_110_353 ();
 FILLCELL_X32 FILLER_110_385 ();
 FILLCELL_X32 FILLER_110_417 ();
 FILLCELL_X32 FILLER_110_449 ();
 FILLCELL_X32 FILLER_110_481 ();
 FILLCELL_X32 FILLER_110_513 ();
 FILLCELL_X32 FILLER_110_545 ();
 FILLCELL_X32 FILLER_110_577 ();
 FILLCELL_X16 FILLER_110_609 ();
 FILLCELL_X4 FILLER_110_625 ();
 FILLCELL_X2 FILLER_110_629 ();
 FILLCELL_X32 FILLER_110_632 ();
 FILLCELL_X32 FILLER_110_664 ();
 FILLCELL_X32 FILLER_110_696 ();
 FILLCELL_X32 FILLER_110_728 ();
 FILLCELL_X32 FILLER_110_760 ();
 FILLCELL_X32 FILLER_110_792 ();
 FILLCELL_X32 FILLER_110_824 ();
 FILLCELL_X32 FILLER_110_856 ();
 FILLCELL_X32 FILLER_110_888 ();
 FILLCELL_X32 FILLER_110_920 ();
 FILLCELL_X32 FILLER_110_952 ();
 FILLCELL_X32 FILLER_110_984 ();
 FILLCELL_X32 FILLER_110_1016 ();
 FILLCELL_X32 FILLER_110_1048 ();
 FILLCELL_X32 FILLER_110_1080 ();
 FILLCELL_X32 FILLER_110_1112 ();
 FILLCELL_X32 FILLER_110_1144 ();
 FILLCELL_X32 FILLER_110_1176 ();
 FILLCELL_X32 FILLER_110_1208 ();
 FILLCELL_X32 FILLER_110_1240 ();
 FILLCELL_X32 FILLER_110_1272 ();
 FILLCELL_X32 FILLER_110_1304 ();
 FILLCELL_X32 FILLER_110_1336 ();
 FILLCELL_X32 FILLER_110_1368 ();
 FILLCELL_X32 FILLER_110_1400 ();
 FILLCELL_X32 FILLER_110_1432 ();
 FILLCELL_X32 FILLER_110_1464 ();
 FILLCELL_X32 FILLER_110_1496 ();
 FILLCELL_X32 FILLER_110_1528 ();
 FILLCELL_X32 FILLER_110_1560 ();
 FILLCELL_X32 FILLER_110_1592 ();
 FILLCELL_X32 FILLER_110_1624 ();
 FILLCELL_X32 FILLER_110_1656 ();
 FILLCELL_X32 FILLER_110_1688 ();
 FILLCELL_X32 FILLER_110_1720 ();
 FILLCELL_X32 FILLER_110_1752 ();
 FILLCELL_X32 FILLER_110_1784 ();
 FILLCELL_X32 FILLER_110_1816 ();
 FILLCELL_X32 FILLER_110_1848 ();
 FILLCELL_X8 FILLER_110_1880 ();
 FILLCELL_X4 FILLER_110_1888 ();
 FILLCELL_X2 FILLER_110_1892 ();
 FILLCELL_X32 FILLER_110_1895 ();
 FILLCELL_X32 FILLER_110_1927 ();
 FILLCELL_X32 FILLER_110_1959 ();
 FILLCELL_X32 FILLER_110_1991 ();
 FILLCELL_X32 FILLER_110_2023 ();
 FILLCELL_X32 FILLER_110_2055 ();
 FILLCELL_X32 FILLER_110_2087 ();
 FILLCELL_X32 FILLER_110_2119 ();
 FILLCELL_X32 FILLER_110_2151 ();
 FILLCELL_X32 FILLER_110_2183 ();
 FILLCELL_X32 FILLER_110_2215 ();
 FILLCELL_X32 FILLER_110_2247 ();
 FILLCELL_X32 FILLER_110_2279 ();
 FILLCELL_X32 FILLER_110_2311 ();
 FILLCELL_X32 FILLER_110_2343 ();
 FILLCELL_X32 FILLER_110_2375 ();
 FILLCELL_X32 FILLER_110_2407 ();
 FILLCELL_X32 FILLER_110_2439 ();
 FILLCELL_X32 FILLER_110_2471 ();
 FILLCELL_X32 FILLER_110_2503 ();
 FILLCELL_X32 FILLER_110_2535 ();
 FILLCELL_X32 FILLER_110_2567 ();
 FILLCELL_X2 FILLER_110_2599 ();
 FILLCELL_X1 FILLER_110_2601 ();
 FILLCELL_X32 FILLER_111_1 ();
 FILLCELL_X32 FILLER_111_33 ();
 FILLCELL_X32 FILLER_111_65 ();
 FILLCELL_X32 FILLER_111_97 ();
 FILLCELL_X32 FILLER_111_129 ();
 FILLCELL_X32 FILLER_111_161 ();
 FILLCELL_X32 FILLER_111_193 ();
 FILLCELL_X32 FILLER_111_225 ();
 FILLCELL_X32 FILLER_111_257 ();
 FILLCELL_X32 FILLER_111_289 ();
 FILLCELL_X32 FILLER_111_321 ();
 FILLCELL_X32 FILLER_111_353 ();
 FILLCELL_X32 FILLER_111_385 ();
 FILLCELL_X32 FILLER_111_417 ();
 FILLCELL_X32 FILLER_111_449 ();
 FILLCELL_X32 FILLER_111_481 ();
 FILLCELL_X32 FILLER_111_513 ();
 FILLCELL_X32 FILLER_111_545 ();
 FILLCELL_X32 FILLER_111_577 ();
 FILLCELL_X32 FILLER_111_609 ();
 FILLCELL_X32 FILLER_111_641 ();
 FILLCELL_X32 FILLER_111_673 ();
 FILLCELL_X32 FILLER_111_705 ();
 FILLCELL_X32 FILLER_111_737 ();
 FILLCELL_X32 FILLER_111_769 ();
 FILLCELL_X32 FILLER_111_801 ();
 FILLCELL_X32 FILLER_111_833 ();
 FILLCELL_X32 FILLER_111_865 ();
 FILLCELL_X32 FILLER_111_897 ();
 FILLCELL_X32 FILLER_111_929 ();
 FILLCELL_X32 FILLER_111_961 ();
 FILLCELL_X32 FILLER_111_993 ();
 FILLCELL_X32 FILLER_111_1025 ();
 FILLCELL_X32 FILLER_111_1057 ();
 FILLCELL_X32 FILLER_111_1089 ();
 FILLCELL_X32 FILLER_111_1121 ();
 FILLCELL_X32 FILLER_111_1153 ();
 FILLCELL_X32 FILLER_111_1185 ();
 FILLCELL_X32 FILLER_111_1217 ();
 FILLCELL_X8 FILLER_111_1249 ();
 FILLCELL_X4 FILLER_111_1257 ();
 FILLCELL_X2 FILLER_111_1261 ();
 FILLCELL_X32 FILLER_111_1264 ();
 FILLCELL_X32 FILLER_111_1296 ();
 FILLCELL_X32 FILLER_111_1328 ();
 FILLCELL_X32 FILLER_111_1360 ();
 FILLCELL_X32 FILLER_111_1392 ();
 FILLCELL_X32 FILLER_111_1424 ();
 FILLCELL_X32 FILLER_111_1456 ();
 FILLCELL_X32 FILLER_111_1488 ();
 FILLCELL_X32 FILLER_111_1520 ();
 FILLCELL_X32 FILLER_111_1552 ();
 FILLCELL_X32 FILLER_111_1584 ();
 FILLCELL_X32 FILLER_111_1616 ();
 FILLCELL_X32 FILLER_111_1648 ();
 FILLCELL_X32 FILLER_111_1680 ();
 FILLCELL_X32 FILLER_111_1712 ();
 FILLCELL_X32 FILLER_111_1744 ();
 FILLCELL_X32 FILLER_111_1776 ();
 FILLCELL_X32 FILLER_111_1808 ();
 FILLCELL_X32 FILLER_111_1840 ();
 FILLCELL_X32 FILLER_111_1872 ();
 FILLCELL_X32 FILLER_111_1904 ();
 FILLCELL_X32 FILLER_111_1936 ();
 FILLCELL_X32 FILLER_111_1968 ();
 FILLCELL_X32 FILLER_111_2000 ();
 FILLCELL_X32 FILLER_111_2032 ();
 FILLCELL_X32 FILLER_111_2064 ();
 FILLCELL_X32 FILLER_111_2096 ();
 FILLCELL_X32 FILLER_111_2128 ();
 FILLCELL_X32 FILLER_111_2160 ();
 FILLCELL_X32 FILLER_111_2192 ();
 FILLCELL_X32 FILLER_111_2224 ();
 FILLCELL_X32 FILLER_111_2256 ();
 FILLCELL_X32 FILLER_111_2288 ();
 FILLCELL_X32 FILLER_111_2320 ();
 FILLCELL_X32 FILLER_111_2352 ();
 FILLCELL_X32 FILLER_111_2384 ();
 FILLCELL_X32 FILLER_111_2416 ();
 FILLCELL_X32 FILLER_111_2448 ();
 FILLCELL_X32 FILLER_111_2480 ();
 FILLCELL_X8 FILLER_111_2512 ();
 FILLCELL_X4 FILLER_111_2520 ();
 FILLCELL_X2 FILLER_111_2524 ();
 FILLCELL_X32 FILLER_111_2527 ();
 FILLCELL_X32 FILLER_111_2559 ();
 FILLCELL_X8 FILLER_111_2591 ();
 FILLCELL_X2 FILLER_111_2599 ();
 FILLCELL_X1 FILLER_111_2601 ();
 FILLCELL_X32 FILLER_112_1 ();
 FILLCELL_X32 FILLER_112_33 ();
 FILLCELL_X32 FILLER_112_65 ();
 FILLCELL_X32 FILLER_112_97 ();
 FILLCELL_X32 FILLER_112_129 ();
 FILLCELL_X32 FILLER_112_161 ();
 FILLCELL_X32 FILLER_112_193 ();
 FILLCELL_X32 FILLER_112_225 ();
 FILLCELL_X32 FILLER_112_257 ();
 FILLCELL_X32 FILLER_112_289 ();
 FILLCELL_X32 FILLER_112_321 ();
 FILLCELL_X32 FILLER_112_353 ();
 FILLCELL_X32 FILLER_112_385 ();
 FILLCELL_X32 FILLER_112_417 ();
 FILLCELL_X32 FILLER_112_449 ();
 FILLCELL_X32 FILLER_112_481 ();
 FILLCELL_X32 FILLER_112_513 ();
 FILLCELL_X32 FILLER_112_545 ();
 FILLCELL_X32 FILLER_112_577 ();
 FILLCELL_X16 FILLER_112_609 ();
 FILLCELL_X4 FILLER_112_625 ();
 FILLCELL_X2 FILLER_112_629 ();
 FILLCELL_X32 FILLER_112_632 ();
 FILLCELL_X32 FILLER_112_664 ();
 FILLCELL_X32 FILLER_112_696 ();
 FILLCELL_X32 FILLER_112_728 ();
 FILLCELL_X32 FILLER_112_760 ();
 FILLCELL_X32 FILLER_112_792 ();
 FILLCELL_X32 FILLER_112_824 ();
 FILLCELL_X32 FILLER_112_856 ();
 FILLCELL_X32 FILLER_112_888 ();
 FILLCELL_X32 FILLER_112_920 ();
 FILLCELL_X32 FILLER_112_952 ();
 FILLCELL_X32 FILLER_112_984 ();
 FILLCELL_X32 FILLER_112_1016 ();
 FILLCELL_X32 FILLER_112_1048 ();
 FILLCELL_X32 FILLER_112_1080 ();
 FILLCELL_X32 FILLER_112_1112 ();
 FILLCELL_X32 FILLER_112_1144 ();
 FILLCELL_X32 FILLER_112_1176 ();
 FILLCELL_X32 FILLER_112_1208 ();
 FILLCELL_X32 FILLER_112_1240 ();
 FILLCELL_X32 FILLER_112_1272 ();
 FILLCELL_X32 FILLER_112_1304 ();
 FILLCELL_X32 FILLER_112_1336 ();
 FILLCELL_X32 FILLER_112_1368 ();
 FILLCELL_X32 FILLER_112_1400 ();
 FILLCELL_X32 FILLER_112_1432 ();
 FILLCELL_X32 FILLER_112_1464 ();
 FILLCELL_X32 FILLER_112_1496 ();
 FILLCELL_X32 FILLER_112_1528 ();
 FILLCELL_X32 FILLER_112_1560 ();
 FILLCELL_X32 FILLER_112_1592 ();
 FILLCELL_X32 FILLER_112_1624 ();
 FILLCELL_X32 FILLER_112_1656 ();
 FILLCELL_X32 FILLER_112_1688 ();
 FILLCELL_X32 FILLER_112_1720 ();
 FILLCELL_X32 FILLER_112_1752 ();
 FILLCELL_X32 FILLER_112_1784 ();
 FILLCELL_X32 FILLER_112_1816 ();
 FILLCELL_X32 FILLER_112_1848 ();
 FILLCELL_X8 FILLER_112_1880 ();
 FILLCELL_X4 FILLER_112_1888 ();
 FILLCELL_X2 FILLER_112_1892 ();
 FILLCELL_X32 FILLER_112_1895 ();
 FILLCELL_X32 FILLER_112_1927 ();
 FILLCELL_X32 FILLER_112_1959 ();
 FILLCELL_X32 FILLER_112_1991 ();
 FILLCELL_X32 FILLER_112_2023 ();
 FILLCELL_X32 FILLER_112_2055 ();
 FILLCELL_X32 FILLER_112_2087 ();
 FILLCELL_X32 FILLER_112_2119 ();
 FILLCELL_X32 FILLER_112_2151 ();
 FILLCELL_X32 FILLER_112_2183 ();
 FILLCELL_X32 FILLER_112_2215 ();
 FILLCELL_X32 FILLER_112_2247 ();
 FILLCELL_X32 FILLER_112_2279 ();
 FILLCELL_X32 FILLER_112_2311 ();
 FILLCELL_X32 FILLER_112_2343 ();
 FILLCELL_X32 FILLER_112_2375 ();
 FILLCELL_X32 FILLER_112_2407 ();
 FILLCELL_X32 FILLER_112_2439 ();
 FILLCELL_X32 FILLER_112_2471 ();
 FILLCELL_X32 FILLER_112_2503 ();
 FILLCELL_X32 FILLER_112_2535 ();
 FILLCELL_X32 FILLER_112_2567 ();
 FILLCELL_X2 FILLER_112_2599 ();
 FILLCELL_X1 FILLER_112_2601 ();
 FILLCELL_X32 FILLER_113_1 ();
 FILLCELL_X32 FILLER_113_33 ();
 FILLCELL_X32 FILLER_113_65 ();
 FILLCELL_X32 FILLER_113_97 ();
 FILLCELL_X32 FILLER_113_129 ();
 FILLCELL_X32 FILLER_113_161 ();
 FILLCELL_X32 FILLER_113_193 ();
 FILLCELL_X32 FILLER_113_225 ();
 FILLCELL_X32 FILLER_113_257 ();
 FILLCELL_X32 FILLER_113_289 ();
 FILLCELL_X32 FILLER_113_321 ();
 FILLCELL_X32 FILLER_113_353 ();
 FILLCELL_X32 FILLER_113_385 ();
 FILLCELL_X32 FILLER_113_417 ();
 FILLCELL_X32 FILLER_113_449 ();
 FILLCELL_X32 FILLER_113_481 ();
 FILLCELL_X32 FILLER_113_513 ();
 FILLCELL_X32 FILLER_113_545 ();
 FILLCELL_X32 FILLER_113_577 ();
 FILLCELL_X32 FILLER_113_609 ();
 FILLCELL_X32 FILLER_113_641 ();
 FILLCELL_X32 FILLER_113_673 ();
 FILLCELL_X32 FILLER_113_705 ();
 FILLCELL_X32 FILLER_113_737 ();
 FILLCELL_X32 FILLER_113_769 ();
 FILLCELL_X32 FILLER_113_801 ();
 FILLCELL_X32 FILLER_113_833 ();
 FILLCELL_X32 FILLER_113_865 ();
 FILLCELL_X32 FILLER_113_897 ();
 FILLCELL_X32 FILLER_113_929 ();
 FILLCELL_X32 FILLER_113_961 ();
 FILLCELL_X32 FILLER_113_993 ();
 FILLCELL_X32 FILLER_113_1025 ();
 FILLCELL_X32 FILLER_113_1057 ();
 FILLCELL_X32 FILLER_113_1089 ();
 FILLCELL_X32 FILLER_113_1121 ();
 FILLCELL_X32 FILLER_113_1153 ();
 FILLCELL_X32 FILLER_113_1185 ();
 FILLCELL_X32 FILLER_113_1217 ();
 FILLCELL_X8 FILLER_113_1249 ();
 FILLCELL_X4 FILLER_113_1257 ();
 FILLCELL_X2 FILLER_113_1261 ();
 FILLCELL_X32 FILLER_113_1264 ();
 FILLCELL_X32 FILLER_113_1296 ();
 FILLCELL_X32 FILLER_113_1328 ();
 FILLCELL_X32 FILLER_113_1360 ();
 FILLCELL_X32 FILLER_113_1392 ();
 FILLCELL_X32 FILLER_113_1424 ();
 FILLCELL_X32 FILLER_113_1456 ();
 FILLCELL_X32 FILLER_113_1488 ();
 FILLCELL_X32 FILLER_113_1520 ();
 FILLCELL_X32 FILLER_113_1552 ();
 FILLCELL_X32 FILLER_113_1584 ();
 FILLCELL_X32 FILLER_113_1616 ();
 FILLCELL_X32 FILLER_113_1648 ();
 FILLCELL_X32 FILLER_113_1680 ();
 FILLCELL_X32 FILLER_113_1712 ();
 FILLCELL_X32 FILLER_113_1744 ();
 FILLCELL_X32 FILLER_113_1776 ();
 FILLCELL_X32 FILLER_113_1808 ();
 FILLCELL_X32 FILLER_113_1840 ();
 FILLCELL_X32 FILLER_113_1872 ();
 FILLCELL_X32 FILLER_113_1904 ();
 FILLCELL_X32 FILLER_113_1936 ();
 FILLCELL_X32 FILLER_113_1968 ();
 FILLCELL_X32 FILLER_113_2000 ();
 FILLCELL_X32 FILLER_113_2032 ();
 FILLCELL_X32 FILLER_113_2064 ();
 FILLCELL_X32 FILLER_113_2096 ();
 FILLCELL_X32 FILLER_113_2128 ();
 FILLCELL_X32 FILLER_113_2160 ();
 FILLCELL_X32 FILLER_113_2192 ();
 FILLCELL_X32 FILLER_113_2224 ();
 FILLCELL_X32 FILLER_113_2256 ();
 FILLCELL_X32 FILLER_113_2288 ();
 FILLCELL_X32 FILLER_113_2320 ();
 FILLCELL_X32 FILLER_113_2352 ();
 FILLCELL_X32 FILLER_113_2384 ();
 FILLCELL_X32 FILLER_113_2416 ();
 FILLCELL_X32 FILLER_113_2448 ();
 FILLCELL_X32 FILLER_113_2480 ();
 FILLCELL_X8 FILLER_113_2512 ();
 FILLCELL_X4 FILLER_113_2520 ();
 FILLCELL_X2 FILLER_113_2524 ();
 FILLCELL_X32 FILLER_113_2527 ();
 FILLCELL_X32 FILLER_113_2559 ();
 FILLCELL_X8 FILLER_113_2591 ();
 FILLCELL_X2 FILLER_113_2599 ();
 FILLCELL_X1 FILLER_113_2601 ();
 FILLCELL_X32 FILLER_114_1 ();
 FILLCELL_X32 FILLER_114_33 ();
 FILLCELL_X32 FILLER_114_65 ();
 FILLCELL_X32 FILLER_114_97 ();
 FILLCELL_X32 FILLER_114_129 ();
 FILLCELL_X32 FILLER_114_161 ();
 FILLCELL_X32 FILLER_114_193 ();
 FILLCELL_X32 FILLER_114_225 ();
 FILLCELL_X32 FILLER_114_257 ();
 FILLCELL_X32 FILLER_114_289 ();
 FILLCELL_X32 FILLER_114_321 ();
 FILLCELL_X32 FILLER_114_353 ();
 FILLCELL_X32 FILLER_114_385 ();
 FILLCELL_X32 FILLER_114_417 ();
 FILLCELL_X32 FILLER_114_449 ();
 FILLCELL_X32 FILLER_114_481 ();
 FILLCELL_X32 FILLER_114_513 ();
 FILLCELL_X32 FILLER_114_545 ();
 FILLCELL_X32 FILLER_114_577 ();
 FILLCELL_X16 FILLER_114_609 ();
 FILLCELL_X4 FILLER_114_625 ();
 FILLCELL_X2 FILLER_114_629 ();
 FILLCELL_X32 FILLER_114_632 ();
 FILLCELL_X32 FILLER_114_664 ();
 FILLCELL_X32 FILLER_114_696 ();
 FILLCELL_X32 FILLER_114_728 ();
 FILLCELL_X32 FILLER_114_760 ();
 FILLCELL_X32 FILLER_114_792 ();
 FILLCELL_X32 FILLER_114_824 ();
 FILLCELL_X32 FILLER_114_856 ();
 FILLCELL_X32 FILLER_114_888 ();
 FILLCELL_X32 FILLER_114_920 ();
 FILLCELL_X32 FILLER_114_952 ();
 FILLCELL_X32 FILLER_114_984 ();
 FILLCELL_X32 FILLER_114_1016 ();
 FILLCELL_X32 FILLER_114_1048 ();
 FILLCELL_X32 FILLER_114_1080 ();
 FILLCELL_X32 FILLER_114_1112 ();
 FILLCELL_X32 FILLER_114_1144 ();
 FILLCELL_X32 FILLER_114_1176 ();
 FILLCELL_X32 FILLER_114_1208 ();
 FILLCELL_X32 FILLER_114_1240 ();
 FILLCELL_X32 FILLER_114_1272 ();
 FILLCELL_X32 FILLER_114_1304 ();
 FILLCELL_X32 FILLER_114_1336 ();
 FILLCELL_X32 FILLER_114_1368 ();
 FILLCELL_X32 FILLER_114_1400 ();
 FILLCELL_X32 FILLER_114_1432 ();
 FILLCELL_X32 FILLER_114_1464 ();
 FILLCELL_X32 FILLER_114_1496 ();
 FILLCELL_X32 FILLER_114_1528 ();
 FILLCELL_X32 FILLER_114_1560 ();
 FILLCELL_X32 FILLER_114_1592 ();
 FILLCELL_X32 FILLER_114_1624 ();
 FILLCELL_X32 FILLER_114_1656 ();
 FILLCELL_X32 FILLER_114_1688 ();
 FILLCELL_X32 FILLER_114_1720 ();
 FILLCELL_X32 FILLER_114_1752 ();
 FILLCELL_X32 FILLER_114_1784 ();
 FILLCELL_X32 FILLER_114_1816 ();
 FILLCELL_X32 FILLER_114_1848 ();
 FILLCELL_X8 FILLER_114_1880 ();
 FILLCELL_X4 FILLER_114_1888 ();
 FILLCELL_X2 FILLER_114_1892 ();
 FILLCELL_X32 FILLER_114_1895 ();
 FILLCELL_X32 FILLER_114_1927 ();
 FILLCELL_X32 FILLER_114_1959 ();
 FILLCELL_X32 FILLER_114_1991 ();
 FILLCELL_X32 FILLER_114_2023 ();
 FILLCELL_X32 FILLER_114_2055 ();
 FILLCELL_X32 FILLER_114_2087 ();
 FILLCELL_X32 FILLER_114_2119 ();
 FILLCELL_X32 FILLER_114_2151 ();
 FILLCELL_X32 FILLER_114_2183 ();
 FILLCELL_X32 FILLER_114_2215 ();
 FILLCELL_X32 FILLER_114_2247 ();
 FILLCELL_X32 FILLER_114_2279 ();
 FILLCELL_X32 FILLER_114_2311 ();
 FILLCELL_X32 FILLER_114_2343 ();
 FILLCELL_X32 FILLER_114_2375 ();
 FILLCELL_X32 FILLER_114_2407 ();
 FILLCELL_X32 FILLER_114_2439 ();
 FILLCELL_X32 FILLER_114_2471 ();
 FILLCELL_X32 FILLER_114_2503 ();
 FILLCELL_X32 FILLER_114_2535 ();
 FILLCELL_X32 FILLER_114_2567 ();
 FILLCELL_X2 FILLER_114_2599 ();
 FILLCELL_X1 FILLER_114_2601 ();
 FILLCELL_X32 FILLER_115_1 ();
 FILLCELL_X32 FILLER_115_33 ();
 FILLCELL_X32 FILLER_115_65 ();
 FILLCELL_X32 FILLER_115_97 ();
 FILLCELL_X32 FILLER_115_129 ();
 FILLCELL_X32 FILLER_115_161 ();
 FILLCELL_X32 FILLER_115_193 ();
 FILLCELL_X32 FILLER_115_225 ();
 FILLCELL_X32 FILLER_115_257 ();
 FILLCELL_X32 FILLER_115_289 ();
 FILLCELL_X32 FILLER_115_321 ();
 FILLCELL_X32 FILLER_115_353 ();
 FILLCELL_X32 FILLER_115_385 ();
 FILLCELL_X32 FILLER_115_417 ();
 FILLCELL_X32 FILLER_115_449 ();
 FILLCELL_X32 FILLER_115_481 ();
 FILLCELL_X32 FILLER_115_513 ();
 FILLCELL_X32 FILLER_115_545 ();
 FILLCELL_X32 FILLER_115_577 ();
 FILLCELL_X32 FILLER_115_609 ();
 FILLCELL_X32 FILLER_115_641 ();
 FILLCELL_X32 FILLER_115_673 ();
 FILLCELL_X32 FILLER_115_705 ();
 FILLCELL_X32 FILLER_115_737 ();
 FILLCELL_X32 FILLER_115_769 ();
 FILLCELL_X32 FILLER_115_801 ();
 FILLCELL_X32 FILLER_115_833 ();
 FILLCELL_X32 FILLER_115_865 ();
 FILLCELL_X32 FILLER_115_897 ();
 FILLCELL_X32 FILLER_115_929 ();
 FILLCELL_X32 FILLER_115_961 ();
 FILLCELL_X32 FILLER_115_993 ();
 FILLCELL_X32 FILLER_115_1025 ();
 FILLCELL_X32 FILLER_115_1057 ();
 FILLCELL_X32 FILLER_115_1089 ();
 FILLCELL_X32 FILLER_115_1121 ();
 FILLCELL_X32 FILLER_115_1153 ();
 FILLCELL_X32 FILLER_115_1185 ();
 FILLCELL_X32 FILLER_115_1217 ();
 FILLCELL_X8 FILLER_115_1249 ();
 FILLCELL_X4 FILLER_115_1257 ();
 FILLCELL_X2 FILLER_115_1261 ();
 FILLCELL_X32 FILLER_115_1264 ();
 FILLCELL_X32 FILLER_115_1296 ();
 FILLCELL_X32 FILLER_115_1328 ();
 FILLCELL_X32 FILLER_115_1360 ();
 FILLCELL_X32 FILLER_115_1392 ();
 FILLCELL_X32 FILLER_115_1424 ();
 FILLCELL_X32 FILLER_115_1456 ();
 FILLCELL_X32 FILLER_115_1488 ();
 FILLCELL_X32 FILLER_115_1520 ();
 FILLCELL_X32 FILLER_115_1552 ();
 FILLCELL_X32 FILLER_115_1584 ();
 FILLCELL_X32 FILLER_115_1616 ();
 FILLCELL_X32 FILLER_115_1648 ();
 FILLCELL_X32 FILLER_115_1680 ();
 FILLCELL_X32 FILLER_115_1712 ();
 FILLCELL_X32 FILLER_115_1744 ();
 FILLCELL_X32 FILLER_115_1776 ();
 FILLCELL_X32 FILLER_115_1808 ();
 FILLCELL_X32 FILLER_115_1840 ();
 FILLCELL_X32 FILLER_115_1872 ();
 FILLCELL_X32 FILLER_115_1904 ();
 FILLCELL_X32 FILLER_115_1936 ();
 FILLCELL_X32 FILLER_115_1968 ();
 FILLCELL_X32 FILLER_115_2000 ();
 FILLCELL_X32 FILLER_115_2032 ();
 FILLCELL_X32 FILLER_115_2064 ();
 FILLCELL_X32 FILLER_115_2096 ();
 FILLCELL_X32 FILLER_115_2128 ();
 FILLCELL_X32 FILLER_115_2160 ();
 FILLCELL_X32 FILLER_115_2192 ();
 FILLCELL_X32 FILLER_115_2224 ();
 FILLCELL_X32 FILLER_115_2256 ();
 FILLCELL_X32 FILLER_115_2288 ();
 FILLCELL_X32 FILLER_115_2320 ();
 FILLCELL_X32 FILLER_115_2352 ();
 FILLCELL_X32 FILLER_115_2384 ();
 FILLCELL_X32 FILLER_115_2416 ();
 FILLCELL_X32 FILLER_115_2448 ();
 FILLCELL_X32 FILLER_115_2480 ();
 FILLCELL_X8 FILLER_115_2512 ();
 FILLCELL_X4 FILLER_115_2520 ();
 FILLCELL_X2 FILLER_115_2524 ();
 FILLCELL_X32 FILLER_115_2527 ();
 FILLCELL_X32 FILLER_115_2559 ();
 FILLCELL_X8 FILLER_115_2591 ();
 FILLCELL_X2 FILLER_115_2599 ();
 FILLCELL_X1 FILLER_115_2601 ();
 FILLCELL_X32 FILLER_116_1 ();
 FILLCELL_X32 FILLER_116_33 ();
 FILLCELL_X32 FILLER_116_65 ();
 FILLCELL_X32 FILLER_116_97 ();
 FILLCELL_X32 FILLER_116_129 ();
 FILLCELL_X32 FILLER_116_161 ();
 FILLCELL_X32 FILLER_116_193 ();
 FILLCELL_X32 FILLER_116_225 ();
 FILLCELL_X32 FILLER_116_257 ();
 FILLCELL_X32 FILLER_116_289 ();
 FILLCELL_X32 FILLER_116_321 ();
 FILLCELL_X32 FILLER_116_353 ();
 FILLCELL_X32 FILLER_116_385 ();
 FILLCELL_X32 FILLER_116_417 ();
 FILLCELL_X32 FILLER_116_449 ();
 FILLCELL_X32 FILLER_116_481 ();
 FILLCELL_X32 FILLER_116_513 ();
 FILLCELL_X32 FILLER_116_545 ();
 FILLCELL_X32 FILLER_116_577 ();
 FILLCELL_X16 FILLER_116_609 ();
 FILLCELL_X4 FILLER_116_625 ();
 FILLCELL_X2 FILLER_116_629 ();
 FILLCELL_X32 FILLER_116_632 ();
 FILLCELL_X32 FILLER_116_664 ();
 FILLCELL_X32 FILLER_116_696 ();
 FILLCELL_X32 FILLER_116_728 ();
 FILLCELL_X32 FILLER_116_760 ();
 FILLCELL_X32 FILLER_116_792 ();
 FILLCELL_X32 FILLER_116_824 ();
 FILLCELL_X32 FILLER_116_856 ();
 FILLCELL_X32 FILLER_116_888 ();
 FILLCELL_X32 FILLER_116_920 ();
 FILLCELL_X32 FILLER_116_952 ();
 FILLCELL_X32 FILLER_116_984 ();
 FILLCELL_X32 FILLER_116_1016 ();
 FILLCELL_X32 FILLER_116_1048 ();
 FILLCELL_X32 FILLER_116_1080 ();
 FILLCELL_X32 FILLER_116_1112 ();
 FILLCELL_X32 FILLER_116_1144 ();
 FILLCELL_X32 FILLER_116_1176 ();
 FILLCELL_X32 FILLER_116_1208 ();
 FILLCELL_X32 FILLER_116_1240 ();
 FILLCELL_X32 FILLER_116_1272 ();
 FILLCELL_X32 FILLER_116_1304 ();
 FILLCELL_X32 FILLER_116_1336 ();
 FILLCELL_X32 FILLER_116_1368 ();
 FILLCELL_X32 FILLER_116_1400 ();
 FILLCELL_X32 FILLER_116_1432 ();
 FILLCELL_X32 FILLER_116_1464 ();
 FILLCELL_X32 FILLER_116_1496 ();
 FILLCELL_X32 FILLER_116_1528 ();
 FILLCELL_X32 FILLER_116_1560 ();
 FILLCELL_X32 FILLER_116_1592 ();
 FILLCELL_X32 FILLER_116_1624 ();
 FILLCELL_X32 FILLER_116_1656 ();
 FILLCELL_X32 FILLER_116_1688 ();
 FILLCELL_X32 FILLER_116_1720 ();
 FILLCELL_X32 FILLER_116_1752 ();
 FILLCELL_X32 FILLER_116_1784 ();
 FILLCELL_X32 FILLER_116_1816 ();
 FILLCELL_X32 FILLER_116_1848 ();
 FILLCELL_X8 FILLER_116_1880 ();
 FILLCELL_X4 FILLER_116_1888 ();
 FILLCELL_X2 FILLER_116_1892 ();
 FILLCELL_X32 FILLER_116_1895 ();
 FILLCELL_X32 FILLER_116_1927 ();
 FILLCELL_X32 FILLER_116_1959 ();
 FILLCELL_X32 FILLER_116_1991 ();
 FILLCELL_X32 FILLER_116_2023 ();
 FILLCELL_X32 FILLER_116_2055 ();
 FILLCELL_X32 FILLER_116_2087 ();
 FILLCELL_X32 FILLER_116_2119 ();
 FILLCELL_X32 FILLER_116_2151 ();
 FILLCELL_X32 FILLER_116_2183 ();
 FILLCELL_X32 FILLER_116_2215 ();
 FILLCELL_X32 FILLER_116_2247 ();
 FILLCELL_X32 FILLER_116_2279 ();
 FILLCELL_X32 FILLER_116_2311 ();
 FILLCELL_X32 FILLER_116_2343 ();
 FILLCELL_X32 FILLER_116_2375 ();
 FILLCELL_X32 FILLER_116_2407 ();
 FILLCELL_X32 FILLER_116_2439 ();
 FILLCELL_X32 FILLER_116_2471 ();
 FILLCELL_X32 FILLER_116_2503 ();
 FILLCELL_X32 FILLER_116_2535 ();
 FILLCELL_X32 FILLER_116_2567 ();
 FILLCELL_X2 FILLER_116_2599 ();
 FILLCELL_X1 FILLER_116_2601 ();
 FILLCELL_X32 FILLER_117_1 ();
 FILLCELL_X32 FILLER_117_33 ();
 FILLCELL_X32 FILLER_117_65 ();
 FILLCELL_X32 FILLER_117_97 ();
 FILLCELL_X32 FILLER_117_129 ();
 FILLCELL_X32 FILLER_117_161 ();
 FILLCELL_X32 FILLER_117_193 ();
 FILLCELL_X32 FILLER_117_225 ();
 FILLCELL_X32 FILLER_117_257 ();
 FILLCELL_X32 FILLER_117_289 ();
 FILLCELL_X32 FILLER_117_321 ();
 FILLCELL_X32 FILLER_117_353 ();
 FILLCELL_X32 FILLER_117_385 ();
 FILLCELL_X32 FILLER_117_417 ();
 FILLCELL_X32 FILLER_117_449 ();
 FILLCELL_X32 FILLER_117_481 ();
 FILLCELL_X32 FILLER_117_513 ();
 FILLCELL_X32 FILLER_117_545 ();
 FILLCELL_X32 FILLER_117_577 ();
 FILLCELL_X32 FILLER_117_609 ();
 FILLCELL_X32 FILLER_117_641 ();
 FILLCELL_X32 FILLER_117_673 ();
 FILLCELL_X32 FILLER_117_705 ();
 FILLCELL_X32 FILLER_117_737 ();
 FILLCELL_X32 FILLER_117_769 ();
 FILLCELL_X32 FILLER_117_801 ();
 FILLCELL_X32 FILLER_117_833 ();
 FILLCELL_X32 FILLER_117_865 ();
 FILLCELL_X32 FILLER_117_897 ();
 FILLCELL_X32 FILLER_117_929 ();
 FILLCELL_X32 FILLER_117_961 ();
 FILLCELL_X32 FILLER_117_993 ();
 FILLCELL_X32 FILLER_117_1025 ();
 FILLCELL_X32 FILLER_117_1057 ();
 FILLCELL_X32 FILLER_117_1089 ();
 FILLCELL_X32 FILLER_117_1121 ();
 FILLCELL_X32 FILLER_117_1153 ();
 FILLCELL_X32 FILLER_117_1185 ();
 FILLCELL_X32 FILLER_117_1217 ();
 FILLCELL_X8 FILLER_117_1249 ();
 FILLCELL_X4 FILLER_117_1257 ();
 FILLCELL_X2 FILLER_117_1261 ();
 FILLCELL_X32 FILLER_117_1264 ();
 FILLCELL_X32 FILLER_117_1296 ();
 FILLCELL_X32 FILLER_117_1328 ();
 FILLCELL_X32 FILLER_117_1360 ();
 FILLCELL_X32 FILLER_117_1392 ();
 FILLCELL_X32 FILLER_117_1424 ();
 FILLCELL_X32 FILLER_117_1456 ();
 FILLCELL_X32 FILLER_117_1488 ();
 FILLCELL_X32 FILLER_117_1520 ();
 FILLCELL_X32 FILLER_117_1552 ();
 FILLCELL_X32 FILLER_117_1584 ();
 FILLCELL_X32 FILLER_117_1616 ();
 FILLCELL_X32 FILLER_117_1648 ();
 FILLCELL_X32 FILLER_117_1680 ();
 FILLCELL_X32 FILLER_117_1712 ();
 FILLCELL_X32 FILLER_117_1744 ();
 FILLCELL_X32 FILLER_117_1776 ();
 FILLCELL_X32 FILLER_117_1808 ();
 FILLCELL_X32 FILLER_117_1840 ();
 FILLCELL_X32 FILLER_117_1872 ();
 FILLCELL_X32 FILLER_117_1904 ();
 FILLCELL_X32 FILLER_117_1936 ();
 FILLCELL_X32 FILLER_117_1968 ();
 FILLCELL_X32 FILLER_117_2000 ();
 FILLCELL_X32 FILLER_117_2032 ();
 FILLCELL_X32 FILLER_117_2064 ();
 FILLCELL_X32 FILLER_117_2096 ();
 FILLCELL_X32 FILLER_117_2128 ();
 FILLCELL_X32 FILLER_117_2160 ();
 FILLCELL_X32 FILLER_117_2192 ();
 FILLCELL_X32 FILLER_117_2224 ();
 FILLCELL_X32 FILLER_117_2256 ();
 FILLCELL_X32 FILLER_117_2288 ();
 FILLCELL_X32 FILLER_117_2320 ();
 FILLCELL_X32 FILLER_117_2352 ();
 FILLCELL_X32 FILLER_117_2384 ();
 FILLCELL_X32 FILLER_117_2416 ();
 FILLCELL_X32 FILLER_117_2448 ();
 FILLCELL_X32 FILLER_117_2480 ();
 FILLCELL_X8 FILLER_117_2512 ();
 FILLCELL_X4 FILLER_117_2520 ();
 FILLCELL_X2 FILLER_117_2524 ();
 FILLCELL_X32 FILLER_117_2527 ();
 FILLCELL_X32 FILLER_117_2559 ();
 FILLCELL_X8 FILLER_117_2591 ();
 FILLCELL_X2 FILLER_117_2599 ();
 FILLCELL_X1 FILLER_117_2601 ();
 FILLCELL_X32 FILLER_118_1 ();
 FILLCELL_X32 FILLER_118_33 ();
 FILLCELL_X32 FILLER_118_65 ();
 FILLCELL_X32 FILLER_118_97 ();
 FILLCELL_X32 FILLER_118_129 ();
 FILLCELL_X32 FILLER_118_161 ();
 FILLCELL_X32 FILLER_118_193 ();
 FILLCELL_X32 FILLER_118_225 ();
 FILLCELL_X32 FILLER_118_257 ();
 FILLCELL_X32 FILLER_118_289 ();
 FILLCELL_X32 FILLER_118_321 ();
 FILLCELL_X32 FILLER_118_353 ();
 FILLCELL_X32 FILLER_118_385 ();
 FILLCELL_X32 FILLER_118_417 ();
 FILLCELL_X32 FILLER_118_449 ();
 FILLCELL_X32 FILLER_118_481 ();
 FILLCELL_X32 FILLER_118_513 ();
 FILLCELL_X32 FILLER_118_545 ();
 FILLCELL_X32 FILLER_118_577 ();
 FILLCELL_X16 FILLER_118_609 ();
 FILLCELL_X4 FILLER_118_625 ();
 FILLCELL_X2 FILLER_118_629 ();
 FILLCELL_X32 FILLER_118_632 ();
 FILLCELL_X32 FILLER_118_664 ();
 FILLCELL_X32 FILLER_118_696 ();
 FILLCELL_X32 FILLER_118_728 ();
 FILLCELL_X32 FILLER_118_760 ();
 FILLCELL_X32 FILLER_118_792 ();
 FILLCELL_X32 FILLER_118_824 ();
 FILLCELL_X32 FILLER_118_856 ();
 FILLCELL_X32 FILLER_118_888 ();
 FILLCELL_X32 FILLER_118_920 ();
 FILLCELL_X32 FILLER_118_952 ();
 FILLCELL_X32 FILLER_118_984 ();
 FILLCELL_X32 FILLER_118_1016 ();
 FILLCELL_X32 FILLER_118_1048 ();
 FILLCELL_X32 FILLER_118_1080 ();
 FILLCELL_X32 FILLER_118_1112 ();
 FILLCELL_X32 FILLER_118_1144 ();
 FILLCELL_X32 FILLER_118_1176 ();
 FILLCELL_X32 FILLER_118_1208 ();
 FILLCELL_X32 FILLER_118_1240 ();
 FILLCELL_X32 FILLER_118_1272 ();
 FILLCELL_X32 FILLER_118_1304 ();
 FILLCELL_X32 FILLER_118_1336 ();
 FILLCELL_X32 FILLER_118_1368 ();
 FILLCELL_X32 FILLER_118_1400 ();
 FILLCELL_X32 FILLER_118_1432 ();
 FILLCELL_X32 FILLER_118_1464 ();
 FILLCELL_X32 FILLER_118_1496 ();
 FILLCELL_X32 FILLER_118_1528 ();
 FILLCELL_X32 FILLER_118_1560 ();
 FILLCELL_X32 FILLER_118_1592 ();
 FILLCELL_X32 FILLER_118_1624 ();
 FILLCELL_X32 FILLER_118_1656 ();
 FILLCELL_X32 FILLER_118_1688 ();
 FILLCELL_X32 FILLER_118_1720 ();
 FILLCELL_X32 FILLER_118_1752 ();
 FILLCELL_X32 FILLER_118_1784 ();
 FILLCELL_X32 FILLER_118_1816 ();
 FILLCELL_X32 FILLER_118_1848 ();
 FILLCELL_X8 FILLER_118_1880 ();
 FILLCELL_X4 FILLER_118_1888 ();
 FILLCELL_X2 FILLER_118_1892 ();
 FILLCELL_X32 FILLER_118_1895 ();
 FILLCELL_X32 FILLER_118_1927 ();
 FILLCELL_X32 FILLER_118_1959 ();
 FILLCELL_X32 FILLER_118_1991 ();
 FILLCELL_X32 FILLER_118_2023 ();
 FILLCELL_X32 FILLER_118_2055 ();
 FILLCELL_X32 FILLER_118_2087 ();
 FILLCELL_X32 FILLER_118_2119 ();
 FILLCELL_X32 FILLER_118_2151 ();
 FILLCELL_X32 FILLER_118_2183 ();
 FILLCELL_X32 FILLER_118_2215 ();
 FILLCELL_X32 FILLER_118_2247 ();
 FILLCELL_X32 FILLER_118_2279 ();
 FILLCELL_X32 FILLER_118_2311 ();
 FILLCELL_X32 FILLER_118_2343 ();
 FILLCELL_X32 FILLER_118_2375 ();
 FILLCELL_X32 FILLER_118_2407 ();
 FILLCELL_X32 FILLER_118_2439 ();
 FILLCELL_X32 FILLER_118_2471 ();
 FILLCELL_X32 FILLER_118_2503 ();
 FILLCELL_X32 FILLER_118_2535 ();
 FILLCELL_X32 FILLER_118_2567 ();
 FILLCELL_X2 FILLER_118_2599 ();
 FILLCELL_X1 FILLER_118_2601 ();
 FILLCELL_X32 FILLER_119_1 ();
 FILLCELL_X32 FILLER_119_33 ();
 FILLCELL_X32 FILLER_119_65 ();
 FILLCELL_X32 FILLER_119_97 ();
 FILLCELL_X32 FILLER_119_129 ();
 FILLCELL_X32 FILLER_119_161 ();
 FILLCELL_X32 FILLER_119_193 ();
 FILLCELL_X32 FILLER_119_225 ();
 FILLCELL_X32 FILLER_119_257 ();
 FILLCELL_X32 FILLER_119_289 ();
 FILLCELL_X32 FILLER_119_321 ();
 FILLCELL_X32 FILLER_119_353 ();
 FILLCELL_X32 FILLER_119_385 ();
 FILLCELL_X32 FILLER_119_417 ();
 FILLCELL_X32 FILLER_119_449 ();
 FILLCELL_X32 FILLER_119_481 ();
 FILLCELL_X32 FILLER_119_513 ();
 FILLCELL_X32 FILLER_119_545 ();
 FILLCELL_X32 FILLER_119_577 ();
 FILLCELL_X32 FILLER_119_609 ();
 FILLCELL_X32 FILLER_119_641 ();
 FILLCELL_X32 FILLER_119_673 ();
 FILLCELL_X32 FILLER_119_705 ();
 FILLCELL_X32 FILLER_119_737 ();
 FILLCELL_X32 FILLER_119_769 ();
 FILLCELL_X32 FILLER_119_801 ();
 FILLCELL_X32 FILLER_119_833 ();
 FILLCELL_X32 FILLER_119_865 ();
 FILLCELL_X32 FILLER_119_897 ();
 FILLCELL_X32 FILLER_119_929 ();
 FILLCELL_X32 FILLER_119_961 ();
 FILLCELL_X32 FILLER_119_993 ();
 FILLCELL_X32 FILLER_119_1025 ();
 FILLCELL_X32 FILLER_119_1057 ();
 FILLCELL_X32 FILLER_119_1089 ();
 FILLCELL_X32 FILLER_119_1121 ();
 FILLCELL_X32 FILLER_119_1153 ();
 FILLCELL_X32 FILLER_119_1185 ();
 FILLCELL_X32 FILLER_119_1217 ();
 FILLCELL_X8 FILLER_119_1249 ();
 FILLCELL_X4 FILLER_119_1257 ();
 FILLCELL_X2 FILLER_119_1261 ();
 FILLCELL_X32 FILLER_119_1264 ();
 FILLCELL_X32 FILLER_119_1296 ();
 FILLCELL_X32 FILLER_119_1328 ();
 FILLCELL_X32 FILLER_119_1360 ();
 FILLCELL_X32 FILLER_119_1392 ();
 FILLCELL_X32 FILLER_119_1424 ();
 FILLCELL_X32 FILLER_119_1456 ();
 FILLCELL_X32 FILLER_119_1488 ();
 FILLCELL_X32 FILLER_119_1520 ();
 FILLCELL_X32 FILLER_119_1552 ();
 FILLCELL_X32 FILLER_119_1584 ();
 FILLCELL_X32 FILLER_119_1616 ();
 FILLCELL_X32 FILLER_119_1648 ();
 FILLCELL_X32 FILLER_119_1680 ();
 FILLCELL_X32 FILLER_119_1712 ();
 FILLCELL_X32 FILLER_119_1744 ();
 FILLCELL_X32 FILLER_119_1776 ();
 FILLCELL_X32 FILLER_119_1808 ();
 FILLCELL_X32 FILLER_119_1840 ();
 FILLCELL_X32 FILLER_119_1872 ();
 FILLCELL_X32 FILLER_119_1904 ();
 FILLCELL_X32 FILLER_119_1936 ();
 FILLCELL_X32 FILLER_119_1968 ();
 FILLCELL_X32 FILLER_119_2000 ();
 FILLCELL_X32 FILLER_119_2032 ();
 FILLCELL_X32 FILLER_119_2064 ();
 FILLCELL_X32 FILLER_119_2096 ();
 FILLCELL_X32 FILLER_119_2128 ();
 FILLCELL_X32 FILLER_119_2160 ();
 FILLCELL_X32 FILLER_119_2192 ();
 FILLCELL_X32 FILLER_119_2224 ();
 FILLCELL_X32 FILLER_119_2256 ();
 FILLCELL_X32 FILLER_119_2288 ();
 FILLCELL_X32 FILLER_119_2320 ();
 FILLCELL_X32 FILLER_119_2352 ();
 FILLCELL_X32 FILLER_119_2384 ();
 FILLCELL_X32 FILLER_119_2416 ();
 FILLCELL_X32 FILLER_119_2448 ();
 FILLCELL_X32 FILLER_119_2480 ();
 FILLCELL_X8 FILLER_119_2512 ();
 FILLCELL_X4 FILLER_119_2520 ();
 FILLCELL_X2 FILLER_119_2524 ();
 FILLCELL_X32 FILLER_119_2527 ();
 FILLCELL_X32 FILLER_119_2559 ();
 FILLCELL_X8 FILLER_119_2591 ();
 FILLCELL_X2 FILLER_119_2599 ();
 FILLCELL_X1 FILLER_119_2601 ();
 FILLCELL_X32 FILLER_120_1 ();
 FILLCELL_X32 FILLER_120_33 ();
 FILLCELL_X32 FILLER_120_65 ();
 FILLCELL_X32 FILLER_120_97 ();
 FILLCELL_X32 FILLER_120_129 ();
 FILLCELL_X32 FILLER_120_161 ();
 FILLCELL_X32 FILLER_120_193 ();
 FILLCELL_X32 FILLER_120_225 ();
 FILLCELL_X32 FILLER_120_257 ();
 FILLCELL_X32 FILLER_120_289 ();
 FILLCELL_X32 FILLER_120_321 ();
 FILLCELL_X32 FILLER_120_353 ();
 FILLCELL_X32 FILLER_120_385 ();
 FILLCELL_X32 FILLER_120_417 ();
 FILLCELL_X32 FILLER_120_449 ();
 FILLCELL_X32 FILLER_120_481 ();
 FILLCELL_X32 FILLER_120_513 ();
 FILLCELL_X32 FILLER_120_545 ();
 FILLCELL_X32 FILLER_120_577 ();
 FILLCELL_X16 FILLER_120_609 ();
 FILLCELL_X4 FILLER_120_625 ();
 FILLCELL_X2 FILLER_120_629 ();
 FILLCELL_X32 FILLER_120_632 ();
 FILLCELL_X32 FILLER_120_664 ();
 FILLCELL_X32 FILLER_120_696 ();
 FILLCELL_X32 FILLER_120_728 ();
 FILLCELL_X32 FILLER_120_760 ();
 FILLCELL_X32 FILLER_120_792 ();
 FILLCELL_X32 FILLER_120_824 ();
 FILLCELL_X32 FILLER_120_856 ();
 FILLCELL_X32 FILLER_120_888 ();
 FILLCELL_X32 FILLER_120_920 ();
 FILLCELL_X32 FILLER_120_952 ();
 FILLCELL_X32 FILLER_120_984 ();
 FILLCELL_X32 FILLER_120_1016 ();
 FILLCELL_X32 FILLER_120_1048 ();
 FILLCELL_X32 FILLER_120_1080 ();
 FILLCELL_X32 FILLER_120_1112 ();
 FILLCELL_X32 FILLER_120_1144 ();
 FILLCELL_X32 FILLER_120_1176 ();
 FILLCELL_X32 FILLER_120_1208 ();
 FILLCELL_X32 FILLER_120_1240 ();
 FILLCELL_X32 FILLER_120_1272 ();
 FILLCELL_X32 FILLER_120_1304 ();
 FILLCELL_X32 FILLER_120_1336 ();
 FILLCELL_X32 FILLER_120_1368 ();
 FILLCELL_X32 FILLER_120_1400 ();
 FILLCELL_X32 FILLER_120_1432 ();
 FILLCELL_X32 FILLER_120_1464 ();
 FILLCELL_X32 FILLER_120_1496 ();
 FILLCELL_X32 FILLER_120_1528 ();
 FILLCELL_X32 FILLER_120_1560 ();
 FILLCELL_X32 FILLER_120_1592 ();
 FILLCELL_X32 FILLER_120_1624 ();
 FILLCELL_X32 FILLER_120_1656 ();
 FILLCELL_X32 FILLER_120_1688 ();
 FILLCELL_X32 FILLER_120_1720 ();
 FILLCELL_X32 FILLER_120_1752 ();
 FILLCELL_X32 FILLER_120_1784 ();
 FILLCELL_X32 FILLER_120_1816 ();
 FILLCELL_X32 FILLER_120_1848 ();
 FILLCELL_X8 FILLER_120_1880 ();
 FILLCELL_X4 FILLER_120_1888 ();
 FILLCELL_X2 FILLER_120_1892 ();
 FILLCELL_X32 FILLER_120_1895 ();
 FILLCELL_X32 FILLER_120_1927 ();
 FILLCELL_X32 FILLER_120_1959 ();
 FILLCELL_X32 FILLER_120_1991 ();
 FILLCELL_X32 FILLER_120_2023 ();
 FILLCELL_X32 FILLER_120_2055 ();
 FILLCELL_X32 FILLER_120_2087 ();
 FILLCELL_X32 FILLER_120_2119 ();
 FILLCELL_X32 FILLER_120_2151 ();
 FILLCELL_X32 FILLER_120_2183 ();
 FILLCELL_X32 FILLER_120_2215 ();
 FILLCELL_X32 FILLER_120_2247 ();
 FILLCELL_X32 FILLER_120_2279 ();
 FILLCELL_X32 FILLER_120_2311 ();
 FILLCELL_X32 FILLER_120_2343 ();
 FILLCELL_X32 FILLER_120_2375 ();
 FILLCELL_X32 FILLER_120_2407 ();
 FILLCELL_X32 FILLER_120_2439 ();
 FILLCELL_X32 FILLER_120_2471 ();
 FILLCELL_X32 FILLER_120_2503 ();
 FILLCELL_X32 FILLER_120_2535 ();
 FILLCELL_X32 FILLER_120_2567 ();
 FILLCELL_X2 FILLER_120_2599 ();
 FILLCELL_X1 FILLER_120_2601 ();
 FILLCELL_X32 FILLER_121_1 ();
 FILLCELL_X32 FILLER_121_33 ();
 FILLCELL_X32 FILLER_121_65 ();
 FILLCELL_X32 FILLER_121_97 ();
 FILLCELL_X32 FILLER_121_129 ();
 FILLCELL_X32 FILLER_121_161 ();
 FILLCELL_X32 FILLER_121_193 ();
 FILLCELL_X32 FILLER_121_225 ();
 FILLCELL_X32 FILLER_121_257 ();
 FILLCELL_X32 FILLER_121_289 ();
 FILLCELL_X32 FILLER_121_321 ();
 FILLCELL_X32 FILLER_121_353 ();
 FILLCELL_X32 FILLER_121_385 ();
 FILLCELL_X32 FILLER_121_417 ();
 FILLCELL_X32 FILLER_121_449 ();
 FILLCELL_X32 FILLER_121_481 ();
 FILLCELL_X32 FILLER_121_513 ();
 FILLCELL_X32 FILLER_121_545 ();
 FILLCELL_X32 FILLER_121_577 ();
 FILLCELL_X32 FILLER_121_609 ();
 FILLCELL_X32 FILLER_121_641 ();
 FILLCELL_X32 FILLER_121_673 ();
 FILLCELL_X32 FILLER_121_705 ();
 FILLCELL_X32 FILLER_121_737 ();
 FILLCELL_X32 FILLER_121_769 ();
 FILLCELL_X32 FILLER_121_801 ();
 FILLCELL_X32 FILLER_121_833 ();
 FILLCELL_X32 FILLER_121_865 ();
 FILLCELL_X32 FILLER_121_897 ();
 FILLCELL_X32 FILLER_121_929 ();
 FILLCELL_X32 FILLER_121_961 ();
 FILLCELL_X32 FILLER_121_993 ();
 FILLCELL_X32 FILLER_121_1025 ();
 FILLCELL_X32 FILLER_121_1057 ();
 FILLCELL_X32 FILLER_121_1089 ();
 FILLCELL_X32 FILLER_121_1121 ();
 FILLCELL_X32 FILLER_121_1153 ();
 FILLCELL_X32 FILLER_121_1185 ();
 FILLCELL_X32 FILLER_121_1217 ();
 FILLCELL_X8 FILLER_121_1249 ();
 FILLCELL_X4 FILLER_121_1257 ();
 FILLCELL_X2 FILLER_121_1261 ();
 FILLCELL_X32 FILLER_121_1264 ();
 FILLCELL_X32 FILLER_121_1296 ();
 FILLCELL_X32 FILLER_121_1328 ();
 FILLCELL_X32 FILLER_121_1360 ();
 FILLCELL_X32 FILLER_121_1392 ();
 FILLCELL_X32 FILLER_121_1424 ();
 FILLCELL_X32 FILLER_121_1456 ();
 FILLCELL_X32 FILLER_121_1488 ();
 FILLCELL_X32 FILLER_121_1520 ();
 FILLCELL_X32 FILLER_121_1552 ();
 FILLCELL_X32 FILLER_121_1584 ();
 FILLCELL_X32 FILLER_121_1616 ();
 FILLCELL_X32 FILLER_121_1648 ();
 FILLCELL_X32 FILLER_121_1680 ();
 FILLCELL_X32 FILLER_121_1712 ();
 FILLCELL_X32 FILLER_121_1744 ();
 FILLCELL_X32 FILLER_121_1776 ();
 FILLCELL_X32 FILLER_121_1808 ();
 FILLCELL_X32 FILLER_121_1840 ();
 FILLCELL_X32 FILLER_121_1872 ();
 FILLCELL_X32 FILLER_121_1904 ();
 FILLCELL_X32 FILLER_121_1936 ();
 FILLCELL_X32 FILLER_121_1968 ();
 FILLCELL_X32 FILLER_121_2000 ();
 FILLCELL_X32 FILLER_121_2032 ();
 FILLCELL_X32 FILLER_121_2064 ();
 FILLCELL_X32 FILLER_121_2096 ();
 FILLCELL_X32 FILLER_121_2128 ();
 FILLCELL_X32 FILLER_121_2160 ();
 FILLCELL_X32 FILLER_121_2192 ();
 FILLCELL_X32 FILLER_121_2224 ();
 FILLCELL_X32 FILLER_121_2256 ();
 FILLCELL_X32 FILLER_121_2288 ();
 FILLCELL_X32 FILLER_121_2320 ();
 FILLCELL_X32 FILLER_121_2352 ();
 FILLCELL_X32 FILLER_121_2384 ();
 FILLCELL_X32 FILLER_121_2416 ();
 FILLCELL_X32 FILLER_121_2448 ();
 FILLCELL_X32 FILLER_121_2480 ();
 FILLCELL_X8 FILLER_121_2512 ();
 FILLCELL_X4 FILLER_121_2520 ();
 FILLCELL_X2 FILLER_121_2524 ();
 FILLCELL_X32 FILLER_121_2527 ();
 FILLCELL_X32 FILLER_121_2559 ();
 FILLCELL_X8 FILLER_121_2591 ();
 FILLCELL_X2 FILLER_121_2599 ();
 FILLCELL_X1 FILLER_121_2601 ();
 FILLCELL_X32 FILLER_122_1 ();
 FILLCELL_X32 FILLER_122_33 ();
 FILLCELL_X32 FILLER_122_65 ();
 FILLCELL_X32 FILLER_122_97 ();
 FILLCELL_X32 FILLER_122_129 ();
 FILLCELL_X32 FILLER_122_161 ();
 FILLCELL_X32 FILLER_122_193 ();
 FILLCELL_X32 FILLER_122_225 ();
 FILLCELL_X32 FILLER_122_257 ();
 FILLCELL_X32 FILLER_122_289 ();
 FILLCELL_X32 FILLER_122_321 ();
 FILLCELL_X32 FILLER_122_353 ();
 FILLCELL_X32 FILLER_122_385 ();
 FILLCELL_X32 FILLER_122_417 ();
 FILLCELL_X32 FILLER_122_449 ();
 FILLCELL_X32 FILLER_122_481 ();
 FILLCELL_X32 FILLER_122_513 ();
 FILLCELL_X32 FILLER_122_545 ();
 FILLCELL_X32 FILLER_122_577 ();
 FILLCELL_X16 FILLER_122_609 ();
 FILLCELL_X4 FILLER_122_625 ();
 FILLCELL_X2 FILLER_122_629 ();
 FILLCELL_X32 FILLER_122_632 ();
 FILLCELL_X32 FILLER_122_664 ();
 FILLCELL_X32 FILLER_122_696 ();
 FILLCELL_X32 FILLER_122_728 ();
 FILLCELL_X32 FILLER_122_760 ();
 FILLCELL_X32 FILLER_122_792 ();
 FILLCELL_X32 FILLER_122_824 ();
 FILLCELL_X32 FILLER_122_856 ();
 FILLCELL_X32 FILLER_122_888 ();
 FILLCELL_X32 FILLER_122_920 ();
 FILLCELL_X32 FILLER_122_952 ();
 FILLCELL_X32 FILLER_122_984 ();
 FILLCELL_X32 FILLER_122_1016 ();
 FILLCELL_X32 FILLER_122_1048 ();
 FILLCELL_X32 FILLER_122_1080 ();
 FILLCELL_X32 FILLER_122_1112 ();
 FILLCELL_X32 FILLER_122_1144 ();
 FILLCELL_X32 FILLER_122_1176 ();
 FILLCELL_X32 FILLER_122_1208 ();
 FILLCELL_X32 FILLER_122_1240 ();
 FILLCELL_X32 FILLER_122_1272 ();
 FILLCELL_X32 FILLER_122_1304 ();
 FILLCELL_X32 FILLER_122_1336 ();
 FILLCELL_X32 FILLER_122_1368 ();
 FILLCELL_X32 FILLER_122_1400 ();
 FILLCELL_X32 FILLER_122_1432 ();
 FILLCELL_X32 FILLER_122_1464 ();
 FILLCELL_X32 FILLER_122_1496 ();
 FILLCELL_X32 FILLER_122_1528 ();
 FILLCELL_X32 FILLER_122_1560 ();
 FILLCELL_X32 FILLER_122_1592 ();
 FILLCELL_X32 FILLER_122_1624 ();
 FILLCELL_X32 FILLER_122_1656 ();
 FILLCELL_X32 FILLER_122_1688 ();
 FILLCELL_X32 FILLER_122_1720 ();
 FILLCELL_X32 FILLER_122_1752 ();
 FILLCELL_X32 FILLER_122_1784 ();
 FILLCELL_X32 FILLER_122_1816 ();
 FILLCELL_X32 FILLER_122_1848 ();
 FILLCELL_X8 FILLER_122_1880 ();
 FILLCELL_X4 FILLER_122_1888 ();
 FILLCELL_X2 FILLER_122_1892 ();
 FILLCELL_X32 FILLER_122_1895 ();
 FILLCELL_X32 FILLER_122_1927 ();
 FILLCELL_X32 FILLER_122_1959 ();
 FILLCELL_X32 FILLER_122_1991 ();
 FILLCELL_X32 FILLER_122_2023 ();
 FILLCELL_X32 FILLER_122_2055 ();
 FILLCELL_X32 FILLER_122_2087 ();
 FILLCELL_X32 FILLER_122_2119 ();
 FILLCELL_X32 FILLER_122_2151 ();
 FILLCELL_X32 FILLER_122_2183 ();
 FILLCELL_X32 FILLER_122_2215 ();
 FILLCELL_X32 FILLER_122_2247 ();
 FILLCELL_X32 FILLER_122_2279 ();
 FILLCELL_X32 FILLER_122_2311 ();
 FILLCELL_X32 FILLER_122_2343 ();
 FILLCELL_X32 FILLER_122_2375 ();
 FILLCELL_X32 FILLER_122_2407 ();
 FILLCELL_X32 FILLER_122_2439 ();
 FILLCELL_X32 FILLER_122_2471 ();
 FILLCELL_X32 FILLER_122_2503 ();
 FILLCELL_X32 FILLER_122_2535 ();
 FILLCELL_X32 FILLER_122_2567 ();
 FILLCELL_X2 FILLER_122_2599 ();
 FILLCELL_X1 FILLER_122_2601 ();
 FILLCELL_X32 FILLER_123_1 ();
 FILLCELL_X32 FILLER_123_33 ();
 FILLCELL_X32 FILLER_123_65 ();
 FILLCELL_X32 FILLER_123_97 ();
 FILLCELL_X32 FILLER_123_129 ();
 FILLCELL_X32 FILLER_123_161 ();
 FILLCELL_X32 FILLER_123_193 ();
 FILLCELL_X32 FILLER_123_225 ();
 FILLCELL_X32 FILLER_123_257 ();
 FILLCELL_X32 FILLER_123_289 ();
 FILLCELL_X32 FILLER_123_321 ();
 FILLCELL_X32 FILLER_123_353 ();
 FILLCELL_X32 FILLER_123_385 ();
 FILLCELL_X32 FILLER_123_417 ();
 FILLCELL_X32 FILLER_123_449 ();
 FILLCELL_X32 FILLER_123_481 ();
 FILLCELL_X32 FILLER_123_513 ();
 FILLCELL_X32 FILLER_123_545 ();
 FILLCELL_X32 FILLER_123_577 ();
 FILLCELL_X32 FILLER_123_609 ();
 FILLCELL_X32 FILLER_123_641 ();
 FILLCELL_X32 FILLER_123_673 ();
 FILLCELL_X32 FILLER_123_705 ();
 FILLCELL_X32 FILLER_123_737 ();
 FILLCELL_X32 FILLER_123_769 ();
 FILLCELL_X32 FILLER_123_801 ();
 FILLCELL_X32 FILLER_123_833 ();
 FILLCELL_X32 FILLER_123_865 ();
 FILLCELL_X32 FILLER_123_897 ();
 FILLCELL_X32 FILLER_123_929 ();
 FILLCELL_X32 FILLER_123_961 ();
 FILLCELL_X32 FILLER_123_993 ();
 FILLCELL_X32 FILLER_123_1025 ();
 FILLCELL_X32 FILLER_123_1057 ();
 FILLCELL_X32 FILLER_123_1089 ();
 FILLCELL_X32 FILLER_123_1121 ();
 FILLCELL_X32 FILLER_123_1153 ();
 FILLCELL_X32 FILLER_123_1185 ();
 FILLCELL_X32 FILLER_123_1217 ();
 FILLCELL_X8 FILLER_123_1249 ();
 FILLCELL_X4 FILLER_123_1257 ();
 FILLCELL_X2 FILLER_123_1261 ();
 FILLCELL_X32 FILLER_123_1264 ();
 FILLCELL_X32 FILLER_123_1296 ();
 FILLCELL_X32 FILLER_123_1328 ();
 FILLCELL_X32 FILLER_123_1360 ();
 FILLCELL_X32 FILLER_123_1392 ();
 FILLCELL_X32 FILLER_123_1424 ();
 FILLCELL_X32 FILLER_123_1456 ();
 FILLCELL_X32 FILLER_123_1488 ();
 FILLCELL_X32 FILLER_123_1520 ();
 FILLCELL_X32 FILLER_123_1552 ();
 FILLCELL_X32 FILLER_123_1584 ();
 FILLCELL_X32 FILLER_123_1616 ();
 FILLCELL_X32 FILLER_123_1648 ();
 FILLCELL_X32 FILLER_123_1680 ();
 FILLCELL_X32 FILLER_123_1712 ();
 FILLCELL_X32 FILLER_123_1744 ();
 FILLCELL_X32 FILLER_123_1776 ();
 FILLCELL_X32 FILLER_123_1808 ();
 FILLCELL_X32 FILLER_123_1840 ();
 FILLCELL_X32 FILLER_123_1872 ();
 FILLCELL_X32 FILLER_123_1904 ();
 FILLCELL_X32 FILLER_123_1936 ();
 FILLCELL_X32 FILLER_123_1968 ();
 FILLCELL_X32 FILLER_123_2000 ();
 FILLCELL_X32 FILLER_123_2032 ();
 FILLCELL_X32 FILLER_123_2064 ();
 FILLCELL_X32 FILLER_123_2096 ();
 FILLCELL_X32 FILLER_123_2128 ();
 FILLCELL_X32 FILLER_123_2160 ();
 FILLCELL_X32 FILLER_123_2192 ();
 FILLCELL_X32 FILLER_123_2224 ();
 FILLCELL_X32 FILLER_123_2256 ();
 FILLCELL_X32 FILLER_123_2288 ();
 FILLCELL_X32 FILLER_123_2320 ();
 FILLCELL_X32 FILLER_123_2352 ();
 FILLCELL_X32 FILLER_123_2384 ();
 FILLCELL_X32 FILLER_123_2416 ();
 FILLCELL_X32 FILLER_123_2448 ();
 FILLCELL_X32 FILLER_123_2480 ();
 FILLCELL_X8 FILLER_123_2512 ();
 FILLCELL_X4 FILLER_123_2520 ();
 FILLCELL_X2 FILLER_123_2524 ();
 FILLCELL_X32 FILLER_123_2527 ();
 FILLCELL_X32 FILLER_123_2559 ();
 FILLCELL_X8 FILLER_123_2591 ();
 FILLCELL_X2 FILLER_123_2599 ();
 FILLCELL_X1 FILLER_123_2601 ();
 FILLCELL_X32 FILLER_124_1 ();
 FILLCELL_X32 FILLER_124_33 ();
 FILLCELL_X32 FILLER_124_65 ();
 FILLCELL_X32 FILLER_124_97 ();
 FILLCELL_X32 FILLER_124_129 ();
 FILLCELL_X32 FILLER_124_161 ();
 FILLCELL_X32 FILLER_124_193 ();
 FILLCELL_X32 FILLER_124_225 ();
 FILLCELL_X32 FILLER_124_257 ();
 FILLCELL_X32 FILLER_124_289 ();
 FILLCELL_X32 FILLER_124_321 ();
 FILLCELL_X32 FILLER_124_353 ();
 FILLCELL_X32 FILLER_124_385 ();
 FILLCELL_X32 FILLER_124_417 ();
 FILLCELL_X32 FILLER_124_449 ();
 FILLCELL_X32 FILLER_124_481 ();
 FILLCELL_X32 FILLER_124_513 ();
 FILLCELL_X32 FILLER_124_545 ();
 FILLCELL_X32 FILLER_124_577 ();
 FILLCELL_X16 FILLER_124_609 ();
 FILLCELL_X4 FILLER_124_625 ();
 FILLCELL_X2 FILLER_124_629 ();
 FILLCELL_X32 FILLER_124_632 ();
 FILLCELL_X32 FILLER_124_664 ();
 FILLCELL_X32 FILLER_124_696 ();
 FILLCELL_X32 FILLER_124_728 ();
 FILLCELL_X32 FILLER_124_760 ();
 FILLCELL_X32 FILLER_124_792 ();
 FILLCELL_X32 FILLER_124_824 ();
 FILLCELL_X32 FILLER_124_856 ();
 FILLCELL_X32 FILLER_124_888 ();
 FILLCELL_X32 FILLER_124_920 ();
 FILLCELL_X32 FILLER_124_952 ();
 FILLCELL_X32 FILLER_124_984 ();
 FILLCELL_X32 FILLER_124_1016 ();
 FILLCELL_X32 FILLER_124_1048 ();
 FILLCELL_X32 FILLER_124_1080 ();
 FILLCELL_X32 FILLER_124_1112 ();
 FILLCELL_X32 FILLER_124_1144 ();
 FILLCELL_X32 FILLER_124_1176 ();
 FILLCELL_X32 FILLER_124_1208 ();
 FILLCELL_X32 FILLER_124_1240 ();
 FILLCELL_X32 FILLER_124_1272 ();
 FILLCELL_X32 FILLER_124_1304 ();
 FILLCELL_X32 FILLER_124_1336 ();
 FILLCELL_X32 FILLER_124_1368 ();
 FILLCELL_X32 FILLER_124_1400 ();
 FILLCELL_X32 FILLER_124_1432 ();
 FILLCELL_X32 FILLER_124_1464 ();
 FILLCELL_X32 FILLER_124_1496 ();
 FILLCELL_X32 FILLER_124_1528 ();
 FILLCELL_X32 FILLER_124_1560 ();
 FILLCELL_X32 FILLER_124_1592 ();
 FILLCELL_X32 FILLER_124_1624 ();
 FILLCELL_X32 FILLER_124_1656 ();
 FILLCELL_X32 FILLER_124_1688 ();
 FILLCELL_X32 FILLER_124_1720 ();
 FILLCELL_X32 FILLER_124_1752 ();
 FILLCELL_X32 FILLER_124_1784 ();
 FILLCELL_X32 FILLER_124_1816 ();
 FILLCELL_X32 FILLER_124_1848 ();
 FILLCELL_X8 FILLER_124_1880 ();
 FILLCELL_X4 FILLER_124_1888 ();
 FILLCELL_X2 FILLER_124_1892 ();
 FILLCELL_X32 FILLER_124_1895 ();
 FILLCELL_X32 FILLER_124_1927 ();
 FILLCELL_X32 FILLER_124_1959 ();
 FILLCELL_X32 FILLER_124_1991 ();
 FILLCELL_X32 FILLER_124_2023 ();
 FILLCELL_X32 FILLER_124_2055 ();
 FILLCELL_X32 FILLER_124_2087 ();
 FILLCELL_X32 FILLER_124_2119 ();
 FILLCELL_X32 FILLER_124_2151 ();
 FILLCELL_X32 FILLER_124_2183 ();
 FILLCELL_X32 FILLER_124_2215 ();
 FILLCELL_X32 FILLER_124_2247 ();
 FILLCELL_X32 FILLER_124_2279 ();
 FILLCELL_X32 FILLER_124_2311 ();
 FILLCELL_X32 FILLER_124_2343 ();
 FILLCELL_X32 FILLER_124_2375 ();
 FILLCELL_X32 FILLER_124_2407 ();
 FILLCELL_X32 FILLER_124_2439 ();
 FILLCELL_X32 FILLER_124_2471 ();
 FILLCELL_X32 FILLER_124_2503 ();
 FILLCELL_X32 FILLER_124_2535 ();
 FILLCELL_X32 FILLER_124_2567 ();
 FILLCELL_X2 FILLER_124_2599 ();
 FILLCELL_X1 FILLER_124_2601 ();
 FILLCELL_X32 FILLER_125_1 ();
 FILLCELL_X32 FILLER_125_33 ();
 FILLCELL_X32 FILLER_125_65 ();
 FILLCELL_X32 FILLER_125_97 ();
 FILLCELL_X32 FILLER_125_129 ();
 FILLCELL_X32 FILLER_125_161 ();
 FILLCELL_X32 FILLER_125_193 ();
 FILLCELL_X32 FILLER_125_225 ();
 FILLCELL_X32 FILLER_125_257 ();
 FILLCELL_X32 FILLER_125_289 ();
 FILLCELL_X32 FILLER_125_321 ();
 FILLCELL_X32 FILLER_125_353 ();
 FILLCELL_X32 FILLER_125_385 ();
 FILLCELL_X32 FILLER_125_417 ();
 FILLCELL_X32 FILLER_125_449 ();
 FILLCELL_X32 FILLER_125_481 ();
 FILLCELL_X32 FILLER_125_513 ();
 FILLCELL_X32 FILLER_125_545 ();
 FILLCELL_X32 FILLER_125_577 ();
 FILLCELL_X32 FILLER_125_609 ();
 FILLCELL_X32 FILLER_125_641 ();
 FILLCELL_X32 FILLER_125_673 ();
 FILLCELL_X32 FILLER_125_705 ();
 FILLCELL_X32 FILLER_125_737 ();
 FILLCELL_X32 FILLER_125_769 ();
 FILLCELL_X32 FILLER_125_801 ();
 FILLCELL_X32 FILLER_125_833 ();
 FILLCELL_X32 FILLER_125_865 ();
 FILLCELL_X32 FILLER_125_897 ();
 FILLCELL_X32 FILLER_125_929 ();
 FILLCELL_X32 FILLER_125_961 ();
 FILLCELL_X32 FILLER_125_993 ();
 FILLCELL_X32 FILLER_125_1025 ();
 FILLCELL_X32 FILLER_125_1057 ();
 FILLCELL_X32 FILLER_125_1089 ();
 FILLCELL_X32 FILLER_125_1121 ();
 FILLCELL_X32 FILLER_125_1153 ();
 FILLCELL_X32 FILLER_125_1185 ();
 FILLCELL_X32 FILLER_125_1217 ();
 FILLCELL_X8 FILLER_125_1249 ();
 FILLCELL_X4 FILLER_125_1257 ();
 FILLCELL_X2 FILLER_125_1261 ();
 FILLCELL_X32 FILLER_125_1264 ();
 FILLCELL_X32 FILLER_125_1296 ();
 FILLCELL_X32 FILLER_125_1328 ();
 FILLCELL_X32 FILLER_125_1360 ();
 FILLCELL_X32 FILLER_125_1392 ();
 FILLCELL_X32 FILLER_125_1424 ();
 FILLCELL_X32 FILLER_125_1456 ();
 FILLCELL_X32 FILLER_125_1488 ();
 FILLCELL_X32 FILLER_125_1520 ();
 FILLCELL_X32 FILLER_125_1552 ();
 FILLCELL_X32 FILLER_125_1584 ();
 FILLCELL_X32 FILLER_125_1616 ();
 FILLCELL_X32 FILLER_125_1648 ();
 FILLCELL_X32 FILLER_125_1680 ();
 FILLCELL_X32 FILLER_125_1712 ();
 FILLCELL_X32 FILLER_125_1744 ();
 FILLCELL_X32 FILLER_125_1776 ();
 FILLCELL_X32 FILLER_125_1808 ();
 FILLCELL_X32 FILLER_125_1840 ();
 FILLCELL_X32 FILLER_125_1872 ();
 FILLCELL_X32 FILLER_125_1904 ();
 FILLCELL_X32 FILLER_125_1936 ();
 FILLCELL_X32 FILLER_125_1968 ();
 FILLCELL_X32 FILLER_125_2000 ();
 FILLCELL_X32 FILLER_125_2032 ();
 FILLCELL_X32 FILLER_125_2064 ();
 FILLCELL_X32 FILLER_125_2096 ();
 FILLCELL_X32 FILLER_125_2128 ();
 FILLCELL_X32 FILLER_125_2160 ();
 FILLCELL_X32 FILLER_125_2192 ();
 FILLCELL_X32 FILLER_125_2224 ();
 FILLCELL_X32 FILLER_125_2256 ();
 FILLCELL_X32 FILLER_125_2288 ();
 FILLCELL_X32 FILLER_125_2320 ();
 FILLCELL_X32 FILLER_125_2352 ();
 FILLCELL_X32 FILLER_125_2384 ();
 FILLCELL_X32 FILLER_125_2416 ();
 FILLCELL_X32 FILLER_125_2448 ();
 FILLCELL_X32 FILLER_125_2480 ();
 FILLCELL_X8 FILLER_125_2512 ();
 FILLCELL_X4 FILLER_125_2520 ();
 FILLCELL_X2 FILLER_125_2524 ();
 FILLCELL_X32 FILLER_125_2527 ();
 FILLCELL_X32 FILLER_125_2559 ();
 FILLCELL_X8 FILLER_125_2591 ();
 FILLCELL_X2 FILLER_125_2599 ();
 FILLCELL_X1 FILLER_125_2601 ();
 FILLCELL_X32 FILLER_126_1 ();
 FILLCELL_X32 FILLER_126_33 ();
 FILLCELL_X32 FILLER_126_65 ();
 FILLCELL_X32 FILLER_126_97 ();
 FILLCELL_X32 FILLER_126_129 ();
 FILLCELL_X32 FILLER_126_161 ();
 FILLCELL_X32 FILLER_126_193 ();
 FILLCELL_X32 FILLER_126_225 ();
 FILLCELL_X32 FILLER_126_257 ();
 FILLCELL_X32 FILLER_126_289 ();
 FILLCELL_X32 FILLER_126_321 ();
 FILLCELL_X32 FILLER_126_353 ();
 FILLCELL_X32 FILLER_126_385 ();
 FILLCELL_X32 FILLER_126_417 ();
 FILLCELL_X32 FILLER_126_449 ();
 FILLCELL_X32 FILLER_126_481 ();
 FILLCELL_X32 FILLER_126_513 ();
 FILLCELL_X32 FILLER_126_545 ();
 FILLCELL_X32 FILLER_126_577 ();
 FILLCELL_X16 FILLER_126_609 ();
 FILLCELL_X4 FILLER_126_625 ();
 FILLCELL_X2 FILLER_126_629 ();
 FILLCELL_X32 FILLER_126_632 ();
 FILLCELL_X32 FILLER_126_664 ();
 FILLCELL_X32 FILLER_126_696 ();
 FILLCELL_X32 FILLER_126_728 ();
 FILLCELL_X32 FILLER_126_760 ();
 FILLCELL_X32 FILLER_126_792 ();
 FILLCELL_X32 FILLER_126_824 ();
 FILLCELL_X32 FILLER_126_856 ();
 FILLCELL_X32 FILLER_126_888 ();
 FILLCELL_X32 FILLER_126_920 ();
 FILLCELL_X32 FILLER_126_952 ();
 FILLCELL_X32 FILLER_126_984 ();
 FILLCELL_X32 FILLER_126_1016 ();
 FILLCELL_X32 FILLER_126_1048 ();
 FILLCELL_X32 FILLER_126_1080 ();
 FILLCELL_X32 FILLER_126_1112 ();
 FILLCELL_X32 FILLER_126_1144 ();
 FILLCELL_X32 FILLER_126_1176 ();
 FILLCELL_X32 FILLER_126_1208 ();
 FILLCELL_X32 FILLER_126_1240 ();
 FILLCELL_X32 FILLER_126_1272 ();
 FILLCELL_X32 FILLER_126_1304 ();
 FILLCELL_X32 FILLER_126_1336 ();
 FILLCELL_X32 FILLER_126_1368 ();
 FILLCELL_X32 FILLER_126_1400 ();
 FILLCELL_X32 FILLER_126_1432 ();
 FILLCELL_X32 FILLER_126_1464 ();
 FILLCELL_X32 FILLER_126_1496 ();
 FILLCELL_X32 FILLER_126_1528 ();
 FILLCELL_X32 FILLER_126_1560 ();
 FILLCELL_X32 FILLER_126_1592 ();
 FILLCELL_X32 FILLER_126_1624 ();
 FILLCELL_X32 FILLER_126_1656 ();
 FILLCELL_X32 FILLER_126_1688 ();
 FILLCELL_X32 FILLER_126_1720 ();
 FILLCELL_X32 FILLER_126_1752 ();
 FILLCELL_X32 FILLER_126_1784 ();
 FILLCELL_X32 FILLER_126_1816 ();
 FILLCELL_X32 FILLER_126_1848 ();
 FILLCELL_X8 FILLER_126_1880 ();
 FILLCELL_X4 FILLER_126_1888 ();
 FILLCELL_X2 FILLER_126_1892 ();
 FILLCELL_X32 FILLER_126_1895 ();
 FILLCELL_X32 FILLER_126_1927 ();
 FILLCELL_X32 FILLER_126_1959 ();
 FILLCELL_X32 FILLER_126_1991 ();
 FILLCELL_X32 FILLER_126_2023 ();
 FILLCELL_X32 FILLER_126_2055 ();
 FILLCELL_X32 FILLER_126_2087 ();
 FILLCELL_X32 FILLER_126_2119 ();
 FILLCELL_X32 FILLER_126_2151 ();
 FILLCELL_X32 FILLER_126_2183 ();
 FILLCELL_X32 FILLER_126_2215 ();
 FILLCELL_X32 FILLER_126_2247 ();
 FILLCELL_X32 FILLER_126_2279 ();
 FILLCELL_X32 FILLER_126_2311 ();
 FILLCELL_X32 FILLER_126_2343 ();
 FILLCELL_X32 FILLER_126_2375 ();
 FILLCELL_X32 FILLER_126_2407 ();
 FILLCELL_X32 FILLER_126_2439 ();
 FILLCELL_X32 FILLER_126_2471 ();
 FILLCELL_X32 FILLER_126_2503 ();
 FILLCELL_X32 FILLER_126_2535 ();
 FILLCELL_X32 FILLER_126_2567 ();
 FILLCELL_X2 FILLER_126_2599 ();
 FILLCELL_X1 FILLER_126_2601 ();
 FILLCELL_X32 FILLER_127_1 ();
 FILLCELL_X32 FILLER_127_33 ();
 FILLCELL_X32 FILLER_127_65 ();
 FILLCELL_X32 FILLER_127_97 ();
 FILLCELL_X32 FILLER_127_129 ();
 FILLCELL_X32 FILLER_127_161 ();
 FILLCELL_X32 FILLER_127_193 ();
 FILLCELL_X32 FILLER_127_225 ();
 FILLCELL_X32 FILLER_127_257 ();
 FILLCELL_X32 FILLER_127_289 ();
 FILLCELL_X32 FILLER_127_321 ();
 FILLCELL_X32 FILLER_127_353 ();
 FILLCELL_X32 FILLER_127_385 ();
 FILLCELL_X32 FILLER_127_417 ();
 FILLCELL_X32 FILLER_127_449 ();
 FILLCELL_X32 FILLER_127_481 ();
 FILLCELL_X32 FILLER_127_513 ();
 FILLCELL_X32 FILLER_127_545 ();
 FILLCELL_X32 FILLER_127_577 ();
 FILLCELL_X32 FILLER_127_609 ();
 FILLCELL_X32 FILLER_127_641 ();
 FILLCELL_X32 FILLER_127_673 ();
 FILLCELL_X32 FILLER_127_705 ();
 FILLCELL_X32 FILLER_127_737 ();
 FILLCELL_X32 FILLER_127_769 ();
 FILLCELL_X32 FILLER_127_801 ();
 FILLCELL_X32 FILLER_127_833 ();
 FILLCELL_X32 FILLER_127_865 ();
 FILLCELL_X32 FILLER_127_897 ();
 FILLCELL_X32 FILLER_127_929 ();
 FILLCELL_X32 FILLER_127_961 ();
 FILLCELL_X32 FILLER_127_993 ();
 FILLCELL_X32 FILLER_127_1025 ();
 FILLCELL_X32 FILLER_127_1057 ();
 FILLCELL_X32 FILLER_127_1089 ();
 FILLCELL_X32 FILLER_127_1121 ();
 FILLCELL_X32 FILLER_127_1153 ();
 FILLCELL_X32 FILLER_127_1185 ();
 FILLCELL_X32 FILLER_127_1217 ();
 FILLCELL_X8 FILLER_127_1249 ();
 FILLCELL_X4 FILLER_127_1257 ();
 FILLCELL_X2 FILLER_127_1261 ();
 FILLCELL_X32 FILLER_127_1264 ();
 FILLCELL_X32 FILLER_127_1296 ();
 FILLCELL_X32 FILLER_127_1328 ();
 FILLCELL_X32 FILLER_127_1360 ();
 FILLCELL_X32 FILLER_127_1392 ();
 FILLCELL_X32 FILLER_127_1424 ();
 FILLCELL_X32 FILLER_127_1456 ();
 FILLCELL_X32 FILLER_127_1488 ();
 FILLCELL_X32 FILLER_127_1520 ();
 FILLCELL_X32 FILLER_127_1552 ();
 FILLCELL_X32 FILLER_127_1584 ();
 FILLCELL_X32 FILLER_127_1616 ();
 FILLCELL_X32 FILLER_127_1648 ();
 FILLCELL_X32 FILLER_127_1680 ();
 FILLCELL_X32 FILLER_127_1712 ();
 FILLCELL_X32 FILLER_127_1744 ();
 FILLCELL_X32 FILLER_127_1776 ();
 FILLCELL_X32 FILLER_127_1808 ();
 FILLCELL_X32 FILLER_127_1840 ();
 FILLCELL_X32 FILLER_127_1872 ();
 FILLCELL_X32 FILLER_127_1904 ();
 FILLCELL_X32 FILLER_127_1936 ();
 FILLCELL_X32 FILLER_127_1968 ();
 FILLCELL_X32 FILLER_127_2000 ();
 FILLCELL_X32 FILLER_127_2032 ();
 FILLCELL_X32 FILLER_127_2064 ();
 FILLCELL_X32 FILLER_127_2096 ();
 FILLCELL_X32 FILLER_127_2128 ();
 FILLCELL_X32 FILLER_127_2160 ();
 FILLCELL_X32 FILLER_127_2192 ();
 FILLCELL_X32 FILLER_127_2224 ();
 FILLCELL_X32 FILLER_127_2256 ();
 FILLCELL_X32 FILLER_127_2288 ();
 FILLCELL_X32 FILLER_127_2320 ();
 FILLCELL_X32 FILLER_127_2352 ();
 FILLCELL_X32 FILLER_127_2384 ();
 FILLCELL_X32 FILLER_127_2416 ();
 FILLCELL_X32 FILLER_127_2448 ();
 FILLCELL_X32 FILLER_127_2480 ();
 FILLCELL_X8 FILLER_127_2512 ();
 FILLCELL_X4 FILLER_127_2520 ();
 FILLCELL_X2 FILLER_127_2524 ();
 FILLCELL_X32 FILLER_127_2527 ();
 FILLCELL_X32 FILLER_127_2559 ();
 FILLCELL_X8 FILLER_127_2591 ();
 FILLCELL_X2 FILLER_127_2599 ();
 FILLCELL_X1 FILLER_127_2601 ();
 FILLCELL_X32 FILLER_128_1 ();
 FILLCELL_X32 FILLER_128_33 ();
 FILLCELL_X32 FILLER_128_65 ();
 FILLCELL_X32 FILLER_128_97 ();
 FILLCELL_X32 FILLER_128_129 ();
 FILLCELL_X32 FILLER_128_161 ();
 FILLCELL_X32 FILLER_128_193 ();
 FILLCELL_X32 FILLER_128_225 ();
 FILLCELL_X32 FILLER_128_257 ();
 FILLCELL_X32 FILLER_128_289 ();
 FILLCELL_X32 FILLER_128_321 ();
 FILLCELL_X32 FILLER_128_353 ();
 FILLCELL_X32 FILLER_128_385 ();
 FILLCELL_X32 FILLER_128_417 ();
 FILLCELL_X32 FILLER_128_449 ();
 FILLCELL_X32 FILLER_128_481 ();
 FILLCELL_X32 FILLER_128_513 ();
 FILLCELL_X32 FILLER_128_545 ();
 FILLCELL_X32 FILLER_128_577 ();
 FILLCELL_X16 FILLER_128_609 ();
 FILLCELL_X4 FILLER_128_625 ();
 FILLCELL_X2 FILLER_128_629 ();
 FILLCELL_X32 FILLER_128_632 ();
 FILLCELL_X32 FILLER_128_664 ();
 FILLCELL_X32 FILLER_128_696 ();
 FILLCELL_X32 FILLER_128_728 ();
 FILLCELL_X32 FILLER_128_760 ();
 FILLCELL_X32 FILLER_128_792 ();
 FILLCELL_X32 FILLER_128_824 ();
 FILLCELL_X32 FILLER_128_856 ();
 FILLCELL_X32 FILLER_128_888 ();
 FILLCELL_X32 FILLER_128_920 ();
 FILLCELL_X32 FILLER_128_952 ();
 FILLCELL_X32 FILLER_128_984 ();
 FILLCELL_X32 FILLER_128_1016 ();
 FILLCELL_X32 FILLER_128_1048 ();
 FILLCELL_X32 FILLER_128_1080 ();
 FILLCELL_X32 FILLER_128_1112 ();
 FILLCELL_X32 FILLER_128_1144 ();
 FILLCELL_X32 FILLER_128_1176 ();
 FILLCELL_X32 FILLER_128_1208 ();
 FILLCELL_X32 FILLER_128_1240 ();
 FILLCELL_X32 FILLER_128_1272 ();
 FILLCELL_X32 FILLER_128_1304 ();
 FILLCELL_X32 FILLER_128_1336 ();
 FILLCELL_X32 FILLER_128_1368 ();
 FILLCELL_X32 FILLER_128_1400 ();
 FILLCELL_X32 FILLER_128_1432 ();
 FILLCELL_X32 FILLER_128_1464 ();
 FILLCELL_X32 FILLER_128_1496 ();
 FILLCELL_X32 FILLER_128_1528 ();
 FILLCELL_X32 FILLER_128_1560 ();
 FILLCELL_X32 FILLER_128_1592 ();
 FILLCELL_X32 FILLER_128_1624 ();
 FILLCELL_X32 FILLER_128_1656 ();
 FILLCELL_X32 FILLER_128_1688 ();
 FILLCELL_X32 FILLER_128_1720 ();
 FILLCELL_X32 FILLER_128_1752 ();
 FILLCELL_X32 FILLER_128_1784 ();
 FILLCELL_X32 FILLER_128_1816 ();
 FILLCELL_X32 FILLER_128_1848 ();
 FILLCELL_X8 FILLER_128_1880 ();
 FILLCELL_X4 FILLER_128_1888 ();
 FILLCELL_X2 FILLER_128_1892 ();
 FILLCELL_X32 FILLER_128_1895 ();
 FILLCELL_X32 FILLER_128_1927 ();
 FILLCELL_X32 FILLER_128_1959 ();
 FILLCELL_X32 FILLER_128_1991 ();
 FILLCELL_X32 FILLER_128_2023 ();
 FILLCELL_X32 FILLER_128_2055 ();
 FILLCELL_X32 FILLER_128_2087 ();
 FILLCELL_X32 FILLER_128_2119 ();
 FILLCELL_X32 FILLER_128_2151 ();
 FILLCELL_X32 FILLER_128_2183 ();
 FILLCELL_X32 FILLER_128_2215 ();
 FILLCELL_X32 FILLER_128_2247 ();
 FILLCELL_X32 FILLER_128_2279 ();
 FILLCELL_X32 FILLER_128_2311 ();
 FILLCELL_X32 FILLER_128_2343 ();
 FILLCELL_X32 FILLER_128_2375 ();
 FILLCELL_X32 FILLER_128_2407 ();
 FILLCELL_X32 FILLER_128_2439 ();
 FILLCELL_X32 FILLER_128_2471 ();
 FILLCELL_X32 FILLER_128_2503 ();
 FILLCELL_X32 FILLER_128_2535 ();
 FILLCELL_X32 FILLER_128_2567 ();
 FILLCELL_X2 FILLER_128_2599 ();
 FILLCELL_X1 FILLER_128_2601 ();
 FILLCELL_X32 FILLER_129_1 ();
 FILLCELL_X32 FILLER_129_33 ();
 FILLCELL_X32 FILLER_129_65 ();
 FILLCELL_X32 FILLER_129_97 ();
 FILLCELL_X32 FILLER_129_129 ();
 FILLCELL_X32 FILLER_129_161 ();
 FILLCELL_X32 FILLER_129_193 ();
 FILLCELL_X32 FILLER_129_225 ();
 FILLCELL_X32 FILLER_129_257 ();
 FILLCELL_X32 FILLER_129_289 ();
 FILLCELL_X32 FILLER_129_321 ();
 FILLCELL_X32 FILLER_129_353 ();
 FILLCELL_X32 FILLER_129_385 ();
 FILLCELL_X32 FILLER_129_417 ();
 FILLCELL_X32 FILLER_129_449 ();
 FILLCELL_X32 FILLER_129_481 ();
 FILLCELL_X32 FILLER_129_513 ();
 FILLCELL_X32 FILLER_129_545 ();
 FILLCELL_X32 FILLER_129_577 ();
 FILLCELL_X32 FILLER_129_609 ();
 FILLCELL_X32 FILLER_129_641 ();
 FILLCELL_X32 FILLER_129_673 ();
 FILLCELL_X32 FILLER_129_705 ();
 FILLCELL_X32 FILLER_129_737 ();
 FILLCELL_X32 FILLER_129_769 ();
 FILLCELL_X32 FILLER_129_801 ();
 FILLCELL_X32 FILLER_129_833 ();
 FILLCELL_X32 FILLER_129_865 ();
 FILLCELL_X32 FILLER_129_897 ();
 FILLCELL_X32 FILLER_129_929 ();
 FILLCELL_X32 FILLER_129_961 ();
 FILLCELL_X32 FILLER_129_993 ();
 FILLCELL_X32 FILLER_129_1025 ();
 FILLCELL_X32 FILLER_129_1057 ();
 FILLCELL_X32 FILLER_129_1089 ();
 FILLCELL_X32 FILLER_129_1121 ();
 FILLCELL_X32 FILLER_129_1153 ();
 FILLCELL_X32 FILLER_129_1185 ();
 FILLCELL_X32 FILLER_129_1217 ();
 FILLCELL_X8 FILLER_129_1249 ();
 FILLCELL_X4 FILLER_129_1257 ();
 FILLCELL_X2 FILLER_129_1261 ();
 FILLCELL_X32 FILLER_129_1264 ();
 FILLCELL_X32 FILLER_129_1296 ();
 FILLCELL_X32 FILLER_129_1328 ();
 FILLCELL_X32 FILLER_129_1360 ();
 FILLCELL_X32 FILLER_129_1392 ();
 FILLCELL_X32 FILLER_129_1424 ();
 FILLCELL_X32 FILLER_129_1456 ();
 FILLCELL_X32 FILLER_129_1488 ();
 FILLCELL_X32 FILLER_129_1520 ();
 FILLCELL_X32 FILLER_129_1552 ();
 FILLCELL_X32 FILLER_129_1584 ();
 FILLCELL_X32 FILLER_129_1616 ();
 FILLCELL_X32 FILLER_129_1648 ();
 FILLCELL_X32 FILLER_129_1680 ();
 FILLCELL_X32 FILLER_129_1712 ();
 FILLCELL_X32 FILLER_129_1744 ();
 FILLCELL_X32 FILLER_129_1776 ();
 FILLCELL_X32 FILLER_129_1808 ();
 FILLCELL_X32 FILLER_129_1840 ();
 FILLCELL_X32 FILLER_129_1872 ();
 FILLCELL_X32 FILLER_129_1904 ();
 FILLCELL_X32 FILLER_129_1936 ();
 FILLCELL_X32 FILLER_129_1968 ();
 FILLCELL_X32 FILLER_129_2000 ();
 FILLCELL_X32 FILLER_129_2032 ();
 FILLCELL_X32 FILLER_129_2064 ();
 FILLCELL_X32 FILLER_129_2096 ();
 FILLCELL_X32 FILLER_129_2128 ();
 FILLCELL_X32 FILLER_129_2160 ();
 FILLCELL_X32 FILLER_129_2192 ();
 FILLCELL_X32 FILLER_129_2224 ();
 FILLCELL_X32 FILLER_129_2256 ();
 FILLCELL_X32 FILLER_129_2288 ();
 FILLCELL_X32 FILLER_129_2320 ();
 FILLCELL_X32 FILLER_129_2352 ();
 FILLCELL_X32 FILLER_129_2384 ();
 FILLCELL_X32 FILLER_129_2416 ();
 FILLCELL_X32 FILLER_129_2448 ();
 FILLCELL_X32 FILLER_129_2480 ();
 FILLCELL_X8 FILLER_129_2512 ();
 FILLCELL_X4 FILLER_129_2520 ();
 FILLCELL_X2 FILLER_129_2524 ();
 FILLCELL_X32 FILLER_129_2527 ();
 FILLCELL_X32 FILLER_129_2559 ();
 FILLCELL_X8 FILLER_129_2591 ();
 FILLCELL_X2 FILLER_129_2599 ();
 FILLCELL_X1 FILLER_129_2601 ();
 FILLCELL_X32 FILLER_130_1 ();
 FILLCELL_X32 FILLER_130_33 ();
 FILLCELL_X32 FILLER_130_65 ();
 FILLCELL_X32 FILLER_130_97 ();
 FILLCELL_X32 FILLER_130_129 ();
 FILLCELL_X32 FILLER_130_161 ();
 FILLCELL_X32 FILLER_130_193 ();
 FILLCELL_X32 FILLER_130_225 ();
 FILLCELL_X32 FILLER_130_257 ();
 FILLCELL_X32 FILLER_130_289 ();
 FILLCELL_X32 FILLER_130_321 ();
 FILLCELL_X32 FILLER_130_353 ();
 FILLCELL_X32 FILLER_130_385 ();
 FILLCELL_X32 FILLER_130_417 ();
 FILLCELL_X32 FILLER_130_449 ();
 FILLCELL_X32 FILLER_130_481 ();
 FILLCELL_X32 FILLER_130_513 ();
 FILLCELL_X32 FILLER_130_545 ();
 FILLCELL_X32 FILLER_130_577 ();
 FILLCELL_X16 FILLER_130_609 ();
 FILLCELL_X4 FILLER_130_625 ();
 FILLCELL_X2 FILLER_130_629 ();
 FILLCELL_X32 FILLER_130_632 ();
 FILLCELL_X32 FILLER_130_664 ();
 FILLCELL_X32 FILLER_130_696 ();
 FILLCELL_X32 FILLER_130_728 ();
 FILLCELL_X32 FILLER_130_760 ();
 FILLCELL_X32 FILLER_130_792 ();
 FILLCELL_X32 FILLER_130_824 ();
 FILLCELL_X32 FILLER_130_856 ();
 FILLCELL_X32 FILLER_130_888 ();
 FILLCELL_X32 FILLER_130_920 ();
 FILLCELL_X32 FILLER_130_952 ();
 FILLCELL_X32 FILLER_130_984 ();
 FILLCELL_X32 FILLER_130_1016 ();
 FILLCELL_X32 FILLER_130_1048 ();
 FILLCELL_X32 FILLER_130_1080 ();
 FILLCELL_X32 FILLER_130_1112 ();
 FILLCELL_X32 FILLER_130_1144 ();
 FILLCELL_X32 FILLER_130_1176 ();
 FILLCELL_X32 FILLER_130_1208 ();
 FILLCELL_X32 FILLER_130_1240 ();
 FILLCELL_X32 FILLER_130_1272 ();
 FILLCELL_X32 FILLER_130_1304 ();
 FILLCELL_X32 FILLER_130_1336 ();
 FILLCELL_X32 FILLER_130_1368 ();
 FILLCELL_X32 FILLER_130_1400 ();
 FILLCELL_X32 FILLER_130_1432 ();
 FILLCELL_X32 FILLER_130_1464 ();
 FILLCELL_X32 FILLER_130_1496 ();
 FILLCELL_X32 FILLER_130_1528 ();
 FILLCELL_X32 FILLER_130_1560 ();
 FILLCELL_X32 FILLER_130_1592 ();
 FILLCELL_X32 FILLER_130_1624 ();
 FILLCELL_X32 FILLER_130_1656 ();
 FILLCELL_X32 FILLER_130_1688 ();
 FILLCELL_X32 FILLER_130_1720 ();
 FILLCELL_X32 FILLER_130_1752 ();
 FILLCELL_X32 FILLER_130_1784 ();
 FILLCELL_X32 FILLER_130_1816 ();
 FILLCELL_X32 FILLER_130_1848 ();
 FILLCELL_X8 FILLER_130_1880 ();
 FILLCELL_X4 FILLER_130_1888 ();
 FILLCELL_X2 FILLER_130_1892 ();
 FILLCELL_X32 FILLER_130_1895 ();
 FILLCELL_X32 FILLER_130_1927 ();
 FILLCELL_X32 FILLER_130_1959 ();
 FILLCELL_X32 FILLER_130_1991 ();
 FILLCELL_X32 FILLER_130_2023 ();
 FILLCELL_X32 FILLER_130_2055 ();
 FILLCELL_X32 FILLER_130_2087 ();
 FILLCELL_X32 FILLER_130_2119 ();
 FILLCELL_X32 FILLER_130_2151 ();
 FILLCELL_X32 FILLER_130_2183 ();
 FILLCELL_X32 FILLER_130_2215 ();
 FILLCELL_X32 FILLER_130_2247 ();
 FILLCELL_X32 FILLER_130_2279 ();
 FILLCELL_X32 FILLER_130_2311 ();
 FILLCELL_X32 FILLER_130_2343 ();
 FILLCELL_X32 FILLER_130_2375 ();
 FILLCELL_X32 FILLER_130_2407 ();
 FILLCELL_X32 FILLER_130_2439 ();
 FILLCELL_X32 FILLER_130_2471 ();
 FILLCELL_X32 FILLER_130_2503 ();
 FILLCELL_X32 FILLER_130_2535 ();
 FILLCELL_X32 FILLER_130_2567 ();
 FILLCELL_X2 FILLER_130_2599 ();
 FILLCELL_X1 FILLER_130_2601 ();
 FILLCELL_X32 FILLER_131_1 ();
 FILLCELL_X32 FILLER_131_33 ();
 FILLCELL_X32 FILLER_131_65 ();
 FILLCELL_X32 FILLER_131_97 ();
 FILLCELL_X32 FILLER_131_129 ();
 FILLCELL_X32 FILLER_131_161 ();
 FILLCELL_X32 FILLER_131_193 ();
 FILLCELL_X32 FILLER_131_225 ();
 FILLCELL_X32 FILLER_131_257 ();
 FILLCELL_X32 FILLER_131_289 ();
 FILLCELL_X32 FILLER_131_321 ();
 FILLCELL_X32 FILLER_131_353 ();
 FILLCELL_X32 FILLER_131_385 ();
 FILLCELL_X32 FILLER_131_417 ();
 FILLCELL_X32 FILLER_131_449 ();
 FILLCELL_X32 FILLER_131_481 ();
 FILLCELL_X32 FILLER_131_513 ();
 FILLCELL_X32 FILLER_131_545 ();
 FILLCELL_X32 FILLER_131_577 ();
 FILLCELL_X32 FILLER_131_609 ();
 FILLCELL_X32 FILLER_131_641 ();
 FILLCELL_X32 FILLER_131_673 ();
 FILLCELL_X32 FILLER_131_705 ();
 FILLCELL_X32 FILLER_131_737 ();
 FILLCELL_X32 FILLER_131_769 ();
 FILLCELL_X32 FILLER_131_801 ();
 FILLCELL_X32 FILLER_131_833 ();
 FILLCELL_X32 FILLER_131_865 ();
 FILLCELL_X32 FILLER_131_897 ();
 FILLCELL_X32 FILLER_131_929 ();
 FILLCELL_X32 FILLER_131_961 ();
 FILLCELL_X32 FILLER_131_993 ();
 FILLCELL_X32 FILLER_131_1025 ();
 FILLCELL_X32 FILLER_131_1057 ();
 FILLCELL_X32 FILLER_131_1089 ();
 FILLCELL_X32 FILLER_131_1121 ();
 FILLCELL_X32 FILLER_131_1153 ();
 FILLCELL_X32 FILLER_131_1185 ();
 FILLCELL_X32 FILLER_131_1217 ();
 FILLCELL_X8 FILLER_131_1249 ();
 FILLCELL_X4 FILLER_131_1257 ();
 FILLCELL_X2 FILLER_131_1261 ();
 FILLCELL_X32 FILLER_131_1264 ();
 FILLCELL_X32 FILLER_131_1296 ();
 FILLCELL_X32 FILLER_131_1328 ();
 FILLCELL_X32 FILLER_131_1360 ();
 FILLCELL_X32 FILLER_131_1392 ();
 FILLCELL_X32 FILLER_131_1424 ();
 FILLCELL_X32 FILLER_131_1456 ();
 FILLCELL_X32 FILLER_131_1488 ();
 FILLCELL_X32 FILLER_131_1520 ();
 FILLCELL_X32 FILLER_131_1552 ();
 FILLCELL_X32 FILLER_131_1584 ();
 FILLCELL_X32 FILLER_131_1616 ();
 FILLCELL_X32 FILLER_131_1648 ();
 FILLCELL_X32 FILLER_131_1680 ();
 FILLCELL_X32 FILLER_131_1712 ();
 FILLCELL_X32 FILLER_131_1744 ();
 FILLCELL_X32 FILLER_131_1776 ();
 FILLCELL_X32 FILLER_131_1808 ();
 FILLCELL_X32 FILLER_131_1840 ();
 FILLCELL_X32 FILLER_131_1872 ();
 FILLCELL_X32 FILLER_131_1904 ();
 FILLCELL_X32 FILLER_131_1936 ();
 FILLCELL_X32 FILLER_131_1968 ();
 FILLCELL_X32 FILLER_131_2000 ();
 FILLCELL_X32 FILLER_131_2032 ();
 FILLCELL_X32 FILLER_131_2064 ();
 FILLCELL_X32 FILLER_131_2096 ();
 FILLCELL_X32 FILLER_131_2128 ();
 FILLCELL_X32 FILLER_131_2160 ();
 FILLCELL_X32 FILLER_131_2192 ();
 FILLCELL_X32 FILLER_131_2224 ();
 FILLCELL_X32 FILLER_131_2256 ();
 FILLCELL_X32 FILLER_131_2288 ();
 FILLCELL_X32 FILLER_131_2320 ();
 FILLCELL_X32 FILLER_131_2352 ();
 FILLCELL_X32 FILLER_131_2384 ();
 FILLCELL_X32 FILLER_131_2416 ();
 FILLCELL_X32 FILLER_131_2448 ();
 FILLCELL_X32 FILLER_131_2480 ();
 FILLCELL_X8 FILLER_131_2512 ();
 FILLCELL_X4 FILLER_131_2520 ();
 FILLCELL_X2 FILLER_131_2524 ();
 FILLCELL_X32 FILLER_131_2527 ();
 FILLCELL_X32 FILLER_131_2559 ();
 FILLCELL_X8 FILLER_131_2591 ();
 FILLCELL_X2 FILLER_131_2599 ();
 FILLCELL_X1 FILLER_131_2601 ();
 FILLCELL_X32 FILLER_132_1 ();
 FILLCELL_X32 FILLER_132_33 ();
 FILLCELL_X32 FILLER_132_65 ();
 FILLCELL_X32 FILLER_132_97 ();
 FILLCELL_X32 FILLER_132_129 ();
 FILLCELL_X32 FILLER_132_161 ();
 FILLCELL_X32 FILLER_132_193 ();
 FILLCELL_X32 FILLER_132_225 ();
 FILLCELL_X32 FILLER_132_257 ();
 FILLCELL_X32 FILLER_132_289 ();
 FILLCELL_X32 FILLER_132_321 ();
 FILLCELL_X32 FILLER_132_353 ();
 FILLCELL_X32 FILLER_132_385 ();
 FILLCELL_X32 FILLER_132_417 ();
 FILLCELL_X32 FILLER_132_449 ();
 FILLCELL_X32 FILLER_132_481 ();
 FILLCELL_X32 FILLER_132_513 ();
 FILLCELL_X32 FILLER_132_545 ();
 FILLCELL_X32 FILLER_132_577 ();
 FILLCELL_X16 FILLER_132_609 ();
 FILLCELL_X4 FILLER_132_625 ();
 FILLCELL_X2 FILLER_132_629 ();
 FILLCELL_X32 FILLER_132_632 ();
 FILLCELL_X32 FILLER_132_664 ();
 FILLCELL_X32 FILLER_132_696 ();
 FILLCELL_X32 FILLER_132_728 ();
 FILLCELL_X32 FILLER_132_760 ();
 FILLCELL_X32 FILLER_132_792 ();
 FILLCELL_X32 FILLER_132_824 ();
 FILLCELL_X32 FILLER_132_856 ();
 FILLCELL_X32 FILLER_132_888 ();
 FILLCELL_X32 FILLER_132_920 ();
 FILLCELL_X32 FILLER_132_952 ();
 FILLCELL_X32 FILLER_132_984 ();
 FILLCELL_X32 FILLER_132_1016 ();
 FILLCELL_X32 FILLER_132_1048 ();
 FILLCELL_X32 FILLER_132_1080 ();
 FILLCELL_X32 FILLER_132_1112 ();
 FILLCELL_X32 FILLER_132_1144 ();
 FILLCELL_X32 FILLER_132_1176 ();
 FILLCELL_X32 FILLER_132_1208 ();
 FILLCELL_X32 FILLER_132_1240 ();
 FILLCELL_X32 FILLER_132_1272 ();
 FILLCELL_X32 FILLER_132_1304 ();
 FILLCELL_X32 FILLER_132_1336 ();
 FILLCELL_X32 FILLER_132_1368 ();
 FILLCELL_X32 FILLER_132_1400 ();
 FILLCELL_X32 FILLER_132_1432 ();
 FILLCELL_X32 FILLER_132_1464 ();
 FILLCELL_X32 FILLER_132_1496 ();
 FILLCELL_X32 FILLER_132_1528 ();
 FILLCELL_X32 FILLER_132_1560 ();
 FILLCELL_X32 FILLER_132_1592 ();
 FILLCELL_X32 FILLER_132_1624 ();
 FILLCELL_X32 FILLER_132_1656 ();
 FILLCELL_X32 FILLER_132_1688 ();
 FILLCELL_X32 FILLER_132_1720 ();
 FILLCELL_X32 FILLER_132_1752 ();
 FILLCELL_X32 FILLER_132_1784 ();
 FILLCELL_X32 FILLER_132_1816 ();
 FILLCELL_X32 FILLER_132_1848 ();
 FILLCELL_X8 FILLER_132_1880 ();
 FILLCELL_X4 FILLER_132_1888 ();
 FILLCELL_X2 FILLER_132_1892 ();
 FILLCELL_X32 FILLER_132_1895 ();
 FILLCELL_X32 FILLER_132_1927 ();
 FILLCELL_X32 FILLER_132_1959 ();
 FILLCELL_X32 FILLER_132_1991 ();
 FILLCELL_X32 FILLER_132_2023 ();
 FILLCELL_X32 FILLER_132_2055 ();
 FILLCELL_X32 FILLER_132_2087 ();
 FILLCELL_X32 FILLER_132_2119 ();
 FILLCELL_X32 FILLER_132_2151 ();
 FILLCELL_X32 FILLER_132_2183 ();
 FILLCELL_X32 FILLER_132_2215 ();
 FILLCELL_X32 FILLER_132_2247 ();
 FILLCELL_X32 FILLER_132_2279 ();
 FILLCELL_X32 FILLER_132_2311 ();
 FILLCELL_X32 FILLER_132_2343 ();
 FILLCELL_X32 FILLER_132_2375 ();
 FILLCELL_X32 FILLER_132_2407 ();
 FILLCELL_X32 FILLER_132_2439 ();
 FILLCELL_X32 FILLER_132_2471 ();
 FILLCELL_X32 FILLER_132_2503 ();
 FILLCELL_X32 FILLER_132_2535 ();
 FILLCELL_X32 FILLER_132_2567 ();
 FILLCELL_X2 FILLER_132_2599 ();
 FILLCELL_X1 FILLER_132_2601 ();
 FILLCELL_X32 FILLER_133_1 ();
 FILLCELL_X32 FILLER_133_33 ();
 FILLCELL_X32 FILLER_133_65 ();
 FILLCELL_X32 FILLER_133_97 ();
 FILLCELL_X32 FILLER_133_129 ();
 FILLCELL_X32 FILLER_133_161 ();
 FILLCELL_X32 FILLER_133_193 ();
 FILLCELL_X32 FILLER_133_225 ();
 FILLCELL_X32 FILLER_133_257 ();
 FILLCELL_X32 FILLER_133_289 ();
 FILLCELL_X32 FILLER_133_321 ();
 FILLCELL_X32 FILLER_133_353 ();
 FILLCELL_X32 FILLER_133_385 ();
 FILLCELL_X32 FILLER_133_417 ();
 FILLCELL_X32 FILLER_133_449 ();
 FILLCELL_X32 FILLER_133_481 ();
 FILLCELL_X32 FILLER_133_513 ();
 FILLCELL_X32 FILLER_133_545 ();
 FILLCELL_X32 FILLER_133_577 ();
 FILLCELL_X32 FILLER_133_609 ();
 FILLCELL_X32 FILLER_133_641 ();
 FILLCELL_X32 FILLER_133_673 ();
 FILLCELL_X32 FILLER_133_705 ();
 FILLCELL_X32 FILLER_133_737 ();
 FILLCELL_X32 FILLER_133_769 ();
 FILLCELL_X32 FILLER_133_801 ();
 FILLCELL_X32 FILLER_133_833 ();
 FILLCELL_X32 FILLER_133_865 ();
 FILLCELL_X32 FILLER_133_897 ();
 FILLCELL_X32 FILLER_133_929 ();
 FILLCELL_X32 FILLER_133_961 ();
 FILLCELL_X32 FILLER_133_993 ();
 FILLCELL_X32 FILLER_133_1025 ();
 FILLCELL_X32 FILLER_133_1057 ();
 FILLCELL_X32 FILLER_133_1089 ();
 FILLCELL_X32 FILLER_133_1121 ();
 FILLCELL_X32 FILLER_133_1153 ();
 FILLCELL_X32 FILLER_133_1185 ();
 FILLCELL_X32 FILLER_133_1217 ();
 FILLCELL_X8 FILLER_133_1249 ();
 FILLCELL_X4 FILLER_133_1257 ();
 FILLCELL_X2 FILLER_133_1261 ();
 FILLCELL_X32 FILLER_133_1264 ();
 FILLCELL_X32 FILLER_133_1296 ();
 FILLCELL_X32 FILLER_133_1328 ();
 FILLCELL_X32 FILLER_133_1360 ();
 FILLCELL_X32 FILLER_133_1392 ();
 FILLCELL_X32 FILLER_133_1424 ();
 FILLCELL_X32 FILLER_133_1456 ();
 FILLCELL_X32 FILLER_133_1488 ();
 FILLCELL_X32 FILLER_133_1520 ();
 FILLCELL_X32 FILLER_133_1552 ();
 FILLCELL_X32 FILLER_133_1584 ();
 FILLCELL_X32 FILLER_133_1616 ();
 FILLCELL_X32 FILLER_133_1648 ();
 FILLCELL_X32 FILLER_133_1680 ();
 FILLCELL_X32 FILLER_133_1712 ();
 FILLCELL_X32 FILLER_133_1744 ();
 FILLCELL_X32 FILLER_133_1776 ();
 FILLCELL_X32 FILLER_133_1808 ();
 FILLCELL_X32 FILLER_133_1840 ();
 FILLCELL_X32 FILLER_133_1872 ();
 FILLCELL_X32 FILLER_133_1904 ();
 FILLCELL_X32 FILLER_133_1936 ();
 FILLCELL_X32 FILLER_133_1968 ();
 FILLCELL_X32 FILLER_133_2000 ();
 FILLCELL_X32 FILLER_133_2032 ();
 FILLCELL_X32 FILLER_133_2064 ();
 FILLCELL_X32 FILLER_133_2096 ();
 FILLCELL_X32 FILLER_133_2128 ();
 FILLCELL_X32 FILLER_133_2160 ();
 FILLCELL_X32 FILLER_133_2192 ();
 FILLCELL_X32 FILLER_133_2224 ();
 FILLCELL_X32 FILLER_133_2256 ();
 FILLCELL_X32 FILLER_133_2288 ();
 FILLCELL_X32 FILLER_133_2320 ();
 FILLCELL_X32 FILLER_133_2352 ();
 FILLCELL_X32 FILLER_133_2384 ();
 FILLCELL_X32 FILLER_133_2416 ();
 FILLCELL_X32 FILLER_133_2448 ();
 FILLCELL_X32 FILLER_133_2480 ();
 FILLCELL_X8 FILLER_133_2512 ();
 FILLCELL_X4 FILLER_133_2520 ();
 FILLCELL_X2 FILLER_133_2524 ();
 FILLCELL_X32 FILLER_133_2527 ();
 FILLCELL_X32 FILLER_133_2559 ();
 FILLCELL_X8 FILLER_133_2591 ();
 FILLCELL_X2 FILLER_133_2599 ();
 FILLCELL_X1 FILLER_133_2601 ();
 FILLCELL_X32 FILLER_134_1 ();
 FILLCELL_X32 FILLER_134_33 ();
 FILLCELL_X32 FILLER_134_65 ();
 FILLCELL_X32 FILLER_134_97 ();
 FILLCELL_X32 FILLER_134_129 ();
 FILLCELL_X32 FILLER_134_161 ();
 FILLCELL_X32 FILLER_134_193 ();
 FILLCELL_X32 FILLER_134_225 ();
 FILLCELL_X32 FILLER_134_257 ();
 FILLCELL_X32 FILLER_134_289 ();
 FILLCELL_X32 FILLER_134_321 ();
 FILLCELL_X32 FILLER_134_353 ();
 FILLCELL_X32 FILLER_134_385 ();
 FILLCELL_X32 FILLER_134_417 ();
 FILLCELL_X32 FILLER_134_449 ();
 FILLCELL_X32 FILLER_134_481 ();
 FILLCELL_X32 FILLER_134_513 ();
 FILLCELL_X32 FILLER_134_545 ();
 FILLCELL_X32 FILLER_134_577 ();
 FILLCELL_X16 FILLER_134_609 ();
 FILLCELL_X4 FILLER_134_625 ();
 FILLCELL_X2 FILLER_134_629 ();
 FILLCELL_X32 FILLER_134_632 ();
 FILLCELL_X32 FILLER_134_664 ();
 FILLCELL_X32 FILLER_134_696 ();
 FILLCELL_X32 FILLER_134_728 ();
 FILLCELL_X32 FILLER_134_760 ();
 FILLCELL_X32 FILLER_134_792 ();
 FILLCELL_X32 FILLER_134_824 ();
 FILLCELL_X32 FILLER_134_856 ();
 FILLCELL_X32 FILLER_134_888 ();
 FILLCELL_X32 FILLER_134_920 ();
 FILLCELL_X32 FILLER_134_952 ();
 FILLCELL_X32 FILLER_134_984 ();
 FILLCELL_X32 FILLER_134_1016 ();
 FILLCELL_X32 FILLER_134_1048 ();
 FILLCELL_X32 FILLER_134_1080 ();
 FILLCELL_X32 FILLER_134_1112 ();
 FILLCELL_X32 FILLER_134_1144 ();
 FILLCELL_X32 FILLER_134_1176 ();
 FILLCELL_X32 FILLER_134_1208 ();
 FILLCELL_X32 FILLER_134_1240 ();
 FILLCELL_X32 FILLER_134_1272 ();
 FILLCELL_X32 FILLER_134_1304 ();
 FILLCELL_X32 FILLER_134_1336 ();
 FILLCELL_X32 FILLER_134_1368 ();
 FILLCELL_X32 FILLER_134_1400 ();
 FILLCELL_X32 FILLER_134_1432 ();
 FILLCELL_X32 FILLER_134_1464 ();
 FILLCELL_X32 FILLER_134_1496 ();
 FILLCELL_X32 FILLER_134_1528 ();
 FILLCELL_X32 FILLER_134_1560 ();
 FILLCELL_X32 FILLER_134_1592 ();
 FILLCELL_X32 FILLER_134_1624 ();
 FILLCELL_X32 FILLER_134_1656 ();
 FILLCELL_X32 FILLER_134_1688 ();
 FILLCELL_X32 FILLER_134_1720 ();
 FILLCELL_X32 FILLER_134_1752 ();
 FILLCELL_X32 FILLER_134_1784 ();
 FILLCELL_X32 FILLER_134_1816 ();
 FILLCELL_X32 FILLER_134_1848 ();
 FILLCELL_X8 FILLER_134_1880 ();
 FILLCELL_X4 FILLER_134_1888 ();
 FILLCELL_X2 FILLER_134_1892 ();
 FILLCELL_X32 FILLER_134_1895 ();
 FILLCELL_X32 FILLER_134_1927 ();
 FILLCELL_X32 FILLER_134_1959 ();
 FILLCELL_X32 FILLER_134_1991 ();
 FILLCELL_X32 FILLER_134_2023 ();
 FILLCELL_X32 FILLER_134_2055 ();
 FILLCELL_X32 FILLER_134_2087 ();
 FILLCELL_X32 FILLER_134_2119 ();
 FILLCELL_X32 FILLER_134_2151 ();
 FILLCELL_X32 FILLER_134_2183 ();
 FILLCELL_X32 FILLER_134_2215 ();
 FILLCELL_X32 FILLER_134_2247 ();
 FILLCELL_X32 FILLER_134_2279 ();
 FILLCELL_X32 FILLER_134_2311 ();
 FILLCELL_X32 FILLER_134_2343 ();
 FILLCELL_X32 FILLER_134_2375 ();
 FILLCELL_X32 FILLER_134_2407 ();
 FILLCELL_X32 FILLER_134_2439 ();
 FILLCELL_X32 FILLER_134_2471 ();
 FILLCELL_X32 FILLER_134_2503 ();
 FILLCELL_X32 FILLER_134_2535 ();
 FILLCELL_X32 FILLER_134_2567 ();
 FILLCELL_X2 FILLER_134_2599 ();
 FILLCELL_X1 FILLER_134_2601 ();
 FILLCELL_X32 FILLER_135_1 ();
 FILLCELL_X32 FILLER_135_33 ();
 FILLCELL_X32 FILLER_135_65 ();
 FILLCELL_X32 FILLER_135_97 ();
 FILLCELL_X32 FILLER_135_129 ();
 FILLCELL_X32 FILLER_135_161 ();
 FILLCELL_X32 FILLER_135_193 ();
 FILLCELL_X32 FILLER_135_225 ();
 FILLCELL_X32 FILLER_135_257 ();
 FILLCELL_X32 FILLER_135_289 ();
 FILLCELL_X32 FILLER_135_321 ();
 FILLCELL_X32 FILLER_135_353 ();
 FILLCELL_X32 FILLER_135_385 ();
 FILLCELL_X32 FILLER_135_417 ();
 FILLCELL_X32 FILLER_135_449 ();
 FILLCELL_X32 FILLER_135_481 ();
 FILLCELL_X32 FILLER_135_513 ();
 FILLCELL_X32 FILLER_135_545 ();
 FILLCELL_X32 FILLER_135_577 ();
 FILLCELL_X32 FILLER_135_609 ();
 FILLCELL_X32 FILLER_135_641 ();
 FILLCELL_X32 FILLER_135_673 ();
 FILLCELL_X32 FILLER_135_705 ();
 FILLCELL_X32 FILLER_135_737 ();
 FILLCELL_X32 FILLER_135_769 ();
 FILLCELL_X32 FILLER_135_801 ();
 FILLCELL_X32 FILLER_135_833 ();
 FILLCELL_X32 FILLER_135_865 ();
 FILLCELL_X32 FILLER_135_897 ();
 FILLCELL_X32 FILLER_135_929 ();
 FILLCELL_X32 FILLER_135_961 ();
 FILLCELL_X32 FILLER_135_993 ();
 FILLCELL_X32 FILLER_135_1025 ();
 FILLCELL_X32 FILLER_135_1057 ();
 FILLCELL_X32 FILLER_135_1089 ();
 FILLCELL_X32 FILLER_135_1121 ();
 FILLCELL_X32 FILLER_135_1153 ();
 FILLCELL_X32 FILLER_135_1185 ();
 FILLCELL_X32 FILLER_135_1217 ();
 FILLCELL_X8 FILLER_135_1249 ();
 FILLCELL_X4 FILLER_135_1257 ();
 FILLCELL_X2 FILLER_135_1261 ();
 FILLCELL_X32 FILLER_135_1264 ();
 FILLCELL_X32 FILLER_135_1296 ();
 FILLCELL_X32 FILLER_135_1328 ();
 FILLCELL_X32 FILLER_135_1360 ();
 FILLCELL_X32 FILLER_135_1392 ();
 FILLCELL_X32 FILLER_135_1424 ();
 FILLCELL_X32 FILLER_135_1456 ();
 FILLCELL_X32 FILLER_135_1488 ();
 FILLCELL_X32 FILLER_135_1520 ();
 FILLCELL_X32 FILLER_135_1552 ();
 FILLCELL_X32 FILLER_135_1584 ();
 FILLCELL_X32 FILLER_135_1616 ();
 FILLCELL_X32 FILLER_135_1648 ();
 FILLCELL_X32 FILLER_135_1680 ();
 FILLCELL_X32 FILLER_135_1712 ();
 FILLCELL_X32 FILLER_135_1744 ();
 FILLCELL_X32 FILLER_135_1776 ();
 FILLCELL_X32 FILLER_135_1808 ();
 FILLCELL_X32 FILLER_135_1840 ();
 FILLCELL_X32 FILLER_135_1872 ();
 FILLCELL_X32 FILLER_135_1904 ();
 FILLCELL_X32 FILLER_135_1936 ();
 FILLCELL_X32 FILLER_135_1968 ();
 FILLCELL_X32 FILLER_135_2000 ();
 FILLCELL_X32 FILLER_135_2032 ();
 FILLCELL_X32 FILLER_135_2064 ();
 FILLCELL_X32 FILLER_135_2096 ();
 FILLCELL_X32 FILLER_135_2128 ();
 FILLCELL_X32 FILLER_135_2160 ();
 FILLCELL_X32 FILLER_135_2192 ();
 FILLCELL_X32 FILLER_135_2224 ();
 FILLCELL_X32 FILLER_135_2256 ();
 FILLCELL_X32 FILLER_135_2288 ();
 FILLCELL_X32 FILLER_135_2320 ();
 FILLCELL_X32 FILLER_135_2352 ();
 FILLCELL_X32 FILLER_135_2384 ();
 FILLCELL_X32 FILLER_135_2416 ();
 FILLCELL_X32 FILLER_135_2448 ();
 FILLCELL_X32 FILLER_135_2480 ();
 FILLCELL_X8 FILLER_135_2512 ();
 FILLCELL_X4 FILLER_135_2520 ();
 FILLCELL_X2 FILLER_135_2524 ();
 FILLCELL_X32 FILLER_135_2527 ();
 FILLCELL_X32 FILLER_135_2559 ();
 FILLCELL_X8 FILLER_135_2591 ();
 FILLCELL_X2 FILLER_135_2599 ();
 FILLCELL_X1 FILLER_135_2601 ();
 FILLCELL_X32 FILLER_136_1 ();
 FILLCELL_X32 FILLER_136_33 ();
 FILLCELL_X32 FILLER_136_65 ();
 FILLCELL_X32 FILLER_136_97 ();
 FILLCELL_X32 FILLER_136_129 ();
 FILLCELL_X32 FILLER_136_161 ();
 FILLCELL_X32 FILLER_136_193 ();
 FILLCELL_X32 FILLER_136_225 ();
 FILLCELL_X32 FILLER_136_257 ();
 FILLCELL_X32 FILLER_136_289 ();
 FILLCELL_X32 FILLER_136_321 ();
 FILLCELL_X32 FILLER_136_353 ();
 FILLCELL_X32 FILLER_136_385 ();
 FILLCELL_X32 FILLER_136_417 ();
 FILLCELL_X32 FILLER_136_449 ();
 FILLCELL_X32 FILLER_136_481 ();
 FILLCELL_X32 FILLER_136_513 ();
 FILLCELL_X32 FILLER_136_545 ();
 FILLCELL_X32 FILLER_136_577 ();
 FILLCELL_X16 FILLER_136_609 ();
 FILLCELL_X4 FILLER_136_625 ();
 FILLCELL_X2 FILLER_136_629 ();
 FILLCELL_X32 FILLER_136_632 ();
 FILLCELL_X32 FILLER_136_664 ();
 FILLCELL_X32 FILLER_136_696 ();
 FILLCELL_X32 FILLER_136_728 ();
 FILLCELL_X32 FILLER_136_760 ();
 FILLCELL_X32 FILLER_136_792 ();
 FILLCELL_X32 FILLER_136_824 ();
 FILLCELL_X32 FILLER_136_856 ();
 FILLCELL_X32 FILLER_136_888 ();
 FILLCELL_X32 FILLER_136_920 ();
 FILLCELL_X32 FILLER_136_952 ();
 FILLCELL_X32 FILLER_136_984 ();
 FILLCELL_X32 FILLER_136_1016 ();
 FILLCELL_X32 FILLER_136_1048 ();
 FILLCELL_X32 FILLER_136_1080 ();
 FILLCELL_X32 FILLER_136_1112 ();
 FILLCELL_X32 FILLER_136_1144 ();
 FILLCELL_X32 FILLER_136_1176 ();
 FILLCELL_X32 FILLER_136_1208 ();
 FILLCELL_X32 FILLER_136_1240 ();
 FILLCELL_X32 FILLER_136_1272 ();
 FILLCELL_X32 FILLER_136_1304 ();
 FILLCELL_X32 FILLER_136_1336 ();
 FILLCELL_X32 FILLER_136_1368 ();
 FILLCELL_X32 FILLER_136_1400 ();
 FILLCELL_X32 FILLER_136_1432 ();
 FILLCELL_X32 FILLER_136_1464 ();
 FILLCELL_X32 FILLER_136_1496 ();
 FILLCELL_X32 FILLER_136_1528 ();
 FILLCELL_X32 FILLER_136_1560 ();
 FILLCELL_X32 FILLER_136_1592 ();
 FILLCELL_X32 FILLER_136_1624 ();
 FILLCELL_X32 FILLER_136_1656 ();
 FILLCELL_X32 FILLER_136_1688 ();
 FILLCELL_X32 FILLER_136_1720 ();
 FILLCELL_X32 FILLER_136_1752 ();
 FILLCELL_X32 FILLER_136_1784 ();
 FILLCELL_X32 FILLER_136_1816 ();
 FILLCELL_X32 FILLER_136_1848 ();
 FILLCELL_X8 FILLER_136_1880 ();
 FILLCELL_X4 FILLER_136_1888 ();
 FILLCELL_X2 FILLER_136_1892 ();
 FILLCELL_X32 FILLER_136_1895 ();
 FILLCELL_X32 FILLER_136_1927 ();
 FILLCELL_X32 FILLER_136_1959 ();
 FILLCELL_X32 FILLER_136_1991 ();
 FILLCELL_X32 FILLER_136_2023 ();
 FILLCELL_X32 FILLER_136_2055 ();
 FILLCELL_X32 FILLER_136_2087 ();
 FILLCELL_X32 FILLER_136_2119 ();
 FILLCELL_X32 FILLER_136_2151 ();
 FILLCELL_X32 FILLER_136_2183 ();
 FILLCELL_X32 FILLER_136_2215 ();
 FILLCELL_X32 FILLER_136_2247 ();
 FILLCELL_X32 FILLER_136_2279 ();
 FILLCELL_X32 FILLER_136_2311 ();
 FILLCELL_X32 FILLER_136_2343 ();
 FILLCELL_X32 FILLER_136_2375 ();
 FILLCELL_X32 FILLER_136_2407 ();
 FILLCELL_X32 FILLER_136_2439 ();
 FILLCELL_X32 FILLER_136_2471 ();
 FILLCELL_X32 FILLER_136_2503 ();
 FILLCELL_X32 FILLER_136_2535 ();
 FILLCELL_X32 FILLER_136_2567 ();
 FILLCELL_X2 FILLER_136_2599 ();
 FILLCELL_X1 FILLER_136_2601 ();
 FILLCELL_X32 FILLER_137_1 ();
 FILLCELL_X32 FILLER_137_33 ();
 FILLCELL_X32 FILLER_137_65 ();
 FILLCELL_X32 FILLER_137_97 ();
 FILLCELL_X32 FILLER_137_129 ();
 FILLCELL_X32 FILLER_137_161 ();
 FILLCELL_X32 FILLER_137_193 ();
 FILLCELL_X32 FILLER_137_225 ();
 FILLCELL_X32 FILLER_137_257 ();
 FILLCELL_X32 FILLER_137_289 ();
 FILLCELL_X32 FILLER_137_321 ();
 FILLCELL_X32 FILLER_137_353 ();
 FILLCELL_X32 FILLER_137_385 ();
 FILLCELL_X32 FILLER_137_417 ();
 FILLCELL_X32 FILLER_137_449 ();
 FILLCELL_X32 FILLER_137_481 ();
 FILLCELL_X32 FILLER_137_513 ();
 FILLCELL_X32 FILLER_137_545 ();
 FILLCELL_X32 FILLER_137_577 ();
 FILLCELL_X32 FILLER_137_609 ();
 FILLCELL_X32 FILLER_137_641 ();
 FILLCELL_X32 FILLER_137_673 ();
 FILLCELL_X32 FILLER_137_705 ();
 FILLCELL_X32 FILLER_137_737 ();
 FILLCELL_X32 FILLER_137_769 ();
 FILLCELL_X32 FILLER_137_801 ();
 FILLCELL_X32 FILLER_137_833 ();
 FILLCELL_X32 FILLER_137_865 ();
 FILLCELL_X32 FILLER_137_897 ();
 FILLCELL_X32 FILLER_137_929 ();
 FILLCELL_X32 FILLER_137_961 ();
 FILLCELL_X32 FILLER_137_993 ();
 FILLCELL_X32 FILLER_137_1025 ();
 FILLCELL_X32 FILLER_137_1057 ();
 FILLCELL_X32 FILLER_137_1089 ();
 FILLCELL_X32 FILLER_137_1121 ();
 FILLCELL_X32 FILLER_137_1153 ();
 FILLCELL_X32 FILLER_137_1185 ();
 FILLCELL_X32 FILLER_137_1217 ();
 FILLCELL_X8 FILLER_137_1249 ();
 FILLCELL_X4 FILLER_137_1257 ();
 FILLCELL_X2 FILLER_137_1261 ();
 FILLCELL_X32 FILLER_137_1264 ();
 FILLCELL_X32 FILLER_137_1296 ();
 FILLCELL_X32 FILLER_137_1328 ();
 FILLCELL_X32 FILLER_137_1360 ();
 FILLCELL_X32 FILLER_137_1392 ();
 FILLCELL_X32 FILLER_137_1424 ();
 FILLCELL_X32 FILLER_137_1456 ();
 FILLCELL_X32 FILLER_137_1488 ();
 FILLCELL_X32 FILLER_137_1520 ();
 FILLCELL_X32 FILLER_137_1552 ();
 FILLCELL_X32 FILLER_137_1584 ();
 FILLCELL_X32 FILLER_137_1616 ();
 FILLCELL_X32 FILLER_137_1648 ();
 FILLCELL_X32 FILLER_137_1680 ();
 FILLCELL_X32 FILLER_137_1712 ();
 FILLCELL_X32 FILLER_137_1744 ();
 FILLCELL_X32 FILLER_137_1776 ();
 FILLCELL_X32 FILLER_137_1808 ();
 FILLCELL_X32 FILLER_137_1840 ();
 FILLCELL_X32 FILLER_137_1872 ();
 FILLCELL_X32 FILLER_137_1904 ();
 FILLCELL_X32 FILLER_137_1936 ();
 FILLCELL_X32 FILLER_137_1968 ();
 FILLCELL_X32 FILLER_137_2000 ();
 FILLCELL_X32 FILLER_137_2032 ();
 FILLCELL_X32 FILLER_137_2064 ();
 FILLCELL_X32 FILLER_137_2096 ();
 FILLCELL_X32 FILLER_137_2128 ();
 FILLCELL_X32 FILLER_137_2160 ();
 FILLCELL_X32 FILLER_137_2192 ();
 FILLCELL_X32 FILLER_137_2224 ();
 FILLCELL_X32 FILLER_137_2256 ();
 FILLCELL_X32 FILLER_137_2288 ();
 FILLCELL_X32 FILLER_137_2320 ();
 FILLCELL_X32 FILLER_137_2352 ();
 FILLCELL_X32 FILLER_137_2384 ();
 FILLCELL_X32 FILLER_137_2416 ();
 FILLCELL_X32 FILLER_137_2448 ();
 FILLCELL_X32 FILLER_137_2480 ();
 FILLCELL_X8 FILLER_137_2512 ();
 FILLCELL_X4 FILLER_137_2520 ();
 FILLCELL_X2 FILLER_137_2524 ();
 FILLCELL_X32 FILLER_137_2527 ();
 FILLCELL_X32 FILLER_137_2559 ();
 FILLCELL_X8 FILLER_137_2591 ();
 FILLCELL_X2 FILLER_137_2599 ();
 FILLCELL_X1 FILLER_137_2601 ();
 FILLCELL_X32 FILLER_138_1 ();
 FILLCELL_X32 FILLER_138_33 ();
 FILLCELL_X32 FILLER_138_65 ();
 FILLCELL_X32 FILLER_138_97 ();
 FILLCELL_X32 FILLER_138_129 ();
 FILLCELL_X32 FILLER_138_161 ();
 FILLCELL_X32 FILLER_138_193 ();
 FILLCELL_X32 FILLER_138_225 ();
 FILLCELL_X32 FILLER_138_257 ();
 FILLCELL_X32 FILLER_138_289 ();
 FILLCELL_X32 FILLER_138_321 ();
 FILLCELL_X32 FILLER_138_353 ();
 FILLCELL_X32 FILLER_138_385 ();
 FILLCELL_X32 FILLER_138_417 ();
 FILLCELL_X32 FILLER_138_449 ();
 FILLCELL_X32 FILLER_138_481 ();
 FILLCELL_X32 FILLER_138_513 ();
 FILLCELL_X32 FILLER_138_545 ();
 FILLCELL_X32 FILLER_138_577 ();
 FILLCELL_X16 FILLER_138_609 ();
 FILLCELL_X4 FILLER_138_625 ();
 FILLCELL_X2 FILLER_138_629 ();
 FILLCELL_X32 FILLER_138_632 ();
 FILLCELL_X32 FILLER_138_664 ();
 FILLCELL_X32 FILLER_138_696 ();
 FILLCELL_X32 FILLER_138_728 ();
 FILLCELL_X32 FILLER_138_760 ();
 FILLCELL_X32 FILLER_138_792 ();
 FILLCELL_X32 FILLER_138_824 ();
 FILLCELL_X32 FILLER_138_856 ();
 FILLCELL_X32 FILLER_138_888 ();
 FILLCELL_X32 FILLER_138_920 ();
 FILLCELL_X32 FILLER_138_952 ();
 FILLCELL_X32 FILLER_138_984 ();
 FILLCELL_X32 FILLER_138_1016 ();
 FILLCELL_X32 FILLER_138_1048 ();
 FILLCELL_X32 FILLER_138_1080 ();
 FILLCELL_X32 FILLER_138_1112 ();
 FILLCELL_X32 FILLER_138_1144 ();
 FILLCELL_X32 FILLER_138_1176 ();
 FILLCELL_X32 FILLER_138_1208 ();
 FILLCELL_X32 FILLER_138_1240 ();
 FILLCELL_X32 FILLER_138_1272 ();
 FILLCELL_X32 FILLER_138_1304 ();
 FILLCELL_X32 FILLER_138_1336 ();
 FILLCELL_X32 FILLER_138_1368 ();
 FILLCELL_X32 FILLER_138_1400 ();
 FILLCELL_X32 FILLER_138_1432 ();
 FILLCELL_X32 FILLER_138_1464 ();
 FILLCELL_X32 FILLER_138_1496 ();
 FILLCELL_X32 FILLER_138_1528 ();
 FILLCELL_X32 FILLER_138_1560 ();
 FILLCELL_X32 FILLER_138_1592 ();
 FILLCELL_X32 FILLER_138_1624 ();
 FILLCELL_X32 FILLER_138_1656 ();
 FILLCELL_X32 FILLER_138_1688 ();
 FILLCELL_X32 FILLER_138_1720 ();
 FILLCELL_X32 FILLER_138_1752 ();
 FILLCELL_X32 FILLER_138_1784 ();
 FILLCELL_X32 FILLER_138_1816 ();
 FILLCELL_X32 FILLER_138_1848 ();
 FILLCELL_X8 FILLER_138_1880 ();
 FILLCELL_X4 FILLER_138_1888 ();
 FILLCELL_X2 FILLER_138_1892 ();
 FILLCELL_X32 FILLER_138_1895 ();
 FILLCELL_X32 FILLER_138_1927 ();
 FILLCELL_X32 FILLER_138_1959 ();
 FILLCELL_X32 FILLER_138_1991 ();
 FILLCELL_X32 FILLER_138_2023 ();
 FILLCELL_X32 FILLER_138_2055 ();
 FILLCELL_X32 FILLER_138_2087 ();
 FILLCELL_X32 FILLER_138_2119 ();
 FILLCELL_X32 FILLER_138_2151 ();
 FILLCELL_X32 FILLER_138_2183 ();
 FILLCELL_X32 FILLER_138_2215 ();
 FILLCELL_X32 FILLER_138_2247 ();
 FILLCELL_X32 FILLER_138_2279 ();
 FILLCELL_X32 FILLER_138_2311 ();
 FILLCELL_X32 FILLER_138_2343 ();
 FILLCELL_X32 FILLER_138_2375 ();
 FILLCELL_X32 FILLER_138_2407 ();
 FILLCELL_X32 FILLER_138_2439 ();
 FILLCELL_X32 FILLER_138_2471 ();
 FILLCELL_X32 FILLER_138_2503 ();
 FILLCELL_X32 FILLER_138_2535 ();
 FILLCELL_X32 FILLER_138_2567 ();
 FILLCELL_X2 FILLER_138_2599 ();
 FILLCELL_X1 FILLER_138_2601 ();
 FILLCELL_X32 FILLER_139_1 ();
 FILLCELL_X32 FILLER_139_33 ();
 FILLCELL_X32 FILLER_139_65 ();
 FILLCELL_X32 FILLER_139_97 ();
 FILLCELL_X32 FILLER_139_129 ();
 FILLCELL_X32 FILLER_139_161 ();
 FILLCELL_X32 FILLER_139_193 ();
 FILLCELL_X32 FILLER_139_225 ();
 FILLCELL_X32 FILLER_139_257 ();
 FILLCELL_X32 FILLER_139_289 ();
 FILLCELL_X32 FILLER_139_321 ();
 FILLCELL_X32 FILLER_139_353 ();
 FILLCELL_X32 FILLER_139_385 ();
 FILLCELL_X32 FILLER_139_417 ();
 FILLCELL_X32 FILLER_139_449 ();
 FILLCELL_X32 FILLER_139_481 ();
 FILLCELL_X32 FILLER_139_513 ();
 FILLCELL_X32 FILLER_139_545 ();
 FILLCELL_X32 FILLER_139_577 ();
 FILLCELL_X32 FILLER_139_609 ();
 FILLCELL_X32 FILLER_139_641 ();
 FILLCELL_X32 FILLER_139_673 ();
 FILLCELL_X32 FILLER_139_705 ();
 FILLCELL_X32 FILLER_139_737 ();
 FILLCELL_X32 FILLER_139_769 ();
 FILLCELL_X32 FILLER_139_801 ();
 FILLCELL_X32 FILLER_139_833 ();
 FILLCELL_X32 FILLER_139_865 ();
 FILLCELL_X32 FILLER_139_897 ();
 FILLCELL_X32 FILLER_139_929 ();
 FILLCELL_X32 FILLER_139_961 ();
 FILLCELL_X32 FILLER_139_993 ();
 FILLCELL_X32 FILLER_139_1025 ();
 FILLCELL_X32 FILLER_139_1057 ();
 FILLCELL_X32 FILLER_139_1089 ();
 FILLCELL_X32 FILLER_139_1121 ();
 FILLCELL_X32 FILLER_139_1153 ();
 FILLCELL_X32 FILLER_139_1185 ();
 FILLCELL_X32 FILLER_139_1217 ();
 FILLCELL_X8 FILLER_139_1249 ();
 FILLCELL_X4 FILLER_139_1257 ();
 FILLCELL_X2 FILLER_139_1261 ();
 FILLCELL_X32 FILLER_139_1264 ();
 FILLCELL_X32 FILLER_139_1296 ();
 FILLCELL_X32 FILLER_139_1328 ();
 FILLCELL_X32 FILLER_139_1360 ();
 FILLCELL_X32 FILLER_139_1392 ();
 FILLCELL_X32 FILLER_139_1424 ();
 FILLCELL_X32 FILLER_139_1456 ();
 FILLCELL_X32 FILLER_139_1488 ();
 FILLCELL_X32 FILLER_139_1520 ();
 FILLCELL_X32 FILLER_139_1552 ();
 FILLCELL_X32 FILLER_139_1584 ();
 FILLCELL_X32 FILLER_139_1616 ();
 FILLCELL_X32 FILLER_139_1648 ();
 FILLCELL_X32 FILLER_139_1680 ();
 FILLCELL_X32 FILLER_139_1712 ();
 FILLCELL_X32 FILLER_139_1744 ();
 FILLCELL_X32 FILLER_139_1776 ();
 FILLCELL_X32 FILLER_139_1808 ();
 FILLCELL_X32 FILLER_139_1840 ();
 FILLCELL_X32 FILLER_139_1872 ();
 FILLCELL_X32 FILLER_139_1904 ();
 FILLCELL_X32 FILLER_139_1936 ();
 FILLCELL_X32 FILLER_139_1968 ();
 FILLCELL_X32 FILLER_139_2000 ();
 FILLCELL_X32 FILLER_139_2032 ();
 FILLCELL_X32 FILLER_139_2064 ();
 FILLCELL_X32 FILLER_139_2096 ();
 FILLCELL_X32 FILLER_139_2128 ();
 FILLCELL_X32 FILLER_139_2160 ();
 FILLCELL_X32 FILLER_139_2192 ();
 FILLCELL_X32 FILLER_139_2224 ();
 FILLCELL_X32 FILLER_139_2256 ();
 FILLCELL_X32 FILLER_139_2288 ();
 FILLCELL_X32 FILLER_139_2320 ();
 FILLCELL_X32 FILLER_139_2352 ();
 FILLCELL_X32 FILLER_139_2384 ();
 FILLCELL_X32 FILLER_139_2416 ();
 FILLCELL_X32 FILLER_139_2448 ();
 FILLCELL_X32 FILLER_139_2480 ();
 FILLCELL_X8 FILLER_139_2512 ();
 FILLCELL_X4 FILLER_139_2520 ();
 FILLCELL_X2 FILLER_139_2524 ();
 FILLCELL_X32 FILLER_139_2527 ();
 FILLCELL_X32 FILLER_139_2559 ();
 FILLCELL_X8 FILLER_139_2591 ();
 FILLCELL_X2 FILLER_139_2599 ();
 FILLCELL_X1 FILLER_139_2601 ();
 FILLCELL_X32 FILLER_140_1 ();
 FILLCELL_X32 FILLER_140_33 ();
 FILLCELL_X32 FILLER_140_65 ();
 FILLCELL_X32 FILLER_140_97 ();
 FILLCELL_X32 FILLER_140_129 ();
 FILLCELL_X32 FILLER_140_161 ();
 FILLCELL_X32 FILLER_140_193 ();
 FILLCELL_X32 FILLER_140_225 ();
 FILLCELL_X32 FILLER_140_257 ();
 FILLCELL_X32 FILLER_140_289 ();
 FILLCELL_X32 FILLER_140_321 ();
 FILLCELL_X32 FILLER_140_353 ();
 FILLCELL_X32 FILLER_140_385 ();
 FILLCELL_X32 FILLER_140_417 ();
 FILLCELL_X32 FILLER_140_449 ();
 FILLCELL_X32 FILLER_140_481 ();
 FILLCELL_X32 FILLER_140_513 ();
 FILLCELL_X32 FILLER_140_545 ();
 FILLCELL_X32 FILLER_140_577 ();
 FILLCELL_X16 FILLER_140_609 ();
 FILLCELL_X4 FILLER_140_625 ();
 FILLCELL_X2 FILLER_140_629 ();
 FILLCELL_X32 FILLER_140_632 ();
 FILLCELL_X32 FILLER_140_664 ();
 FILLCELL_X32 FILLER_140_696 ();
 FILLCELL_X32 FILLER_140_728 ();
 FILLCELL_X32 FILLER_140_760 ();
 FILLCELL_X32 FILLER_140_792 ();
 FILLCELL_X32 FILLER_140_824 ();
 FILLCELL_X32 FILLER_140_856 ();
 FILLCELL_X32 FILLER_140_888 ();
 FILLCELL_X32 FILLER_140_920 ();
 FILLCELL_X32 FILLER_140_952 ();
 FILLCELL_X32 FILLER_140_984 ();
 FILLCELL_X32 FILLER_140_1016 ();
 FILLCELL_X32 FILLER_140_1048 ();
 FILLCELL_X32 FILLER_140_1080 ();
 FILLCELL_X32 FILLER_140_1112 ();
 FILLCELL_X32 FILLER_140_1144 ();
 FILLCELL_X32 FILLER_140_1176 ();
 FILLCELL_X32 FILLER_140_1208 ();
 FILLCELL_X32 FILLER_140_1240 ();
 FILLCELL_X32 FILLER_140_1272 ();
 FILLCELL_X32 FILLER_140_1304 ();
 FILLCELL_X32 FILLER_140_1336 ();
 FILLCELL_X32 FILLER_140_1368 ();
 FILLCELL_X32 FILLER_140_1400 ();
 FILLCELL_X32 FILLER_140_1432 ();
 FILLCELL_X32 FILLER_140_1464 ();
 FILLCELL_X32 FILLER_140_1496 ();
 FILLCELL_X32 FILLER_140_1528 ();
 FILLCELL_X32 FILLER_140_1560 ();
 FILLCELL_X32 FILLER_140_1592 ();
 FILLCELL_X32 FILLER_140_1624 ();
 FILLCELL_X32 FILLER_140_1656 ();
 FILLCELL_X32 FILLER_140_1688 ();
 FILLCELL_X32 FILLER_140_1720 ();
 FILLCELL_X32 FILLER_140_1752 ();
 FILLCELL_X32 FILLER_140_1784 ();
 FILLCELL_X32 FILLER_140_1816 ();
 FILLCELL_X32 FILLER_140_1848 ();
 FILLCELL_X8 FILLER_140_1880 ();
 FILLCELL_X4 FILLER_140_1888 ();
 FILLCELL_X2 FILLER_140_1892 ();
 FILLCELL_X32 FILLER_140_1895 ();
 FILLCELL_X32 FILLER_140_1927 ();
 FILLCELL_X32 FILLER_140_1959 ();
 FILLCELL_X32 FILLER_140_1991 ();
 FILLCELL_X32 FILLER_140_2023 ();
 FILLCELL_X32 FILLER_140_2055 ();
 FILLCELL_X32 FILLER_140_2087 ();
 FILLCELL_X32 FILLER_140_2119 ();
 FILLCELL_X32 FILLER_140_2151 ();
 FILLCELL_X32 FILLER_140_2183 ();
 FILLCELL_X32 FILLER_140_2215 ();
 FILLCELL_X32 FILLER_140_2247 ();
 FILLCELL_X32 FILLER_140_2279 ();
 FILLCELL_X32 FILLER_140_2311 ();
 FILLCELL_X32 FILLER_140_2343 ();
 FILLCELL_X32 FILLER_140_2375 ();
 FILLCELL_X32 FILLER_140_2407 ();
 FILLCELL_X32 FILLER_140_2439 ();
 FILLCELL_X32 FILLER_140_2471 ();
 FILLCELL_X32 FILLER_140_2503 ();
 FILLCELL_X32 FILLER_140_2535 ();
 FILLCELL_X32 FILLER_140_2567 ();
 FILLCELL_X2 FILLER_140_2599 ();
 FILLCELL_X1 FILLER_140_2601 ();
 FILLCELL_X32 FILLER_141_1 ();
 FILLCELL_X32 FILLER_141_33 ();
 FILLCELL_X32 FILLER_141_65 ();
 FILLCELL_X32 FILLER_141_97 ();
 FILLCELL_X32 FILLER_141_129 ();
 FILLCELL_X32 FILLER_141_161 ();
 FILLCELL_X32 FILLER_141_193 ();
 FILLCELL_X32 FILLER_141_225 ();
 FILLCELL_X32 FILLER_141_257 ();
 FILLCELL_X32 FILLER_141_289 ();
 FILLCELL_X32 FILLER_141_321 ();
 FILLCELL_X32 FILLER_141_353 ();
 FILLCELL_X32 FILLER_141_385 ();
 FILLCELL_X32 FILLER_141_417 ();
 FILLCELL_X32 FILLER_141_449 ();
 FILLCELL_X32 FILLER_141_481 ();
 FILLCELL_X32 FILLER_141_513 ();
 FILLCELL_X32 FILLER_141_545 ();
 FILLCELL_X32 FILLER_141_577 ();
 FILLCELL_X32 FILLER_141_609 ();
 FILLCELL_X32 FILLER_141_641 ();
 FILLCELL_X32 FILLER_141_673 ();
 FILLCELL_X32 FILLER_141_705 ();
 FILLCELL_X32 FILLER_141_737 ();
 FILLCELL_X32 FILLER_141_769 ();
 FILLCELL_X32 FILLER_141_801 ();
 FILLCELL_X32 FILLER_141_833 ();
 FILLCELL_X32 FILLER_141_865 ();
 FILLCELL_X32 FILLER_141_897 ();
 FILLCELL_X32 FILLER_141_929 ();
 FILLCELL_X32 FILLER_141_961 ();
 FILLCELL_X32 FILLER_141_993 ();
 FILLCELL_X32 FILLER_141_1025 ();
 FILLCELL_X32 FILLER_141_1057 ();
 FILLCELL_X32 FILLER_141_1089 ();
 FILLCELL_X32 FILLER_141_1121 ();
 FILLCELL_X32 FILLER_141_1153 ();
 FILLCELL_X32 FILLER_141_1185 ();
 FILLCELL_X32 FILLER_141_1217 ();
 FILLCELL_X8 FILLER_141_1249 ();
 FILLCELL_X4 FILLER_141_1257 ();
 FILLCELL_X2 FILLER_141_1261 ();
 FILLCELL_X32 FILLER_141_1264 ();
 FILLCELL_X32 FILLER_141_1296 ();
 FILLCELL_X32 FILLER_141_1328 ();
 FILLCELL_X32 FILLER_141_1360 ();
 FILLCELL_X32 FILLER_141_1392 ();
 FILLCELL_X32 FILLER_141_1424 ();
 FILLCELL_X32 FILLER_141_1456 ();
 FILLCELL_X32 FILLER_141_1488 ();
 FILLCELL_X32 FILLER_141_1520 ();
 FILLCELL_X32 FILLER_141_1552 ();
 FILLCELL_X32 FILLER_141_1584 ();
 FILLCELL_X32 FILLER_141_1616 ();
 FILLCELL_X32 FILLER_141_1648 ();
 FILLCELL_X32 FILLER_141_1680 ();
 FILLCELL_X32 FILLER_141_1712 ();
 FILLCELL_X32 FILLER_141_1744 ();
 FILLCELL_X32 FILLER_141_1776 ();
 FILLCELL_X32 FILLER_141_1808 ();
 FILLCELL_X32 FILLER_141_1840 ();
 FILLCELL_X32 FILLER_141_1872 ();
 FILLCELL_X32 FILLER_141_1904 ();
 FILLCELL_X32 FILLER_141_1936 ();
 FILLCELL_X32 FILLER_141_1968 ();
 FILLCELL_X32 FILLER_141_2000 ();
 FILLCELL_X32 FILLER_141_2032 ();
 FILLCELL_X32 FILLER_141_2064 ();
 FILLCELL_X32 FILLER_141_2096 ();
 FILLCELL_X32 FILLER_141_2128 ();
 FILLCELL_X32 FILLER_141_2160 ();
 FILLCELL_X32 FILLER_141_2192 ();
 FILLCELL_X32 FILLER_141_2224 ();
 FILLCELL_X32 FILLER_141_2256 ();
 FILLCELL_X32 FILLER_141_2288 ();
 FILLCELL_X32 FILLER_141_2320 ();
 FILLCELL_X32 FILLER_141_2352 ();
 FILLCELL_X32 FILLER_141_2384 ();
 FILLCELL_X32 FILLER_141_2416 ();
 FILLCELL_X32 FILLER_141_2448 ();
 FILLCELL_X32 FILLER_141_2480 ();
 FILLCELL_X8 FILLER_141_2512 ();
 FILLCELL_X4 FILLER_141_2520 ();
 FILLCELL_X2 FILLER_141_2524 ();
 FILLCELL_X32 FILLER_141_2527 ();
 FILLCELL_X32 FILLER_141_2559 ();
 FILLCELL_X8 FILLER_141_2591 ();
 FILLCELL_X2 FILLER_141_2599 ();
 FILLCELL_X1 FILLER_141_2601 ();
 FILLCELL_X32 FILLER_142_1 ();
 FILLCELL_X32 FILLER_142_33 ();
 FILLCELL_X32 FILLER_142_65 ();
 FILLCELL_X32 FILLER_142_97 ();
 FILLCELL_X32 FILLER_142_129 ();
 FILLCELL_X32 FILLER_142_161 ();
 FILLCELL_X32 FILLER_142_193 ();
 FILLCELL_X32 FILLER_142_225 ();
 FILLCELL_X32 FILLER_142_257 ();
 FILLCELL_X32 FILLER_142_289 ();
 FILLCELL_X32 FILLER_142_321 ();
 FILLCELL_X32 FILLER_142_353 ();
 FILLCELL_X32 FILLER_142_385 ();
 FILLCELL_X32 FILLER_142_417 ();
 FILLCELL_X32 FILLER_142_449 ();
 FILLCELL_X32 FILLER_142_481 ();
 FILLCELL_X32 FILLER_142_513 ();
 FILLCELL_X32 FILLER_142_545 ();
 FILLCELL_X32 FILLER_142_577 ();
 FILLCELL_X16 FILLER_142_609 ();
 FILLCELL_X4 FILLER_142_625 ();
 FILLCELL_X2 FILLER_142_629 ();
 FILLCELL_X32 FILLER_142_632 ();
 FILLCELL_X32 FILLER_142_664 ();
 FILLCELL_X32 FILLER_142_696 ();
 FILLCELL_X32 FILLER_142_728 ();
 FILLCELL_X32 FILLER_142_760 ();
 FILLCELL_X32 FILLER_142_792 ();
 FILLCELL_X32 FILLER_142_824 ();
 FILLCELL_X32 FILLER_142_856 ();
 FILLCELL_X32 FILLER_142_888 ();
 FILLCELL_X32 FILLER_142_920 ();
 FILLCELL_X32 FILLER_142_952 ();
 FILLCELL_X32 FILLER_142_984 ();
 FILLCELL_X32 FILLER_142_1016 ();
 FILLCELL_X32 FILLER_142_1048 ();
 FILLCELL_X32 FILLER_142_1080 ();
 FILLCELL_X32 FILLER_142_1112 ();
 FILLCELL_X32 FILLER_142_1144 ();
 FILLCELL_X32 FILLER_142_1176 ();
 FILLCELL_X32 FILLER_142_1208 ();
 FILLCELL_X32 FILLER_142_1240 ();
 FILLCELL_X32 FILLER_142_1272 ();
 FILLCELL_X32 FILLER_142_1304 ();
 FILLCELL_X32 FILLER_142_1336 ();
 FILLCELL_X32 FILLER_142_1368 ();
 FILLCELL_X32 FILLER_142_1400 ();
 FILLCELL_X32 FILLER_142_1432 ();
 FILLCELL_X32 FILLER_142_1464 ();
 FILLCELL_X32 FILLER_142_1496 ();
 FILLCELL_X32 FILLER_142_1528 ();
 FILLCELL_X32 FILLER_142_1560 ();
 FILLCELL_X32 FILLER_142_1592 ();
 FILLCELL_X32 FILLER_142_1624 ();
 FILLCELL_X32 FILLER_142_1656 ();
 FILLCELL_X32 FILLER_142_1688 ();
 FILLCELL_X32 FILLER_142_1720 ();
 FILLCELL_X32 FILLER_142_1752 ();
 FILLCELL_X32 FILLER_142_1784 ();
 FILLCELL_X32 FILLER_142_1816 ();
 FILLCELL_X32 FILLER_142_1848 ();
 FILLCELL_X8 FILLER_142_1880 ();
 FILLCELL_X4 FILLER_142_1888 ();
 FILLCELL_X2 FILLER_142_1892 ();
 FILLCELL_X32 FILLER_142_1895 ();
 FILLCELL_X32 FILLER_142_1927 ();
 FILLCELL_X32 FILLER_142_1959 ();
 FILLCELL_X32 FILLER_142_1991 ();
 FILLCELL_X32 FILLER_142_2023 ();
 FILLCELL_X32 FILLER_142_2055 ();
 FILLCELL_X32 FILLER_142_2087 ();
 FILLCELL_X32 FILLER_142_2119 ();
 FILLCELL_X32 FILLER_142_2151 ();
 FILLCELL_X32 FILLER_142_2183 ();
 FILLCELL_X32 FILLER_142_2215 ();
 FILLCELL_X32 FILLER_142_2247 ();
 FILLCELL_X32 FILLER_142_2279 ();
 FILLCELL_X32 FILLER_142_2311 ();
 FILLCELL_X32 FILLER_142_2343 ();
 FILLCELL_X32 FILLER_142_2375 ();
 FILLCELL_X32 FILLER_142_2407 ();
 FILLCELL_X32 FILLER_142_2439 ();
 FILLCELL_X32 FILLER_142_2471 ();
 FILLCELL_X32 FILLER_142_2503 ();
 FILLCELL_X32 FILLER_142_2535 ();
 FILLCELL_X32 FILLER_142_2567 ();
 FILLCELL_X2 FILLER_142_2599 ();
 FILLCELL_X1 FILLER_142_2601 ();
 FILLCELL_X32 FILLER_143_1 ();
 FILLCELL_X32 FILLER_143_33 ();
 FILLCELL_X32 FILLER_143_65 ();
 FILLCELL_X32 FILLER_143_97 ();
 FILLCELL_X32 FILLER_143_129 ();
 FILLCELL_X32 FILLER_143_161 ();
 FILLCELL_X32 FILLER_143_193 ();
 FILLCELL_X32 FILLER_143_225 ();
 FILLCELL_X32 FILLER_143_257 ();
 FILLCELL_X32 FILLER_143_289 ();
 FILLCELL_X32 FILLER_143_321 ();
 FILLCELL_X32 FILLER_143_353 ();
 FILLCELL_X32 FILLER_143_385 ();
 FILLCELL_X32 FILLER_143_417 ();
 FILLCELL_X32 FILLER_143_449 ();
 FILLCELL_X32 FILLER_143_481 ();
 FILLCELL_X32 FILLER_143_513 ();
 FILLCELL_X32 FILLER_143_545 ();
 FILLCELL_X32 FILLER_143_577 ();
 FILLCELL_X32 FILLER_143_609 ();
 FILLCELL_X32 FILLER_143_641 ();
 FILLCELL_X32 FILLER_143_673 ();
 FILLCELL_X32 FILLER_143_705 ();
 FILLCELL_X32 FILLER_143_737 ();
 FILLCELL_X32 FILLER_143_769 ();
 FILLCELL_X32 FILLER_143_801 ();
 FILLCELL_X32 FILLER_143_833 ();
 FILLCELL_X32 FILLER_143_865 ();
 FILLCELL_X32 FILLER_143_897 ();
 FILLCELL_X32 FILLER_143_929 ();
 FILLCELL_X32 FILLER_143_961 ();
 FILLCELL_X32 FILLER_143_993 ();
 FILLCELL_X32 FILLER_143_1025 ();
 FILLCELL_X32 FILLER_143_1057 ();
 FILLCELL_X32 FILLER_143_1089 ();
 FILLCELL_X32 FILLER_143_1121 ();
 FILLCELL_X32 FILLER_143_1153 ();
 FILLCELL_X32 FILLER_143_1185 ();
 FILLCELL_X32 FILLER_143_1217 ();
 FILLCELL_X8 FILLER_143_1249 ();
 FILLCELL_X4 FILLER_143_1257 ();
 FILLCELL_X2 FILLER_143_1261 ();
 FILLCELL_X32 FILLER_143_1264 ();
 FILLCELL_X32 FILLER_143_1296 ();
 FILLCELL_X32 FILLER_143_1328 ();
 FILLCELL_X32 FILLER_143_1360 ();
 FILLCELL_X32 FILLER_143_1392 ();
 FILLCELL_X32 FILLER_143_1424 ();
 FILLCELL_X32 FILLER_143_1456 ();
 FILLCELL_X32 FILLER_143_1488 ();
 FILLCELL_X32 FILLER_143_1520 ();
 FILLCELL_X32 FILLER_143_1552 ();
 FILLCELL_X32 FILLER_143_1584 ();
 FILLCELL_X32 FILLER_143_1616 ();
 FILLCELL_X32 FILLER_143_1648 ();
 FILLCELL_X32 FILLER_143_1680 ();
 FILLCELL_X32 FILLER_143_1712 ();
 FILLCELL_X32 FILLER_143_1744 ();
 FILLCELL_X32 FILLER_143_1776 ();
 FILLCELL_X32 FILLER_143_1808 ();
 FILLCELL_X32 FILLER_143_1840 ();
 FILLCELL_X32 FILLER_143_1872 ();
 FILLCELL_X32 FILLER_143_1904 ();
 FILLCELL_X32 FILLER_143_1936 ();
 FILLCELL_X32 FILLER_143_1968 ();
 FILLCELL_X32 FILLER_143_2000 ();
 FILLCELL_X32 FILLER_143_2032 ();
 FILLCELL_X32 FILLER_143_2064 ();
 FILLCELL_X32 FILLER_143_2096 ();
 FILLCELL_X32 FILLER_143_2128 ();
 FILLCELL_X32 FILLER_143_2160 ();
 FILLCELL_X32 FILLER_143_2192 ();
 FILLCELL_X32 FILLER_143_2224 ();
 FILLCELL_X32 FILLER_143_2256 ();
 FILLCELL_X32 FILLER_143_2288 ();
 FILLCELL_X32 FILLER_143_2320 ();
 FILLCELL_X32 FILLER_143_2352 ();
 FILLCELL_X32 FILLER_143_2384 ();
 FILLCELL_X32 FILLER_143_2416 ();
 FILLCELL_X32 FILLER_143_2448 ();
 FILLCELL_X32 FILLER_143_2480 ();
 FILLCELL_X8 FILLER_143_2512 ();
 FILLCELL_X4 FILLER_143_2520 ();
 FILLCELL_X2 FILLER_143_2524 ();
 FILLCELL_X32 FILLER_143_2527 ();
 FILLCELL_X32 FILLER_143_2559 ();
 FILLCELL_X8 FILLER_143_2591 ();
 FILLCELL_X2 FILLER_143_2599 ();
 FILLCELL_X1 FILLER_143_2601 ();
 FILLCELL_X32 FILLER_144_1 ();
 FILLCELL_X32 FILLER_144_33 ();
 FILLCELL_X32 FILLER_144_65 ();
 FILLCELL_X32 FILLER_144_97 ();
 FILLCELL_X32 FILLER_144_129 ();
 FILLCELL_X32 FILLER_144_161 ();
 FILLCELL_X32 FILLER_144_193 ();
 FILLCELL_X32 FILLER_144_225 ();
 FILLCELL_X32 FILLER_144_257 ();
 FILLCELL_X32 FILLER_144_289 ();
 FILLCELL_X32 FILLER_144_321 ();
 FILLCELL_X32 FILLER_144_353 ();
 FILLCELL_X32 FILLER_144_385 ();
 FILLCELL_X32 FILLER_144_417 ();
 FILLCELL_X32 FILLER_144_449 ();
 FILLCELL_X32 FILLER_144_481 ();
 FILLCELL_X32 FILLER_144_513 ();
 FILLCELL_X32 FILLER_144_545 ();
 FILLCELL_X32 FILLER_144_577 ();
 FILLCELL_X16 FILLER_144_609 ();
 FILLCELL_X4 FILLER_144_625 ();
 FILLCELL_X2 FILLER_144_629 ();
 FILLCELL_X32 FILLER_144_632 ();
 FILLCELL_X32 FILLER_144_664 ();
 FILLCELL_X32 FILLER_144_696 ();
 FILLCELL_X32 FILLER_144_728 ();
 FILLCELL_X32 FILLER_144_760 ();
 FILLCELL_X32 FILLER_144_792 ();
 FILLCELL_X32 FILLER_144_824 ();
 FILLCELL_X32 FILLER_144_856 ();
 FILLCELL_X32 FILLER_144_888 ();
 FILLCELL_X32 FILLER_144_920 ();
 FILLCELL_X32 FILLER_144_952 ();
 FILLCELL_X32 FILLER_144_984 ();
 FILLCELL_X32 FILLER_144_1016 ();
 FILLCELL_X32 FILLER_144_1048 ();
 FILLCELL_X32 FILLER_144_1080 ();
 FILLCELL_X32 FILLER_144_1112 ();
 FILLCELL_X32 FILLER_144_1144 ();
 FILLCELL_X32 FILLER_144_1176 ();
 FILLCELL_X32 FILLER_144_1208 ();
 FILLCELL_X32 FILLER_144_1240 ();
 FILLCELL_X32 FILLER_144_1272 ();
 FILLCELL_X32 FILLER_144_1304 ();
 FILLCELL_X32 FILLER_144_1336 ();
 FILLCELL_X32 FILLER_144_1368 ();
 FILLCELL_X32 FILLER_144_1400 ();
 FILLCELL_X32 FILLER_144_1432 ();
 FILLCELL_X32 FILLER_144_1464 ();
 FILLCELL_X32 FILLER_144_1496 ();
 FILLCELL_X32 FILLER_144_1528 ();
 FILLCELL_X32 FILLER_144_1560 ();
 FILLCELL_X32 FILLER_144_1592 ();
 FILLCELL_X32 FILLER_144_1624 ();
 FILLCELL_X32 FILLER_144_1656 ();
 FILLCELL_X32 FILLER_144_1688 ();
 FILLCELL_X32 FILLER_144_1720 ();
 FILLCELL_X32 FILLER_144_1752 ();
 FILLCELL_X32 FILLER_144_1784 ();
 FILLCELL_X32 FILLER_144_1816 ();
 FILLCELL_X32 FILLER_144_1848 ();
 FILLCELL_X8 FILLER_144_1880 ();
 FILLCELL_X4 FILLER_144_1888 ();
 FILLCELL_X2 FILLER_144_1892 ();
 FILLCELL_X32 FILLER_144_1895 ();
 FILLCELL_X32 FILLER_144_1927 ();
 FILLCELL_X32 FILLER_144_1959 ();
 FILLCELL_X32 FILLER_144_1991 ();
 FILLCELL_X32 FILLER_144_2023 ();
 FILLCELL_X32 FILLER_144_2055 ();
 FILLCELL_X32 FILLER_144_2087 ();
 FILLCELL_X32 FILLER_144_2119 ();
 FILLCELL_X32 FILLER_144_2151 ();
 FILLCELL_X32 FILLER_144_2183 ();
 FILLCELL_X32 FILLER_144_2215 ();
 FILLCELL_X32 FILLER_144_2247 ();
 FILLCELL_X32 FILLER_144_2279 ();
 FILLCELL_X32 FILLER_144_2311 ();
 FILLCELL_X32 FILLER_144_2343 ();
 FILLCELL_X32 FILLER_144_2375 ();
 FILLCELL_X32 FILLER_144_2407 ();
 FILLCELL_X32 FILLER_144_2439 ();
 FILLCELL_X32 FILLER_144_2471 ();
 FILLCELL_X32 FILLER_144_2503 ();
 FILLCELL_X32 FILLER_144_2535 ();
 FILLCELL_X32 FILLER_144_2567 ();
 FILLCELL_X2 FILLER_144_2599 ();
 FILLCELL_X1 FILLER_144_2601 ();
 FILLCELL_X32 FILLER_145_1 ();
 FILLCELL_X32 FILLER_145_33 ();
 FILLCELL_X32 FILLER_145_65 ();
 FILLCELL_X32 FILLER_145_97 ();
 FILLCELL_X32 FILLER_145_129 ();
 FILLCELL_X32 FILLER_145_161 ();
 FILLCELL_X32 FILLER_145_193 ();
 FILLCELL_X32 FILLER_145_225 ();
 FILLCELL_X32 FILLER_145_257 ();
 FILLCELL_X32 FILLER_145_289 ();
 FILLCELL_X32 FILLER_145_321 ();
 FILLCELL_X32 FILLER_145_353 ();
 FILLCELL_X32 FILLER_145_385 ();
 FILLCELL_X32 FILLER_145_417 ();
 FILLCELL_X32 FILLER_145_449 ();
 FILLCELL_X32 FILLER_145_481 ();
 FILLCELL_X32 FILLER_145_513 ();
 FILLCELL_X32 FILLER_145_545 ();
 FILLCELL_X32 FILLER_145_577 ();
 FILLCELL_X32 FILLER_145_609 ();
 FILLCELL_X32 FILLER_145_641 ();
 FILLCELL_X32 FILLER_145_673 ();
 FILLCELL_X32 FILLER_145_705 ();
 FILLCELL_X32 FILLER_145_737 ();
 FILLCELL_X32 FILLER_145_769 ();
 FILLCELL_X32 FILLER_145_801 ();
 FILLCELL_X32 FILLER_145_833 ();
 FILLCELL_X32 FILLER_145_865 ();
 FILLCELL_X32 FILLER_145_897 ();
 FILLCELL_X32 FILLER_145_929 ();
 FILLCELL_X32 FILLER_145_961 ();
 FILLCELL_X32 FILLER_145_993 ();
 FILLCELL_X32 FILLER_145_1025 ();
 FILLCELL_X32 FILLER_145_1057 ();
 FILLCELL_X32 FILLER_145_1089 ();
 FILLCELL_X32 FILLER_145_1121 ();
 FILLCELL_X32 FILLER_145_1153 ();
 FILLCELL_X32 FILLER_145_1185 ();
 FILLCELL_X32 FILLER_145_1217 ();
 FILLCELL_X8 FILLER_145_1249 ();
 FILLCELL_X4 FILLER_145_1257 ();
 FILLCELL_X2 FILLER_145_1261 ();
 FILLCELL_X32 FILLER_145_1264 ();
 FILLCELL_X32 FILLER_145_1296 ();
 FILLCELL_X32 FILLER_145_1328 ();
 FILLCELL_X32 FILLER_145_1360 ();
 FILLCELL_X32 FILLER_145_1392 ();
 FILLCELL_X32 FILLER_145_1424 ();
 FILLCELL_X32 FILLER_145_1456 ();
 FILLCELL_X32 FILLER_145_1488 ();
 FILLCELL_X32 FILLER_145_1520 ();
 FILLCELL_X32 FILLER_145_1552 ();
 FILLCELL_X32 FILLER_145_1584 ();
 FILLCELL_X32 FILLER_145_1616 ();
 FILLCELL_X32 FILLER_145_1648 ();
 FILLCELL_X32 FILLER_145_1680 ();
 FILLCELL_X32 FILLER_145_1712 ();
 FILLCELL_X32 FILLER_145_1744 ();
 FILLCELL_X32 FILLER_145_1776 ();
 FILLCELL_X32 FILLER_145_1808 ();
 FILLCELL_X32 FILLER_145_1840 ();
 FILLCELL_X32 FILLER_145_1872 ();
 FILLCELL_X32 FILLER_145_1904 ();
 FILLCELL_X32 FILLER_145_1936 ();
 FILLCELL_X32 FILLER_145_1968 ();
 FILLCELL_X32 FILLER_145_2000 ();
 FILLCELL_X32 FILLER_145_2032 ();
 FILLCELL_X32 FILLER_145_2064 ();
 FILLCELL_X32 FILLER_145_2096 ();
 FILLCELL_X32 FILLER_145_2128 ();
 FILLCELL_X32 FILLER_145_2160 ();
 FILLCELL_X32 FILLER_145_2192 ();
 FILLCELL_X32 FILLER_145_2224 ();
 FILLCELL_X32 FILLER_145_2256 ();
 FILLCELL_X32 FILLER_145_2288 ();
 FILLCELL_X32 FILLER_145_2320 ();
 FILLCELL_X32 FILLER_145_2352 ();
 FILLCELL_X32 FILLER_145_2384 ();
 FILLCELL_X32 FILLER_145_2416 ();
 FILLCELL_X32 FILLER_145_2448 ();
 FILLCELL_X32 FILLER_145_2480 ();
 FILLCELL_X8 FILLER_145_2512 ();
 FILLCELL_X4 FILLER_145_2520 ();
 FILLCELL_X2 FILLER_145_2524 ();
 FILLCELL_X32 FILLER_145_2527 ();
 FILLCELL_X32 FILLER_145_2559 ();
 FILLCELL_X8 FILLER_145_2591 ();
 FILLCELL_X2 FILLER_145_2599 ();
 FILLCELL_X1 FILLER_145_2601 ();
 FILLCELL_X32 FILLER_146_1 ();
 FILLCELL_X32 FILLER_146_33 ();
 FILLCELL_X32 FILLER_146_65 ();
 FILLCELL_X32 FILLER_146_97 ();
 FILLCELL_X32 FILLER_146_129 ();
 FILLCELL_X32 FILLER_146_161 ();
 FILLCELL_X32 FILLER_146_193 ();
 FILLCELL_X32 FILLER_146_225 ();
 FILLCELL_X32 FILLER_146_257 ();
 FILLCELL_X32 FILLER_146_289 ();
 FILLCELL_X32 FILLER_146_321 ();
 FILLCELL_X32 FILLER_146_353 ();
 FILLCELL_X32 FILLER_146_385 ();
 FILLCELL_X32 FILLER_146_417 ();
 FILLCELL_X32 FILLER_146_449 ();
 FILLCELL_X32 FILLER_146_481 ();
 FILLCELL_X32 FILLER_146_513 ();
 FILLCELL_X32 FILLER_146_545 ();
 FILLCELL_X32 FILLER_146_577 ();
 FILLCELL_X16 FILLER_146_609 ();
 FILLCELL_X4 FILLER_146_625 ();
 FILLCELL_X2 FILLER_146_629 ();
 FILLCELL_X32 FILLER_146_632 ();
 FILLCELL_X32 FILLER_146_664 ();
 FILLCELL_X32 FILLER_146_696 ();
 FILLCELL_X32 FILLER_146_728 ();
 FILLCELL_X32 FILLER_146_760 ();
 FILLCELL_X32 FILLER_146_792 ();
 FILLCELL_X32 FILLER_146_824 ();
 FILLCELL_X32 FILLER_146_856 ();
 FILLCELL_X32 FILLER_146_888 ();
 FILLCELL_X32 FILLER_146_920 ();
 FILLCELL_X32 FILLER_146_952 ();
 FILLCELL_X32 FILLER_146_984 ();
 FILLCELL_X32 FILLER_146_1016 ();
 FILLCELL_X32 FILLER_146_1048 ();
 FILLCELL_X32 FILLER_146_1080 ();
 FILLCELL_X32 FILLER_146_1112 ();
 FILLCELL_X32 FILLER_146_1144 ();
 FILLCELL_X32 FILLER_146_1176 ();
 FILLCELL_X32 FILLER_146_1208 ();
 FILLCELL_X32 FILLER_146_1240 ();
 FILLCELL_X32 FILLER_146_1272 ();
 FILLCELL_X32 FILLER_146_1304 ();
 FILLCELL_X32 FILLER_146_1336 ();
 FILLCELL_X32 FILLER_146_1368 ();
 FILLCELL_X32 FILLER_146_1400 ();
 FILLCELL_X32 FILLER_146_1432 ();
 FILLCELL_X32 FILLER_146_1464 ();
 FILLCELL_X32 FILLER_146_1496 ();
 FILLCELL_X32 FILLER_146_1528 ();
 FILLCELL_X32 FILLER_146_1560 ();
 FILLCELL_X32 FILLER_146_1592 ();
 FILLCELL_X32 FILLER_146_1624 ();
 FILLCELL_X32 FILLER_146_1656 ();
 FILLCELL_X32 FILLER_146_1688 ();
 FILLCELL_X32 FILLER_146_1720 ();
 FILLCELL_X32 FILLER_146_1752 ();
 FILLCELL_X32 FILLER_146_1784 ();
 FILLCELL_X32 FILLER_146_1816 ();
 FILLCELL_X32 FILLER_146_1848 ();
 FILLCELL_X8 FILLER_146_1880 ();
 FILLCELL_X4 FILLER_146_1888 ();
 FILLCELL_X2 FILLER_146_1892 ();
 FILLCELL_X32 FILLER_146_1895 ();
 FILLCELL_X32 FILLER_146_1927 ();
 FILLCELL_X32 FILLER_146_1959 ();
 FILLCELL_X32 FILLER_146_1991 ();
 FILLCELL_X32 FILLER_146_2023 ();
 FILLCELL_X32 FILLER_146_2055 ();
 FILLCELL_X32 FILLER_146_2087 ();
 FILLCELL_X32 FILLER_146_2119 ();
 FILLCELL_X32 FILLER_146_2151 ();
 FILLCELL_X32 FILLER_146_2183 ();
 FILLCELL_X32 FILLER_146_2215 ();
 FILLCELL_X32 FILLER_146_2247 ();
 FILLCELL_X32 FILLER_146_2279 ();
 FILLCELL_X32 FILLER_146_2311 ();
 FILLCELL_X32 FILLER_146_2343 ();
 FILLCELL_X32 FILLER_146_2375 ();
 FILLCELL_X32 FILLER_146_2407 ();
 FILLCELL_X32 FILLER_146_2439 ();
 FILLCELL_X32 FILLER_146_2471 ();
 FILLCELL_X32 FILLER_146_2503 ();
 FILLCELL_X32 FILLER_146_2535 ();
 FILLCELL_X32 FILLER_146_2567 ();
 FILLCELL_X2 FILLER_146_2599 ();
 FILLCELL_X1 FILLER_146_2601 ();
 FILLCELL_X32 FILLER_147_1 ();
 FILLCELL_X32 FILLER_147_33 ();
 FILLCELL_X32 FILLER_147_65 ();
 FILLCELL_X32 FILLER_147_97 ();
 FILLCELL_X32 FILLER_147_129 ();
 FILLCELL_X32 FILLER_147_161 ();
 FILLCELL_X32 FILLER_147_193 ();
 FILLCELL_X32 FILLER_147_225 ();
 FILLCELL_X32 FILLER_147_257 ();
 FILLCELL_X32 FILLER_147_289 ();
 FILLCELL_X32 FILLER_147_321 ();
 FILLCELL_X32 FILLER_147_353 ();
 FILLCELL_X32 FILLER_147_385 ();
 FILLCELL_X32 FILLER_147_417 ();
 FILLCELL_X32 FILLER_147_449 ();
 FILLCELL_X32 FILLER_147_481 ();
 FILLCELL_X32 FILLER_147_513 ();
 FILLCELL_X32 FILLER_147_545 ();
 FILLCELL_X32 FILLER_147_577 ();
 FILLCELL_X32 FILLER_147_609 ();
 FILLCELL_X32 FILLER_147_641 ();
 FILLCELL_X32 FILLER_147_673 ();
 FILLCELL_X32 FILLER_147_705 ();
 FILLCELL_X32 FILLER_147_737 ();
 FILLCELL_X32 FILLER_147_769 ();
 FILLCELL_X32 FILLER_147_801 ();
 FILLCELL_X32 FILLER_147_833 ();
 FILLCELL_X32 FILLER_147_865 ();
 FILLCELL_X32 FILLER_147_897 ();
 FILLCELL_X32 FILLER_147_929 ();
 FILLCELL_X32 FILLER_147_961 ();
 FILLCELL_X32 FILLER_147_993 ();
 FILLCELL_X32 FILLER_147_1025 ();
 FILLCELL_X32 FILLER_147_1057 ();
 FILLCELL_X32 FILLER_147_1089 ();
 FILLCELL_X32 FILLER_147_1121 ();
 FILLCELL_X32 FILLER_147_1153 ();
 FILLCELL_X32 FILLER_147_1185 ();
 FILLCELL_X32 FILLER_147_1217 ();
 FILLCELL_X8 FILLER_147_1249 ();
 FILLCELL_X4 FILLER_147_1257 ();
 FILLCELL_X2 FILLER_147_1261 ();
 FILLCELL_X32 FILLER_147_1264 ();
 FILLCELL_X32 FILLER_147_1296 ();
 FILLCELL_X32 FILLER_147_1328 ();
 FILLCELL_X32 FILLER_147_1360 ();
 FILLCELL_X32 FILLER_147_1392 ();
 FILLCELL_X32 FILLER_147_1424 ();
 FILLCELL_X32 FILLER_147_1456 ();
 FILLCELL_X32 FILLER_147_1488 ();
 FILLCELL_X32 FILLER_147_1520 ();
 FILLCELL_X32 FILLER_147_1552 ();
 FILLCELL_X32 FILLER_147_1584 ();
 FILLCELL_X32 FILLER_147_1616 ();
 FILLCELL_X32 FILLER_147_1648 ();
 FILLCELL_X32 FILLER_147_1680 ();
 FILLCELL_X32 FILLER_147_1712 ();
 FILLCELL_X32 FILLER_147_1744 ();
 FILLCELL_X32 FILLER_147_1776 ();
 FILLCELL_X32 FILLER_147_1808 ();
 FILLCELL_X32 FILLER_147_1840 ();
 FILLCELL_X32 FILLER_147_1872 ();
 FILLCELL_X32 FILLER_147_1904 ();
 FILLCELL_X32 FILLER_147_1936 ();
 FILLCELL_X32 FILLER_147_1968 ();
 FILLCELL_X32 FILLER_147_2000 ();
 FILLCELL_X32 FILLER_147_2032 ();
 FILLCELL_X32 FILLER_147_2064 ();
 FILLCELL_X32 FILLER_147_2096 ();
 FILLCELL_X32 FILLER_147_2128 ();
 FILLCELL_X32 FILLER_147_2160 ();
 FILLCELL_X32 FILLER_147_2192 ();
 FILLCELL_X32 FILLER_147_2224 ();
 FILLCELL_X32 FILLER_147_2256 ();
 FILLCELL_X32 FILLER_147_2288 ();
 FILLCELL_X32 FILLER_147_2320 ();
 FILLCELL_X32 FILLER_147_2352 ();
 FILLCELL_X32 FILLER_147_2384 ();
 FILLCELL_X32 FILLER_147_2416 ();
 FILLCELL_X32 FILLER_147_2448 ();
 FILLCELL_X32 FILLER_147_2480 ();
 FILLCELL_X8 FILLER_147_2512 ();
 FILLCELL_X4 FILLER_147_2520 ();
 FILLCELL_X2 FILLER_147_2524 ();
 FILLCELL_X32 FILLER_147_2527 ();
 FILLCELL_X32 FILLER_147_2559 ();
 FILLCELL_X8 FILLER_147_2591 ();
 FILLCELL_X2 FILLER_147_2599 ();
 FILLCELL_X1 FILLER_147_2601 ();
 FILLCELL_X32 FILLER_148_1 ();
 FILLCELL_X32 FILLER_148_33 ();
 FILLCELL_X32 FILLER_148_65 ();
 FILLCELL_X32 FILLER_148_97 ();
 FILLCELL_X32 FILLER_148_129 ();
 FILLCELL_X32 FILLER_148_161 ();
 FILLCELL_X32 FILLER_148_193 ();
 FILLCELL_X32 FILLER_148_225 ();
 FILLCELL_X32 FILLER_148_257 ();
 FILLCELL_X32 FILLER_148_289 ();
 FILLCELL_X32 FILLER_148_321 ();
 FILLCELL_X32 FILLER_148_353 ();
 FILLCELL_X32 FILLER_148_385 ();
 FILLCELL_X32 FILLER_148_417 ();
 FILLCELL_X32 FILLER_148_449 ();
 FILLCELL_X32 FILLER_148_481 ();
 FILLCELL_X32 FILLER_148_513 ();
 FILLCELL_X32 FILLER_148_545 ();
 FILLCELL_X32 FILLER_148_577 ();
 FILLCELL_X16 FILLER_148_609 ();
 FILLCELL_X4 FILLER_148_625 ();
 FILLCELL_X2 FILLER_148_629 ();
 FILLCELL_X32 FILLER_148_632 ();
 FILLCELL_X32 FILLER_148_664 ();
 FILLCELL_X32 FILLER_148_696 ();
 FILLCELL_X32 FILLER_148_728 ();
 FILLCELL_X32 FILLER_148_760 ();
 FILLCELL_X32 FILLER_148_792 ();
 FILLCELL_X32 FILLER_148_824 ();
 FILLCELL_X32 FILLER_148_856 ();
 FILLCELL_X32 FILLER_148_888 ();
 FILLCELL_X32 FILLER_148_920 ();
 FILLCELL_X32 FILLER_148_952 ();
 FILLCELL_X32 FILLER_148_984 ();
 FILLCELL_X32 FILLER_148_1016 ();
 FILLCELL_X32 FILLER_148_1048 ();
 FILLCELL_X32 FILLER_148_1080 ();
 FILLCELL_X32 FILLER_148_1112 ();
 FILLCELL_X32 FILLER_148_1144 ();
 FILLCELL_X32 FILLER_148_1176 ();
 FILLCELL_X32 FILLER_148_1208 ();
 FILLCELL_X32 FILLER_148_1240 ();
 FILLCELL_X32 FILLER_148_1272 ();
 FILLCELL_X32 FILLER_148_1304 ();
 FILLCELL_X32 FILLER_148_1336 ();
 FILLCELL_X32 FILLER_148_1368 ();
 FILLCELL_X32 FILLER_148_1400 ();
 FILLCELL_X32 FILLER_148_1432 ();
 FILLCELL_X32 FILLER_148_1464 ();
 FILLCELL_X32 FILLER_148_1496 ();
 FILLCELL_X32 FILLER_148_1528 ();
 FILLCELL_X32 FILLER_148_1560 ();
 FILLCELL_X32 FILLER_148_1592 ();
 FILLCELL_X32 FILLER_148_1624 ();
 FILLCELL_X32 FILLER_148_1656 ();
 FILLCELL_X32 FILLER_148_1688 ();
 FILLCELL_X32 FILLER_148_1720 ();
 FILLCELL_X32 FILLER_148_1752 ();
 FILLCELL_X32 FILLER_148_1784 ();
 FILLCELL_X32 FILLER_148_1816 ();
 FILLCELL_X32 FILLER_148_1848 ();
 FILLCELL_X8 FILLER_148_1880 ();
 FILLCELL_X4 FILLER_148_1888 ();
 FILLCELL_X2 FILLER_148_1892 ();
 FILLCELL_X32 FILLER_148_1895 ();
 FILLCELL_X32 FILLER_148_1927 ();
 FILLCELL_X32 FILLER_148_1959 ();
 FILLCELL_X32 FILLER_148_1991 ();
 FILLCELL_X32 FILLER_148_2023 ();
 FILLCELL_X32 FILLER_148_2055 ();
 FILLCELL_X32 FILLER_148_2087 ();
 FILLCELL_X32 FILLER_148_2119 ();
 FILLCELL_X32 FILLER_148_2151 ();
 FILLCELL_X32 FILLER_148_2183 ();
 FILLCELL_X32 FILLER_148_2215 ();
 FILLCELL_X32 FILLER_148_2247 ();
 FILLCELL_X32 FILLER_148_2279 ();
 FILLCELL_X32 FILLER_148_2311 ();
 FILLCELL_X32 FILLER_148_2343 ();
 FILLCELL_X32 FILLER_148_2375 ();
 FILLCELL_X32 FILLER_148_2407 ();
 FILLCELL_X32 FILLER_148_2439 ();
 FILLCELL_X32 FILLER_148_2471 ();
 FILLCELL_X32 FILLER_148_2503 ();
 FILLCELL_X32 FILLER_148_2535 ();
 FILLCELL_X32 FILLER_148_2567 ();
 FILLCELL_X2 FILLER_148_2599 ();
 FILLCELL_X1 FILLER_148_2601 ();
 FILLCELL_X32 FILLER_149_1 ();
 FILLCELL_X32 FILLER_149_33 ();
 FILLCELL_X32 FILLER_149_65 ();
 FILLCELL_X32 FILLER_149_97 ();
 FILLCELL_X32 FILLER_149_129 ();
 FILLCELL_X32 FILLER_149_161 ();
 FILLCELL_X32 FILLER_149_193 ();
 FILLCELL_X32 FILLER_149_225 ();
 FILLCELL_X32 FILLER_149_257 ();
 FILLCELL_X32 FILLER_149_289 ();
 FILLCELL_X32 FILLER_149_321 ();
 FILLCELL_X32 FILLER_149_353 ();
 FILLCELL_X32 FILLER_149_385 ();
 FILLCELL_X32 FILLER_149_417 ();
 FILLCELL_X32 FILLER_149_449 ();
 FILLCELL_X32 FILLER_149_481 ();
 FILLCELL_X32 FILLER_149_513 ();
 FILLCELL_X32 FILLER_149_545 ();
 FILLCELL_X32 FILLER_149_577 ();
 FILLCELL_X32 FILLER_149_609 ();
 FILLCELL_X32 FILLER_149_641 ();
 FILLCELL_X32 FILLER_149_673 ();
 FILLCELL_X32 FILLER_149_705 ();
 FILLCELL_X32 FILLER_149_737 ();
 FILLCELL_X32 FILLER_149_769 ();
 FILLCELL_X32 FILLER_149_801 ();
 FILLCELL_X32 FILLER_149_833 ();
 FILLCELL_X32 FILLER_149_865 ();
 FILLCELL_X32 FILLER_149_897 ();
 FILLCELL_X32 FILLER_149_929 ();
 FILLCELL_X32 FILLER_149_961 ();
 FILLCELL_X32 FILLER_149_993 ();
 FILLCELL_X32 FILLER_149_1025 ();
 FILLCELL_X32 FILLER_149_1057 ();
 FILLCELL_X32 FILLER_149_1089 ();
 FILLCELL_X32 FILLER_149_1121 ();
 FILLCELL_X32 FILLER_149_1153 ();
 FILLCELL_X32 FILLER_149_1185 ();
 FILLCELL_X32 FILLER_149_1217 ();
 FILLCELL_X8 FILLER_149_1249 ();
 FILLCELL_X4 FILLER_149_1257 ();
 FILLCELL_X2 FILLER_149_1261 ();
 FILLCELL_X32 FILLER_149_1264 ();
 FILLCELL_X32 FILLER_149_1296 ();
 FILLCELL_X32 FILLER_149_1328 ();
 FILLCELL_X32 FILLER_149_1360 ();
 FILLCELL_X32 FILLER_149_1392 ();
 FILLCELL_X32 FILLER_149_1424 ();
 FILLCELL_X32 FILLER_149_1456 ();
 FILLCELL_X32 FILLER_149_1488 ();
 FILLCELL_X32 FILLER_149_1520 ();
 FILLCELL_X32 FILLER_149_1552 ();
 FILLCELL_X32 FILLER_149_1584 ();
 FILLCELL_X32 FILLER_149_1616 ();
 FILLCELL_X32 FILLER_149_1648 ();
 FILLCELL_X32 FILLER_149_1680 ();
 FILLCELL_X32 FILLER_149_1712 ();
 FILLCELL_X32 FILLER_149_1744 ();
 FILLCELL_X32 FILLER_149_1776 ();
 FILLCELL_X32 FILLER_149_1808 ();
 FILLCELL_X32 FILLER_149_1840 ();
 FILLCELL_X32 FILLER_149_1872 ();
 FILLCELL_X32 FILLER_149_1904 ();
 FILLCELL_X32 FILLER_149_1936 ();
 FILLCELL_X32 FILLER_149_1968 ();
 FILLCELL_X32 FILLER_149_2000 ();
 FILLCELL_X32 FILLER_149_2032 ();
 FILLCELL_X32 FILLER_149_2064 ();
 FILLCELL_X32 FILLER_149_2096 ();
 FILLCELL_X32 FILLER_149_2128 ();
 FILLCELL_X32 FILLER_149_2160 ();
 FILLCELL_X32 FILLER_149_2192 ();
 FILLCELL_X32 FILLER_149_2224 ();
 FILLCELL_X32 FILLER_149_2256 ();
 FILLCELL_X32 FILLER_149_2288 ();
 FILLCELL_X32 FILLER_149_2320 ();
 FILLCELL_X32 FILLER_149_2352 ();
 FILLCELL_X32 FILLER_149_2384 ();
 FILLCELL_X32 FILLER_149_2416 ();
 FILLCELL_X32 FILLER_149_2448 ();
 FILLCELL_X32 FILLER_149_2480 ();
 FILLCELL_X8 FILLER_149_2512 ();
 FILLCELL_X4 FILLER_149_2520 ();
 FILLCELL_X2 FILLER_149_2524 ();
 FILLCELL_X32 FILLER_149_2527 ();
 FILLCELL_X32 FILLER_149_2559 ();
 FILLCELL_X8 FILLER_149_2591 ();
 FILLCELL_X2 FILLER_149_2599 ();
 FILLCELL_X1 FILLER_149_2601 ();
 FILLCELL_X32 FILLER_150_1 ();
 FILLCELL_X32 FILLER_150_33 ();
 FILLCELL_X32 FILLER_150_65 ();
 FILLCELL_X32 FILLER_150_97 ();
 FILLCELL_X32 FILLER_150_129 ();
 FILLCELL_X32 FILLER_150_161 ();
 FILLCELL_X32 FILLER_150_193 ();
 FILLCELL_X32 FILLER_150_225 ();
 FILLCELL_X32 FILLER_150_257 ();
 FILLCELL_X32 FILLER_150_289 ();
 FILLCELL_X32 FILLER_150_321 ();
 FILLCELL_X32 FILLER_150_353 ();
 FILLCELL_X32 FILLER_150_385 ();
 FILLCELL_X32 FILLER_150_417 ();
 FILLCELL_X32 FILLER_150_449 ();
 FILLCELL_X32 FILLER_150_481 ();
 FILLCELL_X32 FILLER_150_513 ();
 FILLCELL_X32 FILLER_150_545 ();
 FILLCELL_X32 FILLER_150_577 ();
 FILLCELL_X16 FILLER_150_609 ();
 FILLCELL_X4 FILLER_150_625 ();
 FILLCELL_X2 FILLER_150_629 ();
 FILLCELL_X32 FILLER_150_632 ();
 FILLCELL_X32 FILLER_150_664 ();
 FILLCELL_X32 FILLER_150_696 ();
 FILLCELL_X32 FILLER_150_728 ();
 FILLCELL_X32 FILLER_150_760 ();
 FILLCELL_X32 FILLER_150_792 ();
 FILLCELL_X32 FILLER_150_824 ();
 FILLCELL_X32 FILLER_150_856 ();
 FILLCELL_X32 FILLER_150_888 ();
 FILLCELL_X32 FILLER_150_920 ();
 FILLCELL_X32 FILLER_150_952 ();
 FILLCELL_X32 FILLER_150_984 ();
 FILLCELL_X32 FILLER_150_1016 ();
 FILLCELL_X32 FILLER_150_1048 ();
 FILLCELL_X32 FILLER_150_1080 ();
 FILLCELL_X32 FILLER_150_1112 ();
 FILLCELL_X32 FILLER_150_1144 ();
 FILLCELL_X32 FILLER_150_1176 ();
 FILLCELL_X32 FILLER_150_1208 ();
 FILLCELL_X32 FILLER_150_1240 ();
 FILLCELL_X32 FILLER_150_1272 ();
 FILLCELL_X32 FILLER_150_1304 ();
 FILLCELL_X32 FILLER_150_1336 ();
 FILLCELL_X32 FILLER_150_1368 ();
 FILLCELL_X32 FILLER_150_1400 ();
 FILLCELL_X32 FILLER_150_1432 ();
 FILLCELL_X32 FILLER_150_1464 ();
 FILLCELL_X32 FILLER_150_1496 ();
 FILLCELL_X32 FILLER_150_1528 ();
 FILLCELL_X32 FILLER_150_1560 ();
 FILLCELL_X32 FILLER_150_1592 ();
 FILLCELL_X32 FILLER_150_1624 ();
 FILLCELL_X32 FILLER_150_1656 ();
 FILLCELL_X32 FILLER_150_1688 ();
 FILLCELL_X32 FILLER_150_1720 ();
 FILLCELL_X32 FILLER_150_1752 ();
 FILLCELL_X32 FILLER_150_1784 ();
 FILLCELL_X32 FILLER_150_1816 ();
 FILLCELL_X32 FILLER_150_1848 ();
 FILLCELL_X8 FILLER_150_1880 ();
 FILLCELL_X4 FILLER_150_1888 ();
 FILLCELL_X2 FILLER_150_1892 ();
 FILLCELL_X32 FILLER_150_1895 ();
 FILLCELL_X32 FILLER_150_1927 ();
 FILLCELL_X32 FILLER_150_1959 ();
 FILLCELL_X32 FILLER_150_1991 ();
 FILLCELL_X32 FILLER_150_2023 ();
 FILLCELL_X32 FILLER_150_2055 ();
 FILLCELL_X32 FILLER_150_2087 ();
 FILLCELL_X32 FILLER_150_2119 ();
 FILLCELL_X32 FILLER_150_2151 ();
 FILLCELL_X32 FILLER_150_2183 ();
 FILLCELL_X32 FILLER_150_2215 ();
 FILLCELL_X32 FILLER_150_2247 ();
 FILLCELL_X32 FILLER_150_2279 ();
 FILLCELL_X32 FILLER_150_2311 ();
 FILLCELL_X32 FILLER_150_2343 ();
 FILLCELL_X32 FILLER_150_2375 ();
 FILLCELL_X32 FILLER_150_2407 ();
 FILLCELL_X32 FILLER_150_2439 ();
 FILLCELL_X32 FILLER_150_2471 ();
 FILLCELL_X32 FILLER_150_2503 ();
 FILLCELL_X32 FILLER_150_2535 ();
 FILLCELL_X32 FILLER_150_2567 ();
 FILLCELL_X2 FILLER_150_2599 ();
 FILLCELL_X1 FILLER_150_2601 ();
 FILLCELL_X32 FILLER_151_1 ();
 FILLCELL_X32 FILLER_151_33 ();
 FILLCELL_X32 FILLER_151_65 ();
 FILLCELL_X32 FILLER_151_97 ();
 FILLCELL_X32 FILLER_151_129 ();
 FILLCELL_X32 FILLER_151_161 ();
 FILLCELL_X32 FILLER_151_193 ();
 FILLCELL_X32 FILLER_151_225 ();
 FILLCELL_X32 FILLER_151_257 ();
 FILLCELL_X32 FILLER_151_289 ();
 FILLCELL_X32 FILLER_151_321 ();
 FILLCELL_X32 FILLER_151_353 ();
 FILLCELL_X32 FILLER_151_385 ();
 FILLCELL_X32 FILLER_151_417 ();
 FILLCELL_X32 FILLER_151_449 ();
 FILLCELL_X32 FILLER_151_481 ();
 FILLCELL_X32 FILLER_151_513 ();
 FILLCELL_X32 FILLER_151_545 ();
 FILLCELL_X32 FILLER_151_577 ();
 FILLCELL_X32 FILLER_151_609 ();
 FILLCELL_X32 FILLER_151_641 ();
 FILLCELL_X32 FILLER_151_673 ();
 FILLCELL_X32 FILLER_151_705 ();
 FILLCELL_X32 FILLER_151_737 ();
 FILLCELL_X32 FILLER_151_769 ();
 FILLCELL_X32 FILLER_151_801 ();
 FILLCELL_X32 FILLER_151_833 ();
 FILLCELL_X32 FILLER_151_865 ();
 FILLCELL_X32 FILLER_151_897 ();
 FILLCELL_X32 FILLER_151_929 ();
 FILLCELL_X32 FILLER_151_961 ();
 FILLCELL_X32 FILLER_151_993 ();
 FILLCELL_X32 FILLER_151_1025 ();
 FILLCELL_X32 FILLER_151_1057 ();
 FILLCELL_X32 FILLER_151_1089 ();
 FILLCELL_X32 FILLER_151_1121 ();
 FILLCELL_X32 FILLER_151_1153 ();
 FILLCELL_X32 FILLER_151_1185 ();
 FILLCELL_X32 FILLER_151_1217 ();
 FILLCELL_X8 FILLER_151_1249 ();
 FILLCELL_X4 FILLER_151_1257 ();
 FILLCELL_X2 FILLER_151_1261 ();
 FILLCELL_X32 FILLER_151_1264 ();
 FILLCELL_X32 FILLER_151_1296 ();
 FILLCELL_X32 FILLER_151_1328 ();
 FILLCELL_X32 FILLER_151_1360 ();
 FILLCELL_X32 FILLER_151_1392 ();
 FILLCELL_X32 FILLER_151_1424 ();
 FILLCELL_X32 FILLER_151_1456 ();
 FILLCELL_X32 FILLER_151_1488 ();
 FILLCELL_X32 FILLER_151_1520 ();
 FILLCELL_X32 FILLER_151_1552 ();
 FILLCELL_X32 FILLER_151_1584 ();
 FILLCELL_X32 FILLER_151_1616 ();
 FILLCELL_X32 FILLER_151_1648 ();
 FILLCELL_X32 FILLER_151_1680 ();
 FILLCELL_X32 FILLER_151_1712 ();
 FILLCELL_X32 FILLER_151_1744 ();
 FILLCELL_X32 FILLER_151_1776 ();
 FILLCELL_X32 FILLER_151_1808 ();
 FILLCELL_X32 FILLER_151_1840 ();
 FILLCELL_X32 FILLER_151_1872 ();
 FILLCELL_X32 FILLER_151_1904 ();
 FILLCELL_X32 FILLER_151_1936 ();
 FILLCELL_X32 FILLER_151_1968 ();
 FILLCELL_X32 FILLER_151_2000 ();
 FILLCELL_X32 FILLER_151_2032 ();
 FILLCELL_X32 FILLER_151_2064 ();
 FILLCELL_X32 FILLER_151_2096 ();
 FILLCELL_X32 FILLER_151_2128 ();
 FILLCELL_X32 FILLER_151_2160 ();
 FILLCELL_X32 FILLER_151_2192 ();
 FILLCELL_X32 FILLER_151_2224 ();
 FILLCELL_X32 FILLER_151_2256 ();
 FILLCELL_X32 FILLER_151_2288 ();
 FILLCELL_X32 FILLER_151_2320 ();
 FILLCELL_X32 FILLER_151_2352 ();
 FILLCELL_X32 FILLER_151_2384 ();
 FILLCELL_X32 FILLER_151_2416 ();
 FILLCELL_X32 FILLER_151_2448 ();
 FILLCELL_X32 FILLER_151_2480 ();
 FILLCELL_X8 FILLER_151_2512 ();
 FILLCELL_X4 FILLER_151_2520 ();
 FILLCELL_X2 FILLER_151_2524 ();
 FILLCELL_X32 FILLER_151_2527 ();
 FILLCELL_X32 FILLER_151_2559 ();
 FILLCELL_X8 FILLER_151_2591 ();
 FILLCELL_X2 FILLER_151_2599 ();
 FILLCELL_X1 FILLER_151_2601 ();
 FILLCELL_X32 FILLER_152_1 ();
 FILLCELL_X32 FILLER_152_33 ();
 FILLCELL_X32 FILLER_152_65 ();
 FILLCELL_X32 FILLER_152_97 ();
 FILLCELL_X32 FILLER_152_129 ();
 FILLCELL_X32 FILLER_152_161 ();
 FILLCELL_X32 FILLER_152_193 ();
 FILLCELL_X32 FILLER_152_225 ();
 FILLCELL_X32 FILLER_152_257 ();
 FILLCELL_X32 FILLER_152_289 ();
 FILLCELL_X32 FILLER_152_321 ();
 FILLCELL_X32 FILLER_152_353 ();
 FILLCELL_X32 FILLER_152_385 ();
 FILLCELL_X32 FILLER_152_417 ();
 FILLCELL_X32 FILLER_152_449 ();
 FILLCELL_X32 FILLER_152_481 ();
 FILLCELL_X32 FILLER_152_513 ();
 FILLCELL_X32 FILLER_152_545 ();
 FILLCELL_X32 FILLER_152_577 ();
 FILLCELL_X16 FILLER_152_609 ();
 FILLCELL_X4 FILLER_152_625 ();
 FILLCELL_X2 FILLER_152_629 ();
 FILLCELL_X32 FILLER_152_632 ();
 FILLCELL_X32 FILLER_152_664 ();
 FILLCELL_X32 FILLER_152_696 ();
 FILLCELL_X32 FILLER_152_728 ();
 FILLCELL_X32 FILLER_152_760 ();
 FILLCELL_X32 FILLER_152_792 ();
 FILLCELL_X32 FILLER_152_824 ();
 FILLCELL_X32 FILLER_152_856 ();
 FILLCELL_X32 FILLER_152_888 ();
 FILLCELL_X32 FILLER_152_920 ();
 FILLCELL_X32 FILLER_152_952 ();
 FILLCELL_X32 FILLER_152_984 ();
 FILLCELL_X32 FILLER_152_1016 ();
 FILLCELL_X32 FILLER_152_1048 ();
 FILLCELL_X32 FILLER_152_1080 ();
 FILLCELL_X32 FILLER_152_1112 ();
 FILLCELL_X32 FILLER_152_1144 ();
 FILLCELL_X32 FILLER_152_1176 ();
 FILLCELL_X32 FILLER_152_1208 ();
 FILLCELL_X32 FILLER_152_1240 ();
 FILLCELL_X32 FILLER_152_1272 ();
 FILLCELL_X32 FILLER_152_1304 ();
 FILLCELL_X32 FILLER_152_1336 ();
 FILLCELL_X32 FILLER_152_1368 ();
 FILLCELL_X32 FILLER_152_1400 ();
 FILLCELL_X32 FILLER_152_1432 ();
 FILLCELL_X32 FILLER_152_1464 ();
 FILLCELL_X32 FILLER_152_1496 ();
 FILLCELL_X32 FILLER_152_1528 ();
 FILLCELL_X32 FILLER_152_1560 ();
 FILLCELL_X32 FILLER_152_1592 ();
 FILLCELL_X32 FILLER_152_1624 ();
 FILLCELL_X32 FILLER_152_1656 ();
 FILLCELL_X32 FILLER_152_1688 ();
 FILLCELL_X32 FILLER_152_1720 ();
 FILLCELL_X32 FILLER_152_1752 ();
 FILLCELL_X32 FILLER_152_1784 ();
 FILLCELL_X32 FILLER_152_1816 ();
 FILLCELL_X32 FILLER_152_1848 ();
 FILLCELL_X8 FILLER_152_1880 ();
 FILLCELL_X4 FILLER_152_1888 ();
 FILLCELL_X2 FILLER_152_1892 ();
 FILLCELL_X32 FILLER_152_1895 ();
 FILLCELL_X32 FILLER_152_1927 ();
 FILLCELL_X32 FILLER_152_1959 ();
 FILLCELL_X32 FILLER_152_1991 ();
 FILLCELL_X32 FILLER_152_2023 ();
 FILLCELL_X32 FILLER_152_2055 ();
 FILLCELL_X32 FILLER_152_2087 ();
 FILLCELL_X32 FILLER_152_2119 ();
 FILLCELL_X32 FILLER_152_2151 ();
 FILLCELL_X32 FILLER_152_2183 ();
 FILLCELL_X32 FILLER_152_2215 ();
 FILLCELL_X32 FILLER_152_2247 ();
 FILLCELL_X32 FILLER_152_2279 ();
 FILLCELL_X32 FILLER_152_2311 ();
 FILLCELL_X32 FILLER_152_2343 ();
 FILLCELL_X32 FILLER_152_2375 ();
 FILLCELL_X32 FILLER_152_2407 ();
 FILLCELL_X32 FILLER_152_2439 ();
 FILLCELL_X32 FILLER_152_2471 ();
 FILLCELL_X32 FILLER_152_2503 ();
 FILLCELL_X32 FILLER_152_2535 ();
 FILLCELL_X32 FILLER_152_2567 ();
 FILLCELL_X2 FILLER_152_2599 ();
 FILLCELL_X1 FILLER_152_2601 ();
 FILLCELL_X32 FILLER_153_1 ();
 FILLCELL_X32 FILLER_153_33 ();
 FILLCELL_X32 FILLER_153_65 ();
 FILLCELL_X32 FILLER_153_97 ();
 FILLCELL_X32 FILLER_153_129 ();
 FILLCELL_X32 FILLER_153_161 ();
 FILLCELL_X32 FILLER_153_193 ();
 FILLCELL_X32 FILLER_153_225 ();
 FILLCELL_X32 FILLER_153_257 ();
 FILLCELL_X32 FILLER_153_289 ();
 FILLCELL_X32 FILLER_153_321 ();
 FILLCELL_X32 FILLER_153_353 ();
 FILLCELL_X32 FILLER_153_385 ();
 FILLCELL_X32 FILLER_153_417 ();
 FILLCELL_X32 FILLER_153_449 ();
 FILLCELL_X32 FILLER_153_481 ();
 FILLCELL_X32 FILLER_153_513 ();
 FILLCELL_X32 FILLER_153_545 ();
 FILLCELL_X32 FILLER_153_577 ();
 FILLCELL_X32 FILLER_153_609 ();
 FILLCELL_X32 FILLER_153_641 ();
 FILLCELL_X32 FILLER_153_673 ();
 FILLCELL_X32 FILLER_153_705 ();
 FILLCELL_X32 FILLER_153_737 ();
 FILLCELL_X32 FILLER_153_769 ();
 FILLCELL_X32 FILLER_153_801 ();
 FILLCELL_X32 FILLER_153_833 ();
 FILLCELL_X32 FILLER_153_865 ();
 FILLCELL_X32 FILLER_153_897 ();
 FILLCELL_X32 FILLER_153_929 ();
 FILLCELL_X32 FILLER_153_961 ();
 FILLCELL_X32 FILLER_153_993 ();
 FILLCELL_X32 FILLER_153_1025 ();
 FILLCELL_X32 FILLER_153_1057 ();
 FILLCELL_X32 FILLER_153_1089 ();
 FILLCELL_X32 FILLER_153_1121 ();
 FILLCELL_X32 FILLER_153_1153 ();
 FILLCELL_X32 FILLER_153_1185 ();
 FILLCELL_X32 FILLER_153_1217 ();
 FILLCELL_X8 FILLER_153_1249 ();
 FILLCELL_X4 FILLER_153_1257 ();
 FILLCELL_X2 FILLER_153_1261 ();
 FILLCELL_X32 FILLER_153_1264 ();
 FILLCELL_X32 FILLER_153_1296 ();
 FILLCELL_X32 FILLER_153_1328 ();
 FILLCELL_X32 FILLER_153_1360 ();
 FILLCELL_X32 FILLER_153_1392 ();
 FILLCELL_X32 FILLER_153_1424 ();
 FILLCELL_X32 FILLER_153_1456 ();
 FILLCELL_X32 FILLER_153_1488 ();
 FILLCELL_X32 FILLER_153_1520 ();
 FILLCELL_X32 FILLER_153_1552 ();
 FILLCELL_X32 FILLER_153_1584 ();
 FILLCELL_X32 FILLER_153_1616 ();
 FILLCELL_X32 FILLER_153_1648 ();
 FILLCELL_X32 FILLER_153_1680 ();
 FILLCELL_X32 FILLER_153_1712 ();
 FILLCELL_X32 FILLER_153_1744 ();
 FILLCELL_X32 FILLER_153_1776 ();
 FILLCELL_X32 FILLER_153_1808 ();
 FILLCELL_X32 FILLER_153_1840 ();
 FILLCELL_X32 FILLER_153_1872 ();
 FILLCELL_X32 FILLER_153_1904 ();
 FILLCELL_X32 FILLER_153_1936 ();
 FILLCELL_X32 FILLER_153_1968 ();
 FILLCELL_X32 FILLER_153_2000 ();
 FILLCELL_X32 FILLER_153_2032 ();
 FILLCELL_X32 FILLER_153_2064 ();
 FILLCELL_X32 FILLER_153_2096 ();
 FILLCELL_X32 FILLER_153_2128 ();
 FILLCELL_X32 FILLER_153_2160 ();
 FILLCELL_X32 FILLER_153_2192 ();
 FILLCELL_X32 FILLER_153_2224 ();
 FILLCELL_X32 FILLER_153_2256 ();
 FILLCELL_X32 FILLER_153_2288 ();
 FILLCELL_X32 FILLER_153_2320 ();
 FILLCELL_X32 FILLER_153_2352 ();
 FILLCELL_X32 FILLER_153_2384 ();
 FILLCELL_X32 FILLER_153_2416 ();
 FILLCELL_X32 FILLER_153_2448 ();
 FILLCELL_X32 FILLER_153_2480 ();
 FILLCELL_X8 FILLER_153_2512 ();
 FILLCELL_X4 FILLER_153_2520 ();
 FILLCELL_X2 FILLER_153_2524 ();
 FILLCELL_X32 FILLER_153_2527 ();
 FILLCELL_X32 FILLER_153_2559 ();
 FILLCELL_X8 FILLER_153_2591 ();
 FILLCELL_X2 FILLER_153_2599 ();
 FILLCELL_X1 FILLER_153_2601 ();
 FILLCELL_X32 FILLER_154_1 ();
 FILLCELL_X32 FILLER_154_33 ();
 FILLCELL_X32 FILLER_154_65 ();
 FILLCELL_X32 FILLER_154_97 ();
 FILLCELL_X32 FILLER_154_129 ();
 FILLCELL_X32 FILLER_154_161 ();
 FILLCELL_X32 FILLER_154_193 ();
 FILLCELL_X32 FILLER_154_225 ();
 FILLCELL_X32 FILLER_154_257 ();
 FILLCELL_X32 FILLER_154_289 ();
 FILLCELL_X32 FILLER_154_321 ();
 FILLCELL_X32 FILLER_154_353 ();
 FILLCELL_X32 FILLER_154_385 ();
 FILLCELL_X32 FILLER_154_417 ();
 FILLCELL_X32 FILLER_154_449 ();
 FILLCELL_X32 FILLER_154_481 ();
 FILLCELL_X32 FILLER_154_513 ();
 FILLCELL_X32 FILLER_154_545 ();
 FILLCELL_X32 FILLER_154_577 ();
 FILLCELL_X16 FILLER_154_609 ();
 FILLCELL_X4 FILLER_154_625 ();
 FILLCELL_X2 FILLER_154_629 ();
 FILLCELL_X32 FILLER_154_632 ();
 FILLCELL_X32 FILLER_154_664 ();
 FILLCELL_X32 FILLER_154_696 ();
 FILLCELL_X32 FILLER_154_728 ();
 FILLCELL_X32 FILLER_154_760 ();
 FILLCELL_X32 FILLER_154_792 ();
 FILLCELL_X32 FILLER_154_824 ();
 FILLCELL_X32 FILLER_154_856 ();
 FILLCELL_X32 FILLER_154_888 ();
 FILLCELL_X32 FILLER_154_920 ();
 FILLCELL_X32 FILLER_154_952 ();
 FILLCELL_X32 FILLER_154_984 ();
 FILLCELL_X32 FILLER_154_1016 ();
 FILLCELL_X32 FILLER_154_1048 ();
 FILLCELL_X32 FILLER_154_1080 ();
 FILLCELL_X32 FILLER_154_1112 ();
 FILLCELL_X32 FILLER_154_1144 ();
 FILLCELL_X32 FILLER_154_1176 ();
 FILLCELL_X32 FILLER_154_1208 ();
 FILLCELL_X32 FILLER_154_1240 ();
 FILLCELL_X32 FILLER_154_1272 ();
 FILLCELL_X32 FILLER_154_1304 ();
 FILLCELL_X32 FILLER_154_1336 ();
 FILLCELL_X32 FILLER_154_1368 ();
 FILLCELL_X32 FILLER_154_1400 ();
 FILLCELL_X32 FILLER_154_1432 ();
 FILLCELL_X32 FILLER_154_1464 ();
 FILLCELL_X32 FILLER_154_1496 ();
 FILLCELL_X32 FILLER_154_1528 ();
 FILLCELL_X32 FILLER_154_1560 ();
 FILLCELL_X32 FILLER_154_1592 ();
 FILLCELL_X32 FILLER_154_1624 ();
 FILLCELL_X32 FILLER_154_1656 ();
 FILLCELL_X32 FILLER_154_1688 ();
 FILLCELL_X32 FILLER_154_1720 ();
 FILLCELL_X32 FILLER_154_1752 ();
 FILLCELL_X32 FILLER_154_1784 ();
 FILLCELL_X32 FILLER_154_1816 ();
 FILLCELL_X32 FILLER_154_1848 ();
 FILLCELL_X8 FILLER_154_1880 ();
 FILLCELL_X4 FILLER_154_1888 ();
 FILLCELL_X2 FILLER_154_1892 ();
 FILLCELL_X32 FILLER_154_1895 ();
 FILLCELL_X32 FILLER_154_1927 ();
 FILLCELL_X32 FILLER_154_1959 ();
 FILLCELL_X32 FILLER_154_1991 ();
 FILLCELL_X32 FILLER_154_2023 ();
 FILLCELL_X32 FILLER_154_2055 ();
 FILLCELL_X32 FILLER_154_2087 ();
 FILLCELL_X32 FILLER_154_2119 ();
 FILLCELL_X32 FILLER_154_2151 ();
 FILLCELL_X32 FILLER_154_2183 ();
 FILLCELL_X32 FILLER_154_2215 ();
 FILLCELL_X32 FILLER_154_2247 ();
 FILLCELL_X32 FILLER_154_2279 ();
 FILLCELL_X32 FILLER_154_2311 ();
 FILLCELL_X32 FILLER_154_2343 ();
 FILLCELL_X32 FILLER_154_2375 ();
 FILLCELL_X32 FILLER_154_2407 ();
 FILLCELL_X32 FILLER_154_2439 ();
 FILLCELL_X32 FILLER_154_2471 ();
 FILLCELL_X32 FILLER_154_2503 ();
 FILLCELL_X32 FILLER_154_2535 ();
 FILLCELL_X32 FILLER_154_2567 ();
 FILLCELL_X2 FILLER_154_2599 ();
 FILLCELL_X1 FILLER_154_2601 ();
 FILLCELL_X32 FILLER_155_1 ();
 FILLCELL_X32 FILLER_155_33 ();
 FILLCELL_X32 FILLER_155_65 ();
 FILLCELL_X32 FILLER_155_97 ();
 FILLCELL_X32 FILLER_155_129 ();
 FILLCELL_X32 FILLER_155_161 ();
 FILLCELL_X32 FILLER_155_193 ();
 FILLCELL_X32 FILLER_155_225 ();
 FILLCELL_X32 FILLER_155_257 ();
 FILLCELL_X32 FILLER_155_289 ();
 FILLCELL_X32 FILLER_155_321 ();
 FILLCELL_X32 FILLER_155_353 ();
 FILLCELL_X32 FILLER_155_385 ();
 FILLCELL_X32 FILLER_155_417 ();
 FILLCELL_X32 FILLER_155_449 ();
 FILLCELL_X32 FILLER_155_481 ();
 FILLCELL_X32 FILLER_155_513 ();
 FILLCELL_X32 FILLER_155_545 ();
 FILLCELL_X32 FILLER_155_577 ();
 FILLCELL_X32 FILLER_155_609 ();
 FILLCELL_X32 FILLER_155_641 ();
 FILLCELL_X32 FILLER_155_673 ();
 FILLCELL_X32 FILLER_155_705 ();
 FILLCELL_X32 FILLER_155_737 ();
 FILLCELL_X32 FILLER_155_769 ();
 FILLCELL_X32 FILLER_155_801 ();
 FILLCELL_X32 FILLER_155_833 ();
 FILLCELL_X32 FILLER_155_865 ();
 FILLCELL_X32 FILLER_155_897 ();
 FILLCELL_X32 FILLER_155_929 ();
 FILLCELL_X32 FILLER_155_961 ();
 FILLCELL_X32 FILLER_155_993 ();
 FILLCELL_X32 FILLER_155_1025 ();
 FILLCELL_X32 FILLER_155_1057 ();
 FILLCELL_X32 FILLER_155_1089 ();
 FILLCELL_X32 FILLER_155_1121 ();
 FILLCELL_X32 FILLER_155_1153 ();
 FILLCELL_X32 FILLER_155_1185 ();
 FILLCELL_X32 FILLER_155_1217 ();
 FILLCELL_X8 FILLER_155_1249 ();
 FILLCELL_X4 FILLER_155_1257 ();
 FILLCELL_X2 FILLER_155_1261 ();
 FILLCELL_X32 FILLER_155_1264 ();
 FILLCELL_X32 FILLER_155_1296 ();
 FILLCELL_X32 FILLER_155_1328 ();
 FILLCELL_X32 FILLER_155_1360 ();
 FILLCELL_X32 FILLER_155_1392 ();
 FILLCELL_X32 FILLER_155_1424 ();
 FILLCELL_X32 FILLER_155_1456 ();
 FILLCELL_X32 FILLER_155_1488 ();
 FILLCELL_X32 FILLER_155_1520 ();
 FILLCELL_X32 FILLER_155_1552 ();
 FILLCELL_X32 FILLER_155_1584 ();
 FILLCELL_X32 FILLER_155_1616 ();
 FILLCELL_X32 FILLER_155_1648 ();
 FILLCELL_X32 FILLER_155_1680 ();
 FILLCELL_X32 FILLER_155_1712 ();
 FILLCELL_X32 FILLER_155_1744 ();
 FILLCELL_X32 FILLER_155_1776 ();
 FILLCELL_X32 FILLER_155_1808 ();
 FILLCELL_X32 FILLER_155_1840 ();
 FILLCELL_X32 FILLER_155_1872 ();
 FILLCELL_X32 FILLER_155_1904 ();
 FILLCELL_X32 FILLER_155_1936 ();
 FILLCELL_X32 FILLER_155_1968 ();
 FILLCELL_X32 FILLER_155_2000 ();
 FILLCELL_X32 FILLER_155_2032 ();
 FILLCELL_X32 FILLER_155_2064 ();
 FILLCELL_X32 FILLER_155_2096 ();
 FILLCELL_X32 FILLER_155_2128 ();
 FILLCELL_X32 FILLER_155_2160 ();
 FILLCELL_X32 FILLER_155_2192 ();
 FILLCELL_X32 FILLER_155_2224 ();
 FILLCELL_X32 FILLER_155_2256 ();
 FILLCELL_X32 FILLER_155_2288 ();
 FILLCELL_X32 FILLER_155_2320 ();
 FILLCELL_X32 FILLER_155_2352 ();
 FILLCELL_X32 FILLER_155_2384 ();
 FILLCELL_X32 FILLER_155_2416 ();
 FILLCELL_X32 FILLER_155_2448 ();
 FILLCELL_X32 FILLER_155_2480 ();
 FILLCELL_X8 FILLER_155_2512 ();
 FILLCELL_X4 FILLER_155_2520 ();
 FILLCELL_X2 FILLER_155_2524 ();
 FILLCELL_X32 FILLER_155_2527 ();
 FILLCELL_X32 FILLER_155_2559 ();
 FILLCELL_X8 FILLER_155_2591 ();
 FILLCELL_X2 FILLER_155_2599 ();
 FILLCELL_X1 FILLER_155_2601 ();
 FILLCELL_X32 FILLER_156_1 ();
 FILLCELL_X32 FILLER_156_33 ();
 FILLCELL_X32 FILLER_156_65 ();
 FILLCELL_X32 FILLER_156_97 ();
 FILLCELL_X32 FILLER_156_129 ();
 FILLCELL_X32 FILLER_156_161 ();
 FILLCELL_X32 FILLER_156_193 ();
 FILLCELL_X32 FILLER_156_225 ();
 FILLCELL_X32 FILLER_156_257 ();
 FILLCELL_X32 FILLER_156_289 ();
 FILLCELL_X32 FILLER_156_321 ();
 FILLCELL_X32 FILLER_156_353 ();
 FILLCELL_X32 FILLER_156_385 ();
 FILLCELL_X32 FILLER_156_417 ();
 FILLCELL_X32 FILLER_156_449 ();
 FILLCELL_X32 FILLER_156_481 ();
 FILLCELL_X32 FILLER_156_513 ();
 FILLCELL_X32 FILLER_156_545 ();
 FILLCELL_X32 FILLER_156_577 ();
 FILLCELL_X16 FILLER_156_609 ();
 FILLCELL_X4 FILLER_156_625 ();
 FILLCELL_X2 FILLER_156_629 ();
 FILLCELL_X32 FILLER_156_632 ();
 FILLCELL_X32 FILLER_156_664 ();
 FILLCELL_X32 FILLER_156_696 ();
 FILLCELL_X32 FILLER_156_728 ();
 FILLCELL_X32 FILLER_156_760 ();
 FILLCELL_X32 FILLER_156_792 ();
 FILLCELL_X32 FILLER_156_824 ();
 FILLCELL_X32 FILLER_156_856 ();
 FILLCELL_X32 FILLER_156_888 ();
 FILLCELL_X32 FILLER_156_920 ();
 FILLCELL_X32 FILLER_156_952 ();
 FILLCELL_X32 FILLER_156_984 ();
 FILLCELL_X32 FILLER_156_1016 ();
 FILLCELL_X32 FILLER_156_1048 ();
 FILLCELL_X32 FILLER_156_1080 ();
 FILLCELL_X32 FILLER_156_1112 ();
 FILLCELL_X32 FILLER_156_1144 ();
 FILLCELL_X32 FILLER_156_1176 ();
 FILLCELL_X32 FILLER_156_1208 ();
 FILLCELL_X32 FILLER_156_1240 ();
 FILLCELL_X32 FILLER_156_1272 ();
 FILLCELL_X32 FILLER_156_1304 ();
 FILLCELL_X32 FILLER_156_1336 ();
 FILLCELL_X32 FILLER_156_1368 ();
 FILLCELL_X32 FILLER_156_1400 ();
 FILLCELL_X32 FILLER_156_1432 ();
 FILLCELL_X32 FILLER_156_1464 ();
 FILLCELL_X32 FILLER_156_1496 ();
 FILLCELL_X32 FILLER_156_1528 ();
 FILLCELL_X32 FILLER_156_1560 ();
 FILLCELL_X32 FILLER_156_1592 ();
 FILLCELL_X32 FILLER_156_1624 ();
 FILLCELL_X32 FILLER_156_1656 ();
 FILLCELL_X32 FILLER_156_1688 ();
 FILLCELL_X32 FILLER_156_1720 ();
 FILLCELL_X32 FILLER_156_1752 ();
 FILLCELL_X32 FILLER_156_1784 ();
 FILLCELL_X32 FILLER_156_1816 ();
 FILLCELL_X32 FILLER_156_1848 ();
 FILLCELL_X8 FILLER_156_1880 ();
 FILLCELL_X4 FILLER_156_1888 ();
 FILLCELL_X2 FILLER_156_1892 ();
 FILLCELL_X32 FILLER_156_1895 ();
 FILLCELL_X32 FILLER_156_1927 ();
 FILLCELL_X32 FILLER_156_1959 ();
 FILLCELL_X32 FILLER_156_1991 ();
 FILLCELL_X32 FILLER_156_2023 ();
 FILLCELL_X32 FILLER_156_2055 ();
 FILLCELL_X32 FILLER_156_2087 ();
 FILLCELL_X32 FILLER_156_2119 ();
 FILLCELL_X32 FILLER_156_2151 ();
 FILLCELL_X32 FILLER_156_2183 ();
 FILLCELL_X32 FILLER_156_2215 ();
 FILLCELL_X32 FILLER_156_2247 ();
 FILLCELL_X32 FILLER_156_2279 ();
 FILLCELL_X32 FILLER_156_2311 ();
 FILLCELL_X32 FILLER_156_2343 ();
 FILLCELL_X32 FILLER_156_2375 ();
 FILLCELL_X32 FILLER_156_2407 ();
 FILLCELL_X32 FILLER_156_2439 ();
 FILLCELL_X32 FILLER_156_2471 ();
 FILLCELL_X32 FILLER_156_2503 ();
 FILLCELL_X32 FILLER_156_2535 ();
 FILLCELL_X32 FILLER_156_2567 ();
 FILLCELL_X2 FILLER_156_2599 ();
 FILLCELL_X1 FILLER_156_2601 ();
 FILLCELL_X32 FILLER_157_1 ();
 FILLCELL_X32 FILLER_157_33 ();
 FILLCELL_X32 FILLER_157_65 ();
 FILLCELL_X32 FILLER_157_97 ();
 FILLCELL_X32 FILLER_157_129 ();
 FILLCELL_X32 FILLER_157_161 ();
 FILLCELL_X32 FILLER_157_193 ();
 FILLCELL_X32 FILLER_157_225 ();
 FILLCELL_X32 FILLER_157_257 ();
 FILLCELL_X32 FILLER_157_289 ();
 FILLCELL_X32 FILLER_157_321 ();
 FILLCELL_X32 FILLER_157_353 ();
 FILLCELL_X32 FILLER_157_385 ();
 FILLCELL_X32 FILLER_157_417 ();
 FILLCELL_X32 FILLER_157_449 ();
 FILLCELL_X32 FILLER_157_481 ();
 FILLCELL_X32 FILLER_157_513 ();
 FILLCELL_X32 FILLER_157_545 ();
 FILLCELL_X32 FILLER_157_577 ();
 FILLCELL_X32 FILLER_157_609 ();
 FILLCELL_X32 FILLER_157_641 ();
 FILLCELL_X32 FILLER_157_673 ();
 FILLCELL_X32 FILLER_157_705 ();
 FILLCELL_X32 FILLER_157_737 ();
 FILLCELL_X32 FILLER_157_769 ();
 FILLCELL_X32 FILLER_157_801 ();
 FILLCELL_X32 FILLER_157_833 ();
 FILLCELL_X32 FILLER_157_865 ();
 FILLCELL_X32 FILLER_157_897 ();
 FILLCELL_X32 FILLER_157_929 ();
 FILLCELL_X32 FILLER_157_961 ();
 FILLCELL_X32 FILLER_157_993 ();
 FILLCELL_X32 FILLER_157_1025 ();
 FILLCELL_X32 FILLER_157_1057 ();
 FILLCELL_X32 FILLER_157_1089 ();
 FILLCELL_X32 FILLER_157_1121 ();
 FILLCELL_X32 FILLER_157_1153 ();
 FILLCELL_X32 FILLER_157_1185 ();
 FILLCELL_X32 FILLER_157_1217 ();
 FILLCELL_X8 FILLER_157_1249 ();
 FILLCELL_X4 FILLER_157_1257 ();
 FILLCELL_X2 FILLER_157_1261 ();
 FILLCELL_X32 FILLER_157_1264 ();
 FILLCELL_X32 FILLER_157_1296 ();
 FILLCELL_X32 FILLER_157_1328 ();
 FILLCELL_X32 FILLER_157_1360 ();
 FILLCELL_X32 FILLER_157_1392 ();
 FILLCELL_X32 FILLER_157_1424 ();
 FILLCELL_X32 FILLER_157_1456 ();
 FILLCELL_X32 FILLER_157_1488 ();
 FILLCELL_X32 FILLER_157_1520 ();
 FILLCELL_X32 FILLER_157_1552 ();
 FILLCELL_X32 FILLER_157_1584 ();
 FILLCELL_X32 FILLER_157_1616 ();
 FILLCELL_X32 FILLER_157_1648 ();
 FILLCELL_X32 FILLER_157_1680 ();
 FILLCELL_X32 FILLER_157_1712 ();
 FILLCELL_X32 FILLER_157_1744 ();
 FILLCELL_X32 FILLER_157_1776 ();
 FILLCELL_X32 FILLER_157_1808 ();
 FILLCELL_X32 FILLER_157_1840 ();
 FILLCELL_X32 FILLER_157_1872 ();
 FILLCELL_X32 FILLER_157_1904 ();
 FILLCELL_X32 FILLER_157_1936 ();
 FILLCELL_X32 FILLER_157_1968 ();
 FILLCELL_X32 FILLER_157_2000 ();
 FILLCELL_X32 FILLER_157_2032 ();
 FILLCELL_X32 FILLER_157_2064 ();
 FILLCELL_X32 FILLER_157_2096 ();
 FILLCELL_X32 FILLER_157_2128 ();
 FILLCELL_X32 FILLER_157_2160 ();
 FILLCELL_X32 FILLER_157_2192 ();
 FILLCELL_X32 FILLER_157_2224 ();
 FILLCELL_X32 FILLER_157_2256 ();
 FILLCELL_X32 FILLER_157_2288 ();
 FILLCELL_X32 FILLER_157_2320 ();
 FILLCELL_X32 FILLER_157_2352 ();
 FILLCELL_X32 FILLER_157_2384 ();
 FILLCELL_X32 FILLER_157_2416 ();
 FILLCELL_X32 FILLER_157_2448 ();
 FILLCELL_X32 FILLER_157_2480 ();
 FILLCELL_X8 FILLER_157_2512 ();
 FILLCELL_X4 FILLER_157_2520 ();
 FILLCELL_X2 FILLER_157_2524 ();
 FILLCELL_X32 FILLER_157_2527 ();
 FILLCELL_X32 FILLER_157_2559 ();
 FILLCELL_X8 FILLER_157_2591 ();
 FILLCELL_X2 FILLER_157_2599 ();
 FILLCELL_X1 FILLER_157_2601 ();
 FILLCELL_X32 FILLER_158_1 ();
 FILLCELL_X32 FILLER_158_33 ();
 FILLCELL_X32 FILLER_158_65 ();
 FILLCELL_X32 FILLER_158_97 ();
 FILLCELL_X32 FILLER_158_129 ();
 FILLCELL_X32 FILLER_158_161 ();
 FILLCELL_X32 FILLER_158_193 ();
 FILLCELL_X32 FILLER_158_225 ();
 FILLCELL_X32 FILLER_158_257 ();
 FILLCELL_X32 FILLER_158_289 ();
 FILLCELL_X32 FILLER_158_321 ();
 FILLCELL_X32 FILLER_158_353 ();
 FILLCELL_X32 FILLER_158_385 ();
 FILLCELL_X32 FILLER_158_417 ();
 FILLCELL_X32 FILLER_158_449 ();
 FILLCELL_X32 FILLER_158_481 ();
 FILLCELL_X32 FILLER_158_513 ();
 FILLCELL_X32 FILLER_158_545 ();
 FILLCELL_X32 FILLER_158_577 ();
 FILLCELL_X16 FILLER_158_609 ();
 FILLCELL_X4 FILLER_158_625 ();
 FILLCELL_X2 FILLER_158_629 ();
 FILLCELL_X32 FILLER_158_632 ();
 FILLCELL_X32 FILLER_158_664 ();
 FILLCELL_X32 FILLER_158_696 ();
 FILLCELL_X32 FILLER_158_728 ();
 FILLCELL_X32 FILLER_158_760 ();
 FILLCELL_X32 FILLER_158_792 ();
 FILLCELL_X32 FILLER_158_824 ();
 FILLCELL_X32 FILLER_158_856 ();
 FILLCELL_X32 FILLER_158_888 ();
 FILLCELL_X32 FILLER_158_920 ();
 FILLCELL_X32 FILLER_158_952 ();
 FILLCELL_X32 FILLER_158_984 ();
 FILLCELL_X32 FILLER_158_1016 ();
 FILLCELL_X32 FILLER_158_1048 ();
 FILLCELL_X32 FILLER_158_1080 ();
 FILLCELL_X32 FILLER_158_1112 ();
 FILLCELL_X32 FILLER_158_1144 ();
 FILLCELL_X32 FILLER_158_1176 ();
 FILLCELL_X32 FILLER_158_1208 ();
 FILLCELL_X32 FILLER_158_1240 ();
 FILLCELL_X32 FILLER_158_1272 ();
 FILLCELL_X32 FILLER_158_1304 ();
 FILLCELL_X32 FILLER_158_1336 ();
 FILLCELL_X32 FILLER_158_1368 ();
 FILLCELL_X32 FILLER_158_1400 ();
 FILLCELL_X32 FILLER_158_1432 ();
 FILLCELL_X32 FILLER_158_1464 ();
 FILLCELL_X32 FILLER_158_1496 ();
 FILLCELL_X32 FILLER_158_1528 ();
 FILLCELL_X32 FILLER_158_1560 ();
 FILLCELL_X32 FILLER_158_1592 ();
 FILLCELL_X32 FILLER_158_1624 ();
 FILLCELL_X32 FILLER_158_1656 ();
 FILLCELL_X32 FILLER_158_1688 ();
 FILLCELL_X32 FILLER_158_1720 ();
 FILLCELL_X32 FILLER_158_1752 ();
 FILLCELL_X32 FILLER_158_1784 ();
 FILLCELL_X32 FILLER_158_1816 ();
 FILLCELL_X32 FILLER_158_1848 ();
 FILLCELL_X8 FILLER_158_1880 ();
 FILLCELL_X4 FILLER_158_1888 ();
 FILLCELL_X2 FILLER_158_1892 ();
 FILLCELL_X32 FILLER_158_1895 ();
 FILLCELL_X32 FILLER_158_1927 ();
 FILLCELL_X32 FILLER_158_1959 ();
 FILLCELL_X32 FILLER_158_1991 ();
 FILLCELL_X32 FILLER_158_2023 ();
 FILLCELL_X32 FILLER_158_2055 ();
 FILLCELL_X32 FILLER_158_2087 ();
 FILLCELL_X32 FILLER_158_2119 ();
 FILLCELL_X32 FILLER_158_2151 ();
 FILLCELL_X32 FILLER_158_2183 ();
 FILLCELL_X32 FILLER_158_2215 ();
 FILLCELL_X32 FILLER_158_2247 ();
 FILLCELL_X32 FILLER_158_2279 ();
 FILLCELL_X32 FILLER_158_2311 ();
 FILLCELL_X32 FILLER_158_2343 ();
 FILLCELL_X32 FILLER_158_2375 ();
 FILLCELL_X32 FILLER_158_2407 ();
 FILLCELL_X32 FILLER_158_2439 ();
 FILLCELL_X32 FILLER_158_2471 ();
 FILLCELL_X32 FILLER_158_2503 ();
 FILLCELL_X32 FILLER_158_2535 ();
 FILLCELL_X32 FILLER_158_2567 ();
 FILLCELL_X2 FILLER_158_2599 ();
 FILLCELL_X1 FILLER_158_2601 ();
 FILLCELL_X32 FILLER_159_1 ();
 FILLCELL_X32 FILLER_159_33 ();
 FILLCELL_X32 FILLER_159_65 ();
 FILLCELL_X32 FILLER_159_97 ();
 FILLCELL_X32 FILLER_159_129 ();
 FILLCELL_X32 FILLER_159_161 ();
 FILLCELL_X32 FILLER_159_193 ();
 FILLCELL_X32 FILLER_159_225 ();
 FILLCELL_X32 FILLER_159_257 ();
 FILLCELL_X32 FILLER_159_289 ();
 FILLCELL_X32 FILLER_159_321 ();
 FILLCELL_X32 FILLER_159_353 ();
 FILLCELL_X32 FILLER_159_385 ();
 FILLCELL_X32 FILLER_159_417 ();
 FILLCELL_X32 FILLER_159_449 ();
 FILLCELL_X32 FILLER_159_481 ();
 FILLCELL_X32 FILLER_159_513 ();
 FILLCELL_X32 FILLER_159_545 ();
 FILLCELL_X32 FILLER_159_577 ();
 FILLCELL_X32 FILLER_159_609 ();
 FILLCELL_X32 FILLER_159_641 ();
 FILLCELL_X32 FILLER_159_673 ();
 FILLCELL_X32 FILLER_159_705 ();
 FILLCELL_X32 FILLER_159_737 ();
 FILLCELL_X32 FILLER_159_769 ();
 FILLCELL_X32 FILLER_159_801 ();
 FILLCELL_X32 FILLER_159_833 ();
 FILLCELL_X32 FILLER_159_865 ();
 FILLCELL_X32 FILLER_159_897 ();
 FILLCELL_X32 FILLER_159_929 ();
 FILLCELL_X32 FILLER_159_961 ();
 FILLCELL_X32 FILLER_159_993 ();
 FILLCELL_X32 FILLER_159_1025 ();
 FILLCELL_X32 FILLER_159_1057 ();
 FILLCELL_X32 FILLER_159_1089 ();
 FILLCELL_X32 FILLER_159_1121 ();
 FILLCELL_X32 FILLER_159_1153 ();
 FILLCELL_X32 FILLER_159_1185 ();
 FILLCELL_X32 FILLER_159_1217 ();
 FILLCELL_X8 FILLER_159_1249 ();
 FILLCELL_X4 FILLER_159_1257 ();
 FILLCELL_X2 FILLER_159_1261 ();
 FILLCELL_X32 FILLER_159_1264 ();
 FILLCELL_X32 FILLER_159_1296 ();
 FILLCELL_X32 FILLER_159_1328 ();
 FILLCELL_X32 FILLER_159_1360 ();
 FILLCELL_X32 FILLER_159_1392 ();
 FILLCELL_X32 FILLER_159_1424 ();
 FILLCELL_X32 FILLER_159_1456 ();
 FILLCELL_X32 FILLER_159_1488 ();
 FILLCELL_X32 FILLER_159_1520 ();
 FILLCELL_X32 FILLER_159_1552 ();
 FILLCELL_X32 FILLER_159_1584 ();
 FILLCELL_X32 FILLER_159_1616 ();
 FILLCELL_X32 FILLER_159_1648 ();
 FILLCELL_X32 FILLER_159_1680 ();
 FILLCELL_X32 FILLER_159_1712 ();
 FILLCELL_X32 FILLER_159_1744 ();
 FILLCELL_X32 FILLER_159_1776 ();
 FILLCELL_X32 FILLER_159_1808 ();
 FILLCELL_X32 FILLER_159_1840 ();
 FILLCELL_X32 FILLER_159_1872 ();
 FILLCELL_X32 FILLER_159_1904 ();
 FILLCELL_X32 FILLER_159_1936 ();
 FILLCELL_X32 FILLER_159_1968 ();
 FILLCELL_X32 FILLER_159_2000 ();
 FILLCELL_X32 FILLER_159_2032 ();
 FILLCELL_X32 FILLER_159_2064 ();
 FILLCELL_X32 FILLER_159_2096 ();
 FILLCELL_X32 FILLER_159_2128 ();
 FILLCELL_X32 FILLER_159_2160 ();
 FILLCELL_X32 FILLER_159_2192 ();
 FILLCELL_X32 FILLER_159_2224 ();
 FILLCELL_X32 FILLER_159_2256 ();
 FILLCELL_X32 FILLER_159_2288 ();
 FILLCELL_X32 FILLER_159_2320 ();
 FILLCELL_X32 FILLER_159_2352 ();
 FILLCELL_X32 FILLER_159_2384 ();
 FILLCELL_X32 FILLER_159_2416 ();
 FILLCELL_X32 FILLER_159_2448 ();
 FILLCELL_X32 FILLER_159_2480 ();
 FILLCELL_X8 FILLER_159_2512 ();
 FILLCELL_X4 FILLER_159_2520 ();
 FILLCELL_X2 FILLER_159_2524 ();
 FILLCELL_X32 FILLER_159_2527 ();
 FILLCELL_X32 FILLER_159_2559 ();
 FILLCELL_X8 FILLER_159_2591 ();
 FILLCELL_X2 FILLER_159_2599 ();
 FILLCELL_X1 FILLER_159_2601 ();
 FILLCELL_X32 FILLER_160_1 ();
 FILLCELL_X32 FILLER_160_33 ();
 FILLCELL_X32 FILLER_160_65 ();
 FILLCELL_X32 FILLER_160_97 ();
 FILLCELL_X32 FILLER_160_129 ();
 FILLCELL_X32 FILLER_160_161 ();
 FILLCELL_X32 FILLER_160_193 ();
 FILLCELL_X32 FILLER_160_225 ();
 FILLCELL_X32 FILLER_160_257 ();
 FILLCELL_X32 FILLER_160_289 ();
 FILLCELL_X32 FILLER_160_321 ();
 FILLCELL_X32 FILLER_160_353 ();
 FILLCELL_X32 FILLER_160_385 ();
 FILLCELL_X32 FILLER_160_417 ();
 FILLCELL_X32 FILLER_160_449 ();
 FILLCELL_X32 FILLER_160_481 ();
 FILLCELL_X32 FILLER_160_513 ();
 FILLCELL_X32 FILLER_160_545 ();
 FILLCELL_X32 FILLER_160_577 ();
 FILLCELL_X16 FILLER_160_609 ();
 FILLCELL_X4 FILLER_160_625 ();
 FILLCELL_X2 FILLER_160_629 ();
 FILLCELL_X32 FILLER_160_632 ();
 FILLCELL_X32 FILLER_160_664 ();
 FILLCELL_X32 FILLER_160_696 ();
 FILLCELL_X32 FILLER_160_728 ();
 FILLCELL_X32 FILLER_160_760 ();
 FILLCELL_X32 FILLER_160_792 ();
 FILLCELL_X32 FILLER_160_824 ();
 FILLCELL_X32 FILLER_160_856 ();
 FILLCELL_X32 FILLER_160_888 ();
 FILLCELL_X32 FILLER_160_920 ();
 FILLCELL_X32 FILLER_160_952 ();
 FILLCELL_X32 FILLER_160_984 ();
 FILLCELL_X32 FILLER_160_1016 ();
 FILLCELL_X32 FILLER_160_1048 ();
 FILLCELL_X32 FILLER_160_1080 ();
 FILLCELL_X32 FILLER_160_1112 ();
 FILLCELL_X32 FILLER_160_1144 ();
 FILLCELL_X32 FILLER_160_1176 ();
 FILLCELL_X32 FILLER_160_1208 ();
 FILLCELL_X32 FILLER_160_1240 ();
 FILLCELL_X32 FILLER_160_1272 ();
 FILLCELL_X32 FILLER_160_1304 ();
 FILLCELL_X32 FILLER_160_1336 ();
 FILLCELL_X32 FILLER_160_1368 ();
 FILLCELL_X32 FILLER_160_1400 ();
 FILLCELL_X32 FILLER_160_1432 ();
 FILLCELL_X32 FILLER_160_1464 ();
 FILLCELL_X32 FILLER_160_1496 ();
 FILLCELL_X32 FILLER_160_1528 ();
 FILLCELL_X32 FILLER_160_1560 ();
 FILLCELL_X32 FILLER_160_1592 ();
 FILLCELL_X32 FILLER_160_1624 ();
 FILLCELL_X32 FILLER_160_1656 ();
 FILLCELL_X32 FILLER_160_1688 ();
 FILLCELL_X32 FILLER_160_1720 ();
 FILLCELL_X32 FILLER_160_1752 ();
 FILLCELL_X32 FILLER_160_1784 ();
 FILLCELL_X32 FILLER_160_1816 ();
 FILLCELL_X32 FILLER_160_1848 ();
 FILLCELL_X8 FILLER_160_1880 ();
 FILLCELL_X4 FILLER_160_1888 ();
 FILLCELL_X2 FILLER_160_1892 ();
 FILLCELL_X32 FILLER_160_1895 ();
 FILLCELL_X32 FILLER_160_1927 ();
 FILLCELL_X32 FILLER_160_1959 ();
 FILLCELL_X32 FILLER_160_1991 ();
 FILLCELL_X32 FILLER_160_2023 ();
 FILLCELL_X32 FILLER_160_2055 ();
 FILLCELL_X32 FILLER_160_2087 ();
 FILLCELL_X32 FILLER_160_2119 ();
 FILLCELL_X32 FILLER_160_2151 ();
 FILLCELL_X32 FILLER_160_2183 ();
 FILLCELL_X32 FILLER_160_2215 ();
 FILLCELL_X32 FILLER_160_2247 ();
 FILLCELL_X32 FILLER_160_2279 ();
 FILLCELL_X32 FILLER_160_2311 ();
 FILLCELL_X32 FILLER_160_2343 ();
 FILLCELL_X32 FILLER_160_2375 ();
 FILLCELL_X32 FILLER_160_2407 ();
 FILLCELL_X32 FILLER_160_2439 ();
 FILLCELL_X32 FILLER_160_2471 ();
 FILLCELL_X32 FILLER_160_2503 ();
 FILLCELL_X32 FILLER_160_2535 ();
 FILLCELL_X32 FILLER_160_2567 ();
 FILLCELL_X2 FILLER_160_2599 ();
 FILLCELL_X1 FILLER_160_2601 ();
 FILLCELL_X32 FILLER_161_1 ();
 FILLCELL_X32 FILLER_161_33 ();
 FILLCELL_X32 FILLER_161_65 ();
 FILLCELL_X32 FILLER_161_97 ();
 FILLCELL_X32 FILLER_161_129 ();
 FILLCELL_X32 FILLER_161_161 ();
 FILLCELL_X32 FILLER_161_193 ();
 FILLCELL_X32 FILLER_161_225 ();
 FILLCELL_X32 FILLER_161_257 ();
 FILLCELL_X32 FILLER_161_289 ();
 FILLCELL_X32 FILLER_161_321 ();
 FILLCELL_X32 FILLER_161_353 ();
 FILLCELL_X32 FILLER_161_385 ();
 FILLCELL_X32 FILLER_161_417 ();
 FILLCELL_X32 FILLER_161_449 ();
 FILLCELL_X32 FILLER_161_481 ();
 FILLCELL_X32 FILLER_161_513 ();
 FILLCELL_X32 FILLER_161_545 ();
 FILLCELL_X32 FILLER_161_577 ();
 FILLCELL_X32 FILLER_161_609 ();
 FILLCELL_X32 FILLER_161_641 ();
 FILLCELL_X32 FILLER_161_673 ();
 FILLCELL_X32 FILLER_161_705 ();
 FILLCELL_X32 FILLER_161_737 ();
 FILLCELL_X32 FILLER_161_769 ();
 FILLCELL_X32 FILLER_161_801 ();
 FILLCELL_X32 FILLER_161_833 ();
 FILLCELL_X32 FILLER_161_865 ();
 FILLCELL_X32 FILLER_161_897 ();
 FILLCELL_X32 FILLER_161_929 ();
 FILLCELL_X32 FILLER_161_961 ();
 FILLCELL_X32 FILLER_161_993 ();
 FILLCELL_X32 FILLER_161_1025 ();
 FILLCELL_X32 FILLER_161_1057 ();
 FILLCELL_X32 FILLER_161_1089 ();
 FILLCELL_X32 FILLER_161_1121 ();
 FILLCELL_X32 FILLER_161_1153 ();
 FILLCELL_X32 FILLER_161_1185 ();
 FILLCELL_X32 FILLER_161_1217 ();
 FILLCELL_X8 FILLER_161_1249 ();
 FILLCELL_X4 FILLER_161_1257 ();
 FILLCELL_X2 FILLER_161_1261 ();
 FILLCELL_X32 FILLER_161_1264 ();
 FILLCELL_X32 FILLER_161_1296 ();
 FILLCELL_X32 FILLER_161_1328 ();
 FILLCELL_X32 FILLER_161_1360 ();
 FILLCELL_X32 FILLER_161_1392 ();
 FILLCELL_X32 FILLER_161_1424 ();
 FILLCELL_X32 FILLER_161_1456 ();
 FILLCELL_X16 FILLER_161_1488 ();
 FILLCELL_X32 FILLER_161_1521 ();
 FILLCELL_X32 FILLER_161_1553 ();
 FILLCELL_X32 FILLER_161_1585 ();
 FILLCELL_X32 FILLER_161_1617 ();
 FILLCELL_X32 FILLER_161_1649 ();
 FILLCELL_X32 FILLER_161_1681 ();
 FILLCELL_X32 FILLER_161_1713 ();
 FILLCELL_X32 FILLER_161_1745 ();
 FILLCELL_X32 FILLER_161_1777 ();
 FILLCELL_X32 FILLER_161_1809 ();
 FILLCELL_X32 FILLER_161_1841 ();
 FILLCELL_X32 FILLER_161_1873 ();
 FILLCELL_X32 FILLER_161_1905 ();
 FILLCELL_X32 FILLER_161_1937 ();
 FILLCELL_X32 FILLER_161_1969 ();
 FILLCELL_X32 FILLER_161_2001 ();
 FILLCELL_X32 FILLER_161_2033 ();
 FILLCELL_X32 FILLER_161_2065 ();
 FILLCELL_X32 FILLER_161_2097 ();
 FILLCELL_X32 FILLER_161_2129 ();
 FILLCELL_X32 FILLER_161_2161 ();
 FILLCELL_X32 FILLER_161_2193 ();
 FILLCELL_X32 FILLER_161_2225 ();
 FILLCELL_X32 FILLER_161_2257 ();
 FILLCELL_X32 FILLER_161_2289 ();
 FILLCELL_X32 FILLER_161_2321 ();
 FILLCELL_X32 FILLER_161_2353 ();
 FILLCELL_X32 FILLER_161_2385 ();
 FILLCELL_X32 FILLER_161_2417 ();
 FILLCELL_X32 FILLER_161_2449 ();
 FILLCELL_X32 FILLER_161_2481 ();
 FILLCELL_X8 FILLER_161_2513 ();
 FILLCELL_X4 FILLER_161_2521 ();
 FILLCELL_X1 FILLER_161_2525 ();
 FILLCELL_X32 FILLER_161_2527 ();
 FILLCELL_X32 FILLER_161_2559 ();
 FILLCELL_X8 FILLER_161_2591 ();
 FILLCELL_X2 FILLER_161_2599 ();
 FILLCELL_X1 FILLER_161_2601 ();
 FILLCELL_X32 FILLER_162_1 ();
 FILLCELL_X32 FILLER_162_33 ();
 FILLCELL_X32 FILLER_162_65 ();
 FILLCELL_X32 FILLER_162_97 ();
 FILLCELL_X32 FILLER_162_129 ();
 FILLCELL_X32 FILLER_162_161 ();
 FILLCELL_X32 FILLER_162_193 ();
 FILLCELL_X32 FILLER_162_225 ();
 FILLCELL_X32 FILLER_162_257 ();
 FILLCELL_X32 FILLER_162_289 ();
 FILLCELL_X32 FILLER_162_321 ();
 FILLCELL_X32 FILLER_162_353 ();
 FILLCELL_X32 FILLER_162_385 ();
 FILLCELL_X32 FILLER_162_417 ();
 FILLCELL_X32 FILLER_162_449 ();
 FILLCELL_X32 FILLER_162_481 ();
 FILLCELL_X32 FILLER_162_513 ();
 FILLCELL_X32 FILLER_162_545 ();
 FILLCELL_X32 FILLER_162_577 ();
 FILLCELL_X16 FILLER_162_609 ();
 FILLCELL_X4 FILLER_162_625 ();
 FILLCELL_X2 FILLER_162_629 ();
 FILLCELL_X32 FILLER_162_632 ();
 FILLCELL_X32 FILLER_162_664 ();
 FILLCELL_X32 FILLER_162_696 ();
 FILLCELL_X32 FILLER_162_728 ();
 FILLCELL_X32 FILLER_162_760 ();
 FILLCELL_X32 FILLER_162_792 ();
 FILLCELL_X32 FILLER_162_824 ();
 FILLCELL_X32 FILLER_162_856 ();
 FILLCELL_X32 FILLER_162_888 ();
 FILLCELL_X32 FILLER_162_920 ();
 FILLCELL_X32 FILLER_162_952 ();
 FILLCELL_X32 FILLER_162_984 ();
 FILLCELL_X32 FILLER_162_1016 ();
 FILLCELL_X32 FILLER_162_1048 ();
 FILLCELL_X32 FILLER_162_1080 ();
 FILLCELL_X32 FILLER_162_1112 ();
 FILLCELL_X32 FILLER_162_1144 ();
 FILLCELL_X32 FILLER_162_1176 ();
 FILLCELL_X32 FILLER_162_1208 ();
 FILLCELL_X32 FILLER_162_1240 ();
 FILLCELL_X32 FILLER_162_1272 ();
 FILLCELL_X32 FILLER_162_1321 ();
 FILLCELL_X32 FILLER_162_1353 ();
 FILLCELL_X32 FILLER_162_1385 ();
 FILLCELL_X32 FILLER_162_1417 ();
 FILLCELL_X16 FILLER_162_1449 ();
 FILLCELL_X8 FILLER_162_1465 ();
 FILLCELL_X2 FILLER_162_1473 ();
 FILLCELL_X8 FILLER_162_1499 ();
 FILLCELL_X4 FILLER_162_1507 ();
 FILLCELL_X2 FILLER_162_1511 ();
 FILLCELL_X32 FILLER_162_1537 ();
 FILLCELL_X32 FILLER_162_1569 ();
 FILLCELL_X32 FILLER_162_1601 ();
 FILLCELL_X32 FILLER_162_1633 ();
 FILLCELL_X32 FILLER_162_1665 ();
 FILLCELL_X32 FILLER_162_1697 ();
 FILLCELL_X32 FILLER_162_1729 ();
 FILLCELL_X32 FILLER_162_1761 ();
 FILLCELL_X32 FILLER_162_1793 ();
 FILLCELL_X32 FILLER_162_1825 ();
 FILLCELL_X32 FILLER_162_1857 ();
 FILLCELL_X4 FILLER_162_1889 ();
 FILLCELL_X1 FILLER_162_1893 ();
 FILLCELL_X32 FILLER_162_1895 ();
 FILLCELL_X32 FILLER_162_1927 ();
 FILLCELL_X32 FILLER_162_1959 ();
 FILLCELL_X32 FILLER_162_1991 ();
 FILLCELL_X32 FILLER_162_2023 ();
 FILLCELL_X32 FILLER_162_2055 ();
 FILLCELL_X32 FILLER_162_2087 ();
 FILLCELL_X32 FILLER_162_2119 ();
 FILLCELL_X32 FILLER_162_2151 ();
 FILLCELL_X32 FILLER_162_2183 ();
 FILLCELL_X32 FILLER_162_2215 ();
 FILLCELL_X32 FILLER_162_2247 ();
 FILLCELL_X32 FILLER_162_2279 ();
 FILLCELL_X32 FILLER_162_2311 ();
 FILLCELL_X32 FILLER_162_2343 ();
 FILLCELL_X32 FILLER_162_2375 ();
 FILLCELL_X32 FILLER_162_2407 ();
 FILLCELL_X32 FILLER_162_2439 ();
 FILLCELL_X32 FILLER_162_2471 ();
 FILLCELL_X32 FILLER_162_2503 ();
 FILLCELL_X32 FILLER_162_2535 ();
 FILLCELL_X32 FILLER_162_2567 ();
 FILLCELL_X2 FILLER_162_2599 ();
 FILLCELL_X1 FILLER_162_2601 ();
 FILLCELL_X32 FILLER_163_1 ();
 FILLCELL_X32 FILLER_163_33 ();
 FILLCELL_X32 FILLER_163_65 ();
 FILLCELL_X32 FILLER_163_97 ();
 FILLCELL_X32 FILLER_163_129 ();
 FILLCELL_X32 FILLER_163_161 ();
 FILLCELL_X32 FILLER_163_193 ();
 FILLCELL_X32 FILLER_163_225 ();
 FILLCELL_X32 FILLER_163_257 ();
 FILLCELL_X32 FILLER_163_289 ();
 FILLCELL_X32 FILLER_163_321 ();
 FILLCELL_X32 FILLER_163_353 ();
 FILLCELL_X32 FILLER_163_385 ();
 FILLCELL_X32 FILLER_163_417 ();
 FILLCELL_X32 FILLER_163_449 ();
 FILLCELL_X32 FILLER_163_481 ();
 FILLCELL_X32 FILLER_163_513 ();
 FILLCELL_X32 FILLER_163_545 ();
 FILLCELL_X32 FILLER_163_577 ();
 FILLCELL_X32 FILLER_163_609 ();
 FILLCELL_X32 FILLER_163_641 ();
 FILLCELL_X32 FILLER_163_673 ();
 FILLCELL_X32 FILLER_163_705 ();
 FILLCELL_X32 FILLER_163_737 ();
 FILLCELL_X32 FILLER_163_769 ();
 FILLCELL_X32 FILLER_163_801 ();
 FILLCELL_X32 FILLER_163_833 ();
 FILLCELL_X32 FILLER_163_865 ();
 FILLCELL_X32 FILLER_163_897 ();
 FILLCELL_X32 FILLER_163_929 ();
 FILLCELL_X32 FILLER_163_961 ();
 FILLCELL_X32 FILLER_163_993 ();
 FILLCELL_X32 FILLER_163_1025 ();
 FILLCELL_X32 FILLER_163_1057 ();
 FILLCELL_X32 FILLER_163_1089 ();
 FILLCELL_X32 FILLER_163_1121 ();
 FILLCELL_X32 FILLER_163_1153 ();
 FILLCELL_X32 FILLER_163_1185 ();
 FILLCELL_X32 FILLER_163_1217 ();
 FILLCELL_X8 FILLER_163_1249 ();
 FILLCELL_X4 FILLER_163_1257 ();
 FILLCELL_X2 FILLER_163_1261 ();
 FILLCELL_X32 FILLER_163_1264 ();
 FILLCELL_X2 FILLER_163_1296 ();
 FILLCELL_X1 FILLER_163_1298 ();
 FILLCELL_X16 FILLER_163_1330 ();
 FILLCELL_X8 FILLER_163_1346 ();
 FILLCELL_X4 FILLER_163_1354 ();
 FILLCELL_X1 FILLER_163_1358 ();
 FILLCELL_X2 FILLER_163_1376 ();
 FILLCELL_X1 FILLER_163_1378 ();
 FILLCELL_X16 FILLER_163_1386 ();
 FILLCELL_X32 FILLER_163_1426 ();
 FILLCELL_X2 FILLER_163_1458 ();
 FILLCELL_X4 FILLER_163_1477 ();
 FILLCELL_X32 FILLER_163_1488 ();
 FILLCELL_X2 FILLER_163_1520 ();
 FILLCELL_X4 FILLER_163_1529 ();
 FILLCELL_X1 FILLER_163_1533 ();
 FILLCELL_X16 FILLER_163_1541 ();
 FILLCELL_X32 FILLER_163_1581 ();
 FILLCELL_X32 FILLER_163_1613 ();
 FILLCELL_X32 FILLER_163_1645 ();
 FILLCELL_X32 FILLER_163_1677 ();
 FILLCELL_X32 FILLER_163_1709 ();
 FILLCELL_X32 FILLER_163_1741 ();
 FILLCELL_X32 FILLER_163_1773 ();
 FILLCELL_X32 FILLER_163_1805 ();
 FILLCELL_X32 FILLER_163_1837 ();
 FILLCELL_X32 FILLER_163_1869 ();
 FILLCELL_X32 FILLER_163_1901 ();
 FILLCELL_X32 FILLER_163_1933 ();
 FILLCELL_X32 FILLER_163_1965 ();
 FILLCELL_X32 FILLER_163_1997 ();
 FILLCELL_X32 FILLER_163_2029 ();
 FILLCELL_X32 FILLER_163_2061 ();
 FILLCELL_X32 FILLER_163_2093 ();
 FILLCELL_X32 FILLER_163_2125 ();
 FILLCELL_X32 FILLER_163_2157 ();
 FILLCELL_X32 FILLER_163_2189 ();
 FILLCELL_X32 FILLER_163_2221 ();
 FILLCELL_X32 FILLER_163_2253 ();
 FILLCELL_X32 FILLER_163_2285 ();
 FILLCELL_X32 FILLER_163_2317 ();
 FILLCELL_X32 FILLER_163_2349 ();
 FILLCELL_X32 FILLER_163_2381 ();
 FILLCELL_X32 FILLER_163_2413 ();
 FILLCELL_X32 FILLER_163_2445 ();
 FILLCELL_X32 FILLER_163_2477 ();
 FILLCELL_X16 FILLER_163_2509 ();
 FILLCELL_X1 FILLER_163_2525 ();
 FILLCELL_X32 FILLER_163_2527 ();
 FILLCELL_X32 FILLER_163_2559 ();
 FILLCELL_X8 FILLER_163_2591 ();
 FILLCELL_X2 FILLER_163_2599 ();
 FILLCELL_X1 FILLER_163_2601 ();
 FILLCELL_X32 FILLER_164_1 ();
 FILLCELL_X32 FILLER_164_33 ();
 FILLCELL_X32 FILLER_164_65 ();
 FILLCELL_X32 FILLER_164_97 ();
 FILLCELL_X32 FILLER_164_129 ();
 FILLCELL_X32 FILLER_164_161 ();
 FILLCELL_X32 FILLER_164_193 ();
 FILLCELL_X32 FILLER_164_225 ();
 FILLCELL_X32 FILLER_164_257 ();
 FILLCELL_X32 FILLER_164_289 ();
 FILLCELL_X32 FILLER_164_321 ();
 FILLCELL_X32 FILLER_164_353 ();
 FILLCELL_X32 FILLER_164_385 ();
 FILLCELL_X32 FILLER_164_417 ();
 FILLCELL_X32 FILLER_164_449 ();
 FILLCELL_X32 FILLER_164_481 ();
 FILLCELL_X32 FILLER_164_513 ();
 FILLCELL_X32 FILLER_164_545 ();
 FILLCELL_X32 FILLER_164_577 ();
 FILLCELL_X16 FILLER_164_609 ();
 FILLCELL_X4 FILLER_164_625 ();
 FILLCELL_X2 FILLER_164_629 ();
 FILLCELL_X32 FILLER_164_632 ();
 FILLCELL_X32 FILLER_164_664 ();
 FILLCELL_X32 FILLER_164_696 ();
 FILLCELL_X32 FILLER_164_728 ();
 FILLCELL_X32 FILLER_164_760 ();
 FILLCELL_X32 FILLER_164_792 ();
 FILLCELL_X32 FILLER_164_824 ();
 FILLCELL_X32 FILLER_164_856 ();
 FILLCELL_X32 FILLER_164_888 ();
 FILLCELL_X32 FILLER_164_920 ();
 FILLCELL_X32 FILLER_164_952 ();
 FILLCELL_X32 FILLER_164_984 ();
 FILLCELL_X32 FILLER_164_1016 ();
 FILLCELL_X32 FILLER_164_1048 ();
 FILLCELL_X32 FILLER_164_1080 ();
 FILLCELL_X32 FILLER_164_1112 ();
 FILLCELL_X32 FILLER_164_1144 ();
 FILLCELL_X32 FILLER_164_1176 ();
 FILLCELL_X32 FILLER_164_1208 ();
 FILLCELL_X32 FILLER_164_1240 ();
 FILLCELL_X32 FILLER_164_1272 ();
 FILLCELL_X4 FILLER_164_1304 ();
 FILLCELL_X32 FILLER_164_1315 ();
 FILLCELL_X8 FILLER_164_1347 ();
 FILLCELL_X4 FILLER_164_1355 ();
 FILLCELL_X4 FILLER_164_1366 ();
 FILLCELL_X8 FILLER_164_1387 ();
 FILLCELL_X2 FILLER_164_1395 ();
 FILLCELL_X1 FILLER_164_1397 ();
 FILLCELL_X16 FILLER_164_1429 ();
 FILLCELL_X8 FILLER_164_1445 ();
 FILLCELL_X4 FILLER_164_1453 ();
 FILLCELL_X16 FILLER_164_1464 ();
 FILLCELL_X16 FILLER_164_1514 ();
 FILLCELL_X8 FILLER_164_1530 ();
 FILLCELL_X2 FILLER_164_1538 ();
 FILLCELL_X1 FILLER_164_1540 ();
 FILLCELL_X32 FILLER_164_1572 ();
 FILLCELL_X32 FILLER_164_1604 ();
 FILLCELL_X32 FILLER_164_1636 ();
 FILLCELL_X32 FILLER_164_1668 ();
 FILLCELL_X32 FILLER_164_1700 ();
 FILLCELL_X32 FILLER_164_1732 ();
 FILLCELL_X32 FILLER_164_1764 ();
 FILLCELL_X32 FILLER_164_1796 ();
 FILLCELL_X32 FILLER_164_1828 ();
 FILLCELL_X32 FILLER_164_1860 ();
 FILLCELL_X2 FILLER_164_1892 ();
 FILLCELL_X32 FILLER_164_1895 ();
 FILLCELL_X32 FILLER_164_1927 ();
 FILLCELL_X32 FILLER_164_1959 ();
 FILLCELL_X32 FILLER_164_1991 ();
 FILLCELL_X32 FILLER_164_2023 ();
 FILLCELL_X32 FILLER_164_2055 ();
 FILLCELL_X32 FILLER_164_2087 ();
 FILLCELL_X32 FILLER_164_2119 ();
 FILLCELL_X32 FILLER_164_2151 ();
 FILLCELL_X32 FILLER_164_2183 ();
 FILLCELL_X32 FILLER_164_2215 ();
 FILLCELL_X32 FILLER_164_2247 ();
 FILLCELL_X32 FILLER_164_2279 ();
 FILLCELL_X32 FILLER_164_2311 ();
 FILLCELL_X32 FILLER_164_2343 ();
 FILLCELL_X32 FILLER_164_2375 ();
 FILLCELL_X32 FILLER_164_2407 ();
 FILLCELL_X32 FILLER_164_2439 ();
 FILLCELL_X32 FILLER_164_2471 ();
 FILLCELL_X32 FILLER_164_2503 ();
 FILLCELL_X32 FILLER_164_2535 ();
 FILLCELL_X32 FILLER_164_2567 ();
 FILLCELL_X2 FILLER_164_2599 ();
 FILLCELL_X1 FILLER_164_2601 ();
 FILLCELL_X32 FILLER_165_1 ();
 FILLCELL_X32 FILLER_165_33 ();
 FILLCELL_X32 FILLER_165_65 ();
 FILLCELL_X32 FILLER_165_97 ();
 FILLCELL_X32 FILLER_165_129 ();
 FILLCELL_X32 FILLER_165_161 ();
 FILLCELL_X32 FILLER_165_193 ();
 FILLCELL_X32 FILLER_165_225 ();
 FILLCELL_X32 FILLER_165_257 ();
 FILLCELL_X32 FILLER_165_289 ();
 FILLCELL_X32 FILLER_165_321 ();
 FILLCELL_X32 FILLER_165_353 ();
 FILLCELL_X32 FILLER_165_385 ();
 FILLCELL_X32 FILLER_165_417 ();
 FILLCELL_X32 FILLER_165_449 ();
 FILLCELL_X32 FILLER_165_481 ();
 FILLCELL_X32 FILLER_165_513 ();
 FILLCELL_X32 FILLER_165_545 ();
 FILLCELL_X32 FILLER_165_577 ();
 FILLCELL_X32 FILLER_165_609 ();
 FILLCELL_X32 FILLER_165_641 ();
 FILLCELL_X32 FILLER_165_673 ();
 FILLCELL_X32 FILLER_165_705 ();
 FILLCELL_X32 FILLER_165_737 ();
 FILLCELL_X32 FILLER_165_769 ();
 FILLCELL_X32 FILLER_165_801 ();
 FILLCELL_X32 FILLER_165_833 ();
 FILLCELL_X32 FILLER_165_865 ();
 FILLCELL_X32 FILLER_165_897 ();
 FILLCELL_X32 FILLER_165_929 ();
 FILLCELL_X32 FILLER_165_961 ();
 FILLCELL_X32 FILLER_165_993 ();
 FILLCELL_X32 FILLER_165_1025 ();
 FILLCELL_X32 FILLER_165_1057 ();
 FILLCELL_X32 FILLER_165_1089 ();
 FILLCELL_X32 FILLER_165_1121 ();
 FILLCELL_X32 FILLER_165_1153 ();
 FILLCELL_X32 FILLER_165_1185 ();
 FILLCELL_X32 FILLER_165_1217 ();
 FILLCELL_X8 FILLER_165_1249 ();
 FILLCELL_X4 FILLER_165_1257 ();
 FILLCELL_X2 FILLER_165_1261 ();
 FILLCELL_X32 FILLER_165_1264 ();
 FILLCELL_X32 FILLER_165_1296 ();
 FILLCELL_X32 FILLER_165_1328 ();
 FILLCELL_X16 FILLER_165_1360 ();
 FILLCELL_X32 FILLER_165_1383 ();
 FILLCELL_X32 FILLER_165_1415 ();
 FILLCELL_X4 FILLER_165_1447 ();
 FILLCELL_X2 FILLER_165_1451 ();
 FILLCELL_X1 FILLER_165_1470 ();
 FILLCELL_X16 FILLER_165_1478 ();
 FILLCELL_X8 FILLER_165_1501 ();
 FILLCELL_X2 FILLER_165_1509 ();
 FILLCELL_X32 FILLER_165_1518 ();
 FILLCELL_X32 FILLER_165_1550 ();
 FILLCELL_X32 FILLER_165_1582 ();
 FILLCELL_X32 FILLER_165_1614 ();
 FILLCELL_X32 FILLER_165_1646 ();
 FILLCELL_X32 FILLER_165_1678 ();
 FILLCELL_X32 FILLER_165_1710 ();
 FILLCELL_X32 FILLER_165_1742 ();
 FILLCELL_X32 FILLER_165_1774 ();
 FILLCELL_X32 FILLER_165_1806 ();
 FILLCELL_X32 FILLER_165_1838 ();
 FILLCELL_X32 FILLER_165_1870 ();
 FILLCELL_X32 FILLER_165_1902 ();
 FILLCELL_X32 FILLER_165_1934 ();
 FILLCELL_X32 FILLER_165_1966 ();
 FILLCELL_X32 FILLER_165_1998 ();
 FILLCELL_X32 FILLER_165_2030 ();
 FILLCELL_X32 FILLER_165_2062 ();
 FILLCELL_X32 FILLER_165_2094 ();
 FILLCELL_X32 FILLER_165_2126 ();
 FILLCELL_X32 FILLER_165_2158 ();
 FILLCELL_X32 FILLER_165_2190 ();
 FILLCELL_X32 FILLER_165_2222 ();
 FILLCELL_X32 FILLER_165_2254 ();
 FILLCELL_X32 FILLER_165_2286 ();
 FILLCELL_X32 FILLER_165_2318 ();
 FILLCELL_X32 FILLER_165_2350 ();
 FILLCELL_X32 FILLER_165_2382 ();
 FILLCELL_X32 FILLER_165_2414 ();
 FILLCELL_X32 FILLER_165_2446 ();
 FILLCELL_X32 FILLER_165_2478 ();
 FILLCELL_X16 FILLER_165_2510 ();
 FILLCELL_X32 FILLER_165_2527 ();
 FILLCELL_X32 FILLER_165_2559 ();
 FILLCELL_X8 FILLER_165_2591 ();
 FILLCELL_X2 FILLER_165_2599 ();
 FILLCELL_X1 FILLER_165_2601 ();
 FILLCELL_X4 FILLER_166_1 ();
 FILLCELL_X2 FILLER_166_5 ();
 FILLCELL_X1 FILLER_166_7 ();
 FILLCELL_X32 FILLER_166_11 ();
 FILLCELL_X32 FILLER_166_43 ();
 FILLCELL_X32 FILLER_166_75 ();
 FILLCELL_X32 FILLER_166_107 ();
 FILLCELL_X32 FILLER_166_139 ();
 FILLCELL_X32 FILLER_166_171 ();
 FILLCELL_X32 FILLER_166_203 ();
 FILLCELL_X32 FILLER_166_235 ();
 FILLCELL_X32 FILLER_166_267 ();
 FILLCELL_X32 FILLER_166_299 ();
 FILLCELL_X32 FILLER_166_331 ();
 FILLCELL_X32 FILLER_166_363 ();
 FILLCELL_X32 FILLER_166_395 ();
 FILLCELL_X32 FILLER_166_427 ();
 FILLCELL_X32 FILLER_166_459 ();
 FILLCELL_X32 FILLER_166_491 ();
 FILLCELL_X32 FILLER_166_523 ();
 FILLCELL_X32 FILLER_166_555 ();
 FILLCELL_X32 FILLER_166_587 ();
 FILLCELL_X8 FILLER_166_619 ();
 FILLCELL_X4 FILLER_166_627 ();
 FILLCELL_X32 FILLER_166_632 ();
 FILLCELL_X32 FILLER_166_664 ();
 FILLCELL_X32 FILLER_166_696 ();
 FILLCELL_X32 FILLER_166_728 ();
 FILLCELL_X32 FILLER_166_760 ();
 FILLCELL_X32 FILLER_166_792 ();
 FILLCELL_X32 FILLER_166_824 ();
 FILLCELL_X32 FILLER_166_856 ();
 FILLCELL_X32 FILLER_166_888 ();
 FILLCELL_X32 FILLER_166_920 ();
 FILLCELL_X32 FILLER_166_952 ();
 FILLCELL_X32 FILLER_166_984 ();
 FILLCELL_X32 FILLER_166_1016 ();
 FILLCELL_X32 FILLER_166_1048 ();
 FILLCELL_X32 FILLER_166_1080 ();
 FILLCELL_X16 FILLER_166_1112 ();
 FILLCELL_X8 FILLER_166_1128 ();
 FILLCELL_X4 FILLER_166_1136 ();
 FILLCELL_X32 FILLER_166_1147 ();
 FILLCELL_X32 FILLER_166_1179 ();
 FILLCELL_X32 FILLER_166_1211 ();
 FILLCELL_X16 FILLER_166_1243 ();
 FILLCELL_X8 FILLER_166_1259 ();
 FILLCELL_X1 FILLER_166_1267 ();
 FILLCELL_X32 FILLER_166_1292 ();
 FILLCELL_X32 FILLER_166_1324 ();
 FILLCELL_X32 FILLER_166_1356 ();
 FILLCELL_X32 FILLER_166_1388 ();
 FILLCELL_X32 FILLER_166_1420 ();
 FILLCELL_X1 FILLER_166_1452 ();
 FILLCELL_X16 FILLER_166_1460 ();
 FILLCELL_X8 FILLER_166_1476 ();
 FILLCELL_X4 FILLER_166_1484 ();
 FILLCELL_X2 FILLER_166_1488 ();
 FILLCELL_X1 FILLER_166_1490 ();
 FILLCELL_X1 FILLER_166_1498 ();
 FILLCELL_X16 FILLER_166_1506 ();
 FILLCELL_X2 FILLER_166_1522 ();
 FILLCELL_X16 FILLER_166_1531 ();
 FILLCELL_X4 FILLER_166_1547 ();
 FILLCELL_X2 FILLER_166_1551 ();
 FILLCELL_X32 FILLER_166_1560 ();
 FILLCELL_X32 FILLER_166_1592 ();
 FILLCELL_X32 FILLER_166_1624 ();
 FILLCELL_X32 FILLER_166_1656 ();
 FILLCELL_X32 FILLER_166_1688 ();
 FILLCELL_X32 FILLER_166_1720 ();
 FILLCELL_X32 FILLER_166_1752 ();
 FILLCELL_X32 FILLER_166_1784 ();
 FILLCELL_X32 FILLER_166_1816 ();
 FILLCELL_X32 FILLER_166_1848 ();
 FILLCELL_X8 FILLER_166_1880 ();
 FILLCELL_X4 FILLER_166_1888 ();
 FILLCELL_X2 FILLER_166_1892 ();
 FILLCELL_X32 FILLER_166_1895 ();
 FILLCELL_X32 FILLER_166_1927 ();
 FILLCELL_X32 FILLER_166_1959 ();
 FILLCELL_X32 FILLER_166_1991 ();
 FILLCELL_X32 FILLER_166_2023 ();
 FILLCELL_X32 FILLER_166_2055 ();
 FILLCELL_X32 FILLER_166_2087 ();
 FILLCELL_X32 FILLER_166_2119 ();
 FILLCELL_X32 FILLER_166_2151 ();
 FILLCELL_X32 FILLER_166_2183 ();
 FILLCELL_X32 FILLER_166_2215 ();
 FILLCELL_X32 FILLER_166_2247 ();
 FILLCELL_X32 FILLER_166_2279 ();
 FILLCELL_X32 FILLER_166_2311 ();
 FILLCELL_X32 FILLER_166_2343 ();
 FILLCELL_X32 FILLER_166_2375 ();
 FILLCELL_X32 FILLER_166_2407 ();
 FILLCELL_X32 FILLER_166_2439 ();
 FILLCELL_X32 FILLER_166_2471 ();
 FILLCELL_X32 FILLER_166_2503 ();
 FILLCELL_X32 FILLER_166_2535 ();
 FILLCELL_X32 FILLER_166_2567 ();
 FILLCELL_X2 FILLER_166_2599 ();
 FILLCELL_X1 FILLER_166_2601 ();
 FILLCELL_X4 FILLER_167_1 ();
 FILLCELL_X32 FILLER_167_8 ();
 FILLCELL_X32 FILLER_167_40 ();
 FILLCELL_X32 FILLER_167_72 ();
 FILLCELL_X32 FILLER_167_104 ();
 FILLCELL_X32 FILLER_167_136 ();
 FILLCELL_X32 FILLER_167_168 ();
 FILLCELL_X32 FILLER_167_200 ();
 FILLCELL_X32 FILLER_167_232 ();
 FILLCELL_X32 FILLER_167_264 ();
 FILLCELL_X32 FILLER_167_296 ();
 FILLCELL_X32 FILLER_167_328 ();
 FILLCELL_X32 FILLER_167_360 ();
 FILLCELL_X32 FILLER_167_392 ();
 FILLCELL_X32 FILLER_167_424 ();
 FILLCELL_X32 FILLER_167_456 ();
 FILLCELL_X32 FILLER_167_488 ();
 FILLCELL_X32 FILLER_167_520 ();
 FILLCELL_X32 FILLER_167_552 ();
 FILLCELL_X32 FILLER_167_584 ();
 FILLCELL_X32 FILLER_167_616 ();
 FILLCELL_X32 FILLER_167_648 ();
 FILLCELL_X32 FILLER_167_680 ();
 FILLCELL_X32 FILLER_167_712 ();
 FILLCELL_X32 FILLER_167_744 ();
 FILLCELL_X32 FILLER_167_776 ();
 FILLCELL_X32 FILLER_167_808 ();
 FILLCELL_X32 FILLER_167_840 ();
 FILLCELL_X32 FILLER_167_872 ();
 FILLCELL_X32 FILLER_167_904 ();
 FILLCELL_X32 FILLER_167_936 ();
 FILLCELL_X32 FILLER_167_968 ();
 FILLCELL_X32 FILLER_167_1000 ();
 FILLCELL_X32 FILLER_167_1032 ();
 FILLCELL_X32 FILLER_167_1064 ();
 FILLCELL_X32 FILLER_167_1096 ();
 FILLCELL_X4 FILLER_167_1128 ();
 FILLCELL_X2 FILLER_167_1132 ();
 FILLCELL_X32 FILLER_167_1151 ();
 FILLCELL_X32 FILLER_167_1183 ();
 FILLCELL_X32 FILLER_167_1215 ();
 FILLCELL_X16 FILLER_167_1247 ();
 FILLCELL_X4 FILLER_167_1264 ();
 FILLCELL_X2 FILLER_167_1268 ();
 FILLCELL_X1 FILLER_167_1270 ();
 FILLCELL_X4 FILLER_167_1278 ();
 FILLCELL_X2 FILLER_167_1282 ();
 FILLCELL_X8 FILLER_167_1308 ();
 FILLCELL_X4 FILLER_167_1316 ();
 FILLCELL_X2 FILLER_167_1320 ();
 FILLCELL_X16 FILLER_167_1346 ();
 FILLCELL_X4 FILLER_167_1362 ();
 FILLCELL_X1 FILLER_167_1366 ();
 FILLCELL_X32 FILLER_167_1374 ();
 FILLCELL_X32 FILLER_167_1406 ();
 FILLCELL_X32 FILLER_167_1438 ();
 FILLCELL_X16 FILLER_167_1470 ();
 FILLCELL_X1 FILLER_167_1486 ();
 FILLCELL_X16 FILLER_167_1504 ();
 FILLCELL_X8 FILLER_167_1520 ();
 FILLCELL_X4 FILLER_167_1528 ();
 FILLCELL_X1 FILLER_167_1532 ();
 FILLCELL_X2 FILLER_167_1540 ();
 FILLCELL_X1 FILLER_167_1542 ();
 FILLCELL_X32 FILLER_167_1567 ();
 FILLCELL_X32 FILLER_167_1599 ();
 FILLCELL_X32 FILLER_167_1631 ();
 FILLCELL_X32 FILLER_167_1663 ();
 FILLCELL_X32 FILLER_167_1695 ();
 FILLCELL_X32 FILLER_167_1727 ();
 FILLCELL_X32 FILLER_167_1759 ();
 FILLCELL_X32 FILLER_167_1791 ();
 FILLCELL_X32 FILLER_167_1823 ();
 FILLCELL_X32 FILLER_167_1855 ();
 FILLCELL_X32 FILLER_167_1887 ();
 FILLCELL_X32 FILLER_167_1919 ();
 FILLCELL_X32 FILLER_167_1951 ();
 FILLCELL_X32 FILLER_167_1983 ();
 FILLCELL_X32 FILLER_167_2015 ();
 FILLCELL_X32 FILLER_167_2047 ();
 FILLCELL_X32 FILLER_167_2079 ();
 FILLCELL_X32 FILLER_167_2111 ();
 FILLCELL_X32 FILLER_167_2143 ();
 FILLCELL_X32 FILLER_167_2175 ();
 FILLCELL_X32 FILLER_167_2207 ();
 FILLCELL_X32 FILLER_167_2239 ();
 FILLCELL_X32 FILLER_167_2271 ();
 FILLCELL_X32 FILLER_167_2303 ();
 FILLCELL_X32 FILLER_167_2335 ();
 FILLCELL_X32 FILLER_167_2367 ();
 FILLCELL_X32 FILLER_167_2399 ();
 FILLCELL_X32 FILLER_167_2431 ();
 FILLCELL_X32 FILLER_167_2463 ();
 FILLCELL_X16 FILLER_167_2495 ();
 FILLCELL_X8 FILLER_167_2511 ();
 FILLCELL_X4 FILLER_167_2519 ();
 FILLCELL_X2 FILLER_167_2523 ();
 FILLCELL_X1 FILLER_167_2525 ();
 FILLCELL_X32 FILLER_167_2527 ();
 FILLCELL_X32 FILLER_167_2559 ();
 FILLCELL_X8 FILLER_167_2591 ();
 FILLCELL_X2 FILLER_167_2599 ();
 FILLCELL_X1 FILLER_167_2601 ();
 FILLCELL_X1 FILLER_168_1 ();
 FILLCELL_X1 FILLER_168_8 ();
 FILLCELL_X2 FILLER_168_12 ();
 FILLCELL_X1 FILLER_168_14 ();
 FILLCELL_X32 FILLER_168_18 ();
 FILLCELL_X32 FILLER_168_50 ();
 FILLCELL_X32 FILLER_168_82 ();
 FILLCELL_X32 FILLER_168_114 ();
 FILLCELL_X32 FILLER_168_146 ();
 FILLCELL_X32 FILLER_168_178 ();
 FILLCELL_X32 FILLER_168_210 ();
 FILLCELL_X32 FILLER_168_242 ();
 FILLCELL_X32 FILLER_168_274 ();
 FILLCELL_X32 FILLER_168_306 ();
 FILLCELL_X32 FILLER_168_338 ();
 FILLCELL_X32 FILLER_168_370 ();
 FILLCELL_X32 FILLER_168_402 ();
 FILLCELL_X32 FILLER_168_434 ();
 FILLCELL_X32 FILLER_168_466 ();
 FILLCELL_X32 FILLER_168_498 ();
 FILLCELL_X32 FILLER_168_530 ();
 FILLCELL_X32 FILLER_168_562 ();
 FILLCELL_X32 FILLER_168_594 ();
 FILLCELL_X4 FILLER_168_626 ();
 FILLCELL_X1 FILLER_168_630 ();
 FILLCELL_X32 FILLER_168_632 ();
 FILLCELL_X32 FILLER_168_664 ();
 FILLCELL_X32 FILLER_168_696 ();
 FILLCELL_X32 FILLER_168_728 ();
 FILLCELL_X32 FILLER_168_760 ();
 FILLCELL_X32 FILLER_168_792 ();
 FILLCELL_X32 FILLER_168_824 ();
 FILLCELL_X32 FILLER_168_856 ();
 FILLCELL_X32 FILLER_168_888 ();
 FILLCELL_X32 FILLER_168_920 ();
 FILLCELL_X32 FILLER_168_952 ();
 FILLCELL_X32 FILLER_168_984 ();
 FILLCELL_X32 FILLER_168_1016 ();
 FILLCELL_X16 FILLER_168_1048 ();
 FILLCELL_X8 FILLER_168_1064 ();
 FILLCELL_X4 FILLER_168_1072 ();
 FILLCELL_X1 FILLER_168_1076 ();
 FILLCELL_X32 FILLER_168_1093 ();
 FILLCELL_X8 FILLER_168_1125 ();
 FILLCELL_X4 FILLER_168_1133 ();
 FILLCELL_X1 FILLER_168_1141 ();
 FILLCELL_X32 FILLER_168_1145 ();
 FILLCELL_X16 FILLER_168_1177 ();
 FILLCELL_X8 FILLER_168_1193 ();
 FILLCELL_X1 FILLER_168_1201 ();
 FILLCELL_X1 FILLER_168_1212 ();
 FILLCELL_X32 FILLER_168_1232 ();
 FILLCELL_X4 FILLER_168_1264 ();
 FILLCELL_X2 FILLER_168_1268 ();
 FILLCELL_X1 FILLER_168_1270 ();
 FILLCELL_X4 FILLER_168_1288 ();
 FILLCELL_X2 FILLER_168_1292 ();
 FILLCELL_X16 FILLER_168_1301 ();
 FILLCELL_X8 FILLER_168_1317 ();
 FILLCELL_X4 FILLER_168_1325 ();
 FILLCELL_X2 FILLER_168_1329 ();
 FILLCELL_X1 FILLER_168_1331 ();
 FILLCELL_X2 FILLER_168_1353 ();
 FILLCELL_X16 FILLER_168_1386 ();
 FILLCELL_X32 FILLER_168_1426 ();
 FILLCELL_X32 FILLER_168_1458 ();
 FILLCELL_X32 FILLER_168_1490 ();
 FILLCELL_X8 FILLER_168_1522 ();
 FILLCELL_X4 FILLER_168_1547 ();
 FILLCELL_X2 FILLER_168_1551 ();
 FILLCELL_X32 FILLER_168_1560 ();
 FILLCELL_X32 FILLER_168_1592 ();
 FILLCELL_X32 FILLER_168_1624 ();
 FILLCELL_X32 FILLER_168_1656 ();
 FILLCELL_X32 FILLER_168_1688 ();
 FILLCELL_X32 FILLER_168_1720 ();
 FILLCELL_X32 FILLER_168_1752 ();
 FILLCELL_X32 FILLER_168_1784 ();
 FILLCELL_X32 FILLER_168_1816 ();
 FILLCELL_X32 FILLER_168_1848 ();
 FILLCELL_X8 FILLER_168_1880 ();
 FILLCELL_X4 FILLER_168_1888 ();
 FILLCELL_X2 FILLER_168_1892 ();
 FILLCELL_X32 FILLER_168_1895 ();
 FILLCELL_X32 FILLER_168_1927 ();
 FILLCELL_X32 FILLER_168_1959 ();
 FILLCELL_X32 FILLER_168_1991 ();
 FILLCELL_X32 FILLER_168_2023 ();
 FILLCELL_X32 FILLER_168_2055 ();
 FILLCELL_X32 FILLER_168_2087 ();
 FILLCELL_X32 FILLER_168_2119 ();
 FILLCELL_X32 FILLER_168_2151 ();
 FILLCELL_X32 FILLER_168_2183 ();
 FILLCELL_X32 FILLER_168_2215 ();
 FILLCELL_X32 FILLER_168_2247 ();
 FILLCELL_X32 FILLER_168_2279 ();
 FILLCELL_X32 FILLER_168_2311 ();
 FILLCELL_X32 FILLER_168_2343 ();
 FILLCELL_X32 FILLER_168_2375 ();
 FILLCELL_X32 FILLER_168_2407 ();
 FILLCELL_X32 FILLER_168_2439 ();
 FILLCELL_X32 FILLER_168_2471 ();
 FILLCELL_X32 FILLER_168_2503 ();
 FILLCELL_X32 FILLER_168_2535 ();
 FILLCELL_X32 FILLER_168_2567 ();
 FILLCELL_X2 FILLER_168_2599 ();
 FILLCELL_X1 FILLER_168_2601 ();
 FILLCELL_X16 FILLER_169_1 ();
 FILLCELL_X32 FILLER_169_22 ();
 FILLCELL_X32 FILLER_169_54 ();
 FILLCELL_X32 FILLER_169_86 ();
 FILLCELL_X32 FILLER_169_118 ();
 FILLCELL_X32 FILLER_169_150 ();
 FILLCELL_X32 FILLER_169_182 ();
 FILLCELL_X32 FILLER_169_214 ();
 FILLCELL_X32 FILLER_169_246 ();
 FILLCELL_X32 FILLER_169_278 ();
 FILLCELL_X32 FILLER_169_310 ();
 FILLCELL_X32 FILLER_169_342 ();
 FILLCELL_X32 FILLER_169_374 ();
 FILLCELL_X32 FILLER_169_406 ();
 FILLCELL_X32 FILLER_169_438 ();
 FILLCELL_X32 FILLER_169_470 ();
 FILLCELL_X32 FILLER_169_502 ();
 FILLCELL_X32 FILLER_169_534 ();
 FILLCELL_X32 FILLER_169_566 ();
 FILLCELL_X32 FILLER_169_598 ();
 FILLCELL_X32 FILLER_169_630 ();
 FILLCELL_X32 FILLER_169_662 ();
 FILLCELL_X32 FILLER_169_694 ();
 FILLCELL_X32 FILLER_169_726 ();
 FILLCELL_X32 FILLER_169_758 ();
 FILLCELL_X32 FILLER_169_790 ();
 FILLCELL_X32 FILLER_169_822 ();
 FILLCELL_X32 FILLER_169_854 ();
 FILLCELL_X32 FILLER_169_886 ();
 FILLCELL_X32 FILLER_169_918 ();
 FILLCELL_X32 FILLER_169_950 ();
 FILLCELL_X32 FILLER_169_982 ();
 FILLCELL_X32 FILLER_169_1014 ();
 FILLCELL_X8 FILLER_169_1046 ();
 FILLCELL_X2 FILLER_169_1054 ();
 FILLCELL_X4 FILLER_169_1065 ();
 FILLCELL_X2 FILLER_169_1069 ();
 FILLCELL_X1 FILLER_169_1071 ();
 FILLCELL_X2 FILLER_169_1082 ();
 FILLCELL_X1 FILLER_169_1094 ();
 FILLCELL_X32 FILLER_169_1115 ();
 FILLCELL_X4 FILLER_169_1147 ();
 FILLCELL_X1 FILLER_169_1151 ();
 FILLCELL_X8 FILLER_169_1161 ();
 FILLCELL_X2 FILLER_169_1169 ();
 FILLCELL_X1 FILLER_169_1171 ();
 FILLCELL_X8 FILLER_169_1191 ();
 FILLCELL_X4 FILLER_169_1199 ();
 FILLCELL_X2 FILLER_169_1210 ();
 FILLCELL_X1 FILLER_169_1215 ();
 FILLCELL_X32 FILLER_169_1229 ();
 FILLCELL_X2 FILLER_169_1261 ();
 FILLCELL_X16 FILLER_169_1264 ();
 FILLCELL_X8 FILLER_169_1280 ();
 FILLCELL_X4 FILLER_169_1288 ();
 FILLCELL_X2 FILLER_169_1292 ();
 FILLCELL_X1 FILLER_169_1294 ();
 FILLCELL_X8 FILLER_169_1316 ();
 FILLCELL_X4 FILLER_169_1324 ();
 FILLCELL_X16 FILLER_169_1345 ();
 FILLCELL_X2 FILLER_169_1361 ();
 FILLCELL_X1 FILLER_169_1363 ();
 FILLCELL_X16 FILLER_169_1381 ();
 FILLCELL_X1 FILLER_169_1397 ();
 FILLCELL_X1 FILLER_169_1422 ();
 FILLCELL_X8 FILLER_169_1430 ();
 FILLCELL_X2 FILLER_169_1438 ();
 FILLCELL_X8 FILLER_169_1464 ();
 FILLCELL_X4 FILLER_169_1472 ();
 FILLCELL_X2 FILLER_169_1476 ();
 FILLCELL_X8 FILLER_169_1485 ();
 FILLCELL_X4 FILLER_169_1493 ();
 FILLCELL_X1 FILLER_169_1497 ();
 FILLCELL_X8 FILLER_169_1505 ();
 FILLCELL_X4 FILLER_169_1513 ();
 FILLCELL_X2 FILLER_169_1517 ();
 FILLCELL_X32 FILLER_169_1524 ();
 FILLCELL_X32 FILLER_169_1556 ();
 FILLCELL_X32 FILLER_169_1588 ();
 FILLCELL_X32 FILLER_169_1620 ();
 FILLCELL_X32 FILLER_169_1652 ();
 FILLCELL_X32 FILLER_169_1684 ();
 FILLCELL_X32 FILLER_169_1716 ();
 FILLCELL_X32 FILLER_169_1748 ();
 FILLCELL_X32 FILLER_169_1780 ();
 FILLCELL_X32 FILLER_169_1812 ();
 FILLCELL_X32 FILLER_169_1844 ();
 FILLCELL_X32 FILLER_169_1876 ();
 FILLCELL_X32 FILLER_169_1908 ();
 FILLCELL_X32 FILLER_169_1940 ();
 FILLCELL_X32 FILLER_169_1972 ();
 FILLCELL_X32 FILLER_169_2004 ();
 FILLCELL_X32 FILLER_169_2036 ();
 FILLCELL_X32 FILLER_169_2068 ();
 FILLCELL_X32 FILLER_169_2100 ();
 FILLCELL_X32 FILLER_169_2132 ();
 FILLCELL_X32 FILLER_169_2164 ();
 FILLCELL_X32 FILLER_169_2196 ();
 FILLCELL_X32 FILLER_169_2228 ();
 FILLCELL_X32 FILLER_169_2260 ();
 FILLCELL_X32 FILLER_169_2292 ();
 FILLCELL_X32 FILLER_169_2324 ();
 FILLCELL_X32 FILLER_169_2356 ();
 FILLCELL_X32 FILLER_169_2388 ();
 FILLCELL_X32 FILLER_169_2420 ();
 FILLCELL_X32 FILLER_169_2452 ();
 FILLCELL_X32 FILLER_169_2484 ();
 FILLCELL_X8 FILLER_169_2516 ();
 FILLCELL_X2 FILLER_169_2524 ();
 FILLCELL_X32 FILLER_169_2527 ();
 FILLCELL_X32 FILLER_169_2559 ();
 FILLCELL_X8 FILLER_169_2591 ();
 FILLCELL_X2 FILLER_169_2599 ();
 FILLCELL_X1 FILLER_169_2601 ();
 FILLCELL_X32 FILLER_170_1 ();
 FILLCELL_X32 FILLER_170_33 ();
 FILLCELL_X32 FILLER_170_65 ();
 FILLCELL_X32 FILLER_170_97 ();
 FILLCELL_X32 FILLER_170_129 ();
 FILLCELL_X32 FILLER_170_161 ();
 FILLCELL_X32 FILLER_170_193 ();
 FILLCELL_X32 FILLER_170_225 ();
 FILLCELL_X32 FILLER_170_257 ();
 FILLCELL_X32 FILLER_170_289 ();
 FILLCELL_X32 FILLER_170_321 ();
 FILLCELL_X32 FILLER_170_353 ();
 FILLCELL_X32 FILLER_170_385 ();
 FILLCELL_X32 FILLER_170_417 ();
 FILLCELL_X32 FILLER_170_449 ();
 FILLCELL_X32 FILLER_170_481 ();
 FILLCELL_X32 FILLER_170_513 ();
 FILLCELL_X32 FILLER_170_545 ();
 FILLCELL_X32 FILLER_170_577 ();
 FILLCELL_X16 FILLER_170_609 ();
 FILLCELL_X4 FILLER_170_625 ();
 FILLCELL_X2 FILLER_170_629 ();
 FILLCELL_X32 FILLER_170_632 ();
 FILLCELL_X32 FILLER_170_664 ();
 FILLCELL_X32 FILLER_170_696 ();
 FILLCELL_X32 FILLER_170_728 ();
 FILLCELL_X32 FILLER_170_760 ();
 FILLCELL_X32 FILLER_170_792 ();
 FILLCELL_X32 FILLER_170_824 ();
 FILLCELL_X32 FILLER_170_856 ();
 FILLCELL_X32 FILLER_170_888 ();
 FILLCELL_X32 FILLER_170_920 ();
 FILLCELL_X32 FILLER_170_952 ();
 FILLCELL_X32 FILLER_170_984 ();
 FILLCELL_X32 FILLER_170_1016 ();
 FILLCELL_X16 FILLER_170_1048 ();
 FILLCELL_X8 FILLER_170_1064 ();
 FILLCELL_X4 FILLER_170_1072 ();
 FILLCELL_X2 FILLER_170_1092 ();
 FILLCELL_X1 FILLER_170_1094 ();
 FILLCELL_X16 FILLER_170_1105 ();
 FILLCELL_X8 FILLER_170_1121 ();
 FILLCELL_X2 FILLER_170_1129 ();
 FILLCELL_X2 FILLER_170_1134 ();
 FILLCELL_X1 FILLER_170_1136 ();
 FILLCELL_X1 FILLER_170_1141 ();
 FILLCELL_X4 FILLER_170_1149 ();
 FILLCELL_X1 FILLER_170_1153 ();
 FILLCELL_X8 FILLER_170_1164 ();
 FILLCELL_X1 FILLER_170_1172 ();
 FILLCELL_X4 FILLER_170_1183 ();
 FILLCELL_X1 FILLER_170_1187 ();
 FILLCELL_X8 FILLER_170_1191 ();
 FILLCELL_X1 FILLER_170_1199 ();
 FILLCELL_X4 FILLER_170_1208 ();
 FILLCELL_X2 FILLER_170_1212 ();
 FILLCELL_X4 FILLER_170_1219 ();
 FILLCELL_X2 FILLER_170_1223 ();
 FILLCELL_X1 FILLER_170_1225 ();
 FILLCELL_X8 FILLER_170_1239 ();
 FILLCELL_X4 FILLER_170_1247 ();
 FILLCELL_X16 FILLER_170_1267 ();
 FILLCELL_X8 FILLER_170_1283 ();
 FILLCELL_X32 FILLER_170_1308 ();
 FILLCELL_X32 FILLER_170_1340 ();
 FILLCELL_X4 FILLER_170_1372 ();
 FILLCELL_X1 FILLER_170_1376 ();
 FILLCELL_X16 FILLER_170_1384 ();
 FILLCELL_X2 FILLER_170_1400 ();
 FILLCELL_X1 FILLER_170_1402 ();
 FILLCELL_X16 FILLER_170_1410 ();
 FILLCELL_X2 FILLER_170_1426 ();
 FILLCELL_X1 FILLER_170_1428 ();
 FILLCELL_X1 FILLER_170_1453 ();
 FILLCELL_X8 FILLER_170_1461 ();
 FILLCELL_X2 FILLER_170_1469 ();
 FILLCELL_X1 FILLER_170_1478 ();
 FILLCELL_X1 FILLER_170_1496 ();
 FILLCELL_X16 FILLER_170_1521 ();
 FILLCELL_X8 FILLER_170_1537 ();
 FILLCELL_X2 FILLER_170_1545 ();
 FILLCELL_X1 FILLER_170_1547 ();
 FILLCELL_X32 FILLER_170_1555 ();
 FILLCELL_X32 FILLER_170_1587 ();
 FILLCELL_X32 FILLER_170_1619 ();
 FILLCELL_X32 FILLER_170_1651 ();
 FILLCELL_X32 FILLER_170_1683 ();
 FILLCELL_X32 FILLER_170_1715 ();
 FILLCELL_X32 FILLER_170_1747 ();
 FILLCELL_X32 FILLER_170_1779 ();
 FILLCELL_X32 FILLER_170_1811 ();
 FILLCELL_X32 FILLER_170_1843 ();
 FILLCELL_X16 FILLER_170_1875 ();
 FILLCELL_X2 FILLER_170_1891 ();
 FILLCELL_X1 FILLER_170_1893 ();
 FILLCELL_X32 FILLER_170_1895 ();
 FILLCELL_X32 FILLER_170_1927 ();
 FILLCELL_X32 FILLER_170_1959 ();
 FILLCELL_X32 FILLER_170_1991 ();
 FILLCELL_X32 FILLER_170_2023 ();
 FILLCELL_X32 FILLER_170_2055 ();
 FILLCELL_X32 FILLER_170_2087 ();
 FILLCELL_X32 FILLER_170_2119 ();
 FILLCELL_X32 FILLER_170_2151 ();
 FILLCELL_X32 FILLER_170_2183 ();
 FILLCELL_X32 FILLER_170_2215 ();
 FILLCELL_X32 FILLER_170_2247 ();
 FILLCELL_X32 FILLER_170_2279 ();
 FILLCELL_X32 FILLER_170_2311 ();
 FILLCELL_X32 FILLER_170_2343 ();
 FILLCELL_X32 FILLER_170_2375 ();
 FILLCELL_X32 FILLER_170_2407 ();
 FILLCELL_X32 FILLER_170_2439 ();
 FILLCELL_X32 FILLER_170_2471 ();
 FILLCELL_X32 FILLER_170_2503 ();
 FILLCELL_X32 FILLER_170_2535 ();
 FILLCELL_X32 FILLER_170_2567 ();
 FILLCELL_X2 FILLER_170_2599 ();
 FILLCELL_X1 FILLER_170_2601 ();
 FILLCELL_X16 FILLER_171_1 ();
 FILLCELL_X4 FILLER_171_17 ();
 FILLCELL_X2 FILLER_171_21 ();
 FILLCELL_X1 FILLER_171_23 ();
 FILLCELL_X32 FILLER_171_27 ();
 FILLCELL_X32 FILLER_171_59 ();
 FILLCELL_X32 FILLER_171_91 ();
 FILLCELL_X32 FILLER_171_123 ();
 FILLCELL_X32 FILLER_171_155 ();
 FILLCELL_X32 FILLER_171_187 ();
 FILLCELL_X32 FILLER_171_219 ();
 FILLCELL_X32 FILLER_171_251 ();
 FILLCELL_X32 FILLER_171_283 ();
 FILLCELL_X32 FILLER_171_315 ();
 FILLCELL_X32 FILLER_171_347 ();
 FILLCELL_X32 FILLER_171_379 ();
 FILLCELL_X32 FILLER_171_411 ();
 FILLCELL_X32 FILLER_171_443 ();
 FILLCELL_X32 FILLER_171_475 ();
 FILLCELL_X32 FILLER_171_507 ();
 FILLCELL_X32 FILLER_171_539 ();
 FILLCELL_X32 FILLER_171_571 ();
 FILLCELL_X32 FILLER_171_603 ();
 FILLCELL_X32 FILLER_171_635 ();
 FILLCELL_X32 FILLER_171_667 ();
 FILLCELL_X32 FILLER_171_699 ();
 FILLCELL_X32 FILLER_171_731 ();
 FILLCELL_X32 FILLER_171_763 ();
 FILLCELL_X32 FILLER_171_795 ();
 FILLCELL_X32 FILLER_171_827 ();
 FILLCELL_X32 FILLER_171_859 ();
 FILLCELL_X32 FILLER_171_891 ();
 FILLCELL_X32 FILLER_171_923 ();
 FILLCELL_X32 FILLER_171_955 ();
 FILLCELL_X32 FILLER_171_987 ();
 FILLCELL_X32 FILLER_171_1019 ();
 FILLCELL_X32 FILLER_171_1051 ();
 FILLCELL_X2 FILLER_171_1083 ();
 FILLCELL_X1 FILLER_171_1085 ();
 FILLCELL_X2 FILLER_171_1096 ();
 FILLCELL_X1 FILLER_171_1098 ();
 FILLCELL_X4 FILLER_171_1126 ();
 FILLCELL_X16 FILLER_171_1151 ();
 FILLCELL_X8 FILLER_171_1167 ();
 FILLCELL_X4 FILLER_171_1184 ();
 FILLCELL_X1 FILLER_171_1188 ();
 FILLCELL_X8 FILLER_171_1199 ();
 FILLCELL_X1 FILLER_171_1207 ();
 FILLCELL_X16 FILLER_171_1228 ();
 FILLCELL_X4 FILLER_171_1244 ();
 FILLCELL_X2 FILLER_171_1248 ();
 FILLCELL_X8 FILLER_171_1253 ();
 FILLCELL_X2 FILLER_171_1261 ();
 FILLCELL_X32 FILLER_171_1277 ();
 FILLCELL_X32 FILLER_171_1309 ();
 FILLCELL_X32 FILLER_171_1341 ();
 FILLCELL_X32 FILLER_171_1373 ();
 FILLCELL_X16 FILLER_171_1405 ();
 FILLCELL_X8 FILLER_171_1421 ();
 FILLCELL_X4 FILLER_171_1429 ();
 FILLCELL_X32 FILLER_171_1438 ();
 FILLCELL_X32 FILLER_171_1470 ();
 FILLCELL_X16 FILLER_171_1502 ();
 FILLCELL_X4 FILLER_171_1518 ();
 FILLCELL_X2 FILLER_171_1522 ();
 FILLCELL_X1 FILLER_171_1531 ();
 FILLCELL_X32 FILLER_171_1537 ();
 FILLCELL_X4 FILLER_171_1569 ();
 FILLCELL_X2 FILLER_171_1573 ();
 FILLCELL_X1 FILLER_171_1575 ();
 FILLCELL_X32 FILLER_171_1583 ();
 FILLCELL_X32 FILLER_171_1615 ();
 FILLCELL_X32 FILLER_171_1647 ();
 FILLCELL_X32 FILLER_171_1679 ();
 FILLCELL_X32 FILLER_171_1711 ();
 FILLCELL_X32 FILLER_171_1743 ();
 FILLCELL_X32 FILLER_171_1775 ();
 FILLCELL_X32 FILLER_171_1807 ();
 FILLCELL_X32 FILLER_171_1839 ();
 FILLCELL_X32 FILLER_171_1871 ();
 FILLCELL_X32 FILLER_171_1903 ();
 FILLCELL_X32 FILLER_171_1935 ();
 FILLCELL_X32 FILLER_171_1967 ();
 FILLCELL_X32 FILLER_171_1999 ();
 FILLCELL_X32 FILLER_171_2031 ();
 FILLCELL_X32 FILLER_171_2063 ();
 FILLCELL_X32 FILLER_171_2095 ();
 FILLCELL_X32 FILLER_171_2127 ();
 FILLCELL_X32 FILLER_171_2159 ();
 FILLCELL_X32 FILLER_171_2191 ();
 FILLCELL_X32 FILLER_171_2223 ();
 FILLCELL_X32 FILLER_171_2255 ();
 FILLCELL_X32 FILLER_171_2287 ();
 FILLCELL_X32 FILLER_171_2319 ();
 FILLCELL_X32 FILLER_171_2351 ();
 FILLCELL_X32 FILLER_171_2383 ();
 FILLCELL_X32 FILLER_171_2415 ();
 FILLCELL_X32 FILLER_171_2447 ();
 FILLCELL_X32 FILLER_171_2479 ();
 FILLCELL_X8 FILLER_171_2511 ();
 FILLCELL_X4 FILLER_171_2519 ();
 FILLCELL_X2 FILLER_171_2523 ();
 FILLCELL_X1 FILLER_171_2525 ();
 FILLCELL_X32 FILLER_171_2527 ();
 FILLCELL_X32 FILLER_171_2559 ();
 FILLCELL_X8 FILLER_171_2591 ();
 FILLCELL_X2 FILLER_171_2599 ();
 FILLCELL_X1 FILLER_171_2601 ();
 FILLCELL_X32 FILLER_172_1 ();
 FILLCELL_X32 FILLER_172_33 ();
 FILLCELL_X32 FILLER_172_65 ();
 FILLCELL_X32 FILLER_172_97 ();
 FILLCELL_X32 FILLER_172_129 ();
 FILLCELL_X32 FILLER_172_161 ();
 FILLCELL_X32 FILLER_172_193 ();
 FILLCELL_X32 FILLER_172_225 ();
 FILLCELL_X32 FILLER_172_257 ();
 FILLCELL_X32 FILLER_172_289 ();
 FILLCELL_X32 FILLER_172_321 ();
 FILLCELL_X32 FILLER_172_353 ();
 FILLCELL_X32 FILLER_172_385 ();
 FILLCELL_X32 FILLER_172_417 ();
 FILLCELL_X32 FILLER_172_449 ();
 FILLCELL_X32 FILLER_172_481 ();
 FILLCELL_X32 FILLER_172_513 ();
 FILLCELL_X32 FILLER_172_545 ();
 FILLCELL_X32 FILLER_172_577 ();
 FILLCELL_X16 FILLER_172_609 ();
 FILLCELL_X4 FILLER_172_625 ();
 FILLCELL_X2 FILLER_172_629 ();
 FILLCELL_X32 FILLER_172_632 ();
 FILLCELL_X32 FILLER_172_664 ();
 FILLCELL_X32 FILLER_172_696 ();
 FILLCELL_X32 FILLER_172_728 ();
 FILLCELL_X32 FILLER_172_760 ();
 FILLCELL_X32 FILLER_172_792 ();
 FILLCELL_X32 FILLER_172_824 ();
 FILLCELL_X32 FILLER_172_856 ();
 FILLCELL_X32 FILLER_172_888 ();
 FILLCELL_X32 FILLER_172_920 ();
 FILLCELL_X32 FILLER_172_952 ();
 FILLCELL_X32 FILLER_172_984 ();
 FILLCELL_X32 FILLER_172_1016 ();
 FILLCELL_X32 FILLER_172_1048 ();
 FILLCELL_X8 FILLER_172_1080 ();
 FILLCELL_X4 FILLER_172_1088 ();
 FILLCELL_X2 FILLER_172_1092 ();
 FILLCELL_X4 FILLER_172_1101 ();
 FILLCELL_X1 FILLER_172_1109 ();
 FILLCELL_X16 FILLER_172_1120 ();
 FILLCELL_X8 FILLER_172_1136 ();
 FILLCELL_X4 FILLER_172_1144 ();
 FILLCELL_X2 FILLER_172_1148 ();
 FILLCELL_X1 FILLER_172_1150 ();
 FILLCELL_X2 FILLER_172_1166 ();
 FILLCELL_X16 FILLER_172_1181 ();
 FILLCELL_X4 FILLER_172_1197 ();
 FILLCELL_X4 FILLER_172_1214 ();
 FILLCELL_X2 FILLER_172_1218 ();
 FILLCELL_X1 FILLER_172_1220 ();
 FILLCELL_X16 FILLER_172_1228 ();
 FILLCELL_X4 FILLER_172_1244 ();
 FILLCELL_X2 FILLER_172_1248 ();
 FILLCELL_X1 FILLER_172_1250 ();
 FILLCELL_X1 FILLER_172_1270 ();
 FILLCELL_X8 FILLER_172_1284 ();
 FILLCELL_X2 FILLER_172_1292 ();
 FILLCELL_X16 FILLER_172_1301 ();
 FILLCELL_X8 FILLER_172_1317 ();
 FILLCELL_X4 FILLER_172_1325 ();
 FILLCELL_X1 FILLER_172_1329 ();
 FILLCELL_X32 FILLER_172_1337 ();
 FILLCELL_X32 FILLER_172_1369 ();
 FILLCELL_X32 FILLER_172_1401 ();
 FILLCELL_X4 FILLER_172_1433 ();
 FILLCELL_X32 FILLER_172_1452 ();
 FILLCELL_X32 FILLER_172_1484 ();
 FILLCELL_X32 FILLER_172_1533 ();
 FILLCELL_X2 FILLER_172_1565 ();
 FILLCELL_X1 FILLER_172_1567 ();
 FILLCELL_X32 FILLER_172_1592 ();
 FILLCELL_X32 FILLER_172_1624 ();
 FILLCELL_X32 FILLER_172_1656 ();
 FILLCELL_X32 FILLER_172_1688 ();
 FILLCELL_X32 FILLER_172_1720 ();
 FILLCELL_X32 FILLER_172_1752 ();
 FILLCELL_X32 FILLER_172_1784 ();
 FILLCELL_X32 FILLER_172_1816 ();
 FILLCELL_X32 FILLER_172_1848 ();
 FILLCELL_X8 FILLER_172_1880 ();
 FILLCELL_X4 FILLER_172_1888 ();
 FILLCELL_X2 FILLER_172_1892 ();
 FILLCELL_X32 FILLER_172_1895 ();
 FILLCELL_X32 FILLER_172_1927 ();
 FILLCELL_X32 FILLER_172_1959 ();
 FILLCELL_X32 FILLER_172_1991 ();
 FILLCELL_X32 FILLER_172_2023 ();
 FILLCELL_X32 FILLER_172_2055 ();
 FILLCELL_X32 FILLER_172_2087 ();
 FILLCELL_X32 FILLER_172_2119 ();
 FILLCELL_X32 FILLER_172_2151 ();
 FILLCELL_X32 FILLER_172_2183 ();
 FILLCELL_X32 FILLER_172_2215 ();
 FILLCELL_X32 FILLER_172_2247 ();
 FILLCELL_X32 FILLER_172_2279 ();
 FILLCELL_X32 FILLER_172_2311 ();
 FILLCELL_X32 FILLER_172_2343 ();
 FILLCELL_X32 FILLER_172_2375 ();
 FILLCELL_X32 FILLER_172_2407 ();
 FILLCELL_X32 FILLER_172_2439 ();
 FILLCELL_X32 FILLER_172_2471 ();
 FILLCELL_X32 FILLER_172_2503 ();
 FILLCELL_X32 FILLER_172_2535 ();
 FILLCELL_X32 FILLER_172_2567 ();
 FILLCELL_X2 FILLER_172_2599 ();
 FILLCELL_X1 FILLER_172_2601 ();
 FILLCELL_X32 FILLER_173_1 ();
 FILLCELL_X32 FILLER_173_33 ();
 FILLCELL_X32 FILLER_173_65 ();
 FILLCELL_X32 FILLER_173_97 ();
 FILLCELL_X32 FILLER_173_129 ();
 FILLCELL_X32 FILLER_173_161 ();
 FILLCELL_X32 FILLER_173_193 ();
 FILLCELL_X32 FILLER_173_225 ();
 FILLCELL_X32 FILLER_173_257 ();
 FILLCELL_X32 FILLER_173_289 ();
 FILLCELL_X32 FILLER_173_321 ();
 FILLCELL_X32 FILLER_173_353 ();
 FILLCELL_X32 FILLER_173_385 ();
 FILLCELL_X32 FILLER_173_417 ();
 FILLCELL_X32 FILLER_173_449 ();
 FILLCELL_X32 FILLER_173_481 ();
 FILLCELL_X32 FILLER_173_513 ();
 FILLCELL_X32 FILLER_173_545 ();
 FILLCELL_X32 FILLER_173_577 ();
 FILLCELL_X32 FILLER_173_609 ();
 FILLCELL_X32 FILLER_173_641 ();
 FILLCELL_X32 FILLER_173_673 ();
 FILLCELL_X32 FILLER_173_705 ();
 FILLCELL_X32 FILLER_173_737 ();
 FILLCELL_X32 FILLER_173_769 ();
 FILLCELL_X32 FILLER_173_801 ();
 FILLCELL_X32 FILLER_173_833 ();
 FILLCELL_X32 FILLER_173_865 ();
 FILLCELL_X32 FILLER_173_897 ();
 FILLCELL_X32 FILLER_173_929 ();
 FILLCELL_X32 FILLER_173_961 ();
 FILLCELL_X32 FILLER_173_993 ();
 FILLCELL_X32 FILLER_173_1025 ();
 FILLCELL_X32 FILLER_173_1057 ();
 FILLCELL_X16 FILLER_173_1089 ();
 FILLCELL_X8 FILLER_173_1105 ();
 FILLCELL_X4 FILLER_173_1113 ();
 FILLCELL_X1 FILLER_173_1117 ();
 FILLCELL_X8 FILLER_173_1120 ();
 FILLCELL_X2 FILLER_173_1128 ();
 FILLCELL_X32 FILLER_173_1143 ();
 FILLCELL_X32 FILLER_173_1175 ();
 FILLCELL_X16 FILLER_173_1207 ();
 FILLCELL_X16 FILLER_173_1226 ();
 FILLCELL_X4 FILLER_173_1242 ();
 FILLCELL_X2 FILLER_173_1246 ();
 FILLCELL_X1 FILLER_173_1248 ();
 FILLCELL_X8 FILLER_173_1252 ();
 FILLCELL_X2 FILLER_173_1260 ();
 FILLCELL_X1 FILLER_173_1262 ();
 FILLCELL_X16 FILLER_173_1264 ();
 FILLCELL_X8 FILLER_173_1280 ();
 FILLCELL_X2 FILLER_173_1288 ();
 FILLCELL_X8 FILLER_173_1307 ();
 FILLCELL_X4 FILLER_173_1315 ();
 FILLCELL_X16 FILLER_173_1343 ();
 FILLCELL_X4 FILLER_173_1359 ();
 FILLCELL_X2 FILLER_173_1363 ();
 FILLCELL_X4 FILLER_173_1372 ();
 FILLCELL_X1 FILLER_173_1376 ();
 FILLCELL_X16 FILLER_173_1384 ();
 FILLCELL_X1 FILLER_173_1400 ();
 FILLCELL_X1 FILLER_173_1408 ();
 FILLCELL_X16 FILLER_173_1416 ();
 FILLCELL_X8 FILLER_173_1432 ();
 FILLCELL_X32 FILLER_173_1457 ();
 FILLCELL_X8 FILLER_173_1489 ();
 FILLCELL_X4 FILLER_173_1497 ();
 FILLCELL_X2 FILLER_173_1501 ();
 FILLCELL_X16 FILLER_173_1510 ();
 FILLCELL_X1 FILLER_173_1550 ();
 FILLCELL_X4 FILLER_173_1558 ();
 FILLCELL_X2 FILLER_173_1562 ();
 FILLCELL_X4 FILLER_173_1581 ();
 FILLCELL_X1 FILLER_173_1585 ();
 FILLCELL_X32 FILLER_173_1593 ();
 FILLCELL_X32 FILLER_173_1625 ();
 FILLCELL_X32 FILLER_173_1657 ();
 FILLCELL_X32 FILLER_173_1689 ();
 FILLCELL_X32 FILLER_173_1721 ();
 FILLCELL_X32 FILLER_173_1753 ();
 FILLCELL_X32 FILLER_173_1785 ();
 FILLCELL_X32 FILLER_173_1817 ();
 FILLCELL_X32 FILLER_173_1849 ();
 FILLCELL_X32 FILLER_173_1881 ();
 FILLCELL_X32 FILLER_173_1913 ();
 FILLCELL_X32 FILLER_173_1945 ();
 FILLCELL_X32 FILLER_173_1977 ();
 FILLCELL_X32 FILLER_173_2009 ();
 FILLCELL_X32 FILLER_173_2041 ();
 FILLCELL_X32 FILLER_173_2073 ();
 FILLCELL_X32 FILLER_173_2105 ();
 FILLCELL_X32 FILLER_173_2137 ();
 FILLCELL_X32 FILLER_173_2169 ();
 FILLCELL_X32 FILLER_173_2201 ();
 FILLCELL_X32 FILLER_173_2233 ();
 FILLCELL_X32 FILLER_173_2265 ();
 FILLCELL_X32 FILLER_173_2297 ();
 FILLCELL_X32 FILLER_173_2329 ();
 FILLCELL_X32 FILLER_173_2361 ();
 FILLCELL_X32 FILLER_173_2393 ();
 FILLCELL_X32 FILLER_173_2425 ();
 FILLCELL_X32 FILLER_173_2457 ();
 FILLCELL_X32 FILLER_173_2489 ();
 FILLCELL_X4 FILLER_173_2521 ();
 FILLCELL_X1 FILLER_173_2525 ();
 FILLCELL_X32 FILLER_173_2527 ();
 FILLCELL_X32 FILLER_173_2559 ();
 FILLCELL_X8 FILLER_173_2591 ();
 FILLCELL_X2 FILLER_173_2599 ();
 FILLCELL_X1 FILLER_173_2601 ();
 FILLCELL_X32 FILLER_174_1 ();
 FILLCELL_X32 FILLER_174_33 ();
 FILLCELL_X32 FILLER_174_65 ();
 FILLCELL_X32 FILLER_174_97 ();
 FILLCELL_X32 FILLER_174_129 ();
 FILLCELL_X32 FILLER_174_161 ();
 FILLCELL_X32 FILLER_174_193 ();
 FILLCELL_X32 FILLER_174_225 ();
 FILLCELL_X32 FILLER_174_257 ();
 FILLCELL_X32 FILLER_174_289 ();
 FILLCELL_X32 FILLER_174_321 ();
 FILLCELL_X32 FILLER_174_353 ();
 FILLCELL_X32 FILLER_174_385 ();
 FILLCELL_X32 FILLER_174_417 ();
 FILLCELL_X32 FILLER_174_449 ();
 FILLCELL_X32 FILLER_174_481 ();
 FILLCELL_X32 FILLER_174_513 ();
 FILLCELL_X32 FILLER_174_545 ();
 FILLCELL_X32 FILLER_174_577 ();
 FILLCELL_X16 FILLER_174_609 ();
 FILLCELL_X4 FILLER_174_625 ();
 FILLCELL_X2 FILLER_174_629 ();
 FILLCELL_X32 FILLER_174_632 ();
 FILLCELL_X32 FILLER_174_664 ();
 FILLCELL_X32 FILLER_174_696 ();
 FILLCELL_X32 FILLER_174_728 ();
 FILLCELL_X32 FILLER_174_760 ();
 FILLCELL_X32 FILLER_174_792 ();
 FILLCELL_X32 FILLER_174_824 ();
 FILLCELL_X32 FILLER_174_856 ();
 FILLCELL_X32 FILLER_174_888 ();
 FILLCELL_X32 FILLER_174_920 ();
 FILLCELL_X32 FILLER_174_952 ();
 FILLCELL_X32 FILLER_174_984 ();
 FILLCELL_X32 FILLER_174_1016 ();
 FILLCELL_X32 FILLER_174_1048 ();
 FILLCELL_X16 FILLER_174_1080 ();
 FILLCELL_X4 FILLER_174_1096 ();
 FILLCELL_X1 FILLER_174_1100 ();
 FILLCELL_X4 FILLER_174_1105 ();
 FILLCELL_X2 FILLER_174_1109 ();
 FILLCELL_X32 FILLER_174_1121 ();
 FILLCELL_X2 FILLER_174_1153 ();
 FILLCELL_X1 FILLER_174_1155 ();
 FILLCELL_X8 FILLER_174_1179 ();
 FILLCELL_X4 FILLER_174_1187 ();
 FILLCELL_X2 FILLER_174_1191 ();
 FILLCELL_X1 FILLER_174_1193 ();
 FILLCELL_X16 FILLER_174_1204 ();
 FILLCELL_X8 FILLER_174_1220 ();
 FILLCELL_X2 FILLER_174_1228 ();
 FILLCELL_X8 FILLER_174_1239 ();
 FILLCELL_X2 FILLER_174_1247 ();
 FILLCELL_X1 FILLER_174_1249 ();
 FILLCELL_X1 FILLER_174_1253 ();
 FILLCELL_X8 FILLER_174_1267 ();
 FILLCELL_X4 FILLER_174_1275 ();
 FILLCELL_X2 FILLER_174_1279 ();
 FILLCELL_X1 FILLER_174_1281 ();
 FILLCELL_X4 FILLER_174_1289 ();
 FILLCELL_X1 FILLER_174_1293 ();
 FILLCELL_X8 FILLER_174_1302 ();
 FILLCELL_X4 FILLER_174_1310 ();
 FILLCELL_X16 FILLER_174_1331 ();
 FILLCELL_X8 FILLER_174_1347 ();
 FILLCELL_X1 FILLER_174_1389 ();
 FILLCELL_X16 FILLER_174_1424 ();
 FILLCELL_X4 FILLER_174_1440 ();
 FILLCELL_X2 FILLER_174_1444 ();
 FILLCELL_X32 FILLER_174_1463 ();
 FILLCELL_X2 FILLER_174_1495 ();
 FILLCELL_X1 FILLER_174_1497 ();
 FILLCELL_X1 FILLER_174_1522 ();
 FILLCELL_X32 FILLER_174_1537 ();
 FILLCELL_X4 FILLER_174_1569 ();
 FILLCELL_X2 FILLER_174_1573 ();
 FILLCELL_X1 FILLER_174_1575 ();
 FILLCELL_X8 FILLER_174_1593 ();
 FILLCELL_X2 FILLER_174_1601 ();
 FILLCELL_X32 FILLER_174_1607 ();
 FILLCELL_X32 FILLER_174_1639 ();
 FILLCELL_X32 FILLER_174_1671 ();
 FILLCELL_X32 FILLER_174_1703 ();
 FILLCELL_X32 FILLER_174_1735 ();
 FILLCELL_X32 FILLER_174_1767 ();
 FILLCELL_X32 FILLER_174_1799 ();
 FILLCELL_X32 FILLER_174_1831 ();
 FILLCELL_X16 FILLER_174_1863 ();
 FILLCELL_X8 FILLER_174_1879 ();
 FILLCELL_X4 FILLER_174_1887 ();
 FILLCELL_X2 FILLER_174_1891 ();
 FILLCELL_X1 FILLER_174_1893 ();
 FILLCELL_X32 FILLER_174_1895 ();
 FILLCELL_X32 FILLER_174_1927 ();
 FILLCELL_X32 FILLER_174_1959 ();
 FILLCELL_X32 FILLER_174_1991 ();
 FILLCELL_X32 FILLER_174_2023 ();
 FILLCELL_X32 FILLER_174_2055 ();
 FILLCELL_X32 FILLER_174_2087 ();
 FILLCELL_X32 FILLER_174_2119 ();
 FILLCELL_X32 FILLER_174_2151 ();
 FILLCELL_X32 FILLER_174_2183 ();
 FILLCELL_X32 FILLER_174_2215 ();
 FILLCELL_X32 FILLER_174_2247 ();
 FILLCELL_X32 FILLER_174_2279 ();
 FILLCELL_X32 FILLER_174_2311 ();
 FILLCELL_X32 FILLER_174_2343 ();
 FILLCELL_X32 FILLER_174_2375 ();
 FILLCELL_X32 FILLER_174_2407 ();
 FILLCELL_X32 FILLER_174_2439 ();
 FILLCELL_X32 FILLER_174_2471 ();
 FILLCELL_X32 FILLER_174_2503 ();
 FILLCELL_X32 FILLER_174_2535 ();
 FILLCELL_X32 FILLER_174_2567 ();
 FILLCELL_X2 FILLER_174_2599 ();
 FILLCELL_X1 FILLER_174_2601 ();
 FILLCELL_X16 FILLER_175_1 ();
 FILLCELL_X8 FILLER_175_17 ();
 FILLCELL_X4 FILLER_175_25 ();
 FILLCELL_X32 FILLER_175_36 ();
 FILLCELL_X32 FILLER_175_68 ();
 FILLCELL_X32 FILLER_175_100 ();
 FILLCELL_X32 FILLER_175_132 ();
 FILLCELL_X32 FILLER_175_164 ();
 FILLCELL_X32 FILLER_175_196 ();
 FILLCELL_X32 FILLER_175_228 ();
 FILLCELL_X32 FILLER_175_260 ();
 FILLCELL_X32 FILLER_175_292 ();
 FILLCELL_X32 FILLER_175_324 ();
 FILLCELL_X32 FILLER_175_356 ();
 FILLCELL_X32 FILLER_175_388 ();
 FILLCELL_X32 FILLER_175_420 ();
 FILLCELL_X32 FILLER_175_452 ();
 FILLCELL_X32 FILLER_175_484 ();
 FILLCELL_X32 FILLER_175_516 ();
 FILLCELL_X32 FILLER_175_548 ();
 FILLCELL_X32 FILLER_175_580 ();
 FILLCELL_X32 FILLER_175_612 ();
 FILLCELL_X32 FILLER_175_644 ();
 FILLCELL_X32 FILLER_175_676 ();
 FILLCELL_X32 FILLER_175_708 ();
 FILLCELL_X32 FILLER_175_740 ();
 FILLCELL_X32 FILLER_175_772 ();
 FILLCELL_X32 FILLER_175_804 ();
 FILLCELL_X32 FILLER_175_836 ();
 FILLCELL_X32 FILLER_175_868 ();
 FILLCELL_X32 FILLER_175_900 ();
 FILLCELL_X32 FILLER_175_932 ();
 FILLCELL_X32 FILLER_175_964 ();
 FILLCELL_X32 FILLER_175_996 ();
 FILLCELL_X32 FILLER_175_1028 ();
 FILLCELL_X32 FILLER_175_1060 ();
 FILLCELL_X32 FILLER_175_1092 ();
 FILLCELL_X32 FILLER_175_1124 ();
 FILLCELL_X4 FILLER_175_1156 ();
 FILLCELL_X2 FILLER_175_1160 ();
 FILLCELL_X2 FILLER_175_1166 ();
 FILLCELL_X8 FILLER_175_1179 ();
 FILLCELL_X4 FILLER_175_1187 ();
 FILLCELL_X2 FILLER_175_1191 ();
 FILLCELL_X1 FILLER_175_1193 ();
 FILLCELL_X4 FILLER_175_1204 ();
 FILLCELL_X32 FILLER_175_1218 ();
 FILLCELL_X8 FILLER_175_1264 ();
 FILLCELL_X1 FILLER_175_1272 ();
 FILLCELL_X8 FILLER_175_1290 ();
 FILLCELL_X32 FILLER_175_1313 ();
 FILLCELL_X32 FILLER_175_1345 ();
 FILLCELL_X16 FILLER_175_1377 ();
 FILLCELL_X8 FILLER_175_1393 ();
 FILLCELL_X4 FILLER_175_1401 ();
 FILLCELL_X1 FILLER_175_1405 ();
 FILLCELL_X4 FILLER_175_1413 ();
 FILLCELL_X2 FILLER_175_1417 ();
 FILLCELL_X1 FILLER_175_1419 ();
 FILLCELL_X16 FILLER_175_1427 ();
 FILLCELL_X8 FILLER_175_1443 ();
 FILLCELL_X32 FILLER_175_1458 ();
 FILLCELL_X4 FILLER_175_1490 ();
 FILLCELL_X8 FILLER_175_1511 ();
 FILLCELL_X2 FILLER_175_1519 ();
 FILLCELL_X16 FILLER_175_1538 ();
 FILLCELL_X2 FILLER_175_1554 ();
 FILLCELL_X8 FILLER_175_1563 ();
 FILLCELL_X4 FILLER_175_1571 ();
 FILLCELL_X2 FILLER_175_1575 ();
 FILLCELL_X1 FILLER_175_1577 ();
 FILLCELL_X4 FILLER_175_1616 ();
 FILLCELL_X32 FILLER_175_1624 ();
 FILLCELL_X32 FILLER_175_1656 ();
 FILLCELL_X32 FILLER_175_1688 ();
 FILLCELL_X32 FILLER_175_1720 ();
 FILLCELL_X32 FILLER_175_1752 ();
 FILLCELL_X32 FILLER_175_1784 ();
 FILLCELL_X32 FILLER_175_1816 ();
 FILLCELL_X32 FILLER_175_1848 ();
 FILLCELL_X32 FILLER_175_1880 ();
 FILLCELL_X32 FILLER_175_1912 ();
 FILLCELL_X32 FILLER_175_1944 ();
 FILLCELL_X32 FILLER_175_1976 ();
 FILLCELL_X32 FILLER_175_2008 ();
 FILLCELL_X32 FILLER_175_2040 ();
 FILLCELL_X32 FILLER_175_2072 ();
 FILLCELL_X32 FILLER_175_2104 ();
 FILLCELL_X32 FILLER_175_2136 ();
 FILLCELL_X32 FILLER_175_2168 ();
 FILLCELL_X32 FILLER_175_2200 ();
 FILLCELL_X32 FILLER_175_2232 ();
 FILLCELL_X32 FILLER_175_2264 ();
 FILLCELL_X32 FILLER_175_2296 ();
 FILLCELL_X32 FILLER_175_2328 ();
 FILLCELL_X32 FILLER_175_2360 ();
 FILLCELL_X32 FILLER_175_2392 ();
 FILLCELL_X32 FILLER_175_2424 ();
 FILLCELL_X32 FILLER_175_2456 ();
 FILLCELL_X32 FILLER_175_2488 ();
 FILLCELL_X4 FILLER_175_2520 ();
 FILLCELL_X2 FILLER_175_2524 ();
 FILLCELL_X32 FILLER_175_2527 ();
 FILLCELL_X32 FILLER_175_2559 ();
 FILLCELL_X8 FILLER_175_2591 ();
 FILLCELL_X2 FILLER_175_2599 ();
 FILLCELL_X1 FILLER_175_2601 ();
 FILLCELL_X8 FILLER_176_1 ();
 FILLCELL_X4 FILLER_176_9 ();
 FILLCELL_X32 FILLER_176_16 ();
 FILLCELL_X32 FILLER_176_48 ();
 FILLCELL_X32 FILLER_176_80 ();
 FILLCELL_X32 FILLER_176_112 ();
 FILLCELL_X32 FILLER_176_144 ();
 FILLCELL_X32 FILLER_176_176 ();
 FILLCELL_X32 FILLER_176_208 ();
 FILLCELL_X32 FILLER_176_240 ();
 FILLCELL_X32 FILLER_176_272 ();
 FILLCELL_X32 FILLER_176_304 ();
 FILLCELL_X32 FILLER_176_336 ();
 FILLCELL_X32 FILLER_176_368 ();
 FILLCELL_X32 FILLER_176_400 ();
 FILLCELL_X32 FILLER_176_432 ();
 FILLCELL_X32 FILLER_176_464 ();
 FILLCELL_X32 FILLER_176_496 ();
 FILLCELL_X32 FILLER_176_528 ();
 FILLCELL_X32 FILLER_176_560 ();
 FILLCELL_X32 FILLER_176_592 ();
 FILLCELL_X4 FILLER_176_624 ();
 FILLCELL_X2 FILLER_176_628 ();
 FILLCELL_X1 FILLER_176_630 ();
 FILLCELL_X32 FILLER_176_632 ();
 FILLCELL_X32 FILLER_176_664 ();
 FILLCELL_X32 FILLER_176_696 ();
 FILLCELL_X32 FILLER_176_728 ();
 FILLCELL_X32 FILLER_176_760 ();
 FILLCELL_X32 FILLER_176_792 ();
 FILLCELL_X32 FILLER_176_824 ();
 FILLCELL_X32 FILLER_176_856 ();
 FILLCELL_X32 FILLER_176_888 ();
 FILLCELL_X32 FILLER_176_920 ();
 FILLCELL_X32 FILLER_176_952 ();
 FILLCELL_X32 FILLER_176_984 ();
 FILLCELL_X32 FILLER_176_1016 ();
 FILLCELL_X32 FILLER_176_1048 ();
 FILLCELL_X32 FILLER_176_1080 ();
 FILLCELL_X16 FILLER_176_1112 ();
 FILLCELL_X1 FILLER_176_1128 ();
 FILLCELL_X32 FILLER_176_1235 ();
 FILLCELL_X16 FILLER_176_1267 ();
 FILLCELL_X4 FILLER_176_1283 ();
 FILLCELL_X4 FILLER_176_1294 ();
 FILLCELL_X32 FILLER_176_1305 ();
 FILLCELL_X1 FILLER_176_1337 ();
 FILLCELL_X32 FILLER_176_1345 ();
 FILLCELL_X16 FILLER_176_1377 ();
 FILLCELL_X4 FILLER_176_1393 ();
 FILLCELL_X2 FILLER_176_1397 ();
 FILLCELL_X1 FILLER_176_1399 ();
 FILLCELL_X2 FILLER_176_1407 ();
 FILLCELL_X2 FILLER_176_1423 ();
 FILLCELL_X16 FILLER_176_1432 ();
 FILLCELL_X8 FILLER_176_1448 ();
 FILLCELL_X4 FILLER_176_1456 ();
 FILLCELL_X32 FILLER_176_1467 ();
 FILLCELL_X32 FILLER_176_1499 ();
 FILLCELL_X8 FILLER_176_1531 ();
 FILLCELL_X2 FILLER_176_1539 ();
 FILLCELL_X2 FILLER_176_1548 ();
 FILLCELL_X1 FILLER_176_1550 ();
 FILLCELL_X32 FILLER_176_1558 ();
 FILLCELL_X32 FILLER_176_1590 ();
 FILLCELL_X32 FILLER_176_1622 ();
 FILLCELL_X32 FILLER_176_1654 ();
 FILLCELL_X32 FILLER_176_1686 ();
 FILLCELL_X32 FILLER_176_1718 ();
 FILLCELL_X32 FILLER_176_1750 ();
 FILLCELL_X32 FILLER_176_1782 ();
 FILLCELL_X32 FILLER_176_1814 ();
 FILLCELL_X32 FILLER_176_1846 ();
 FILLCELL_X16 FILLER_176_1878 ();
 FILLCELL_X32 FILLER_176_1895 ();
 FILLCELL_X32 FILLER_176_1927 ();
 FILLCELL_X32 FILLER_176_1959 ();
 FILLCELL_X32 FILLER_176_1991 ();
 FILLCELL_X32 FILLER_176_2023 ();
 FILLCELL_X32 FILLER_176_2055 ();
 FILLCELL_X32 FILLER_176_2087 ();
 FILLCELL_X32 FILLER_176_2119 ();
 FILLCELL_X32 FILLER_176_2151 ();
 FILLCELL_X32 FILLER_176_2183 ();
 FILLCELL_X32 FILLER_176_2215 ();
 FILLCELL_X32 FILLER_176_2247 ();
 FILLCELL_X32 FILLER_176_2279 ();
 FILLCELL_X32 FILLER_176_2311 ();
 FILLCELL_X32 FILLER_176_2343 ();
 FILLCELL_X32 FILLER_176_2375 ();
 FILLCELL_X32 FILLER_176_2407 ();
 FILLCELL_X32 FILLER_176_2439 ();
 FILLCELL_X32 FILLER_176_2471 ();
 FILLCELL_X32 FILLER_176_2503 ();
 FILLCELL_X32 FILLER_176_2535 ();
 FILLCELL_X16 FILLER_176_2567 ();
 FILLCELL_X4 FILLER_176_2583 ();
 FILLCELL_X2 FILLER_176_2587 ();
 FILLCELL_X1 FILLER_176_2589 ();
 FILLCELL_X2 FILLER_176_2593 ();
 FILLCELL_X1 FILLER_176_2595 ();
 FILLCELL_X32 FILLER_177_1 ();
 FILLCELL_X32 FILLER_177_33 ();
 FILLCELL_X32 FILLER_177_65 ();
 FILLCELL_X32 FILLER_177_97 ();
 FILLCELL_X32 FILLER_177_129 ();
 FILLCELL_X32 FILLER_177_161 ();
 FILLCELL_X32 FILLER_177_193 ();
 FILLCELL_X32 FILLER_177_225 ();
 FILLCELL_X32 FILLER_177_257 ();
 FILLCELL_X32 FILLER_177_289 ();
 FILLCELL_X32 FILLER_177_321 ();
 FILLCELL_X32 FILLER_177_353 ();
 FILLCELL_X32 FILLER_177_385 ();
 FILLCELL_X32 FILLER_177_417 ();
 FILLCELL_X32 FILLER_177_449 ();
 FILLCELL_X32 FILLER_177_481 ();
 FILLCELL_X32 FILLER_177_513 ();
 FILLCELL_X32 FILLER_177_545 ();
 FILLCELL_X32 FILLER_177_577 ();
 FILLCELL_X32 FILLER_177_609 ();
 FILLCELL_X32 FILLER_177_641 ();
 FILLCELL_X32 FILLER_177_673 ();
 FILLCELL_X32 FILLER_177_705 ();
 FILLCELL_X32 FILLER_177_737 ();
 FILLCELL_X32 FILLER_177_769 ();
 FILLCELL_X32 FILLER_177_801 ();
 FILLCELL_X32 FILLER_177_833 ();
 FILLCELL_X32 FILLER_177_865 ();
 FILLCELL_X32 FILLER_177_897 ();
 FILLCELL_X32 FILLER_177_929 ();
 FILLCELL_X32 FILLER_177_961 ();
 FILLCELL_X32 FILLER_177_993 ();
 FILLCELL_X32 FILLER_177_1025 ();
 FILLCELL_X32 FILLER_177_1057 ();
 FILLCELL_X32 FILLER_177_1089 ();
 FILLCELL_X8 FILLER_177_1121 ();
 FILLCELL_X4 FILLER_177_1129 ();
 FILLCELL_X2 FILLER_177_1133 ();
 FILLCELL_X32 FILLER_177_1139 ();
 FILLCELL_X32 FILLER_177_1171 ();
 FILLCELL_X16 FILLER_177_1203 ();
 FILLCELL_X16 FILLER_177_1245 ();
 FILLCELL_X2 FILLER_177_1261 ();
 FILLCELL_X32 FILLER_177_1264 ();
 FILLCELL_X4 FILLER_177_1296 ();
 FILLCELL_X2 FILLER_177_1300 ();
 FILLCELL_X1 FILLER_177_1302 ();
 FILLCELL_X16 FILLER_177_1310 ();
 FILLCELL_X1 FILLER_177_1326 ();
 FILLCELL_X1 FILLER_177_1334 ();
 FILLCELL_X32 FILLER_177_1349 ();
 FILLCELL_X1 FILLER_177_1381 ();
 FILLCELL_X32 FILLER_177_1389 ();
 FILLCELL_X32 FILLER_177_1421 ();
 FILLCELL_X2 FILLER_177_1453 ();
 FILLCELL_X1 FILLER_177_1455 ();
 FILLCELL_X32 FILLER_177_1477 ();
 FILLCELL_X2 FILLER_177_1509 ();
 FILLCELL_X8 FILLER_177_1518 ();
 FILLCELL_X4 FILLER_177_1526 ();
 FILLCELL_X1 FILLER_177_1530 ();
 FILLCELL_X16 FILLER_177_1538 ();
 FILLCELL_X2 FILLER_177_1554 ();
 FILLCELL_X1 FILLER_177_1556 ();
 FILLCELL_X32 FILLER_177_1564 ();
 FILLCELL_X32 FILLER_177_1596 ();
 FILLCELL_X32 FILLER_177_1628 ();
 FILLCELL_X32 FILLER_177_1660 ();
 FILLCELL_X32 FILLER_177_1692 ();
 FILLCELL_X32 FILLER_177_1724 ();
 FILLCELL_X32 FILLER_177_1756 ();
 FILLCELL_X32 FILLER_177_1788 ();
 FILLCELL_X32 FILLER_177_1820 ();
 FILLCELL_X32 FILLER_177_1852 ();
 FILLCELL_X32 FILLER_177_1884 ();
 FILLCELL_X32 FILLER_177_1916 ();
 FILLCELL_X32 FILLER_177_1948 ();
 FILLCELL_X32 FILLER_177_1980 ();
 FILLCELL_X32 FILLER_177_2012 ();
 FILLCELL_X32 FILLER_177_2044 ();
 FILLCELL_X32 FILLER_177_2076 ();
 FILLCELL_X32 FILLER_177_2108 ();
 FILLCELL_X32 FILLER_177_2140 ();
 FILLCELL_X32 FILLER_177_2172 ();
 FILLCELL_X32 FILLER_177_2204 ();
 FILLCELL_X32 FILLER_177_2236 ();
 FILLCELL_X32 FILLER_177_2268 ();
 FILLCELL_X32 FILLER_177_2300 ();
 FILLCELL_X32 FILLER_177_2332 ();
 FILLCELL_X32 FILLER_177_2364 ();
 FILLCELL_X32 FILLER_177_2396 ();
 FILLCELL_X32 FILLER_177_2428 ();
 FILLCELL_X32 FILLER_177_2460 ();
 FILLCELL_X32 FILLER_177_2492 ();
 FILLCELL_X2 FILLER_177_2524 ();
 FILLCELL_X32 FILLER_177_2527 ();
 FILLCELL_X16 FILLER_177_2559 ();
 FILLCELL_X1 FILLER_177_2575 ();
 FILLCELL_X1 FILLER_177_2579 ();
 FILLCELL_X2 FILLER_177_2583 ();
 FILLCELL_X8 FILLER_177_2591 ();
 FILLCELL_X2 FILLER_177_2599 ();
 FILLCELL_X1 FILLER_177_2601 ();
 FILLCELL_X32 FILLER_178_1 ();
 FILLCELL_X32 FILLER_178_33 ();
 FILLCELL_X32 FILLER_178_65 ();
 FILLCELL_X32 FILLER_178_97 ();
 FILLCELL_X32 FILLER_178_129 ();
 FILLCELL_X32 FILLER_178_161 ();
 FILLCELL_X32 FILLER_178_193 ();
 FILLCELL_X32 FILLER_178_225 ();
 FILLCELL_X32 FILLER_178_257 ();
 FILLCELL_X32 FILLER_178_289 ();
 FILLCELL_X32 FILLER_178_321 ();
 FILLCELL_X32 FILLER_178_353 ();
 FILLCELL_X32 FILLER_178_385 ();
 FILLCELL_X32 FILLER_178_417 ();
 FILLCELL_X32 FILLER_178_449 ();
 FILLCELL_X32 FILLER_178_481 ();
 FILLCELL_X32 FILLER_178_513 ();
 FILLCELL_X32 FILLER_178_545 ();
 FILLCELL_X32 FILLER_178_577 ();
 FILLCELL_X16 FILLER_178_609 ();
 FILLCELL_X4 FILLER_178_625 ();
 FILLCELL_X2 FILLER_178_629 ();
 FILLCELL_X32 FILLER_178_632 ();
 FILLCELL_X32 FILLER_178_664 ();
 FILLCELL_X32 FILLER_178_696 ();
 FILLCELL_X32 FILLER_178_728 ();
 FILLCELL_X32 FILLER_178_760 ();
 FILLCELL_X32 FILLER_178_792 ();
 FILLCELL_X32 FILLER_178_824 ();
 FILLCELL_X32 FILLER_178_856 ();
 FILLCELL_X32 FILLER_178_888 ();
 FILLCELL_X32 FILLER_178_920 ();
 FILLCELL_X32 FILLER_178_952 ();
 FILLCELL_X32 FILLER_178_984 ();
 FILLCELL_X32 FILLER_178_1016 ();
 FILLCELL_X32 FILLER_178_1048 ();
 FILLCELL_X32 FILLER_178_1080 ();
 FILLCELL_X8 FILLER_178_1112 ();
 FILLCELL_X32 FILLER_178_1124 ();
 FILLCELL_X32 FILLER_178_1156 ();
 FILLCELL_X16 FILLER_178_1188 ();
 FILLCELL_X8 FILLER_178_1204 ();
 FILLCELL_X2 FILLER_178_1212 ();
 FILLCELL_X1 FILLER_178_1214 ();
 FILLCELL_X4 FILLER_178_1218 ();
 FILLCELL_X1 FILLER_178_1222 ();
 FILLCELL_X32 FILLER_178_1226 ();
 FILLCELL_X4 FILLER_178_1258 ();
 FILLCELL_X4 FILLER_178_1279 ();
 FILLCELL_X1 FILLER_178_1283 ();
 FILLCELL_X2 FILLER_178_1301 ();
 FILLCELL_X1 FILLER_178_1303 ();
 FILLCELL_X32 FILLER_178_1318 ();
 FILLCELL_X8 FILLER_178_1350 ();
 FILLCELL_X4 FILLER_178_1358 ();
 FILLCELL_X2 FILLER_178_1362 ();
 FILLCELL_X4 FILLER_178_1378 ();
 FILLCELL_X2 FILLER_178_1382 ();
 FILLCELL_X16 FILLER_178_1391 ();
 FILLCELL_X1 FILLER_178_1407 ();
 FILLCELL_X16 FILLER_178_1425 ();
 FILLCELL_X4 FILLER_178_1441 ();
 FILLCELL_X2 FILLER_178_1445 ();
 FILLCELL_X1 FILLER_178_1447 ();
 FILLCELL_X16 FILLER_178_1465 ();
 FILLCELL_X8 FILLER_178_1481 ();
 FILLCELL_X4 FILLER_178_1489 ();
 FILLCELL_X1 FILLER_178_1493 ();
 FILLCELL_X1 FILLER_178_1525 ();
 FILLCELL_X16 FILLER_178_1550 ();
 FILLCELL_X1 FILLER_178_1566 ();
 FILLCELL_X32 FILLER_178_1591 ();
 FILLCELL_X32 FILLER_178_1623 ();
 FILLCELL_X32 FILLER_178_1655 ();
 FILLCELL_X32 FILLER_178_1687 ();
 FILLCELL_X32 FILLER_178_1719 ();
 FILLCELL_X32 FILLER_178_1751 ();
 FILLCELL_X32 FILLER_178_1783 ();
 FILLCELL_X32 FILLER_178_1815 ();
 FILLCELL_X32 FILLER_178_1847 ();
 FILLCELL_X8 FILLER_178_1879 ();
 FILLCELL_X4 FILLER_178_1887 ();
 FILLCELL_X2 FILLER_178_1891 ();
 FILLCELL_X1 FILLER_178_1893 ();
 FILLCELL_X32 FILLER_178_1895 ();
 FILLCELL_X32 FILLER_178_1927 ();
 FILLCELL_X32 FILLER_178_1959 ();
 FILLCELL_X32 FILLER_178_1991 ();
 FILLCELL_X32 FILLER_178_2023 ();
 FILLCELL_X32 FILLER_178_2055 ();
 FILLCELL_X32 FILLER_178_2087 ();
 FILLCELL_X32 FILLER_178_2119 ();
 FILLCELL_X32 FILLER_178_2151 ();
 FILLCELL_X32 FILLER_178_2183 ();
 FILLCELL_X32 FILLER_178_2215 ();
 FILLCELL_X32 FILLER_178_2247 ();
 FILLCELL_X32 FILLER_178_2279 ();
 FILLCELL_X32 FILLER_178_2311 ();
 FILLCELL_X32 FILLER_178_2343 ();
 FILLCELL_X32 FILLER_178_2375 ();
 FILLCELL_X32 FILLER_178_2407 ();
 FILLCELL_X32 FILLER_178_2439 ();
 FILLCELL_X32 FILLER_178_2471 ();
 FILLCELL_X32 FILLER_178_2503 ();
 FILLCELL_X16 FILLER_178_2535 ();
 FILLCELL_X4 FILLER_178_2551 ();
 FILLCELL_X2 FILLER_178_2555 ();
 FILLCELL_X8 FILLER_178_2563 ();
 FILLCELL_X4 FILLER_178_2571 ();
 FILLCELL_X2 FILLER_178_2575 ();
 FILLCELL_X1 FILLER_178_2577 ();
 FILLCELL_X1 FILLER_178_2581 ();
 FILLCELL_X4 FILLER_178_2585 ();
 FILLCELL_X1 FILLER_178_2589 ();
 FILLCELL_X4 FILLER_178_2593 ();
 FILLCELL_X2 FILLER_178_2597 ();
 FILLCELL_X32 FILLER_179_1 ();
 FILLCELL_X32 FILLER_179_33 ();
 FILLCELL_X32 FILLER_179_65 ();
 FILLCELL_X32 FILLER_179_97 ();
 FILLCELL_X32 FILLER_179_129 ();
 FILLCELL_X32 FILLER_179_161 ();
 FILLCELL_X32 FILLER_179_193 ();
 FILLCELL_X32 FILLER_179_225 ();
 FILLCELL_X32 FILLER_179_257 ();
 FILLCELL_X32 FILLER_179_289 ();
 FILLCELL_X32 FILLER_179_321 ();
 FILLCELL_X32 FILLER_179_353 ();
 FILLCELL_X32 FILLER_179_385 ();
 FILLCELL_X32 FILLER_179_417 ();
 FILLCELL_X32 FILLER_179_449 ();
 FILLCELL_X32 FILLER_179_481 ();
 FILLCELL_X32 FILLER_179_513 ();
 FILLCELL_X32 FILLER_179_545 ();
 FILLCELL_X32 FILLER_179_577 ();
 FILLCELL_X32 FILLER_179_609 ();
 FILLCELL_X32 FILLER_179_641 ();
 FILLCELL_X32 FILLER_179_673 ();
 FILLCELL_X32 FILLER_179_705 ();
 FILLCELL_X32 FILLER_179_737 ();
 FILLCELL_X32 FILLER_179_769 ();
 FILLCELL_X32 FILLER_179_801 ();
 FILLCELL_X32 FILLER_179_833 ();
 FILLCELL_X32 FILLER_179_865 ();
 FILLCELL_X32 FILLER_179_897 ();
 FILLCELL_X32 FILLER_179_929 ();
 FILLCELL_X32 FILLER_179_961 ();
 FILLCELL_X32 FILLER_179_993 ();
 FILLCELL_X32 FILLER_179_1025 ();
 FILLCELL_X32 FILLER_179_1057 ();
 FILLCELL_X8 FILLER_179_1089 ();
 FILLCELL_X1 FILLER_179_1097 ();
 FILLCELL_X1 FILLER_179_1123 ();
 FILLCELL_X32 FILLER_179_1134 ();
 FILLCELL_X32 FILLER_179_1166 ();
 FILLCELL_X32 FILLER_179_1198 ();
 FILLCELL_X32 FILLER_179_1230 ();
 FILLCELL_X1 FILLER_179_1262 ();
 FILLCELL_X2 FILLER_179_1264 ();
 FILLCELL_X8 FILLER_179_1273 ();
 FILLCELL_X2 FILLER_179_1281 ();
 FILLCELL_X16 FILLER_179_1290 ();
 FILLCELL_X8 FILLER_179_1306 ();
 FILLCELL_X2 FILLER_179_1314 ();
 FILLCELL_X1 FILLER_179_1316 ();
 FILLCELL_X16 FILLER_179_1334 ();
 FILLCELL_X16 FILLER_179_1367 ();
 FILLCELL_X1 FILLER_179_1383 ();
 FILLCELL_X8 FILLER_179_1393 ();
 FILLCELL_X4 FILLER_179_1401 ();
 FILLCELL_X1 FILLER_179_1429 ();
 FILLCELL_X4 FILLER_179_1439 ();
 FILLCELL_X2 FILLER_179_1443 ();
 FILLCELL_X1 FILLER_179_1445 ();
 FILLCELL_X4 FILLER_179_1470 ();
 FILLCELL_X2 FILLER_179_1474 ();
 FILLCELL_X1 FILLER_179_1476 ();
 FILLCELL_X16 FILLER_179_1486 ();
 FILLCELL_X2 FILLER_179_1502 ();
 FILLCELL_X32 FILLER_179_1511 ();
 FILLCELL_X8 FILLER_179_1543 ();
 FILLCELL_X2 FILLER_179_1551 ();
 FILLCELL_X32 FILLER_179_1588 ();
 FILLCELL_X32 FILLER_179_1620 ();
 FILLCELL_X32 FILLER_179_1652 ();
 FILLCELL_X32 FILLER_179_1684 ();
 FILLCELL_X32 FILLER_179_1716 ();
 FILLCELL_X32 FILLER_179_1748 ();
 FILLCELL_X32 FILLER_179_1780 ();
 FILLCELL_X32 FILLER_179_1812 ();
 FILLCELL_X32 FILLER_179_1844 ();
 FILLCELL_X32 FILLER_179_1876 ();
 FILLCELL_X32 FILLER_179_1908 ();
 FILLCELL_X32 FILLER_179_1940 ();
 FILLCELL_X32 FILLER_179_1972 ();
 FILLCELL_X32 FILLER_179_2004 ();
 FILLCELL_X32 FILLER_179_2036 ();
 FILLCELL_X32 FILLER_179_2068 ();
 FILLCELL_X32 FILLER_179_2100 ();
 FILLCELL_X32 FILLER_179_2132 ();
 FILLCELL_X32 FILLER_179_2164 ();
 FILLCELL_X32 FILLER_179_2196 ();
 FILLCELL_X32 FILLER_179_2228 ();
 FILLCELL_X32 FILLER_179_2260 ();
 FILLCELL_X32 FILLER_179_2292 ();
 FILLCELL_X32 FILLER_179_2324 ();
 FILLCELL_X32 FILLER_179_2356 ();
 FILLCELL_X32 FILLER_179_2388 ();
 FILLCELL_X32 FILLER_179_2420 ();
 FILLCELL_X32 FILLER_179_2452 ();
 FILLCELL_X32 FILLER_179_2484 ();
 FILLCELL_X8 FILLER_179_2516 ();
 FILLCELL_X2 FILLER_179_2524 ();
 FILLCELL_X32 FILLER_179_2527 ();
 FILLCELL_X32 FILLER_179_2559 ();
 FILLCELL_X8 FILLER_179_2591 ();
 FILLCELL_X2 FILLER_179_2599 ();
 FILLCELL_X1 FILLER_179_2601 ();
 FILLCELL_X32 FILLER_180_8 ();
 FILLCELL_X32 FILLER_180_40 ();
 FILLCELL_X32 FILLER_180_72 ();
 FILLCELL_X32 FILLER_180_104 ();
 FILLCELL_X32 FILLER_180_136 ();
 FILLCELL_X32 FILLER_180_168 ();
 FILLCELL_X32 FILLER_180_200 ();
 FILLCELL_X32 FILLER_180_232 ();
 FILLCELL_X32 FILLER_180_264 ();
 FILLCELL_X32 FILLER_180_296 ();
 FILLCELL_X32 FILLER_180_328 ();
 FILLCELL_X32 FILLER_180_360 ();
 FILLCELL_X32 FILLER_180_392 ();
 FILLCELL_X32 FILLER_180_424 ();
 FILLCELL_X32 FILLER_180_456 ();
 FILLCELL_X32 FILLER_180_488 ();
 FILLCELL_X32 FILLER_180_520 ();
 FILLCELL_X32 FILLER_180_552 ();
 FILLCELL_X32 FILLER_180_584 ();
 FILLCELL_X8 FILLER_180_616 ();
 FILLCELL_X4 FILLER_180_624 ();
 FILLCELL_X2 FILLER_180_628 ();
 FILLCELL_X1 FILLER_180_630 ();
 FILLCELL_X32 FILLER_180_632 ();
 FILLCELL_X32 FILLER_180_664 ();
 FILLCELL_X32 FILLER_180_696 ();
 FILLCELL_X32 FILLER_180_728 ();
 FILLCELL_X32 FILLER_180_760 ();
 FILLCELL_X32 FILLER_180_792 ();
 FILLCELL_X32 FILLER_180_824 ();
 FILLCELL_X32 FILLER_180_856 ();
 FILLCELL_X32 FILLER_180_888 ();
 FILLCELL_X32 FILLER_180_920 ();
 FILLCELL_X32 FILLER_180_952 ();
 FILLCELL_X32 FILLER_180_984 ();
 FILLCELL_X32 FILLER_180_1016 ();
 FILLCELL_X32 FILLER_180_1048 ();
 FILLCELL_X16 FILLER_180_1080 ();
 FILLCELL_X8 FILLER_180_1096 ();
 FILLCELL_X4 FILLER_180_1104 ();
 FILLCELL_X1 FILLER_180_1108 ();
 FILLCELL_X4 FILLER_180_1111 ();
 FILLCELL_X1 FILLER_180_1115 ();
 FILLCELL_X8 FILLER_180_1123 ();
 FILLCELL_X2 FILLER_180_1131 ();
 FILLCELL_X1 FILLER_180_1133 ();
 FILLCELL_X2 FILLER_180_1144 ();
 FILLCELL_X8 FILLER_180_1166 ();
 FILLCELL_X2 FILLER_180_1174 ();
 FILLCELL_X8 FILLER_180_1181 ();
 FILLCELL_X2 FILLER_180_1189 ();
 FILLCELL_X4 FILLER_180_1208 ();
 FILLCELL_X2 FILLER_180_1212 ();
 FILLCELL_X1 FILLER_180_1214 ();
 FILLCELL_X8 FILLER_180_1218 ();
 FILLCELL_X4 FILLER_180_1229 ();
 FILLCELL_X2 FILLER_180_1233 ();
 FILLCELL_X1 FILLER_180_1235 ();
 FILLCELL_X32 FILLER_180_1265 ();
 FILLCELL_X16 FILLER_180_1297 ();
 FILLCELL_X4 FILLER_180_1313 ();
 FILLCELL_X2 FILLER_180_1317 ();
 FILLCELL_X2 FILLER_180_1326 ();
 FILLCELL_X4 FILLER_180_1345 ();
 FILLCELL_X2 FILLER_180_1349 ();
 FILLCELL_X1 FILLER_180_1351 ();
 FILLCELL_X2 FILLER_180_1359 ();
 FILLCELL_X1 FILLER_180_1361 ();
 FILLCELL_X16 FILLER_180_1386 ();
 FILLCELL_X8 FILLER_180_1402 ();
 FILLCELL_X2 FILLER_180_1410 ();
 FILLCELL_X1 FILLER_180_1412 ();
 FILLCELL_X32 FILLER_180_1420 ();
 FILLCELL_X1 FILLER_180_1452 ();
 FILLCELL_X32 FILLER_180_1460 ();
 FILLCELL_X2 FILLER_180_1492 ();
 FILLCELL_X1 FILLER_180_1494 ();
 FILLCELL_X16 FILLER_180_1519 ();
 FILLCELL_X2 FILLER_180_1535 ();
 FILLCELL_X1 FILLER_180_1537 ();
 FILLCELL_X16 FILLER_180_1551 ();
 FILLCELL_X8 FILLER_180_1567 ();
 FILLCELL_X4 FILLER_180_1575 ();
 FILLCELL_X32 FILLER_180_1593 ();
 FILLCELL_X32 FILLER_180_1625 ();
 FILLCELL_X32 FILLER_180_1657 ();
 FILLCELL_X32 FILLER_180_1689 ();
 FILLCELL_X32 FILLER_180_1721 ();
 FILLCELL_X32 FILLER_180_1753 ();
 FILLCELL_X32 FILLER_180_1785 ();
 FILLCELL_X32 FILLER_180_1817 ();
 FILLCELL_X32 FILLER_180_1849 ();
 FILLCELL_X8 FILLER_180_1881 ();
 FILLCELL_X4 FILLER_180_1889 ();
 FILLCELL_X1 FILLER_180_1893 ();
 FILLCELL_X32 FILLER_180_1895 ();
 FILLCELL_X32 FILLER_180_1927 ();
 FILLCELL_X32 FILLER_180_1959 ();
 FILLCELL_X32 FILLER_180_1991 ();
 FILLCELL_X32 FILLER_180_2023 ();
 FILLCELL_X32 FILLER_180_2055 ();
 FILLCELL_X32 FILLER_180_2087 ();
 FILLCELL_X32 FILLER_180_2119 ();
 FILLCELL_X32 FILLER_180_2151 ();
 FILLCELL_X32 FILLER_180_2183 ();
 FILLCELL_X32 FILLER_180_2215 ();
 FILLCELL_X32 FILLER_180_2247 ();
 FILLCELL_X32 FILLER_180_2279 ();
 FILLCELL_X32 FILLER_180_2311 ();
 FILLCELL_X32 FILLER_180_2343 ();
 FILLCELL_X32 FILLER_180_2375 ();
 FILLCELL_X32 FILLER_180_2407 ();
 FILLCELL_X32 FILLER_180_2439 ();
 FILLCELL_X32 FILLER_180_2471 ();
 FILLCELL_X32 FILLER_180_2503 ();
 FILLCELL_X32 FILLER_180_2535 ();
 FILLCELL_X32 FILLER_180_2567 ();
 FILLCELL_X2 FILLER_180_2599 ();
 FILLCELL_X1 FILLER_180_2601 ();
 FILLCELL_X32 FILLER_181_1 ();
 FILLCELL_X32 FILLER_181_33 ();
 FILLCELL_X32 FILLER_181_65 ();
 FILLCELL_X32 FILLER_181_97 ();
 FILLCELL_X32 FILLER_181_129 ();
 FILLCELL_X32 FILLER_181_161 ();
 FILLCELL_X32 FILLER_181_193 ();
 FILLCELL_X32 FILLER_181_225 ();
 FILLCELL_X32 FILLER_181_257 ();
 FILLCELL_X32 FILLER_181_289 ();
 FILLCELL_X32 FILLER_181_321 ();
 FILLCELL_X32 FILLER_181_353 ();
 FILLCELL_X32 FILLER_181_385 ();
 FILLCELL_X32 FILLER_181_417 ();
 FILLCELL_X32 FILLER_181_449 ();
 FILLCELL_X32 FILLER_181_481 ();
 FILLCELL_X32 FILLER_181_513 ();
 FILLCELL_X32 FILLER_181_545 ();
 FILLCELL_X32 FILLER_181_577 ();
 FILLCELL_X32 FILLER_181_609 ();
 FILLCELL_X32 FILLER_181_641 ();
 FILLCELL_X32 FILLER_181_673 ();
 FILLCELL_X32 FILLER_181_705 ();
 FILLCELL_X32 FILLER_181_737 ();
 FILLCELL_X32 FILLER_181_769 ();
 FILLCELL_X32 FILLER_181_801 ();
 FILLCELL_X32 FILLER_181_833 ();
 FILLCELL_X32 FILLER_181_865 ();
 FILLCELL_X32 FILLER_181_897 ();
 FILLCELL_X32 FILLER_181_929 ();
 FILLCELL_X32 FILLER_181_961 ();
 FILLCELL_X32 FILLER_181_993 ();
 FILLCELL_X32 FILLER_181_1025 ();
 FILLCELL_X32 FILLER_181_1057 ();
 FILLCELL_X16 FILLER_181_1089 ();
 FILLCELL_X4 FILLER_181_1105 ();
 FILLCELL_X1 FILLER_181_1109 ();
 FILLCELL_X32 FILLER_181_1117 ();
 FILLCELL_X2 FILLER_181_1153 ();
 FILLCELL_X2 FILLER_181_1162 ();
 FILLCELL_X8 FILLER_181_1168 ();
 FILLCELL_X16 FILLER_181_1201 ();
 FILLCELL_X4 FILLER_181_1217 ();
 FILLCELL_X2 FILLER_181_1221 ();
 FILLCELL_X1 FILLER_181_1223 ();
 FILLCELL_X1 FILLER_181_1227 ();
 FILLCELL_X8 FILLER_181_1241 ();
 FILLCELL_X1 FILLER_181_1249 ();
 FILLCELL_X16 FILLER_181_1277 ();
 FILLCELL_X4 FILLER_181_1293 ();
 FILLCELL_X16 FILLER_181_1301 ();
 FILLCELL_X8 FILLER_181_1317 ();
 FILLCELL_X1 FILLER_181_1325 ();
 FILLCELL_X16 FILLER_181_1333 ();
 FILLCELL_X8 FILLER_181_1349 ();
 FILLCELL_X2 FILLER_181_1357 ();
 FILLCELL_X1 FILLER_181_1359 ();
 FILLCELL_X32 FILLER_181_1365 ();
 FILLCELL_X32 FILLER_181_1397 ();
 FILLCELL_X32 FILLER_181_1429 ();
 FILLCELL_X32 FILLER_181_1461 ();
 FILLCELL_X32 FILLER_181_1493 ();
 FILLCELL_X16 FILLER_181_1525 ();
 FILLCELL_X4 FILLER_181_1541 ();
 FILLCELL_X2 FILLER_181_1545 ();
 FILLCELL_X8 FILLER_181_1554 ();
 FILLCELL_X2 FILLER_181_1562 ();
 FILLCELL_X1 FILLER_181_1564 ();
 FILLCELL_X2 FILLER_181_1603 ();
 FILLCELL_X1 FILLER_181_1605 ();
 FILLCELL_X32 FILLER_181_1630 ();
 FILLCELL_X32 FILLER_181_1662 ();
 FILLCELL_X32 FILLER_181_1694 ();
 FILLCELL_X32 FILLER_181_1726 ();
 FILLCELL_X32 FILLER_181_1758 ();
 FILLCELL_X32 FILLER_181_1790 ();
 FILLCELL_X32 FILLER_181_1822 ();
 FILLCELL_X32 FILLER_181_1854 ();
 FILLCELL_X32 FILLER_181_1886 ();
 FILLCELL_X32 FILLER_181_1918 ();
 FILLCELL_X32 FILLER_181_1950 ();
 FILLCELL_X32 FILLER_181_1982 ();
 FILLCELL_X32 FILLER_181_2014 ();
 FILLCELL_X32 FILLER_181_2046 ();
 FILLCELL_X32 FILLER_181_2078 ();
 FILLCELL_X32 FILLER_181_2110 ();
 FILLCELL_X32 FILLER_181_2142 ();
 FILLCELL_X32 FILLER_181_2174 ();
 FILLCELL_X32 FILLER_181_2206 ();
 FILLCELL_X32 FILLER_181_2238 ();
 FILLCELL_X32 FILLER_181_2270 ();
 FILLCELL_X32 FILLER_181_2302 ();
 FILLCELL_X32 FILLER_181_2334 ();
 FILLCELL_X32 FILLER_181_2366 ();
 FILLCELL_X32 FILLER_181_2398 ();
 FILLCELL_X32 FILLER_181_2430 ();
 FILLCELL_X32 FILLER_181_2462 ();
 FILLCELL_X32 FILLER_181_2494 ();
 FILLCELL_X32 FILLER_181_2527 ();
 FILLCELL_X32 FILLER_181_2559 ();
 FILLCELL_X8 FILLER_181_2591 ();
 FILLCELL_X2 FILLER_181_2599 ();
 FILLCELL_X1 FILLER_181_2601 ();
 FILLCELL_X32 FILLER_182_1 ();
 FILLCELL_X32 FILLER_182_33 ();
 FILLCELL_X32 FILLER_182_65 ();
 FILLCELL_X32 FILLER_182_97 ();
 FILLCELL_X32 FILLER_182_129 ();
 FILLCELL_X32 FILLER_182_161 ();
 FILLCELL_X32 FILLER_182_193 ();
 FILLCELL_X32 FILLER_182_225 ();
 FILLCELL_X32 FILLER_182_257 ();
 FILLCELL_X32 FILLER_182_289 ();
 FILLCELL_X32 FILLER_182_321 ();
 FILLCELL_X32 FILLER_182_353 ();
 FILLCELL_X32 FILLER_182_385 ();
 FILLCELL_X32 FILLER_182_417 ();
 FILLCELL_X32 FILLER_182_449 ();
 FILLCELL_X32 FILLER_182_481 ();
 FILLCELL_X32 FILLER_182_513 ();
 FILLCELL_X32 FILLER_182_545 ();
 FILLCELL_X32 FILLER_182_577 ();
 FILLCELL_X16 FILLER_182_609 ();
 FILLCELL_X4 FILLER_182_625 ();
 FILLCELL_X2 FILLER_182_629 ();
 FILLCELL_X32 FILLER_182_632 ();
 FILLCELL_X32 FILLER_182_664 ();
 FILLCELL_X32 FILLER_182_696 ();
 FILLCELL_X32 FILLER_182_728 ();
 FILLCELL_X32 FILLER_182_760 ();
 FILLCELL_X32 FILLER_182_792 ();
 FILLCELL_X32 FILLER_182_824 ();
 FILLCELL_X32 FILLER_182_856 ();
 FILLCELL_X32 FILLER_182_888 ();
 FILLCELL_X32 FILLER_182_920 ();
 FILLCELL_X32 FILLER_182_952 ();
 FILLCELL_X32 FILLER_182_984 ();
 FILLCELL_X32 FILLER_182_1016 ();
 FILLCELL_X32 FILLER_182_1048 ();
 FILLCELL_X16 FILLER_182_1080 ();
 FILLCELL_X8 FILLER_182_1096 ();
 FILLCELL_X1 FILLER_182_1104 ();
 FILLCELL_X2 FILLER_182_1124 ();
 FILLCELL_X1 FILLER_182_1126 ();
 FILLCELL_X8 FILLER_182_1134 ();
 FILLCELL_X4 FILLER_182_1142 ();
 FILLCELL_X2 FILLER_182_1146 ();
 FILLCELL_X1 FILLER_182_1148 ();
 FILLCELL_X1 FILLER_182_1156 ();
 FILLCELL_X32 FILLER_182_1164 ();
 FILLCELL_X16 FILLER_182_1196 ();
 FILLCELL_X2 FILLER_182_1212 ();
 FILLCELL_X16 FILLER_182_1240 ();
 FILLCELL_X8 FILLER_182_1256 ();
 FILLCELL_X1 FILLER_182_1264 ();
 FILLCELL_X32 FILLER_182_1272 ();
 FILLCELL_X32 FILLER_182_1304 ();
 FILLCELL_X32 FILLER_182_1336 ();
 FILLCELL_X32 FILLER_182_1368 ();
 FILLCELL_X4 FILLER_182_1400 ();
 FILLCELL_X1 FILLER_182_1404 ();
 FILLCELL_X32 FILLER_182_1419 ();
 FILLCELL_X4 FILLER_182_1451 ();
 FILLCELL_X1 FILLER_182_1455 ();
 FILLCELL_X32 FILLER_182_1460 ();
 FILLCELL_X32 FILLER_182_1492 ();
 FILLCELL_X32 FILLER_182_1524 ();
 FILLCELL_X32 FILLER_182_1556 ();
 FILLCELL_X32 FILLER_182_1588 ();
 FILLCELL_X32 FILLER_182_1620 ();
 FILLCELL_X32 FILLER_182_1652 ();
 FILLCELL_X32 FILLER_182_1684 ();
 FILLCELL_X32 FILLER_182_1716 ();
 FILLCELL_X32 FILLER_182_1748 ();
 FILLCELL_X32 FILLER_182_1780 ();
 FILLCELL_X32 FILLER_182_1812 ();
 FILLCELL_X32 FILLER_182_1844 ();
 FILLCELL_X16 FILLER_182_1876 ();
 FILLCELL_X2 FILLER_182_1892 ();
 FILLCELL_X32 FILLER_182_1895 ();
 FILLCELL_X32 FILLER_182_1927 ();
 FILLCELL_X32 FILLER_182_1959 ();
 FILLCELL_X32 FILLER_182_1991 ();
 FILLCELL_X32 FILLER_182_2023 ();
 FILLCELL_X32 FILLER_182_2055 ();
 FILLCELL_X32 FILLER_182_2087 ();
 FILLCELL_X32 FILLER_182_2119 ();
 FILLCELL_X32 FILLER_182_2151 ();
 FILLCELL_X32 FILLER_182_2183 ();
 FILLCELL_X32 FILLER_182_2215 ();
 FILLCELL_X32 FILLER_182_2247 ();
 FILLCELL_X32 FILLER_182_2279 ();
 FILLCELL_X32 FILLER_182_2311 ();
 FILLCELL_X32 FILLER_182_2343 ();
 FILLCELL_X32 FILLER_182_2375 ();
 FILLCELL_X32 FILLER_182_2407 ();
 FILLCELL_X32 FILLER_182_2439 ();
 FILLCELL_X32 FILLER_182_2471 ();
 FILLCELL_X32 FILLER_182_2503 ();
 FILLCELL_X32 FILLER_182_2535 ();
 FILLCELL_X32 FILLER_182_2567 ();
 FILLCELL_X2 FILLER_182_2599 ();
 FILLCELL_X1 FILLER_182_2601 ();
 FILLCELL_X32 FILLER_183_1 ();
 FILLCELL_X32 FILLER_183_33 ();
 FILLCELL_X32 FILLER_183_65 ();
 FILLCELL_X32 FILLER_183_97 ();
 FILLCELL_X32 FILLER_183_129 ();
 FILLCELL_X32 FILLER_183_161 ();
 FILLCELL_X32 FILLER_183_193 ();
 FILLCELL_X32 FILLER_183_225 ();
 FILLCELL_X32 FILLER_183_257 ();
 FILLCELL_X32 FILLER_183_289 ();
 FILLCELL_X32 FILLER_183_321 ();
 FILLCELL_X32 FILLER_183_353 ();
 FILLCELL_X32 FILLER_183_385 ();
 FILLCELL_X32 FILLER_183_417 ();
 FILLCELL_X32 FILLER_183_449 ();
 FILLCELL_X32 FILLER_183_481 ();
 FILLCELL_X32 FILLER_183_513 ();
 FILLCELL_X32 FILLER_183_545 ();
 FILLCELL_X32 FILLER_183_577 ();
 FILLCELL_X32 FILLER_183_609 ();
 FILLCELL_X32 FILLER_183_641 ();
 FILLCELL_X32 FILLER_183_673 ();
 FILLCELL_X32 FILLER_183_705 ();
 FILLCELL_X32 FILLER_183_737 ();
 FILLCELL_X32 FILLER_183_769 ();
 FILLCELL_X32 FILLER_183_801 ();
 FILLCELL_X32 FILLER_183_833 ();
 FILLCELL_X32 FILLER_183_865 ();
 FILLCELL_X32 FILLER_183_897 ();
 FILLCELL_X32 FILLER_183_929 ();
 FILLCELL_X32 FILLER_183_961 ();
 FILLCELL_X32 FILLER_183_993 ();
 FILLCELL_X32 FILLER_183_1025 ();
 FILLCELL_X32 FILLER_183_1057 ();
 FILLCELL_X16 FILLER_183_1089 ();
 FILLCELL_X8 FILLER_183_1105 ();
 FILLCELL_X4 FILLER_183_1113 ();
 FILLCELL_X2 FILLER_183_1117 ();
 FILLCELL_X1 FILLER_183_1126 ();
 FILLCELL_X16 FILLER_183_1158 ();
 FILLCELL_X8 FILLER_183_1174 ();
 FILLCELL_X2 FILLER_183_1182 ();
 FILLCELL_X1 FILLER_183_1184 ();
 FILLCELL_X4 FILLER_183_1202 ();
 FILLCELL_X1 FILLER_183_1206 ();
 FILLCELL_X32 FILLER_183_1212 ();
 FILLCELL_X16 FILLER_183_1244 ();
 FILLCELL_X2 FILLER_183_1260 ();
 FILLCELL_X1 FILLER_183_1262 ();
 FILLCELL_X2 FILLER_183_1264 ();
 FILLCELL_X16 FILLER_183_1283 ();
 FILLCELL_X8 FILLER_183_1299 ();
 FILLCELL_X1 FILLER_183_1307 ();
 FILLCELL_X4 FILLER_183_1315 ();
 FILLCELL_X2 FILLER_183_1319 ();
 FILLCELL_X1 FILLER_183_1321 ();
 FILLCELL_X16 FILLER_183_1329 ();
 FILLCELL_X4 FILLER_183_1345 ();
 FILLCELL_X1 FILLER_183_1349 ();
 FILLCELL_X32 FILLER_183_1357 ();
 FILLCELL_X8 FILLER_183_1389 ();
 FILLCELL_X4 FILLER_183_1397 ();
 FILLCELL_X16 FILLER_183_1418 ();
 FILLCELL_X4 FILLER_183_1434 ();
 FILLCELL_X1 FILLER_183_1438 ();
 FILLCELL_X8 FILLER_183_1446 ();
 FILLCELL_X2 FILLER_183_1454 ();
 FILLCELL_X32 FILLER_183_1463 ();
 FILLCELL_X4 FILLER_183_1495 ();
 FILLCELL_X2 FILLER_183_1499 ();
 FILLCELL_X8 FILLER_183_1508 ();
 FILLCELL_X4 FILLER_183_1516 ();
 FILLCELL_X1 FILLER_183_1520 ();
 FILLCELL_X8 FILLER_183_1528 ();
 FILLCELL_X2 FILLER_183_1536 ();
 FILLCELL_X32 FILLER_183_1545 ();
 FILLCELL_X16 FILLER_183_1577 ();
 FILLCELL_X8 FILLER_183_1593 ();
 FILLCELL_X32 FILLER_183_1608 ();
 FILLCELL_X32 FILLER_183_1640 ();
 FILLCELL_X32 FILLER_183_1672 ();
 FILLCELL_X32 FILLER_183_1704 ();
 FILLCELL_X32 FILLER_183_1736 ();
 FILLCELL_X32 FILLER_183_1768 ();
 FILLCELL_X32 FILLER_183_1800 ();
 FILLCELL_X32 FILLER_183_1832 ();
 FILLCELL_X32 FILLER_183_1864 ();
 FILLCELL_X32 FILLER_183_1896 ();
 FILLCELL_X32 FILLER_183_1928 ();
 FILLCELL_X32 FILLER_183_1960 ();
 FILLCELL_X32 FILLER_183_1992 ();
 FILLCELL_X32 FILLER_183_2024 ();
 FILLCELL_X32 FILLER_183_2056 ();
 FILLCELL_X32 FILLER_183_2088 ();
 FILLCELL_X32 FILLER_183_2120 ();
 FILLCELL_X32 FILLER_183_2152 ();
 FILLCELL_X32 FILLER_183_2184 ();
 FILLCELL_X32 FILLER_183_2216 ();
 FILLCELL_X32 FILLER_183_2248 ();
 FILLCELL_X32 FILLER_183_2280 ();
 FILLCELL_X32 FILLER_183_2312 ();
 FILLCELL_X32 FILLER_183_2344 ();
 FILLCELL_X32 FILLER_183_2376 ();
 FILLCELL_X32 FILLER_183_2408 ();
 FILLCELL_X32 FILLER_183_2440 ();
 FILLCELL_X32 FILLER_183_2472 ();
 FILLCELL_X16 FILLER_183_2504 ();
 FILLCELL_X4 FILLER_183_2520 ();
 FILLCELL_X2 FILLER_183_2524 ();
 FILLCELL_X32 FILLER_183_2527 ();
 FILLCELL_X32 FILLER_183_2559 ();
 FILLCELL_X8 FILLER_183_2591 ();
 FILLCELL_X2 FILLER_183_2599 ();
 FILLCELL_X1 FILLER_183_2601 ();
 FILLCELL_X32 FILLER_184_1 ();
 FILLCELL_X32 FILLER_184_33 ();
 FILLCELL_X32 FILLER_184_65 ();
 FILLCELL_X32 FILLER_184_97 ();
 FILLCELL_X32 FILLER_184_129 ();
 FILLCELL_X32 FILLER_184_161 ();
 FILLCELL_X32 FILLER_184_193 ();
 FILLCELL_X32 FILLER_184_225 ();
 FILLCELL_X32 FILLER_184_257 ();
 FILLCELL_X32 FILLER_184_289 ();
 FILLCELL_X32 FILLER_184_321 ();
 FILLCELL_X32 FILLER_184_353 ();
 FILLCELL_X32 FILLER_184_385 ();
 FILLCELL_X32 FILLER_184_417 ();
 FILLCELL_X32 FILLER_184_449 ();
 FILLCELL_X32 FILLER_184_481 ();
 FILLCELL_X32 FILLER_184_513 ();
 FILLCELL_X32 FILLER_184_545 ();
 FILLCELL_X32 FILLER_184_577 ();
 FILLCELL_X16 FILLER_184_609 ();
 FILLCELL_X4 FILLER_184_625 ();
 FILLCELL_X2 FILLER_184_629 ();
 FILLCELL_X32 FILLER_184_632 ();
 FILLCELL_X32 FILLER_184_664 ();
 FILLCELL_X32 FILLER_184_696 ();
 FILLCELL_X32 FILLER_184_728 ();
 FILLCELL_X32 FILLER_184_760 ();
 FILLCELL_X32 FILLER_184_792 ();
 FILLCELL_X32 FILLER_184_824 ();
 FILLCELL_X32 FILLER_184_856 ();
 FILLCELL_X32 FILLER_184_888 ();
 FILLCELL_X32 FILLER_184_920 ();
 FILLCELL_X32 FILLER_184_952 ();
 FILLCELL_X32 FILLER_184_984 ();
 FILLCELL_X32 FILLER_184_1016 ();
 FILLCELL_X32 FILLER_184_1048 ();
 FILLCELL_X32 FILLER_184_1080 ();
 FILLCELL_X32 FILLER_184_1112 ();
 FILLCELL_X16 FILLER_184_1144 ();
 FILLCELL_X2 FILLER_184_1160 ();
 FILLCELL_X32 FILLER_184_1179 ();
 FILLCELL_X2 FILLER_184_1211 ();
 FILLCELL_X1 FILLER_184_1230 ();
 FILLCELL_X32 FILLER_184_1238 ();
 FILLCELL_X8 FILLER_184_1277 ();
 FILLCELL_X1 FILLER_184_1285 ();
 FILLCELL_X8 FILLER_184_1293 ();
 FILLCELL_X2 FILLER_184_1301 ();
 FILLCELL_X8 FILLER_184_1327 ();
 FILLCELL_X4 FILLER_184_1335 ();
 FILLCELL_X8 FILLER_184_1356 ();
 FILLCELL_X16 FILLER_184_1388 ();
 FILLCELL_X4 FILLER_184_1404 ();
 FILLCELL_X16 FILLER_184_1415 ();
 FILLCELL_X2 FILLER_184_1431 ();
 FILLCELL_X1 FILLER_184_1433 ();
 FILLCELL_X8 FILLER_184_1468 ();
 FILLCELL_X4 FILLER_184_1476 ();
 FILLCELL_X2 FILLER_184_1480 ();
 FILLCELL_X1 FILLER_184_1482 ();
 FILLCELL_X8 FILLER_184_1507 ();
 FILLCELL_X2 FILLER_184_1515 ();
 FILLCELL_X32 FILLER_184_1551 ();
 FILLCELL_X8 FILLER_184_1583 ();
 FILLCELL_X4 FILLER_184_1591 ();
 FILLCELL_X1 FILLER_184_1595 ();
 FILLCELL_X32 FILLER_184_1613 ();
 FILLCELL_X32 FILLER_184_1645 ();
 FILLCELL_X32 FILLER_184_1677 ();
 FILLCELL_X32 FILLER_184_1709 ();
 FILLCELL_X32 FILLER_184_1741 ();
 FILLCELL_X32 FILLER_184_1773 ();
 FILLCELL_X32 FILLER_184_1805 ();
 FILLCELL_X32 FILLER_184_1837 ();
 FILLCELL_X16 FILLER_184_1869 ();
 FILLCELL_X8 FILLER_184_1885 ();
 FILLCELL_X1 FILLER_184_1893 ();
 FILLCELL_X32 FILLER_184_1895 ();
 FILLCELL_X32 FILLER_184_1927 ();
 FILLCELL_X32 FILLER_184_1959 ();
 FILLCELL_X32 FILLER_184_1991 ();
 FILLCELL_X32 FILLER_184_2023 ();
 FILLCELL_X32 FILLER_184_2055 ();
 FILLCELL_X32 FILLER_184_2087 ();
 FILLCELL_X32 FILLER_184_2119 ();
 FILLCELL_X32 FILLER_184_2151 ();
 FILLCELL_X32 FILLER_184_2183 ();
 FILLCELL_X32 FILLER_184_2215 ();
 FILLCELL_X32 FILLER_184_2247 ();
 FILLCELL_X32 FILLER_184_2279 ();
 FILLCELL_X32 FILLER_184_2311 ();
 FILLCELL_X32 FILLER_184_2343 ();
 FILLCELL_X32 FILLER_184_2375 ();
 FILLCELL_X32 FILLER_184_2407 ();
 FILLCELL_X32 FILLER_184_2439 ();
 FILLCELL_X32 FILLER_184_2471 ();
 FILLCELL_X32 FILLER_184_2503 ();
 FILLCELL_X32 FILLER_184_2535 ();
 FILLCELL_X32 FILLER_184_2567 ();
 FILLCELL_X2 FILLER_184_2599 ();
 FILLCELL_X1 FILLER_184_2601 ();
 FILLCELL_X32 FILLER_185_1 ();
 FILLCELL_X32 FILLER_185_33 ();
 FILLCELL_X32 FILLER_185_65 ();
 FILLCELL_X32 FILLER_185_97 ();
 FILLCELL_X32 FILLER_185_129 ();
 FILLCELL_X32 FILLER_185_161 ();
 FILLCELL_X32 FILLER_185_193 ();
 FILLCELL_X32 FILLER_185_225 ();
 FILLCELL_X32 FILLER_185_257 ();
 FILLCELL_X32 FILLER_185_289 ();
 FILLCELL_X32 FILLER_185_321 ();
 FILLCELL_X32 FILLER_185_353 ();
 FILLCELL_X32 FILLER_185_385 ();
 FILLCELL_X32 FILLER_185_417 ();
 FILLCELL_X32 FILLER_185_449 ();
 FILLCELL_X32 FILLER_185_481 ();
 FILLCELL_X32 FILLER_185_513 ();
 FILLCELL_X32 FILLER_185_545 ();
 FILLCELL_X32 FILLER_185_577 ();
 FILLCELL_X32 FILLER_185_609 ();
 FILLCELL_X32 FILLER_185_641 ();
 FILLCELL_X32 FILLER_185_673 ();
 FILLCELL_X32 FILLER_185_705 ();
 FILLCELL_X32 FILLER_185_737 ();
 FILLCELL_X32 FILLER_185_769 ();
 FILLCELL_X32 FILLER_185_801 ();
 FILLCELL_X32 FILLER_185_833 ();
 FILLCELL_X32 FILLER_185_865 ();
 FILLCELL_X32 FILLER_185_897 ();
 FILLCELL_X32 FILLER_185_929 ();
 FILLCELL_X32 FILLER_185_961 ();
 FILLCELL_X32 FILLER_185_993 ();
 FILLCELL_X32 FILLER_185_1025 ();
 FILLCELL_X32 FILLER_185_1057 ();
 FILLCELL_X32 FILLER_185_1089 ();
 FILLCELL_X32 FILLER_185_1121 ();
 FILLCELL_X32 FILLER_185_1153 ();
 FILLCELL_X4 FILLER_185_1185 ();
 FILLCELL_X2 FILLER_185_1189 ();
 FILLCELL_X32 FILLER_185_1196 ();
 FILLCELL_X8 FILLER_185_1228 ();
 FILLCELL_X2 FILLER_185_1236 ();
 FILLCELL_X1 FILLER_185_1238 ();
 FILLCELL_X4 FILLER_185_1256 ();
 FILLCELL_X2 FILLER_185_1260 ();
 FILLCELL_X1 FILLER_185_1262 ();
 FILLCELL_X4 FILLER_185_1264 ();
 FILLCELL_X2 FILLER_185_1268 ();
 FILLCELL_X16 FILLER_185_1287 ();
 FILLCELL_X2 FILLER_185_1303 ();
 FILLCELL_X16 FILLER_185_1336 ();
 FILLCELL_X8 FILLER_185_1352 ();
 FILLCELL_X4 FILLER_185_1360 ();
 FILLCELL_X2 FILLER_185_1364 ();
 FILLCELL_X16 FILLER_185_1373 ();
 FILLCELL_X4 FILLER_185_1389 ();
 FILLCELL_X2 FILLER_185_1393 ();
 FILLCELL_X32 FILLER_185_1419 ();
 FILLCELL_X8 FILLER_185_1451 ();
 FILLCELL_X4 FILLER_185_1459 ();
 FILLCELL_X1 FILLER_185_1463 ();
 FILLCELL_X8 FILLER_185_1471 ();
 FILLCELL_X4 FILLER_185_1479 ();
 FILLCELL_X1 FILLER_185_1483 ();
 FILLCELL_X1 FILLER_185_1501 ();
 FILLCELL_X16 FILLER_185_1509 ();
 FILLCELL_X4 FILLER_185_1525 ();
 FILLCELL_X2 FILLER_185_1529 ();
 FILLCELL_X1 FILLER_185_1531 ();
 FILLCELL_X16 FILLER_185_1539 ();
 FILLCELL_X2 FILLER_185_1555 ();
 FILLCELL_X8 FILLER_185_1564 ();
 FILLCELL_X2 FILLER_185_1572 ();
 FILLCELL_X4 FILLER_185_1605 ();
 FILLCELL_X32 FILLER_185_1616 ();
 FILLCELL_X32 FILLER_185_1648 ();
 FILLCELL_X32 FILLER_185_1680 ();
 FILLCELL_X32 FILLER_185_1712 ();
 FILLCELL_X32 FILLER_185_1744 ();
 FILLCELL_X32 FILLER_185_1776 ();
 FILLCELL_X32 FILLER_185_1808 ();
 FILLCELL_X32 FILLER_185_1840 ();
 FILLCELL_X32 FILLER_185_1872 ();
 FILLCELL_X32 FILLER_185_1904 ();
 FILLCELL_X32 FILLER_185_1936 ();
 FILLCELL_X32 FILLER_185_1968 ();
 FILLCELL_X32 FILLER_185_2000 ();
 FILLCELL_X32 FILLER_185_2032 ();
 FILLCELL_X32 FILLER_185_2064 ();
 FILLCELL_X32 FILLER_185_2096 ();
 FILLCELL_X32 FILLER_185_2128 ();
 FILLCELL_X32 FILLER_185_2160 ();
 FILLCELL_X32 FILLER_185_2192 ();
 FILLCELL_X32 FILLER_185_2224 ();
 FILLCELL_X32 FILLER_185_2256 ();
 FILLCELL_X32 FILLER_185_2288 ();
 FILLCELL_X32 FILLER_185_2320 ();
 FILLCELL_X32 FILLER_185_2352 ();
 FILLCELL_X32 FILLER_185_2384 ();
 FILLCELL_X32 FILLER_185_2416 ();
 FILLCELL_X32 FILLER_185_2448 ();
 FILLCELL_X32 FILLER_185_2480 ();
 FILLCELL_X8 FILLER_185_2512 ();
 FILLCELL_X4 FILLER_185_2520 ();
 FILLCELL_X2 FILLER_185_2524 ();
 FILLCELL_X32 FILLER_185_2527 ();
 FILLCELL_X32 FILLER_185_2559 ();
 FILLCELL_X8 FILLER_185_2591 ();
 FILLCELL_X2 FILLER_185_2599 ();
 FILLCELL_X1 FILLER_185_2601 ();
 FILLCELL_X32 FILLER_186_1 ();
 FILLCELL_X32 FILLER_186_33 ();
 FILLCELL_X32 FILLER_186_65 ();
 FILLCELL_X32 FILLER_186_97 ();
 FILLCELL_X32 FILLER_186_129 ();
 FILLCELL_X32 FILLER_186_161 ();
 FILLCELL_X32 FILLER_186_193 ();
 FILLCELL_X32 FILLER_186_225 ();
 FILLCELL_X32 FILLER_186_257 ();
 FILLCELL_X32 FILLER_186_289 ();
 FILLCELL_X32 FILLER_186_321 ();
 FILLCELL_X32 FILLER_186_353 ();
 FILLCELL_X32 FILLER_186_385 ();
 FILLCELL_X32 FILLER_186_417 ();
 FILLCELL_X32 FILLER_186_449 ();
 FILLCELL_X32 FILLER_186_481 ();
 FILLCELL_X32 FILLER_186_513 ();
 FILLCELL_X32 FILLER_186_545 ();
 FILLCELL_X32 FILLER_186_577 ();
 FILLCELL_X16 FILLER_186_609 ();
 FILLCELL_X4 FILLER_186_625 ();
 FILLCELL_X2 FILLER_186_629 ();
 FILLCELL_X32 FILLER_186_632 ();
 FILLCELL_X32 FILLER_186_664 ();
 FILLCELL_X32 FILLER_186_696 ();
 FILLCELL_X32 FILLER_186_728 ();
 FILLCELL_X32 FILLER_186_760 ();
 FILLCELL_X32 FILLER_186_792 ();
 FILLCELL_X32 FILLER_186_824 ();
 FILLCELL_X32 FILLER_186_856 ();
 FILLCELL_X32 FILLER_186_888 ();
 FILLCELL_X32 FILLER_186_920 ();
 FILLCELL_X32 FILLER_186_952 ();
 FILLCELL_X32 FILLER_186_984 ();
 FILLCELL_X32 FILLER_186_1016 ();
 FILLCELL_X32 FILLER_186_1048 ();
 FILLCELL_X32 FILLER_186_1080 ();
 FILLCELL_X32 FILLER_186_1112 ();
 FILLCELL_X32 FILLER_186_1144 ();
 FILLCELL_X32 FILLER_186_1176 ();
 FILLCELL_X32 FILLER_186_1208 ();
 FILLCELL_X4 FILLER_186_1240 ();
 FILLCELL_X2 FILLER_186_1244 ();
 FILLCELL_X1 FILLER_186_1253 ();
 FILLCELL_X32 FILLER_186_1259 ();
 FILLCELL_X32 FILLER_186_1291 ();
 FILLCELL_X16 FILLER_186_1323 ();
 FILLCELL_X1 FILLER_186_1339 ();
 FILLCELL_X16 FILLER_186_1347 ();
 FILLCELL_X8 FILLER_186_1363 ();
 FILLCELL_X32 FILLER_186_1385 ();
 FILLCELL_X1 FILLER_186_1417 ();
 FILLCELL_X16 FILLER_186_1432 ();
 FILLCELL_X8 FILLER_186_1448 ();
 FILLCELL_X4 FILLER_186_1456 ();
 FILLCELL_X2 FILLER_186_1460 ();
 FILLCELL_X1 FILLER_186_1462 ();
 FILLCELL_X2 FILLER_186_1470 ();
 FILLCELL_X32 FILLER_186_1479 ();
 FILLCELL_X16 FILLER_186_1511 ();
 FILLCELL_X4 FILLER_186_1527 ();
 FILLCELL_X2 FILLER_186_1531 ();
 FILLCELL_X8 FILLER_186_1540 ();
 FILLCELL_X1 FILLER_186_1548 ();
 FILLCELL_X4 FILLER_186_1573 ();
 FILLCELL_X2 FILLER_186_1584 ();
 FILLCELL_X4 FILLER_186_1593 ();
 FILLCELL_X1 FILLER_186_1597 ();
 FILLCELL_X32 FILLER_186_1615 ();
 FILLCELL_X32 FILLER_186_1647 ();
 FILLCELL_X32 FILLER_186_1679 ();
 FILLCELL_X32 FILLER_186_1711 ();
 FILLCELL_X32 FILLER_186_1743 ();
 FILLCELL_X32 FILLER_186_1775 ();
 FILLCELL_X32 FILLER_186_1807 ();
 FILLCELL_X32 FILLER_186_1839 ();
 FILLCELL_X16 FILLER_186_1871 ();
 FILLCELL_X4 FILLER_186_1887 ();
 FILLCELL_X2 FILLER_186_1891 ();
 FILLCELL_X1 FILLER_186_1893 ();
 FILLCELL_X32 FILLER_186_1895 ();
 FILLCELL_X32 FILLER_186_1927 ();
 FILLCELL_X32 FILLER_186_1959 ();
 FILLCELL_X32 FILLER_186_1991 ();
 FILLCELL_X32 FILLER_186_2023 ();
 FILLCELL_X32 FILLER_186_2055 ();
 FILLCELL_X32 FILLER_186_2087 ();
 FILLCELL_X32 FILLER_186_2119 ();
 FILLCELL_X32 FILLER_186_2151 ();
 FILLCELL_X32 FILLER_186_2183 ();
 FILLCELL_X32 FILLER_186_2215 ();
 FILLCELL_X32 FILLER_186_2247 ();
 FILLCELL_X32 FILLER_186_2279 ();
 FILLCELL_X32 FILLER_186_2311 ();
 FILLCELL_X32 FILLER_186_2343 ();
 FILLCELL_X32 FILLER_186_2375 ();
 FILLCELL_X32 FILLER_186_2407 ();
 FILLCELL_X32 FILLER_186_2439 ();
 FILLCELL_X32 FILLER_186_2471 ();
 FILLCELL_X32 FILLER_186_2503 ();
 FILLCELL_X32 FILLER_186_2535 ();
 FILLCELL_X32 FILLER_186_2567 ();
 FILLCELL_X2 FILLER_186_2599 ();
 FILLCELL_X1 FILLER_186_2601 ();
 FILLCELL_X32 FILLER_187_1 ();
 FILLCELL_X32 FILLER_187_33 ();
 FILLCELL_X32 FILLER_187_65 ();
 FILLCELL_X32 FILLER_187_97 ();
 FILLCELL_X32 FILLER_187_129 ();
 FILLCELL_X32 FILLER_187_161 ();
 FILLCELL_X32 FILLER_187_193 ();
 FILLCELL_X32 FILLER_187_225 ();
 FILLCELL_X32 FILLER_187_257 ();
 FILLCELL_X32 FILLER_187_289 ();
 FILLCELL_X32 FILLER_187_321 ();
 FILLCELL_X32 FILLER_187_353 ();
 FILLCELL_X32 FILLER_187_385 ();
 FILLCELL_X32 FILLER_187_417 ();
 FILLCELL_X32 FILLER_187_449 ();
 FILLCELL_X32 FILLER_187_481 ();
 FILLCELL_X32 FILLER_187_513 ();
 FILLCELL_X32 FILLER_187_545 ();
 FILLCELL_X32 FILLER_187_577 ();
 FILLCELL_X32 FILLER_187_609 ();
 FILLCELL_X32 FILLER_187_641 ();
 FILLCELL_X32 FILLER_187_673 ();
 FILLCELL_X32 FILLER_187_705 ();
 FILLCELL_X32 FILLER_187_737 ();
 FILLCELL_X32 FILLER_187_769 ();
 FILLCELL_X32 FILLER_187_801 ();
 FILLCELL_X32 FILLER_187_833 ();
 FILLCELL_X32 FILLER_187_865 ();
 FILLCELL_X32 FILLER_187_897 ();
 FILLCELL_X32 FILLER_187_929 ();
 FILLCELL_X32 FILLER_187_961 ();
 FILLCELL_X32 FILLER_187_993 ();
 FILLCELL_X32 FILLER_187_1025 ();
 FILLCELL_X32 FILLER_187_1057 ();
 FILLCELL_X32 FILLER_187_1089 ();
 FILLCELL_X32 FILLER_187_1121 ();
 FILLCELL_X32 FILLER_187_1153 ();
 FILLCELL_X32 FILLER_187_1185 ();
 FILLCELL_X4 FILLER_187_1227 ();
 FILLCELL_X1 FILLER_187_1231 ();
 FILLCELL_X2 FILLER_187_1249 ();
 FILLCELL_X1 FILLER_187_1251 ();
 FILLCELL_X1 FILLER_187_1262 ();
 FILLCELL_X8 FILLER_187_1264 ();
 FILLCELL_X2 FILLER_187_1272 ();
 FILLCELL_X32 FILLER_187_1281 ();
 FILLCELL_X16 FILLER_187_1313 ();
 FILLCELL_X8 FILLER_187_1329 ();
 FILLCELL_X4 FILLER_187_1337 ();
 FILLCELL_X4 FILLER_187_1358 ();
 FILLCELL_X2 FILLER_187_1362 ();
 FILLCELL_X32 FILLER_187_1371 ();
 FILLCELL_X32 FILLER_187_1403 ();
 FILLCELL_X16 FILLER_187_1435 ();
 FILLCELL_X4 FILLER_187_1451 ();
 FILLCELL_X2 FILLER_187_1455 ();
 FILLCELL_X1 FILLER_187_1457 ();
 FILLCELL_X32 FILLER_187_1465 ();
 FILLCELL_X32 FILLER_187_1497 ();
 FILLCELL_X4 FILLER_187_1529 ();
 FILLCELL_X8 FILLER_187_1540 ();
 FILLCELL_X2 FILLER_187_1548 ();
 FILLCELL_X16 FILLER_187_1553 ();
 FILLCELL_X4 FILLER_187_1569 ();
 FILLCELL_X2 FILLER_187_1573 ();
 FILLCELL_X1 FILLER_187_1575 ();
 FILLCELL_X32 FILLER_187_1583 ();
 FILLCELL_X32 FILLER_187_1615 ();
 FILLCELL_X32 FILLER_187_1647 ();
 FILLCELL_X32 FILLER_187_1679 ();
 FILLCELL_X32 FILLER_187_1711 ();
 FILLCELL_X32 FILLER_187_1743 ();
 FILLCELL_X32 FILLER_187_1775 ();
 FILLCELL_X32 FILLER_187_1807 ();
 FILLCELL_X32 FILLER_187_1839 ();
 FILLCELL_X32 FILLER_187_1871 ();
 FILLCELL_X32 FILLER_187_1903 ();
 FILLCELL_X32 FILLER_187_1935 ();
 FILLCELL_X32 FILLER_187_1967 ();
 FILLCELL_X32 FILLER_187_1999 ();
 FILLCELL_X32 FILLER_187_2031 ();
 FILLCELL_X32 FILLER_187_2063 ();
 FILLCELL_X32 FILLER_187_2095 ();
 FILLCELL_X32 FILLER_187_2127 ();
 FILLCELL_X32 FILLER_187_2159 ();
 FILLCELL_X32 FILLER_187_2191 ();
 FILLCELL_X32 FILLER_187_2223 ();
 FILLCELL_X32 FILLER_187_2255 ();
 FILLCELL_X32 FILLER_187_2287 ();
 FILLCELL_X32 FILLER_187_2319 ();
 FILLCELL_X32 FILLER_187_2351 ();
 FILLCELL_X32 FILLER_187_2383 ();
 FILLCELL_X32 FILLER_187_2415 ();
 FILLCELL_X32 FILLER_187_2447 ();
 FILLCELL_X32 FILLER_187_2479 ();
 FILLCELL_X8 FILLER_187_2511 ();
 FILLCELL_X4 FILLER_187_2519 ();
 FILLCELL_X2 FILLER_187_2523 ();
 FILLCELL_X1 FILLER_187_2525 ();
 FILLCELL_X32 FILLER_187_2527 ();
 FILLCELL_X32 FILLER_187_2559 ();
 FILLCELL_X8 FILLER_187_2591 ();
 FILLCELL_X2 FILLER_187_2599 ();
 FILLCELL_X1 FILLER_187_2601 ();
 FILLCELL_X32 FILLER_188_1 ();
 FILLCELL_X32 FILLER_188_33 ();
 FILLCELL_X32 FILLER_188_65 ();
 FILLCELL_X32 FILLER_188_97 ();
 FILLCELL_X32 FILLER_188_129 ();
 FILLCELL_X32 FILLER_188_161 ();
 FILLCELL_X32 FILLER_188_193 ();
 FILLCELL_X32 FILLER_188_225 ();
 FILLCELL_X32 FILLER_188_257 ();
 FILLCELL_X32 FILLER_188_289 ();
 FILLCELL_X32 FILLER_188_321 ();
 FILLCELL_X32 FILLER_188_353 ();
 FILLCELL_X32 FILLER_188_385 ();
 FILLCELL_X32 FILLER_188_417 ();
 FILLCELL_X32 FILLER_188_449 ();
 FILLCELL_X32 FILLER_188_481 ();
 FILLCELL_X32 FILLER_188_513 ();
 FILLCELL_X32 FILLER_188_545 ();
 FILLCELL_X32 FILLER_188_577 ();
 FILLCELL_X16 FILLER_188_609 ();
 FILLCELL_X4 FILLER_188_625 ();
 FILLCELL_X2 FILLER_188_629 ();
 FILLCELL_X32 FILLER_188_632 ();
 FILLCELL_X32 FILLER_188_664 ();
 FILLCELL_X32 FILLER_188_696 ();
 FILLCELL_X32 FILLER_188_728 ();
 FILLCELL_X32 FILLER_188_760 ();
 FILLCELL_X32 FILLER_188_792 ();
 FILLCELL_X32 FILLER_188_824 ();
 FILLCELL_X32 FILLER_188_856 ();
 FILLCELL_X32 FILLER_188_888 ();
 FILLCELL_X32 FILLER_188_920 ();
 FILLCELL_X32 FILLER_188_952 ();
 FILLCELL_X32 FILLER_188_984 ();
 FILLCELL_X32 FILLER_188_1016 ();
 FILLCELL_X32 FILLER_188_1048 ();
 FILLCELL_X32 FILLER_188_1080 ();
 FILLCELL_X32 FILLER_188_1112 ();
 FILLCELL_X32 FILLER_188_1144 ();
 FILLCELL_X32 FILLER_188_1176 ();
 FILLCELL_X32 FILLER_188_1208 ();
 FILLCELL_X4 FILLER_188_1240 ();
 FILLCELL_X1 FILLER_188_1244 ();
 FILLCELL_X8 FILLER_188_1252 ();
 FILLCELL_X4 FILLER_188_1260 ();
 FILLCELL_X2 FILLER_188_1264 ();
 FILLCELL_X16 FILLER_188_1282 ();
 FILLCELL_X8 FILLER_188_1298 ();
 FILLCELL_X1 FILLER_188_1306 ();
 FILLCELL_X1 FILLER_188_1314 ();
 FILLCELL_X2 FILLER_188_1322 ();
 FILLCELL_X1 FILLER_188_1324 ();
 FILLCELL_X16 FILLER_188_1334 ();
 FILLCELL_X4 FILLER_188_1350 ();
 FILLCELL_X16 FILLER_188_1378 ();
 FILLCELL_X4 FILLER_188_1394 ();
 FILLCELL_X2 FILLER_188_1398 ();
 FILLCELL_X1 FILLER_188_1400 ();
 FILLCELL_X8 FILLER_188_1408 ();
 FILLCELL_X4 FILLER_188_1416 ();
 FILLCELL_X1 FILLER_188_1420 ();
 FILLCELL_X4 FILLER_188_1445 ();
 FILLCELL_X2 FILLER_188_1449 ();
 FILLCELL_X32 FILLER_188_1468 ();
 FILLCELL_X16 FILLER_188_1500 ();
 FILLCELL_X4 FILLER_188_1516 ();
 FILLCELL_X16 FILLER_188_1527 ();
 FILLCELL_X1 FILLER_188_1543 ();
 FILLCELL_X2 FILLER_188_1548 ();
 FILLCELL_X2 FILLER_188_1560 ();
 FILLCELL_X1 FILLER_188_1562 ();
 FILLCELL_X32 FILLER_188_1570 ();
 FILLCELL_X32 FILLER_188_1602 ();
 FILLCELL_X32 FILLER_188_1634 ();
 FILLCELL_X32 FILLER_188_1666 ();
 FILLCELL_X32 FILLER_188_1698 ();
 FILLCELL_X32 FILLER_188_1730 ();
 FILLCELL_X32 FILLER_188_1762 ();
 FILLCELL_X32 FILLER_188_1794 ();
 FILLCELL_X32 FILLER_188_1826 ();
 FILLCELL_X32 FILLER_188_1858 ();
 FILLCELL_X4 FILLER_188_1890 ();
 FILLCELL_X32 FILLER_188_1895 ();
 FILLCELL_X32 FILLER_188_1927 ();
 FILLCELL_X32 FILLER_188_1959 ();
 FILLCELL_X32 FILLER_188_1991 ();
 FILLCELL_X32 FILLER_188_2023 ();
 FILLCELL_X32 FILLER_188_2055 ();
 FILLCELL_X32 FILLER_188_2087 ();
 FILLCELL_X32 FILLER_188_2119 ();
 FILLCELL_X32 FILLER_188_2151 ();
 FILLCELL_X32 FILLER_188_2183 ();
 FILLCELL_X32 FILLER_188_2215 ();
 FILLCELL_X32 FILLER_188_2247 ();
 FILLCELL_X32 FILLER_188_2279 ();
 FILLCELL_X32 FILLER_188_2311 ();
 FILLCELL_X32 FILLER_188_2343 ();
 FILLCELL_X32 FILLER_188_2375 ();
 FILLCELL_X32 FILLER_188_2407 ();
 FILLCELL_X32 FILLER_188_2439 ();
 FILLCELL_X32 FILLER_188_2471 ();
 FILLCELL_X32 FILLER_188_2503 ();
 FILLCELL_X32 FILLER_188_2535 ();
 FILLCELL_X32 FILLER_188_2567 ();
 FILLCELL_X2 FILLER_188_2599 ();
 FILLCELL_X1 FILLER_188_2601 ();
 FILLCELL_X32 FILLER_189_1 ();
 FILLCELL_X32 FILLER_189_33 ();
 FILLCELL_X32 FILLER_189_65 ();
 FILLCELL_X32 FILLER_189_97 ();
 FILLCELL_X32 FILLER_189_129 ();
 FILLCELL_X32 FILLER_189_161 ();
 FILLCELL_X32 FILLER_189_193 ();
 FILLCELL_X32 FILLER_189_225 ();
 FILLCELL_X32 FILLER_189_257 ();
 FILLCELL_X32 FILLER_189_289 ();
 FILLCELL_X32 FILLER_189_321 ();
 FILLCELL_X32 FILLER_189_353 ();
 FILLCELL_X32 FILLER_189_385 ();
 FILLCELL_X32 FILLER_189_417 ();
 FILLCELL_X32 FILLER_189_449 ();
 FILLCELL_X32 FILLER_189_481 ();
 FILLCELL_X32 FILLER_189_513 ();
 FILLCELL_X32 FILLER_189_545 ();
 FILLCELL_X32 FILLER_189_577 ();
 FILLCELL_X32 FILLER_189_609 ();
 FILLCELL_X32 FILLER_189_641 ();
 FILLCELL_X32 FILLER_189_673 ();
 FILLCELL_X32 FILLER_189_705 ();
 FILLCELL_X32 FILLER_189_737 ();
 FILLCELL_X32 FILLER_189_769 ();
 FILLCELL_X32 FILLER_189_801 ();
 FILLCELL_X32 FILLER_189_833 ();
 FILLCELL_X32 FILLER_189_865 ();
 FILLCELL_X32 FILLER_189_897 ();
 FILLCELL_X32 FILLER_189_929 ();
 FILLCELL_X32 FILLER_189_961 ();
 FILLCELL_X32 FILLER_189_993 ();
 FILLCELL_X32 FILLER_189_1025 ();
 FILLCELL_X32 FILLER_189_1057 ();
 FILLCELL_X32 FILLER_189_1089 ();
 FILLCELL_X32 FILLER_189_1121 ();
 FILLCELL_X32 FILLER_189_1153 ();
 FILLCELL_X32 FILLER_189_1185 ();
 FILLCELL_X32 FILLER_189_1217 ();
 FILLCELL_X4 FILLER_189_1249 ();
 FILLCELL_X1 FILLER_189_1253 ();
 FILLCELL_X4 FILLER_189_1258 ();
 FILLCELL_X1 FILLER_189_1262 ();
 FILLCELL_X16 FILLER_189_1264 ();
 FILLCELL_X8 FILLER_189_1280 ();
 FILLCELL_X2 FILLER_189_1288 ();
 FILLCELL_X32 FILLER_189_1329 ();
 FILLCELL_X16 FILLER_189_1361 ();
 FILLCELL_X8 FILLER_189_1377 ();
 FILLCELL_X4 FILLER_189_1385 ();
 FILLCELL_X4 FILLER_189_1406 ();
 FILLCELL_X2 FILLER_189_1410 ();
 FILLCELL_X32 FILLER_189_1419 ();
 FILLCELL_X4 FILLER_189_1451 ();
 FILLCELL_X2 FILLER_189_1455 ();
 FILLCELL_X1 FILLER_189_1457 ();
 FILLCELL_X16 FILLER_189_1465 ();
 FILLCELL_X8 FILLER_189_1481 ();
 FILLCELL_X4 FILLER_189_1489 ();
 FILLCELL_X1 FILLER_189_1517 ();
 FILLCELL_X8 FILLER_189_1552 ();
 FILLCELL_X1 FILLER_189_1560 ();
 FILLCELL_X32 FILLER_189_1585 ();
 FILLCELL_X32 FILLER_189_1617 ();
 FILLCELL_X32 FILLER_189_1649 ();
 FILLCELL_X32 FILLER_189_1681 ();
 FILLCELL_X32 FILLER_189_1713 ();
 FILLCELL_X32 FILLER_189_1745 ();
 FILLCELL_X32 FILLER_189_1777 ();
 FILLCELL_X32 FILLER_189_1809 ();
 FILLCELL_X32 FILLER_189_1841 ();
 FILLCELL_X32 FILLER_189_1873 ();
 FILLCELL_X32 FILLER_189_1905 ();
 FILLCELL_X32 FILLER_189_1937 ();
 FILLCELL_X32 FILLER_189_1969 ();
 FILLCELL_X32 FILLER_189_2001 ();
 FILLCELL_X32 FILLER_189_2033 ();
 FILLCELL_X32 FILLER_189_2065 ();
 FILLCELL_X32 FILLER_189_2097 ();
 FILLCELL_X32 FILLER_189_2129 ();
 FILLCELL_X32 FILLER_189_2161 ();
 FILLCELL_X32 FILLER_189_2193 ();
 FILLCELL_X32 FILLER_189_2225 ();
 FILLCELL_X32 FILLER_189_2257 ();
 FILLCELL_X32 FILLER_189_2289 ();
 FILLCELL_X32 FILLER_189_2321 ();
 FILLCELL_X32 FILLER_189_2353 ();
 FILLCELL_X32 FILLER_189_2385 ();
 FILLCELL_X32 FILLER_189_2417 ();
 FILLCELL_X32 FILLER_189_2449 ();
 FILLCELL_X32 FILLER_189_2481 ();
 FILLCELL_X8 FILLER_189_2513 ();
 FILLCELL_X4 FILLER_189_2521 ();
 FILLCELL_X1 FILLER_189_2525 ();
 FILLCELL_X32 FILLER_189_2527 ();
 FILLCELL_X32 FILLER_189_2559 ();
 FILLCELL_X8 FILLER_189_2591 ();
 FILLCELL_X2 FILLER_189_2599 ();
 FILLCELL_X1 FILLER_189_2601 ();
 FILLCELL_X32 FILLER_190_1 ();
 FILLCELL_X32 FILLER_190_33 ();
 FILLCELL_X32 FILLER_190_65 ();
 FILLCELL_X32 FILLER_190_97 ();
 FILLCELL_X32 FILLER_190_129 ();
 FILLCELL_X32 FILLER_190_161 ();
 FILLCELL_X32 FILLER_190_193 ();
 FILLCELL_X32 FILLER_190_225 ();
 FILLCELL_X32 FILLER_190_257 ();
 FILLCELL_X32 FILLER_190_289 ();
 FILLCELL_X32 FILLER_190_321 ();
 FILLCELL_X32 FILLER_190_353 ();
 FILLCELL_X32 FILLER_190_385 ();
 FILLCELL_X32 FILLER_190_417 ();
 FILLCELL_X32 FILLER_190_449 ();
 FILLCELL_X32 FILLER_190_481 ();
 FILLCELL_X32 FILLER_190_513 ();
 FILLCELL_X32 FILLER_190_545 ();
 FILLCELL_X32 FILLER_190_577 ();
 FILLCELL_X16 FILLER_190_609 ();
 FILLCELL_X4 FILLER_190_625 ();
 FILLCELL_X2 FILLER_190_629 ();
 FILLCELL_X32 FILLER_190_632 ();
 FILLCELL_X32 FILLER_190_664 ();
 FILLCELL_X32 FILLER_190_696 ();
 FILLCELL_X32 FILLER_190_728 ();
 FILLCELL_X32 FILLER_190_760 ();
 FILLCELL_X32 FILLER_190_792 ();
 FILLCELL_X32 FILLER_190_824 ();
 FILLCELL_X32 FILLER_190_856 ();
 FILLCELL_X32 FILLER_190_888 ();
 FILLCELL_X32 FILLER_190_920 ();
 FILLCELL_X32 FILLER_190_952 ();
 FILLCELL_X32 FILLER_190_984 ();
 FILLCELL_X32 FILLER_190_1016 ();
 FILLCELL_X32 FILLER_190_1048 ();
 FILLCELL_X32 FILLER_190_1080 ();
 FILLCELL_X32 FILLER_190_1112 ();
 FILLCELL_X32 FILLER_190_1144 ();
 FILLCELL_X32 FILLER_190_1176 ();
 FILLCELL_X32 FILLER_190_1208 ();
 FILLCELL_X8 FILLER_190_1240 ();
 FILLCELL_X4 FILLER_190_1248 ();
 FILLCELL_X2 FILLER_190_1252 ();
 FILLCELL_X4 FILLER_190_1278 ();
 FILLCELL_X1 FILLER_190_1282 ();
 FILLCELL_X32 FILLER_190_1321 ();
 FILLCELL_X32 FILLER_190_1353 ();
 FILLCELL_X16 FILLER_190_1385 ();
 FILLCELL_X4 FILLER_190_1401 ();
 FILLCELL_X1 FILLER_190_1405 ();
 FILLCELL_X16 FILLER_190_1430 ();
 FILLCELL_X4 FILLER_190_1446 ();
 FILLCELL_X2 FILLER_190_1450 ();
 FILLCELL_X16 FILLER_190_1465 ();
 FILLCELL_X16 FILLER_190_1512 ();
 FILLCELL_X2 FILLER_190_1528 ();
 FILLCELL_X1 FILLER_190_1530 ();
 FILLCELL_X16 FILLER_190_1555 ();
 FILLCELL_X4 FILLER_190_1571 ();
 FILLCELL_X2 FILLER_190_1575 ();
 FILLCELL_X1 FILLER_190_1577 ();
 FILLCELL_X32 FILLER_190_1602 ();
 FILLCELL_X32 FILLER_190_1634 ();
 FILLCELL_X32 FILLER_190_1666 ();
 FILLCELL_X32 FILLER_190_1698 ();
 FILLCELL_X32 FILLER_190_1730 ();
 FILLCELL_X32 FILLER_190_1762 ();
 FILLCELL_X32 FILLER_190_1794 ();
 FILLCELL_X32 FILLER_190_1826 ();
 FILLCELL_X32 FILLER_190_1858 ();
 FILLCELL_X4 FILLER_190_1890 ();
 FILLCELL_X32 FILLER_190_1895 ();
 FILLCELL_X32 FILLER_190_1927 ();
 FILLCELL_X32 FILLER_190_1959 ();
 FILLCELL_X32 FILLER_190_1991 ();
 FILLCELL_X32 FILLER_190_2023 ();
 FILLCELL_X32 FILLER_190_2055 ();
 FILLCELL_X32 FILLER_190_2087 ();
 FILLCELL_X32 FILLER_190_2119 ();
 FILLCELL_X32 FILLER_190_2151 ();
 FILLCELL_X32 FILLER_190_2183 ();
 FILLCELL_X32 FILLER_190_2215 ();
 FILLCELL_X32 FILLER_190_2247 ();
 FILLCELL_X32 FILLER_190_2279 ();
 FILLCELL_X32 FILLER_190_2311 ();
 FILLCELL_X32 FILLER_190_2343 ();
 FILLCELL_X32 FILLER_190_2375 ();
 FILLCELL_X32 FILLER_190_2407 ();
 FILLCELL_X32 FILLER_190_2439 ();
 FILLCELL_X32 FILLER_190_2471 ();
 FILLCELL_X32 FILLER_190_2503 ();
 FILLCELL_X32 FILLER_190_2535 ();
 FILLCELL_X32 FILLER_190_2567 ();
 FILLCELL_X2 FILLER_190_2599 ();
 FILLCELL_X1 FILLER_190_2601 ();
 FILLCELL_X32 FILLER_191_1 ();
 FILLCELL_X32 FILLER_191_33 ();
 FILLCELL_X32 FILLER_191_65 ();
 FILLCELL_X32 FILLER_191_97 ();
 FILLCELL_X32 FILLER_191_129 ();
 FILLCELL_X32 FILLER_191_161 ();
 FILLCELL_X32 FILLER_191_193 ();
 FILLCELL_X32 FILLER_191_225 ();
 FILLCELL_X32 FILLER_191_257 ();
 FILLCELL_X32 FILLER_191_289 ();
 FILLCELL_X32 FILLER_191_321 ();
 FILLCELL_X32 FILLER_191_353 ();
 FILLCELL_X32 FILLER_191_385 ();
 FILLCELL_X32 FILLER_191_417 ();
 FILLCELL_X32 FILLER_191_449 ();
 FILLCELL_X32 FILLER_191_481 ();
 FILLCELL_X32 FILLER_191_513 ();
 FILLCELL_X32 FILLER_191_545 ();
 FILLCELL_X32 FILLER_191_577 ();
 FILLCELL_X32 FILLER_191_609 ();
 FILLCELL_X32 FILLER_191_641 ();
 FILLCELL_X32 FILLER_191_673 ();
 FILLCELL_X32 FILLER_191_705 ();
 FILLCELL_X32 FILLER_191_737 ();
 FILLCELL_X32 FILLER_191_769 ();
 FILLCELL_X32 FILLER_191_801 ();
 FILLCELL_X32 FILLER_191_833 ();
 FILLCELL_X32 FILLER_191_865 ();
 FILLCELL_X32 FILLER_191_897 ();
 FILLCELL_X32 FILLER_191_929 ();
 FILLCELL_X32 FILLER_191_961 ();
 FILLCELL_X32 FILLER_191_993 ();
 FILLCELL_X32 FILLER_191_1025 ();
 FILLCELL_X32 FILLER_191_1057 ();
 FILLCELL_X32 FILLER_191_1089 ();
 FILLCELL_X32 FILLER_191_1121 ();
 FILLCELL_X32 FILLER_191_1153 ();
 FILLCELL_X32 FILLER_191_1185 ();
 FILLCELL_X16 FILLER_191_1217 ();
 FILLCELL_X2 FILLER_191_1233 ();
 FILLCELL_X1 FILLER_191_1235 ();
 FILLCELL_X16 FILLER_191_1243 ();
 FILLCELL_X4 FILLER_191_1259 ();
 FILLCELL_X32 FILLER_191_1264 ();
 FILLCELL_X32 FILLER_191_1296 ();
 FILLCELL_X16 FILLER_191_1328 ();
 FILLCELL_X8 FILLER_191_1344 ();
 FILLCELL_X4 FILLER_191_1352 ();
 FILLCELL_X2 FILLER_191_1356 ();
 FILLCELL_X1 FILLER_191_1358 ();
 FILLCELL_X32 FILLER_191_1363 ();
 FILLCELL_X8 FILLER_191_1395 ();
 FILLCELL_X4 FILLER_191_1403 ();
 FILLCELL_X2 FILLER_191_1407 ();
 FILLCELL_X1 FILLER_191_1409 ();
 FILLCELL_X32 FILLER_191_1414 ();
 FILLCELL_X8 FILLER_191_1446 ();
 FILLCELL_X1 FILLER_191_1454 ();
 FILLCELL_X32 FILLER_191_1469 ();
 FILLCELL_X32 FILLER_191_1501 ();
 FILLCELL_X32 FILLER_191_1533 ();
 FILLCELL_X32 FILLER_191_1565 ();
 FILLCELL_X32 FILLER_191_1597 ();
 FILLCELL_X32 FILLER_191_1629 ();
 FILLCELL_X32 FILLER_191_1661 ();
 FILLCELL_X32 FILLER_191_1693 ();
 FILLCELL_X32 FILLER_191_1725 ();
 FILLCELL_X32 FILLER_191_1757 ();
 FILLCELL_X32 FILLER_191_1789 ();
 FILLCELL_X32 FILLER_191_1821 ();
 FILLCELL_X32 FILLER_191_1853 ();
 FILLCELL_X32 FILLER_191_1885 ();
 FILLCELL_X32 FILLER_191_1917 ();
 FILLCELL_X32 FILLER_191_1949 ();
 FILLCELL_X32 FILLER_191_1981 ();
 FILLCELL_X32 FILLER_191_2013 ();
 FILLCELL_X32 FILLER_191_2045 ();
 FILLCELL_X32 FILLER_191_2077 ();
 FILLCELL_X32 FILLER_191_2109 ();
 FILLCELL_X32 FILLER_191_2141 ();
 FILLCELL_X32 FILLER_191_2173 ();
 FILLCELL_X32 FILLER_191_2205 ();
 FILLCELL_X32 FILLER_191_2237 ();
 FILLCELL_X32 FILLER_191_2269 ();
 FILLCELL_X32 FILLER_191_2301 ();
 FILLCELL_X32 FILLER_191_2333 ();
 FILLCELL_X32 FILLER_191_2365 ();
 FILLCELL_X32 FILLER_191_2397 ();
 FILLCELL_X32 FILLER_191_2429 ();
 FILLCELL_X32 FILLER_191_2461 ();
 FILLCELL_X32 FILLER_191_2493 ();
 FILLCELL_X1 FILLER_191_2525 ();
 FILLCELL_X32 FILLER_191_2527 ();
 FILLCELL_X32 FILLER_191_2559 ();
 FILLCELL_X8 FILLER_191_2591 ();
 FILLCELL_X2 FILLER_191_2599 ();
 FILLCELL_X1 FILLER_191_2601 ();
 FILLCELL_X32 FILLER_192_1 ();
 FILLCELL_X32 FILLER_192_33 ();
 FILLCELL_X32 FILLER_192_65 ();
 FILLCELL_X32 FILLER_192_97 ();
 FILLCELL_X32 FILLER_192_129 ();
 FILLCELL_X32 FILLER_192_161 ();
 FILLCELL_X32 FILLER_192_193 ();
 FILLCELL_X32 FILLER_192_225 ();
 FILLCELL_X32 FILLER_192_257 ();
 FILLCELL_X32 FILLER_192_289 ();
 FILLCELL_X32 FILLER_192_321 ();
 FILLCELL_X32 FILLER_192_353 ();
 FILLCELL_X32 FILLER_192_385 ();
 FILLCELL_X32 FILLER_192_417 ();
 FILLCELL_X32 FILLER_192_449 ();
 FILLCELL_X32 FILLER_192_481 ();
 FILLCELL_X32 FILLER_192_513 ();
 FILLCELL_X32 FILLER_192_545 ();
 FILLCELL_X32 FILLER_192_577 ();
 FILLCELL_X16 FILLER_192_609 ();
 FILLCELL_X4 FILLER_192_625 ();
 FILLCELL_X2 FILLER_192_629 ();
 FILLCELL_X32 FILLER_192_632 ();
 FILLCELL_X32 FILLER_192_664 ();
 FILLCELL_X32 FILLER_192_696 ();
 FILLCELL_X32 FILLER_192_728 ();
 FILLCELL_X32 FILLER_192_760 ();
 FILLCELL_X32 FILLER_192_792 ();
 FILLCELL_X32 FILLER_192_824 ();
 FILLCELL_X32 FILLER_192_856 ();
 FILLCELL_X32 FILLER_192_888 ();
 FILLCELL_X32 FILLER_192_920 ();
 FILLCELL_X32 FILLER_192_952 ();
 FILLCELL_X32 FILLER_192_984 ();
 FILLCELL_X32 FILLER_192_1016 ();
 FILLCELL_X32 FILLER_192_1048 ();
 FILLCELL_X32 FILLER_192_1080 ();
 FILLCELL_X32 FILLER_192_1112 ();
 FILLCELL_X32 FILLER_192_1144 ();
 FILLCELL_X32 FILLER_192_1176 ();
 FILLCELL_X16 FILLER_192_1208 ();
 FILLCELL_X2 FILLER_192_1224 ();
 FILLCELL_X1 FILLER_192_1226 ();
 FILLCELL_X8 FILLER_192_1251 ();
 FILLCELL_X1 FILLER_192_1259 ();
 FILLCELL_X16 FILLER_192_1274 ();
 FILLCELL_X8 FILLER_192_1290 ();
 FILLCELL_X2 FILLER_192_1298 ();
 FILLCELL_X2 FILLER_192_1307 ();
 FILLCELL_X1 FILLER_192_1309 ();
 FILLCELL_X16 FILLER_192_1317 ();
 FILLCELL_X8 FILLER_192_1333 ();
 FILLCELL_X4 FILLER_192_1341 ();
 FILLCELL_X1 FILLER_192_1345 ();
 FILLCELL_X4 FILLER_192_1353 ();
 FILLCELL_X4 FILLER_192_1364 ();
 FILLCELL_X1 FILLER_192_1368 ();
 FILLCELL_X16 FILLER_192_1376 ();
 FILLCELL_X8 FILLER_192_1392 ();
 FILLCELL_X4 FILLER_192_1400 ();
 FILLCELL_X2 FILLER_192_1404 ();
 FILLCELL_X1 FILLER_192_1406 ();
 FILLCELL_X32 FILLER_192_1414 ();
 FILLCELL_X4 FILLER_192_1446 ();
 FILLCELL_X32 FILLER_192_1467 ();
 FILLCELL_X32 FILLER_192_1499 ();
 FILLCELL_X16 FILLER_192_1531 ();
 FILLCELL_X8 FILLER_192_1547 ();
 FILLCELL_X4 FILLER_192_1562 ();
 FILLCELL_X2 FILLER_192_1566 ();
 FILLCELL_X1 FILLER_192_1568 ();
 FILLCELL_X8 FILLER_192_1576 ();
 FILLCELL_X32 FILLER_192_1601 ();
 FILLCELL_X32 FILLER_192_1633 ();
 FILLCELL_X32 FILLER_192_1665 ();
 FILLCELL_X32 FILLER_192_1697 ();
 FILLCELL_X32 FILLER_192_1729 ();
 FILLCELL_X32 FILLER_192_1761 ();
 FILLCELL_X32 FILLER_192_1793 ();
 FILLCELL_X32 FILLER_192_1825 ();
 FILLCELL_X32 FILLER_192_1857 ();
 FILLCELL_X4 FILLER_192_1889 ();
 FILLCELL_X1 FILLER_192_1893 ();
 FILLCELL_X32 FILLER_192_1895 ();
 FILLCELL_X32 FILLER_192_1927 ();
 FILLCELL_X32 FILLER_192_1959 ();
 FILLCELL_X32 FILLER_192_1991 ();
 FILLCELL_X32 FILLER_192_2023 ();
 FILLCELL_X32 FILLER_192_2055 ();
 FILLCELL_X32 FILLER_192_2087 ();
 FILLCELL_X32 FILLER_192_2119 ();
 FILLCELL_X32 FILLER_192_2151 ();
 FILLCELL_X32 FILLER_192_2183 ();
 FILLCELL_X32 FILLER_192_2215 ();
 FILLCELL_X32 FILLER_192_2247 ();
 FILLCELL_X32 FILLER_192_2279 ();
 FILLCELL_X32 FILLER_192_2311 ();
 FILLCELL_X32 FILLER_192_2343 ();
 FILLCELL_X32 FILLER_192_2375 ();
 FILLCELL_X32 FILLER_192_2407 ();
 FILLCELL_X32 FILLER_192_2439 ();
 FILLCELL_X32 FILLER_192_2471 ();
 FILLCELL_X32 FILLER_192_2503 ();
 FILLCELL_X32 FILLER_192_2535 ();
 FILLCELL_X32 FILLER_192_2567 ();
 FILLCELL_X2 FILLER_192_2599 ();
 FILLCELL_X1 FILLER_192_2601 ();
 FILLCELL_X32 FILLER_193_1 ();
 FILLCELL_X32 FILLER_193_33 ();
 FILLCELL_X32 FILLER_193_65 ();
 FILLCELL_X32 FILLER_193_97 ();
 FILLCELL_X32 FILLER_193_129 ();
 FILLCELL_X32 FILLER_193_161 ();
 FILLCELL_X32 FILLER_193_193 ();
 FILLCELL_X32 FILLER_193_225 ();
 FILLCELL_X32 FILLER_193_257 ();
 FILLCELL_X32 FILLER_193_289 ();
 FILLCELL_X32 FILLER_193_321 ();
 FILLCELL_X32 FILLER_193_353 ();
 FILLCELL_X32 FILLER_193_385 ();
 FILLCELL_X32 FILLER_193_417 ();
 FILLCELL_X32 FILLER_193_449 ();
 FILLCELL_X32 FILLER_193_481 ();
 FILLCELL_X32 FILLER_193_513 ();
 FILLCELL_X32 FILLER_193_545 ();
 FILLCELL_X32 FILLER_193_577 ();
 FILLCELL_X32 FILLER_193_609 ();
 FILLCELL_X32 FILLER_193_641 ();
 FILLCELL_X32 FILLER_193_673 ();
 FILLCELL_X32 FILLER_193_705 ();
 FILLCELL_X32 FILLER_193_737 ();
 FILLCELL_X32 FILLER_193_769 ();
 FILLCELL_X32 FILLER_193_801 ();
 FILLCELL_X32 FILLER_193_833 ();
 FILLCELL_X32 FILLER_193_865 ();
 FILLCELL_X32 FILLER_193_897 ();
 FILLCELL_X32 FILLER_193_929 ();
 FILLCELL_X32 FILLER_193_961 ();
 FILLCELL_X32 FILLER_193_993 ();
 FILLCELL_X32 FILLER_193_1025 ();
 FILLCELL_X32 FILLER_193_1057 ();
 FILLCELL_X32 FILLER_193_1089 ();
 FILLCELL_X32 FILLER_193_1121 ();
 FILLCELL_X32 FILLER_193_1153 ();
 FILLCELL_X32 FILLER_193_1185 ();
 FILLCELL_X32 FILLER_193_1217 ();
 FILLCELL_X8 FILLER_193_1249 ();
 FILLCELL_X4 FILLER_193_1257 ();
 FILLCELL_X2 FILLER_193_1261 ();
 FILLCELL_X32 FILLER_193_1264 ();
 FILLCELL_X16 FILLER_193_1296 ();
 FILLCELL_X2 FILLER_193_1312 ();
 FILLCELL_X16 FILLER_193_1321 ();
 FILLCELL_X2 FILLER_193_1337 ();
 FILLCELL_X1 FILLER_193_1339 ();
 FILLCELL_X4 FILLER_193_1357 ();
 FILLCELL_X2 FILLER_193_1361 ();
 FILLCELL_X8 FILLER_193_1387 ();
 FILLCELL_X2 FILLER_193_1395 ();
 FILLCELL_X1 FILLER_193_1397 ();
 FILLCELL_X8 FILLER_193_1405 ();
 FILLCELL_X4 FILLER_193_1413 ();
 FILLCELL_X1 FILLER_193_1417 ();
 FILLCELL_X16 FILLER_193_1425 ();
 FILLCELL_X8 FILLER_193_1441 ();
 FILLCELL_X2 FILLER_193_1449 ();
 FILLCELL_X32 FILLER_193_1482 ();
 FILLCELL_X8 FILLER_193_1514 ();
 FILLCELL_X4 FILLER_193_1522 ();
 FILLCELL_X2 FILLER_193_1526 ();
 FILLCELL_X8 FILLER_193_1535 ();
 FILLCELL_X1 FILLER_193_1543 ();
 FILLCELL_X8 FILLER_193_1548 ();
 FILLCELL_X4 FILLER_193_1556 ();
 FILLCELL_X16 FILLER_193_1577 ();
 FILLCELL_X2 FILLER_193_1593 ();
 FILLCELL_X32 FILLER_193_1602 ();
 FILLCELL_X32 FILLER_193_1634 ();
 FILLCELL_X32 FILLER_193_1666 ();
 FILLCELL_X32 FILLER_193_1698 ();
 FILLCELL_X32 FILLER_193_1730 ();
 FILLCELL_X32 FILLER_193_1762 ();
 FILLCELL_X32 FILLER_193_1794 ();
 FILLCELL_X32 FILLER_193_1826 ();
 FILLCELL_X32 FILLER_193_1858 ();
 FILLCELL_X32 FILLER_193_1890 ();
 FILLCELL_X32 FILLER_193_1922 ();
 FILLCELL_X32 FILLER_193_1954 ();
 FILLCELL_X32 FILLER_193_1986 ();
 FILLCELL_X32 FILLER_193_2018 ();
 FILLCELL_X32 FILLER_193_2050 ();
 FILLCELL_X32 FILLER_193_2082 ();
 FILLCELL_X32 FILLER_193_2114 ();
 FILLCELL_X32 FILLER_193_2146 ();
 FILLCELL_X32 FILLER_193_2178 ();
 FILLCELL_X32 FILLER_193_2210 ();
 FILLCELL_X32 FILLER_193_2242 ();
 FILLCELL_X32 FILLER_193_2274 ();
 FILLCELL_X32 FILLER_193_2306 ();
 FILLCELL_X32 FILLER_193_2338 ();
 FILLCELL_X32 FILLER_193_2370 ();
 FILLCELL_X32 FILLER_193_2402 ();
 FILLCELL_X32 FILLER_193_2434 ();
 FILLCELL_X32 FILLER_193_2466 ();
 FILLCELL_X16 FILLER_193_2498 ();
 FILLCELL_X8 FILLER_193_2514 ();
 FILLCELL_X4 FILLER_193_2522 ();
 FILLCELL_X32 FILLER_193_2527 ();
 FILLCELL_X32 FILLER_193_2559 ();
 FILLCELL_X8 FILLER_193_2591 ();
 FILLCELL_X2 FILLER_193_2599 ();
 FILLCELL_X1 FILLER_193_2601 ();
 FILLCELL_X32 FILLER_194_1 ();
 FILLCELL_X32 FILLER_194_33 ();
 FILLCELL_X32 FILLER_194_65 ();
 FILLCELL_X32 FILLER_194_97 ();
 FILLCELL_X32 FILLER_194_129 ();
 FILLCELL_X32 FILLER_194_161 ();
 FILLCELL_X32 FILLER_194_193 ();
 FILLCELL_X32 FILLER_194_225 ();
 FILLCELL_X32 FILLER_194_257 ();
 FILLCELL_X32 FILLER_194_289 ();
 FILLCELL_X32 FILLER_194_321 ();
 FILLCELL_X32 FILLER_194_353 ();
 FILLCELL_X32 FILLER_194_385 ();
 FILLCELL_X32 FILLER_194_417 ();
 FILLCELL_X32 FILLER_194_449 ();
 FILLCELL_X32 FILLER_194_481 ();
 FILLCELL_X32 FILLER_194_513 ();
 FILLCELL_X32 FILLER_194_545 ();
 FILLCELL_X32 FILLER_194_577 ();
 FILLCELL_X16 FILLER_194_609 ();
 FILLCELL_X4 FILLER_194_625 ();
 FILLCELL_X2 FILLER_194_629 ();
 FILLCELL_X32 FILLER_194_632 ();
 FILLCELL_X32 FILLER_194_664 ();
 FILLCELL_X32 FILLER_194_696 ();
 FILLCELL_X32 FILLER_194_728 ();
 FILLCELL_X32 FILLER_194_760 ();
 FILLCELL_X32 FILLER_194_792 ();
 FILLCELL_X32 FILLER_194_824 ();
 FILLCELL_X32 FILLER_194_856 ();
 FILLCELL_X32 FILLER_194_888 ();
 FILLCELL_X32 FILLER_194_920 ();
 FILLCELL_X32 FILLER_194_952 ();
 FILLCELL_X32 FILLER_194_984 ();
 FILLCELL_X32 FILLER_194_1016 ();
 FILLCELL_X32 FILLER_194_1048 ();
 FILLCELL_X32 FILLER_194_1080 ();
 FILLCELL_X32 FILLER_194_1112 ();
 FILLCELL_X32 FILLER_194_1144 ();
 FILLCELL_X32 FILLER_194_1176 ();
 FILLCELL_X16 FILLER_194_1208 ();
 FILLCELL_X8 FILLER_194_1224 ();
 FILLCELL_X4 FILLER_194_1232 ();
 FILLCELL_X2 FILLER_194_1236 ();
 FILLCELL_X8 FILLER_194_1245 ();
 FILLCELL_X1 FILLER_194_1253 ();
 FILLCELL_X16 FILLER_194_1271 ();
 FILLCELL_X8 FILLER_194_1287 ();
 FILLCELL_X2 FILLER_194_1295 ();
 FILLCELL_X8 FILLER_194_1304 ();
 FILLCELL_X1 FILLER_194_1312 ();
 FILLCELL_X32 FILLER_194_1337 ();
 FILLCELL_X1 FILLER_194_1369 ();
 FILLCELL_X8 FILLER_194_1377 ();
 FILLCELL_X1 FILLER_194_1402 ();
 FILLCELL_X4 FILLER_194_1410 ();
 FILLCELL_X1 FILLER_194_1414 ();
 FILLCELL_X1 FILLER_194_1422 ();
 FILLCELL_X32 FILLER_194_1430 ();
 FILLCELL_X2 FILLER_194_1462 ();
 FILLCELL_X1 FILLER_194_1464 ();
 FILLCELL_X8 FILLER_194_1472 ();
 FILLCELL_X4 FILLER_194_1480 ();
 FILLCELL_X2 FILLER_194_1484 ();
 FILLCELL_X1 FILLER_194_1486 ();
 FILLCELL_X16 FILLER_194_1494 ();
 FILLCELL_X8 FILLER_194_1510 ();
 FILLCELL_X2 FILLER_194_1518 ();
 FILLCELL_X1 FILLER_194_1520 ();
 FILLCELL_X4 FILLER_194_1528 ();
 FILLCELL_X1 FILLER_194_1532 ();
 FILLCELL_X32 FILLER_194_1540 ();
 FILLCELL_X32 FILLER_194_1572 ();
 FILLCELL_X32 FILLER_194_1604 ();
 FILLCELL_X32 FILLER_194_1636 ();
 FILLCELL_X32 FILLER_194_1668 ();
 FILLCELL_X32 FILLER_194_1700 ();
 FILLCELL_X32 FILLER_194_1732 ();
 FILLCELL_X32 FILLER_194_1764 ();
 FILLCELL_X32 FILLER_194_1796 ();
 FILLCELL_X32 FILLER_194_1828 ();
 FILLCELL_X32 FILLER_194_1860 ();
 FILLCELL_X2 FILLER_194_1892 ();
 FILLCELL_X32 FILLER_194_1895 ();
 FILLCELL_X32 FILLER_194_1927 ();
 FILLCELL_X32 FILLER_194_1959 ();
 FILLCELL_X32 FILLER_194_1991 ();
 FILLCELL_X32 FILLER_194_2023 ();
 FILLCELL_X32 FILLER_194_2055 ();
 FILLCELL_X32 FILLER_194_2087 ();
 FILLCELL_X32 FILLER_194_2119 ();
 FILLCELL_X32 FILLER_194_2151 ();
 FILLCELL_X32 FILLER_194_2183 ();
 FILLCELL_X32 FILLER_194_2215 ();
 FILLCELL_X32 FILLER_194_2247 ();
 FILLCELL_X32 FILLER_194_2279 ();
 FILLCELL_X32 FILLER_194_2311 ();
 FILLCELL_X32 FILLER_194_2343 ();
 FILLCELL_X32 FILLER_194_2375 ();
 FILLCELL_X32 FILLER_194_2407 ();
 FILLCELL_X32 FILLER_194_2439 ();
 FILLCELL_X32 FILLER_194_2471 ();
 FILLCELL_X32 FILLER_194_2503 ();
 FILLCELL_X32 FILLER_194_2535 ();
 FILLCELL_X32 FILLER_194_2567 ();
 FILLCELL_X2 FILLER_194_2599 ();
 FILLCELL_X1 FILLER_194_2601 ();
 FILLCELL_X32 FILLER_195_1 ();
 FILLCELL_X32 FILLER_195_33 ();
 FILLCELL_X32 FILLER_195_65 ();
 FILLCELL_X32 FILLER_195_97 ();
 FILLCELL_X32 FILLER_195_129 ();
 FILLCELL_X32 FILLER_195_161 ();
 FILLCELL_X32 FILLER_195_193 ();
 FILLCELL_X32 FILLER_195_225 ();
 FILLCELL_X32 FILLER_195_257 ();
 FILLCELL_X32 FILLER_195_289 ();
 FILLCELL_X32 FILLER_195_321 ();
 FILLCELL_X32 FILLER_195_353 ();
 FILLCELL_X32 FILLER_195_385 ();
 FILLCELL_X32 FILLER_195_417 ();
 FILLCELL_X32 FILLER_195_449 ();
 FILLCELL_X32 FILLER_195_481 ();
 FILLCELL_X32 FILLER_195_513 ();
 FILLCELL_X32 FILLER_195_545 ();
 FILLCELL_X32 FILLER_195_577 ();
 FILLCELL_X32 FILLER_195_609 ();
 FILLCELL_X32 FILLER_195_641 ();
 FILLCELL_X32 FILLER_195_673 ();
 FILLCELL_X32 FILLER_195_705 ();
 FILLCELL_X32 FILLER_195_737 ();
 FILLCELL_X32 FILLER_195_769 ();
 FILLCELL_X32 FILLER_195_801 ();
 FILLCELL_X32 FILLER_195_833 ();
 FILLCELL_X32 FILLER_195_865 ();
 FILLCELL_X32 FILLER_195_897 ();
 FILLCELL_X32 FILLER_195_929 ();
 FILLCELL_X32 FILLER_195_961 ();
 FILLCELL_X32 FILLER_195_993 ();
 FILLCELL_X32 FILLER_195_1025 ();
 FILLCELL_X32 FILLER_195_1057 ();
 FILLCELL_X32 FILLER_195_1089 ();
 FILLCELL_X32 FILLER_195_1121 ();
 FILLCELL_X32 FILLER_195_1153 ();
 FILLCELL_X32 FILLER_195_1185 ();
 FILLCELL_X8 FILLER_195_1217 ();
 FILLCELL_X4 FILLER_195_1225 ();
 FILLCELL_X2 FILLER_195_1229 ();
 FILLCELL_X1 FILLER_195_1231 ();
 FILLCELL_X4 FILLER_195_1249 ();
 FILLCELL_X2 FILLER_195_1253 ();
 FILLCELL_X1 FILLER_195_1255 ();
 FILLCELL_X16 FILLER_195_1264 ();
 FILLCELL_X8 FILLER_195_1280 ();
 FILLCELL_X32 FILLER_195_1312 ();
 FILLCELL_X8 FILLER_195_1344 ();
 FILLCELL_X4 FILLER_195_1352 ();
 FILLCELL_X2 FILLER_195_1356 ();
 FILLCELL_X1 FILLER_195_1358 ();
 FILLCELL_X32 FILLER_195_1366 ();
 FILLCELL_X16 FILLER_195_1398 ();
 FILLCELL_X2 FILLER_195_1414 ();
 FILLCELL_X1 FILLER_195_1416 ();
 FILLCELL_X8 FILLER_195_1434 ();
 FILLCELL_X4 FILLER_195_1442 ();
 FILLCELL_X1 FILLER_195_1446 ();
 FILLCELL_X8 FILLER_195_1451 ();
 FILLCELL_X2 FILLER_195_1459 ();
 FILLCELL_X8 FILLER_195_1478 ();
 FILLCELL_X4 FILLER_195_1486 ();
 FILLCELL_X8 FILLER_195_1514 ();
 FILLCELL_X4 FILLER_195_1522 ();
 FILLCELL_X2 FILLER_195_1526 ();
 FILLCELL_X32 FILLER_195_1545 ();
 FILLCELL_X32 FILLER_195_1577 ();
 FILLCELL_X4 FILLER_195_1609 ();
 FILLCELL_X32 FILLER_195_1617 ();
 FILLCELL_X32 FILLER_195_1649 ();
 FILLCELL_X32 FILLER_195_1681 ();
 FILLCELL_X32 FILLER_195_1713 ();
 FILLCELL_X32 FILLER_195_1745 ();
 FILLCELL_X32 FILLER_195_1777 ();
 FILLCELL_X32 FILLER_195_1809 ();
 FILLCELL_X32 FILLER_195_1841 ();
 FILLCELL_X32 FILLER_195_1873 ();
 FILLCELL_X32 FILLER_195_1905 ();
 FILLCELL_X32 FILLER_195_1937 ();
 FILLCELL_X32 FILLER_195_1969 ();
 FILLCELL_X32 FILLER_195_2001 ();
 FILLCELL_X32 FILLER_195_2033 ();
 FILLCELL_X32 FILLER_195_2065 ();
 FILLCELL_X32 FILLER_195_2097 ();
 FILLCELL_X32 FILLER_195_2129 ();
 FILLCELL_X32 FILLER_195_2161 ();
 FILLCELL_X32 FILLER_195_2193 ();
 FILLCELL_X32 FILLER_195_2225 ();
 FILLCELL_X32 FILLER_195_2257 ();
 FILLCELL_X32 FILLER_195_2289 ();
 FILLCELL_X32 FILLER_195_2321 ();
 FILLCELL_X32 FILLER_195_2353 ();
 FILLCELL_X32 FILLER_195_2385 ();
 FILLCELL_X32 FILLER_195_2417 ();
 FILLCELL_X32 FILLER_195_2449 ();
 FILLCELL_X32 FILLER_195_2481 ();
 FILLCELL_X8 FILLER_195_2513 ();
 FILLCELL_X4 FILLER_195_2521 ();
 FILLCELL_X1 FILLER_195_2525 ();
 FILLCELL_X32 FILLER_195_2527 ();
 FILLCELL_X32 FILLER_195_2559 ();
 FILLCELL_X8 FILLER_195_2591 ();
 FILLCELL_X2 FILLER_195_2599 ();
 FILLCELL_X1 FILLER_195_2601 ();
 FILLCELL_X32 FILLER_196_1 ();
 FILLCELL_X32 FILLER_196_33 ();
 FILLCELL_X32 FILLER_196_65 ();
 FILLCELL_X32 FILLER_196_97 ();
 FILLCELL_X32 FILLER_196_129 ();
 FILLCELL_X32 FILLER_196_161 ();
 FILLCELL_X32 FILLER_196_193 ();
 FILLCELL_X32 FILLER_196_225 ();
 FILLCELL_X32 FILLER_196_257 ();
 FILLCELL_X32 FILLER_196_289 ();
 FILLCELL_X32 FILLER_196_321 ();
 FILLCELL_X32 FILLER_196_353 ();
 FILLCELL_X32 FILLER_196_385 ();
 FILLCELL_X32 FILLER_196_417 ();
 FILLCELL_X32 FILLER_196_449 ();
 FILLCELL_X32 FILLER_196_481 ();
 FILLCELL_X32 FILLER_196_513 ();
 FILLCELL_X32 FILLER_196_545 ();
 FILLCELL_X32 FILLER_196_577 ();
 FILLCELL_X16 FILLER_196_609 ();
 FILLCELL_X4 FILLER_196_625 ();
 FILLCELL_X2 FILLER_196_629 ();
 FILLCELL_X32 FILLER_196_632 ();
 FILLCELL_X32 FILLER_196_664 ();
 FILLCELL_X32 FILLER_196_696 ();
 FILLCELL_X32 FILLER_196_728 ();
 FILLCELL_X32 FILLER_196_760 ();
 FILLCELL_X32 FILLER_196_792 ();
 FILLCELL_X32 FILLER_196_824 ();
 FILLCELL_X32 FILLER_196_856 ();
 FILLCELL_X32 FILLER_196_888 ();
 FILLCELL_X32 FILLER_196_920 ();
 FILLCELL_X32 FILLER_196_952 ();
 FILLCELL_X32 FILLER_196_984 ();
 FILLCELL_X32 FILLER_196_1016 ();
 FILLCELL_X32 FILLER_196_1048 ();
 FILLCELL_X32 FILLER_196_1080 ();
 FILLCELL_X32 FILLER_196_1112 ();
 FILLCELL_X32 FILLER_196_1144 ();
 FILLCELL_X32 FILLER_196_1176 ();
 FILLCELL_X32 FILLER_196_1208 ();
 FILLCELL_X32 FILLER_196_1240 ();
 FILLCELL_X16 FILLER_196_1272 ();
 FILLCELL_X2 FILLER_196_1288 ();
 FILLCELL_X1 FILLER_196_1290 ();
 FILLCELL_X16 FILLER_196_1332 ();
 FILLCELL_X4 FILLER_196_1348 ();
 FILLCELL_X1 FILLER_196_1359 ();
 FILLCELL_X8 FILLER_196_1377 ();
 FILLCELL_X4 FILLER_196_1385 ();
 FILLCELL_X2 FILLER_196_1389 ();
 FILLCELL_X4 FILLER_196_1415 ();
 FILLCELL_X1 FILLER_196_1419 ();
 FILLCELL_X32 FILLER_196_1427 ();
 FILLCELL_X4 FILLER_196_1459 ();
 FILLCELL_X2 FILLER_196_1463 ();
 FILLCELL_X1 FILLER_196_1465 ();
 FILLCELL_X4 FILLER_196_1473 ();
 FILLCELL_X2 FILLER_196_1477 ();
 FILLCELL_X8 FILLER_196_1483 ();
 FILLCELL_X4 FILLER_196_1491 ();
 FILLCELL_X2 FILLER_196_1495 ();
 FILLCELL_X1 FILLER_196_1497 ();
 FILLCELL_X16 FILLER_196_1505 ();
 FILLCELL_X32 FILLER_196_1545 ();
 FILLCELL_X32 FILLER_196_1577 ();
 FILLCELL_X32 FILLER_196_1609 ();
 FILLCELL_X32 FILLER_196_1641 ();
 FILLCELL_X32 FILLER_196_1673 ();
 FILLCELL_X32 FILLER_196_1705 ();
 FILLCELL_X32 FILLER_196_1737 ();
 FILLCELL_X32 FILLER_196_1769 ();
 FILLCELL_X32 FILLER_196_1801 ();
 FILLCELL_X32 FILLER_196_1833 ();
 FILLCELL_X16 FILLER_196_1865 ();
 FILLCELL_X8 FILLER_196_1881 ();
 FILLCELL_X4 FILLER_196_1889 ();
 FILLCELL_X1 FILLER_196_1893 ();
 FILLCELL_X32 FILLER_196_1895 ();
 FILLCELL_X32 FILLER_196_1927 ();
 FILLCELL_X32 FILLER_196_1959 ();
 FILLCELL_X32 FILLER_196_1991 ();
 FILLCELL_X32 FILLER_196_2023 ();
 FILLCELL_X32 FILLER_196_2055 ();
 FILLCELL_X32 FILLER_196_2087 ();
 FILLCELL_X32 FILLER_196_2119 ();
 FILLCELL_X32 FILLER_196_2151 ();
 FILLCELL_X32 FILLER_196_2183 ();
 FILLCELL_X32 FILLER_196_2215 ();
 FILLCELL_X32 FILLER_196_2247 ();
 FILLCELL_X32 FILLER_196_2279 ();
 FILLCELL_X32 FILLER_196_2311 ();
 FILLCELL_X32 FILLER_196_2343 ();
 FILLCELL_X32 FILLER_196_2375 ();
 FILLCELL_X32 FILLER_196_2407 ();
 FILLCELL_X32 FILLER_196_2439 ();
 FILLCELL_X32 FILLER_196_2471 ();
 FILLCELL_X32 FILLER_196_2503 ();
 FILLCELL_X32 FILLER_196_2535 ();
 FILLCELL_X32 FILLER_196_2567 ();
 FILLCELL_X2 FILLER_196_2599 ();
 FILLCELL_X1 FILLER_196_2601 ();
 FILLCELL_X32 FILLER_197_1 ();
 FILLCELL_X32 FILLER_197_33 ();
 FILLCELL_X32 FILLER_197_65 ();
 FILLCELL_X32 FILLER_197_97 ();
 FILLCELL_X32 FILLER_197_129 ();
 FILLCELL_X32 FILLER_197_161 ();
 FILLCELL_X32 FILLER_197_193 ();
 FILLCELL_X32 FILLER_197_225 ();
 FILLCELL_X32 FILLER_197_257 ();
 FILLCELL_X32 FILLER_197_289 ();
 FILLCELL_X32 FILLER_197_321 ();
 FILLCELL_X32 FILLER_197_353 ();
 FILLCELL_X32 FILLER_197_385 ();
 FILLCELL_X32 FILLER_197_417 ();
 FILLCELL_X32 FILLER_197_449 ();
 FILLCELL_X32 FILLER_197_481 ();
 FILLCELL_X32 FILLER_197_513 ();
 FILLCELL_X32 FILLER_197_545 ();
 FILLCELL_X32 FILLER_197_577 ();
 FILLCELL_X32 FILLER_197_609 ();
 FILLCELL_X32 FILLER_197_641 ();
 FILLCELL_X32 FILLER_197_673 ();
 FILLCELL_X32 FILLER_197_705 ();
 FILLCELL_X32 FILLER_197_737 ();
 FILLCELL_X32 FILLER_197_769 ();
 FILLCELL_X32 FILLER_197_801 ();
 FILLCELL_X32 FILLER_197_833 ();
 FILLCELL_X32 FILLER_197_865 ();
 FILLCELL_X32 FILLER_197_897 ();
 FILLCELL_X32 FILLER_197_929 ();
 FILLCELL_X32 FILLER_197_961 ();
 FILLCELL_X32 FILLER_197_993 ();
 FILLCELL_X32 FILLER_197_1025 ();
 FILLCELL_X32 FILLER_197_1057 ();
 FILLCELL_X32 FILLER_197_1089 ();
 FILLCELL_X32 FILLER_197_1121 ();
 FILLCELL_X32 FILLER_197_1153 ();
 FILLCELL_X32 FILLER_197_1185 ();
 FILLCELL_X32 FILLER_197_1217 ();
 FILLCELL_X8 FILLER_197_1249 ();
 FILLCELL_X4 FILLER_197_1257 ();
 FILLCELL_X2 FILLER_197_1261 ();
 FILLCELL_X16 FILLER_197_1264 ();
 FILLCELL_X8 FILLER_197_1280 ();
 FILLCELL_X2 FILLER_197_1288 ();
 FILLCELL_X32 FILLER_197_1297 ();
 FILLCELL_X16 FILLER_197_1329 ();
 FILLCELL_X2 FILLER_197_1345 ();
 FILLCELL_X32 FILLER_197_1364 ();
 FILLCELL_X16 FILLER_197_1396 ();
 FILLCELL_X2 FILLER_197_1412 ();
 FILLCELL_X1 FILLER_197_1414 ();
 FILLCELL_X16 FILLER_197_1432 ();
 FILLCELL_X4 FILLER_197_1448 ();
 FILLCELL_X16 FILLER_197_1476 ();
 FILLCELL_X1 FILLER_197_1492 ();
 FILLCELL_X32 FILLER_197_1510 ();
 FILLCELL_X32 FILLER_197_1542 ();
 FILLCELL_X32 FILLER_197_1574 ();
 FILLCELL_X32 FILLER_197_1606 ();
 FILLCELL_X32 FILLER_197_1638 ();
 FILLCELL_X32 FILLER_197_1670 ();
 FILLCELL_X32 FILLER_197_1702 ();
 FILLCELL_X32 FILLER_197_1734 ();
 FILLCELL_X32 FILLER_197_1766 ();
 FILLCELL_X32 FILLER_197_1798 ();
 FILLCELL_X32 FILLER_197_1830 ();
 FILLCELL_X32 FILLER_197_1862 ();
 FILLCELL_X32 FILLER_197_1894 ();
 FILLCELL_X32 FILLER_197_1926 ();
 FILLCELL_X32 FILLER_197_1958 ();
 FILLCELL_X32 FILLER_197_1990 ();
 FILLCELL_X32 FILLER_197_2022 ();
 FILLCELL_X32 FILLER_197_2054 ();
 FILLCELL_X32 FILLER_197_2086 ();
 FILLCELL_X32 FILLER_197_2118 ();
 FILLCELL_X32 FILLER_197_2150 ();
 FILLCELL_X32 FILLER_197_2182 ();
 FILLCELL_X32 FILLER_197_2214 ();
 FILLCELL_X32 FILLER_197_2246 ();
 FILLCELL_X32 FILLER_197_2278 ();
 FILLCELL_X32 FILLER_197_2310 ();
 FILLCELL_X32 FILLER_197_2342 ();
 FILLCELL_X32 FILLER_197_2374 ();
 FILLCELL_X32 FILLER_197_2406 ();
 FILLCELL_X32 FILLER_197_2438 ();
 FILLCELL_X32 FILLER_197_2470 ();
 FILLCELL_X16 FILLER_197_2502 ();
 FILLCELL_X8 FILLER_197_2518 ();
 FILLCELL_X32 FILLER_197_2527 ();
 FILLCELL_X32 FILLER_197_2559 ();
 FILLCELL_X8 FILLER_197_2591 ();
 FILLCELL_X2 FILLER_197_2599 ();
 FILLCELL_X1 FILLER_197_2601 ();
 FILLCELL_X32 FILLER_198_1 ();
 FILLCELL_X32 FILLER_198_33 ();
 FILLCELL_X32 FILLER_198_65 ();
 FILLCELL_X32 FILLER_198_97 ();
 FILLCELL_X32 FILLER_198_129 ();
 FILLCELL_X32 FILLER_198_161 ();
 FILLCELL_X32 FILLER_198_193 ();
 FILLCELL_X32 FILLER_198_225 ();
 FILLCELL_X32 FILLER_198_257 ();
 FILLCELL_X32 FILLER_198_289 ();
 FILLCELL_X32 FILLER_198_321 ();
 FILLCELL_X32 FILLER_198_353 ();
 FILLCELL_X32 FILLER_198_385 ();
 FILLCELL_X32 FILLER_198_417 ();
 FILLCELL_X32 FILLER_198_449 ();
 FILLCELL_X32 FILLER_198_481 ();
 FILLCELL_X32 FILLER_198_513 ();
 FILLCELL_X32 FILLER_198_545 ();
 FILLCELL_X32 FILLER_198_577 ();
 FILLCELL_X16 FILLER_198_609 ();
 FILLCELL_X4 FILLER_198_625 ();
 FILLCELL_X2 FILLER_198_629 ();
 FILLCELL_X32 FILLER_198_632 ();
 FILLCELL_X32 FILLER_198_664 ();
 FILLCELL_X32 FILLER_198_696 ();
 FILLCELL_X32 FILLER_198_728 ();
 FILLCELL_X32 FILLER_198_760 ();
 FILLCELL_X32 FILLER_198_792 ();
 FILLCELL_X32 FILLER_198_824 ();
 FILLCELL_X32 FILLER_198_856 ();
 FILLCELL_X32 FILLER_198_888 ();
 FILLCELL_X32 FILLER_198_920 ();
 FILLCELL_X32 FILLER_198_952 ();
 FILLCELL_X32 FILLER_198_984 ();
 FILLCELL_X32 FILLER_198_1016 ();
 FILLCELL_X32 FILLER_198_1048 ();
 FILLCELL_X32 FILLER_198_1080 ();
 FILLCELL_X32 FILLER_198_1112 ();
 FILLCELL_X32 FILLER_198_1144 ();
 FILLCELL_X32 FILLER_198_1176 ();
 FILLCELL_X8 FILLER_198_1208 ();
 FILLCELL_X4 FILLER_198_1216 ();
 FILLCELL_X32 FILLER_198_1224 ();
 FILLCELL_X32 FILLER_198_1256 ();
 FILLCELL_X32 FILLER_198_1288 ();
 FILLCELL_X32 FILLER_198_1320 ();
 FILLCELL_X32 FILLER_198_1352 ();
 FILLCELL_X32 FILLER_198_1384 ();
 FILLCELL_X32 FILLER_198_1416 ();
 FILLCELL_X32 FILLER_198_1448 ();
 FILLCELL_X32 FILLER_198_1480 ();
 FILLCELL_X32 FILLER_198_1512 ();
 FILLCELL_X32 FILLER_198_1544 ();
 FILLCELL_X32 FILLER_198_1576 ();
 FILLCELL_X32 FILLER_198_1608 ();
 FILLCELL_X32 FILLER_198_1640 ();
 FILLCELL_X32 FILLER_198_1672 ();
 FILLCELL_X32 FILLER_198_1704 ();
 FILLCELL_X32 FILLER_198_1736 ();
 FILLCELL_X32 FILLER_198_1768 ();
 FILLCELL_X32 FILLER_198_1800 ();
 FILLCELL_X32 FILLER_198_1832 ();
 FILLCELL_X16 FILLER_198_1864 ();
 FILLCELL_X8 FILLER_198_1880 ();
 FILLCELL_X4 FILLER_198_1888 ();
 FILLCELL_X2 FILLER_198_1892 ();
 FILLCELL_X32 FILLER_198_1895 ();
 FILLCELL_X32 FILLER_198_1927 ();
 FILLCELL_X32 FILLER_198_1959 ();
 FILLCELL_X32 FILLER_198_1991 ();
 FILLCELL_X32 FILLER_198_2023 ();
 FILLCELL_X32 FILLER_198_2055 ();
 FILLCELL_X32 FILLER_198_2087 ();
 FILLCELL_X32 FILLER_198_2119 ();
 FILLCELL_X32 FILLER_198_2151 ();
 FILLCELL_X32 FILLER_198_2183 ();
 FILLCELL_X32 FILLER_198_2215 ();
 FILLCELL_X32 FILLER_198_2247 ();
 FILLCELL_X32 FILLER_198_2279 ();
 FILLCELL_X32 FILLER_198_2311 ();
 FILLCELL_X32 FILLER_198_2343 ();
 FILLCELL_X32 FILLER_198_2375 ();
 FILLCELL_X32 FILLER_198_2407 ();
 FILLCELL_X32 FILLER_198_2439 ();
 FILLCELL_X32 FILLER_198_2471 ();
 FILLCELL_X32 FILLER_198_2503 ();
 FILLCELL_X32 FILLER_198_2535 ();
 FILLCELL_X32 FILLER_198_2567 ();
 FILLCELL_X2 FILLER_198_2599 ();
 FILLCELL_X1 FILLER_198_2601 ();
 FILLCELL_X32 FILLER_199_1 ();
 FILLCELL_X32 FILLER_199_33 ();
 FILLCELL_X32 FILLER_199_65 ();
 FILLCELL_X32 FILLER_199_97 ();
 FILLCELL_X32 FILLER_199_129 ();
 FILLCELL_X32 FILLER_199_161 ();
 FILLCELL_X32 FILLER_199_193 ();
 FILLCELL_X32 FILLER_199_225 ();
 FILLCELL_X32 FILLER_199_257 ();
 FILLCELL_X32 FILLER_199_289 ();
 FILLCELL_X32 FILLER_199_321 ();
 FILLCELL_X32 FILLER_199_353 ();
 FILLCELL_X32 FILLER_199_385 ();
 FILLCELL_X32 FILLER_199_417 ();
 FILLCELL_X32 FILLER_199_449 ();
 FILLCELL_X32 FILLER_199_481 ();
 FILLCELL_X32 FILLER_199_513 ();
 FILLCELL_X32 FILLER_199_545 ();
 FILLCELL_X32 FILLER_199_577 ();
 FILLCELL_X32 FILLER_199_609 ();
 FILLCELL_X32 FILLER_199_641 ();
 FILLCELL_X32 FILLER_199_673 ();
 FILLCELL_X32 FILLER_199_705 ();
 FILLCELL_X32 FILLER_199_737 ();
 FILLCELL_X32 FILLER_199_769 ();
 FILLCELL_X32 FILLER_199_801 ();
 FILLCELL_X32 FILLER_199_833 ();
 FILLCELL_X32 FILLER_199_865 ();
 FILLCELL_X32 FILLER_199_897 ();
 FILLCELL_X32 FILLER_199_929 ();
 FILLCELL_X32 FILLER_199_961 ();
 FILLCELL_X32 FILLER_199_993 ();
 FILLCELL_X32 FILLER_199_1025 ();
 FILLCELL_X32 FILLER_199_1057 ();
 FILLCELL_X32 FILLER_199_1089 ();
 FILLCELL_X32 FILLER_199_1121 ();
 FILLCELL_X32 FILLER_199_1153 ();
 FILLCELL_X32 FILLER_199_1185 ();
 FILLCELL_X32 FILLER_199_1217 ();
 FILLCELL_X8 FILLER_199_1249 ();
 FILLCELL_X4 FILLER_199_1257 ();
 FILLCELL_X2 FILLER_199_1261 ();
 FILLCELL_X8 FILLER_199_1264 ();
 FILLCELL_X4 FILLER_199_1272 ();
 FILLCELL_X1 FILLER_199_1276 ();
 FILLCELL_X32 FILLER_199_1281 ();
 FILLCELL_X32 FILLER_199_1313 ();
 FILLCELL_X32 FILLER_199_1345 ();
 FILLCELL_X32 FILLER_199_1377 ();
 FILLCELL_X32 FILLER_199_1409 ();
 FILLCELL_X32 FILLER_199_1441 ();
 FILLCELL_X32 FILLER_199_1473 ();
 FILLCELL_X32 FILLER_199_1505 ();
 FILLCELL_X32 FILLER_199_1537 ();
 FILLCELL_X32 FILLER_199_1569 ();
 FILLCELL_X32 FILLER_199_1601 ();
 FILLCELL_X32 FILLER_199_1633 ();
 FILLCELL_X32 FILLER_199_1665 ();
 FILLCELL_X32 FILLER_199_1697 ();
 FILLCELL_X32 FILLER_199_1729 ();
 FILLCELL_X32 FILLER_199_1761 ();
 FILLCELL_X32 FILLER_199_1793 ();
 FILLCELL_X32 FILLER_199_1825 ();
 FILLCELL_X32 FILLER_199_1857 ();
 FILLCELL_X32 FILLER_199_1889 ();
 FILLCELL_X32 FILLER_199_1921 ();
 FILLCELL_X32 FILLER_199_1953 ();
 FILLCELL_X32 FILLER_199_1985 ();
 FILLCELL_X32 FILLER_199_2017 ();
 FILLCELL_X32 FILLER_199_2049 ();
 FILLCELL_X32 FILLER_199_2081 ();
 FILLCELL_X32 FILLER_199_2113 ();
 FILLCELL_X32 FILLER_199_2145 ();
 FILLCELL_X32 FILLER_199_2177 ();
 FILLCELL_X32 FILLER_199_2209 ();
 FILLCELL_X32 FILLER_199_2241 ();
 FILLCELL_X32 FILLER_199_2273 ();
 FILLCELL_X32 FILLER_199_2305 ();
 FILLCELL_X32 FILLER_199_2337 ();
 FILLCELL_X32 FILLER_199_2369 ();
 FILLCELL_X32 FILLER_199_2401 ();
 FILLCELL_X32 FILLER_199_2433 ();
 FILLCELL_X32 FILLER_199_2465 ();
 FILLCELL_X16 FILLER_199_2497 ();
 FILLCELL_X8 FILLER_199_2513 ();
 FILLCELL_X4 FILLER_199_2521 ();
 FILLCELL_X1 FILLER_199_2525 ();
 FILLCELL_X32 FILLER_199_2527 ();
 FILLCELL_X32 FILLER_199_2559 ();
 FILLCELL_X8 FILLER_199_2591 ();
 FILLCELL_X2 FILLER_199_2599 ();
 FILLCELL_X1 FILLER_199_2601 ();
 FILLCELL_X32 FILLER_200_1 ();
 FILLCELL_X32 FILLER_200_33 ();
 FILLCELL_X32 FILLER_200_65 ();
 FILLCELL_X32 FILLER_200_97 ();
 FILLCELL_X32 FILLER_200_129 ();
 FILLCELL_X32 FILLER_200_161 ();
 FILLCELL_X32 FILLER_200_193 ();
 FILLCELL_X32 FILLER_200_225 ();
 FILLCELL_X32 FILLER_200_257 ();
 FILLCELL_X32 FILLER_200_289 ();
 FILLCELL_X32 FILLER_200_321 ();
 FILLCELL_X32 FILLER_200_353 ();
 FILLCELL_X32 FILLER_200_385 ();
 FILLCELL_X32 FILLER_200_417 ();
 FILLCELL_X32 FILLER_200_449 ();
 FILLCELL_X32 FILLER_200_481 ();
 FILLCELL_X32 FILLER_200_513 ();
 FILLCELL_X32 FILLER_200_545 ();
 FILLCELL_X32 FILLER_200_577 ();
 FILLCELL_X16 FILLER_200_609 ();
 FILLCELL_X4 FILLER_200_625 ();
 FILLCELL_X2 FILLER_200_629 ();
 FILLCELL_X32 FILLER_200_632 ();
 FILLCELL_X32 FILLER_200_664 ();
 FILLCELL_X32 FILLER_200_696 ();
 FILLCELL_X32 FILLER_200_728 ();
 FILLCELL_X32 FILLER_200_760 ();
 FILLCELL_X32 FILLER_200_792 ();
 FILLCELL_X32 FILLER_200_824 ();
 FILLCELL_X32 FILLER_200_856 ();
 FILLCELL_X32 FILLER_200_888 ();
 FILLCELL_X32 FILLER_200_920 ();
 FILLCELL_X32 FILLER_200_952 ();
 FILLCELL_X32 FILLER_200_984 ();
 FILLCELL_X32 FILLER_200_1016 ();
 FILLCELL_X32 FILLER_200_1048 ();
 FILLCELL_X32 FILLER_200_1080 ();
 FILLCELL_X32 FILLER_200_1112 ();
 FILLCELL_X32 FILLER_200_1144 ();
 FILLCELL_X32 FILLER_200_1176 ();
 FILLCELL_X32 FILLER_200_1208 ();
 FILLCELL_X32 FILLER_200_1240 ();
 FILLCELL_X32 FILLER_200_1272 ();
 FILLCELL_X16 FILLER_200_1304 ();
 FILLCELL_X8 FILLER_200_1320 ();
 FILLCELL_X2 FILLER_200_1328 ();
 FILLCELL_X1 FILLER_200_1330 ();
 FILLCELL_X32 FILLER_200_1335 ();
 FILLCELL_X32 FILLER_200_1367 ();
 FILLCELL_X32 FILLER_200_1399 ();
 FILLCELL_X32 FILLER_200_1431 ();
 FILLCELL_X32 FILLER_200_1463 ();
 FILLCELL_X32 FILLER_200_1495 ();
 FILLCELL_X32 FILLER_200_1527 ();
 FILLCELL_X32 FILLER_200_1559 ();
 FILLCELL_X32 FILLER_200_1591 ();
 FILLCELL_X32 FILLER_200_1623 ();
 FILLCELL_X32 FILLER_200_1655 ();
 FILLCELL_X32 FILLER_200_1687 ();
 FILLCELL_X32 FILLER_200_1719 ();
 FILLCELL_X32 FILLER_200_1751 ();
 FILLCELL_X32 FILLER_200_1783 ();
 FILLCELL_X32 FILLER_200_1815 ();
 FILLCELL_X32 FILLER_200_1847 ();
 FILLCELL_X8 FILLER_200_1879 ();
 FILLCELL_X4 FILLER_200_1887 ();
 FILLCELL_X2 FILLER_200_1891 ();
 FILLCELL_X1 FILLER_200_1893 ();
 FILLCELL_X32 FILLER_200_1895 ();
 FILLCELL_X32 FILLER_200_1927 ();
 FILLCELL_X32 FILLER_200_1959 ();
 FILLCELL_X32 FILLER_200_1991 ();
 FILLCELL_X32 FILLER_200_2023 ();
 FILLCELL_X32 FILLER_200_2055 ();
 FILLCELL_X32 FILLER_200_2087 ();
 FILLCELL_X32 FILLER_200_2119 ();
 FILLCELL_X32 FILLER_200_2151 ();
 FILLCELL_X32 FILLER_200_2183 ();
 FILLCELL_X32 FILLER_200_2215 ();
 FILLCELL_X32 FILLER_200_2247 ();
 FILLCELL_X32 FILLER_200_2279 ();
 FILLCELL_X32 FILLER_200_2311 ();
 FILLCELL_X32 FILLER_200_2343 ();
 FILLCELL_X32 FILLER_200_2375 ();
 FILLCELL_X32 FILLER_200_2407 ();
 FILLCELL_X32 FILLER_200_2439 ();
 FILLCELL_X32 FILLER_200_2471 ();
 FILLCELL_X32 FILLER_200_2503 ();
 FILLCELL_X32 FILLER_200_2535 ();
 FILLCELL_X32 FILLER_200_2567 ();
 FILLCELL_X2 FILLER_200_2599 ();
 FILLCELL_X1 FILLER_200_2601 ();
 FILLCELL_X32 FILLER_201_1 ();
 FILLCELL_X32 FILLER_201_33 ();
 FILLCELL_X32 FILLER_201_65 ();
 FILLCELL_X32 FILLER_201_97 ();
 FILLCELL_X32 FILLER_201_129 ();
 FILLCELL_X32 FILLER_201_161 ();
 FILLCELL_X32 FILLER_201_193 ();
 FILLCELL_X32 FILLER_201_225 ();
 FILLCELL_X32 FILLER_201_257 ();
 FILLCELL_X32 FILLER_201_289 ();
 FILLCELL_X32 FILLER_201_321 ();
 FILLCELL_X32 FILLER_201_353 ();
 FILLCELL_X32 FILLER_201_385 ();
 FILLCELL_X32 FILLER_201_417 ();
 FILLCELL_X32 FILLER_201_449 ();
 FILLCELL_X32 FILLER_201_481 ();
 FILLCELL_X32 FILLER_201_513 ();
 FILLCELL_X32 FILLER_201_545 ();
 FILLCELL_X32 FILLER_201_577 ();
 FILLCELL_X32 FILLER_201_609 ();
 FILLCELL_X32 FILLER_201_641 ();
 FILLCELL_X32 FILLER_201_673 ();
 FILLCELL_X32 FILLER_201_705 ();
 FILLCELL_X32 FILLER_201_737 ();
 FILLCELL_X32 FILLER_201_769 ();
 FILLCELL_X32 FILLER_201_801 ();
 FILLCELL_X32 FILLER_201_833 ();
 FILLCELL_X32 FILLER_201_865 ();
 FILLCELL_X32 FILLER_201_897 ();
 FILLCELL_X32 FILLER_201_929 ();
 FILLCELL_X32 FILLER_201_961 ();
 FILLCELL_X32 FILLER_201_993 ();
 FILLCELL_X32 FILLER_201_1025 ();
 FILLCELL_X32 FILLER_201_1057 ();
 FILLCELL_X32 FILLER_201_1089 ();
 FILLCELL_X32 FILLER_201_1121 ();
 FILLCELL_X32 FILLER_201_1153 ();
 FILLCELL_X32 FILLER_201_1185 ();
 FILLCELL_X32 FILLER_201_1217 ();
 FILLCELL_X8 FILLER_201_1249 ();
 FILLCELL_X4 FILLER_201_1257 ();
 FILLCELL_X2 FILLER_201_1261 ();
 FILLCELL_X32 FILLER_201_1264 ();
 FILLCELL_X32 FILLER_201_1296 ();
 FILLCELL_X32 FILLER_201_1328 ();
 FILLCELL_X32 FILLER_201_1360 ();
 FILLCELL_X32 FILLER_201_1392 ();
 FILLCELL_X32 FILLER_201_1424 ();
 FILLCELL_X32 FILLER_201_1456 ();
 FILLCELL_X32 FILLER_201_1488 ();
 FILLCELL_X32 FILLER_201_1520 ();
 FILLCELL_X32 FILLER_201_1552 ();
 FILLCELL_X32 FILLER_201_1584 ();
 FILLCELL_X32 FILLER_201_1616 ();
 FILLCELL_X32 FILLER_201_1648 ();
 FILLCELL_X32 FILLER_201_1680 ();
 FILLCELL_X32 FILLER_201_1712 ();
 FILLCELL_X32 FILLER_201_1744 ();
 FILLCELL_X32 FILLER_201_1776 ();
 FILLCELL_X32 FILLER_201_1808 ();
 FILLCELL_X32 FILLER_201_1840 ();
 FILLCELL_X32 FILLER_201_1872 ();
 FILLCELL_X32 FILLER_201_1904 ();
 FILLCELL_X32 FILLER_201_1936 ();
 FILLCELL_X32 FILLER_201_1968 ();
 FILLCELL_X32 FILLER_201_2000 ();
 FILLCELL_X32 FILLER_201_2032 ();
 FILLCELL_X32 FILLER_201_2064 ();
 FILLCELL_X32 FILLER_201_2096 ();
 FILLCELL_X32 FILLER_201_2128 ();
 FILLCELL_X32 FILLER_201_2160 ();
 FILLCELL_X32 FILLER_201_2192 ();
 FILLCELL_X32 FILLER_201_2224 ();
 FILLCELL_X32 FILLER_201_2256 ();
 FILLCELL_X32 FILLER_201_2288 ();
 FILLCELL_X32 FILLER_201_2320 ();
 FILLCELL_X32 FILLER_201_2352 ();
 FILLCELL_X32 FILLER_201_2384 ();
 FILLCELL_X32 FILLER_201_2416 ();
 FILLCELL_X32 FILLER_201_2448 ();
 FILLCELL_X32 FILLER_201_2480 ();
 FILLCELL_X8 FILLER_201_2512 ();
 FILLCELL_X4 FILLER_201_2520 ();
 FILLCELL_X2 FILLER_201_2524 ();
 FILLCELL_X32 FILLER_201_2527 ();
 FILLCELL_X32 FILLER_201_2559 ();
 FILLCELL_X8 FILLER_201_2591 ();
 FILLCELL_X2 FILLER_201_2599 ();
 FILLCELL_X1 FILLER_201_2601 ();
 FILLCELL_X32 FILLER_202_1 ();
 FILLCELL_X32 FILLER_202_33 ();
 FILLCELL_X32 FILLER_202_65 ();
 FILLCELL_X32 FILLER_202_97 ();
 FILLCELL_X32 FILLER_202_129 ();
 FILLCELL_X32 FILLER_202_161 ();
 FILLCELL_X32 FILLER_202_193 ();
 FILLCELL_X32 FILLER_202_225 ();
 FILLCELL_X32 FILLER_202_257 ();
 FILLCELL_X32 FILLER_202_289 ();
 FILLCELL_X32 FILLER_202_321 ();
 FILLCELL_X32 FILLER_202_353 ();
 FILLCELL_X32 FILLER_202_385 ();
 FILLCELL_X32 FILLER_202_417 ();
 FILLCELL_X32 FILLER_202_449 ();
 FILLCELL_X32 FILLER_202_481 ();
 FILLCELL_X32 FILLER_202_513 ();
 FILLCELL_X32 FILLER_202_545 ();
 FILLCELL_X32 FILLER_202_577 ();
 FILLCELL_X16 FILLER_202_609 ();
 FILLCELL_X4 FILLER_202_625 ();
 FILLCELL_X2 FILLER_202_629 ();
 FILLCELL_X32 FILLER_202_632 ();
 FILLCELL_X32 FILLER_202_664 ();
 FILLCELL_X32 FILLER_202_696 ();
 FILLCELL_X32 FILLER_202_728 ();
 FILLCELL_X32 FILLER_202_760 ();
 FILLCELL_X32 FILLER_202_792 ();
 FILLCELL_X32 FILLER_202_824 ();
 FILLCELL_X32 FILLER_202_856 ();
 FILLCELL_X32 FILLER_202_888 ();
 FILLCELL_X32 FILLER_202_920 ();
 FILLCELL_X32 FILLER_202_952 ();
 FILLCELL_X32 FILLER_202_984 ();
 FILLCELL_X32 FILLER_202_1016 ();
 FILLCELL_X32 FILLER_202_1048 ();
 FILLCELL_X32 FILLER_202_1080 ();
 FILLCELL_X32 FILLER_202_1112 ();
 FILLCELL_X32 FILLER_202_1144 ();
 FILLCELL_X32 FILLER_202_1176 ();
 FILLCELL_X32 FILLER_202_1208 ();
 FILLCELL_X32 FILLER_202_1240 ();
 FILLCELL_X32 FILLER_202_1272 ();
 FILLCELL_X32 FILLER_202_1304 ();
 FILLCELL_X32 FILLER_202_1336 ();
 FILLCELL_X32 FILLER_202_1368 ();
 FILLCELL_X32 FILLER_202_1400 ();
 FILLCELL_X32 FILLER_202_1432 ();
 FILLCELL_X32 FILLER_202_1464 ();
 FILLCELL_X32 FILLER_202_1496 ();
 FILLCELL_X32 FILLER_202_1528 ();
 FILLCELL_X32 FILLER_202_1560 ();
 FILLCELL_X32 FILLER_202_1592 ();
 FILLCELL_X32 FILLER_202_1624 ();
 FILLCELL_X32 FILLER_202_1656 ();
 FILLCELL_X32 FILLER_202_1688 ();
 FILLCELL_X32 FILLER_202_1720 ();
 FILLCELL_X32 FILLER_202_1752 ();
 FILLCELL_X32 FILLER_202_1784 ();
 FILLCELL_X32 FILLER_202_1816 ();
 FILLCELL_X32 FILLER_202_1848 ();
 FILLCELL_X8 FILLER_202_1880 ();
 FILLCELL_X4 FILLER_202_1888 ();
 FILLCELL_X2 FILLER_202_1892 ();
 FILLCELL_X32 FILLER_202_1895 ();
 FILLCELL_X32 FILLER_202_1927 ();
 FILLCELL_X32 FILLER_202_1959 ();
 FILLCELL_X32 FILLER_202_1991 ();
 FILLCELL_X32 FILLER_202_2023 ();
 FILLCELL_X32 FILLER_202_2055 ();
 FILLCELL_X32 FILLER_202_2087 ();
 FILLCELL_X32 FILLER_202_2119 ();
 FILLCELL_X32 FILLER_202_2151 ();
 FILLCELL_X32 FILLER_202_2183 ();
 FILLCELL_X32 FILLER_202_2215 ();
 FILLCELL_X32 FILLER_202_2247 ();
 FILLCELL_X32 FILLER_202_2279 ();
 FILLCELL_X32 FILLER_202_2311 ();
 FILLCELL_X32 FILLER_202_2343 ();
 FILLCELL_X32 FILLER_202_2375 ();
 FILLCELL_X32 FILLER_202_2407 ();
 FILLCELL_X32 FILLER_202_2439 ();
 FILLCELL_X32 FILLER_202_2471 ();
 FILLCELL_X32 FILLER_202_2503 ();
 FILLCELL_X32 FILLER_202_2535 ();
 FILLCELL_X32 FILLER_202_2567 ();
 FILLCELL_X2 FILLER_202_2599 ();
 FILLCELL_X1 FILLER_202_2601 ();
 FILLCELL_X32 FILLER_203_1 ();
 FILLCELL_X32 FILLER_203_33 ();
 FILLCELL_X32 FILLER_203_65 ();
 FILLCELL_X32 FILLER_203_97 ();
 FILLCELL_X32 FILLER_203_129 ();
 FILLCELL_X32 FILLER_203_161 ();
 FILLCELL_X32 FILLER_203_193 ();
 FILLCELL_X32 FILLER_203_225 ();
 FILLCELL_X32 FILLER_203_257 ();
 FILLCELL_X32 FILLER_203_289 ();
 FILLCELL_X32 FILLER_203_321 ();
 FILLCELL_X32 FILLER_203_353 ();
 FILLCELL_X32 FILLER_203_385 ();
 FILLCELL_X32 FILLER_203_417 ();
 FILLCELL_X32 FILLER_203_449 ();
 FILLCELL_X32 FILLER_203_481 ();
 FILLCELL_X32 FILLER_203_513 ();
 FILLCELL_X32 FILLER_203_545 ();
 FILLCELL_X32 FILLER_203_577 ();
 FILLCELL_X32 FILLER_203_609 ();
 FILLCELL_X32 FILLER_203_641 ();
 FILLCELL_X32 FILLER_203_673 ();
 FILLCELL_X32 FILLER_203_705 ();
 FILLCELL_X32 FILLER_203_737 ();
 FILLCELL_X32 FILLER_203_769 ();
 FILLCELL_X32 FILLER_203_801 ();
 FILLCELL_X32 FILLER_203_833 ();
 FILLCELL_X32 FILLER_203_865 ();
 FILLCELL_X32 FILLER_203_897 ();
 FILLCELL_X32 FILLER_203_929 ();
 FILLCELL_X32 FILLER_203_961 ();
 FILLCELL_X32 FILLER_203_993 ();
 FILLCELL_X32 FILLER_203_1025 ();
 FILLCELL_X32 FILLER_203_1057 ();
 FILLCELL_X32 FILLER_203_1089 ();
 FILLCELL_X32 FILLER_203_1121 ();
 FILLCELL_X32 FILLER_203_1153 ();
 FILLCELL_X32 FILLER_203_1185 ();
 FILLCELL_X32 FILLER_203_1217 ();
 FILLCELL_X8 FILLER_203_1249 ();
 FILLCELL_X4 FILLER_203_1257 ();
 FILLCELL_X2 FILLER_203_1261 ();
 FILLCELL_X32 FILLER_203_1264 ();
 FILLCELL_X32 FILLER_203_1296 ();
 FILLCELL_X32 FILLER_203_1328 ();
 FILLCELL_X32 FILLER_203_1360 ();
 FILLCELL_X32 FILLER_203_1392 ();
 FILLCELL_X32 FILLER_203_1424 ();
 FILLCELL_X32 FILLER_203_1456 ();
 FILLCELL_X32 FILLER_203_1488 ();
 FILLCELL_X32 FILLER_203_1520 ();
 FILLCELL_X32 FILLER_203_1552 ();
 FILLCELL_X32 FILLER_203_1584 ();
 FILLCELL_X32 FILLER_203_1616 ();
 FILLCELL_X32 FILLER_203_1648 ();
 FILLCELL_X32 FILLER_203_1680 ();
 FILLCELL_X32 FILLER_203_1712 ();
 FILLCELL_X32 FILLER_203_1744 ();
 FILLCELL_X32 FILLER_203_1776 ();
 FILLCELL_X32 FILLER_203_1808 ();
 FILLCELL_X32 FILLER_203_1840 ();
 FILLCELL_X32 FILLER_203_1872 ();
 FILLCELL_X32 FILLER_203_1904 ();
 FILLCELL_X32 FILLER_203_1936 ();
 FILLCELL_X32 FILLER_203_1968 ();
 FILLCELL_X32 FILLER_203_2000 ();
 FILLCELL_X32 FILLER_203_2032 ();
 FILLCELL_X32 FILLER_203_2064 ();
 FILLCELL_X32 FILLER_203_2096 ();
 FILLCELL_X32 FILLER_203_2128 ();
 FILLCELL_X32 FILLER_203_2160 ();
 FILLCELL_X32 FILLER_203_2192 ();
 FILLCELL_X32 FILLER_203_2224 ();
 FILLCELL_X32 FILLER_203_2256 ();
 FILLCELL_X32 FILLER_203_2288 ();
 FILLCELL_X32 FILLER_203_2320 ();
 FILLCELL_X32 FILLER_203_2352 ();
 FILLCELL_X32 FILLER_203_2384 ();
 FILLCELL_X32 FILLER_203_2416 ();
 FILLCELL_X32 FILLER_203_2448 ();
 FILLCELL_X32 FILLER_203_2480 ();
 FILLCELL_X8 FILLER_203_2512 ();
 FILLCELL_X4 FILLER_203_2520 ();
 FILLCELL_X2 FILLER_203_2524 ();
 FILLCELL_X32 FILLER_203_2527 ();
 FILLCELL_X32 FILLER_203_2559 ();
 FILLCELL_X8 FILLER_203_2591 ();
 FILLCELL_X2 FILLER_203_2599 ();
 FILLCELL_X1 FILLER_203_2601 ();
 FILLCELL_X32 FILLER_204_1 ();
 FILLCELL_X32 FILLER_204_33 ();
 FILLCELL_X32 FILLER_204_65 ();
 FILLCELL_X32 FILLER_204_97 ();
 FILLCELL_X32 FILLER_204_129 ();
 FILLCELL_X32 FILLER_204_161 ();
 FILLCELL_X32 FILLER_204_193 ();
 FILLCELL_X32 FILLER_204_225 ();
 FILLCELL_X32 FILLER_204_257 ();
 FILLCELL_X32 FILLER_204_289 ();
 FILLCELL_X32 FILLER_204_321 ();
 FILLCELL_X32 FILLER_204_353 ();
 FILLCELL_X32 FILLER_204_385 ();
 FILLCELL_X32 FILLER_204_417 ();
 FILLCELL_X32 FILLER_204_449 ();
 FILLCELL_X32 FILLER_204_481 ();
 FILLCELL_X32 FILLER_204_513 ();
 FILLCELL_X32 FILLER_204_545 ();
 FILLCELL_X32 FILLER_204_577 ();
 FILLCELL_X16 FILLER_204_609 ();
 FILLCELL_X4 FILLER_204_625 ();
 FILLCELL_X2 FILLER_204_629 ();
 FILLCELL_X32 FILLER_204_632 ();
 FILLCELL_X32 FILLER_204_664 ();
 FILLCELL_X32 FILLER_204_696 ();
 FILLCELL_X32 FILLER_204_728 ();
 FILLCELL_X32 FILLER_204_760 ();
 FILLCELL_X32 FILLER_204_792 ();
 FILLCELL_X32 FILLER_204_824 ();
 FILLCELL_X32 FILLER_204_856 ();
 FILLCELL_X32 FILLER_204_888 ();
 FILLCELL_X32 FILLER_204_920 ();
 FILLCELL_X32 FILLER_204_952 ();
 FILLCELL_X32 FILLER_204_984 ();
 FILLCELL_X32 FILLER_204_1016 ();
 FILLCELL_X32 FILLER_204_1048 ();
 FILLCELL_X32 FILLER_204_1080 ();
 FILLCELL_X32 FILLER_204_1112 ();
 FILLCELL_X32 FILLER_204_1144 ();
 FILLCELL_X32 FILLER_204_1176 ();
 FILLCELL_X32 FILLER_204_1208 ();
 FILLCELL_X32 FILLER_204_1240 ();
 FILLCELL_X32 FILLER_204_1272 ();
 FILLCELL_X32 FILLER_204_1304 ();
 FILLCELL_X32 FILLER_204_1336 ();
 FILLCELL_X32 FILLER_204_1368 ();
 FILLCELL_X32 FILLER_204_1400 ();
 FILLCELL_X32 FILLER_204_1432 ();
 FILLCELL_X32 FILLER_204_1464 ();
 FILLCELL_X32 FILLER_204_1496 ();
 FILLCELL_X32 FILLER_204_1528 ();
 FILLCELL_X32 FILLER_204_1560 ();
 FILLCELL_X32 FILLER_204_1592 ();
 FILLCELL_X32 FILLER_204_1624 ();
 FILLCELL_X32 FILLER_204_1656 ();
 FILLCELL_X32 FILLER_204_1688 ();
 FILLCELL_X32 FILLER_204_1720 ();
 FILLCELL_X32 FILLER_204_1752 ();
 FILLCELL_X32 FILLER_204_1784 ();
 FILLCELL_X32 FILLER_204_1816 ();
 FILLCELL_X32 FILLER_204_1848 ();
 FILLCELL_X8 FILLER_204_1880 ();
 FILLCELL_X4 FILLER_204_1888 ();
 FILLCELL_X2 FILLER_204_1892 ();
 FILLCELL_X32 FILLER_204_1895 ();
 FILLCELL_X32 FILLER_204_1927 ();
 FILLCELL_X32 FILLER_204_1959 ();
 FILLCELL_X32 FILLER_204_1991 ();
 FILLCELL_X32 FILLER_204_2023 ();
 FILLCELL_X32 FILLER_204_2055 ();
 FILLCELL_X32 FILLER_204_2087 ();
 FILLCELL_X32 FILLER_204_2119 ();
 FILLCELL_X32 FILLER_204_2151 ();
 FILLCELL_X32 FILLER_204_2183 ();
 FILLCELL_X32 FILLER_204_2215 ();
 FILLCELL_X32 FILLER_204_2247 ();
 FILLCELL_X32 FILLER_204_2279 ();
 FILLCELL_X32 FILLER_204_2311 ();
 FILLCELL_X32 FILLER_204_2343 ();
 FILLCELL_X32 FILLER_204_2375 ();
 FILLCELL_X32 FILLER_204_2407 ();
 FILLCELL_X32 FILLER_204_2439 ();
 FILLCELL_X32 FILLER_204_2471 ();
 FILLCELL_X32 FILLER_204_2503 ();
 FILLCELL_X32 FILLER_204_2535 ();
 FILLCELL_X32 FILLER_204_2567 ();
 FILLCELL_X2 FILLER_204_2599 ();
 FILLCELL_X1 FILLER_204_2601 ();
 FILLCELL_X32 FILLER_205_1 ();
 FILLCELL_X32 FILLER_205_33 ();
 FILLCELL_X32 FILLER_205_65 ();
 FILLCELL_X32 FILLER_205_97 ();
 FILLCELL_X32 FILLER_205_129 ();
 FILLCELL_X32 FILLER_205_161 ();
 FILLCELL_X32 FILLER_205_193 ();
 FILLCELL_X32 FILLER_205_225 ();
 FILLCELL_X32 FILLER_205_257 ();
 FILLCELL_X32 FILLER_205_289 ();
 FILLCELL_X32 FILLER_205_321 ();
 FILLCELL_X32 FILLER_205_353 ();
 FILLCELL_X32 FILLER_205_385 ();
 FILLCELL_X32 FILLER_205_417 ();
 FILLCELL_X32 FILLER_205_449 ();
 FILLCELL_X32 FILLER_205_481 ();
 FILLCELL_X32 FILLER_205_513 ();
 FILLCELL_X32 FILLER_205_545 ();
 FILLCELL_X32 FILLER_205_577 ();
 FILLCELL_X32 FILLER_205_609 ();
 FILLCELL_X32 FILLER_205_641 ();
 FILLCELL_X32 FILLER_205_673 ();
 FILLCELL_X32 FILLER_205_705 ();
 FILLCELL_X32 FILLER_205_737 ();
 FILLCELL_X32 FILLER_205_769 ();
 FILLCELL_X32 FILLER_205_801 ();
 FILLCELL_X32 FILLER_205_833 ();
 FILLCELL_X32 FILLER_205_865 ();
 FILLCELL_X32 FILLER_205_897 ();
 FILLCELL_X32 FILLER_205_929 ();
 FILLCELL_X32 FILLER_205_961 ();
 FILLCELL_X32 FILLER_205_993 ();
 FILLCELL_X32 FILLER_205_1025 ();
 FILLCELL_X32 FILLER_205_1057 ();
 FILLCELL_X32 FILLER_205_1089 ();
 FILLCELL_X32 FILLER_205_1121 ();
 FILLCELL_X32 FILLER_205_1153 ();
 FILLCELL_X32 FILLER_205_1185 ();
 FILLCELL_X32 FILLER_205_1217 ();
 FILLCELL_X8 FILLER_205_1249 ();
 FILLCELL_X4 FILLER_205_1257 ();
 FILLCELL_X2 FILLER_205_1261 ();
 FILLCELL_X32 FILLER_205_1264 ();
 FILLCELL_X32 FILLER_205_1296 ();
 FILLCELL_X32 FILLER_205_1328 ();
 FILLCELL_X32 FILLER_205_1360 ();
 FILLCELL_X32 FILLER_205_1392 ();
 FILLCELL_X32 FILLER_205_1424 ();
 FILLCELL_X32 FILLER_205_1456 ();
 FILLCELL_X32 FILLER_205_1488 ();
 FILLCELL_X32 FILLER_205_1520 ();
 FILLCELL_X32 FILLER_205_1552 ();
 FILLCELL_X32 FILLER_205_1584 ();
 FILLCELL_X32 FILLER_205_1616 ();
 FILLCELL_X32 FILLER_205_1648 ();
 FILLCELL_X32 FILLER_205_1680 ();
 FILLCELL_X32 FILLER_205_1712 ();
 FILLCELL_X32 FILLER_205_1744 ();
 FILLCELL_X32 FILLER_205_1776 ();
 FILLCELL_X32 FILLER_205_1808 ();
 FILLCELL_X32 FILLER_205_1840 ();
 FILLCELL_X32 FILLER_205_1872 ();
 FILLCELL_X32 FILLER_205_1904 ();
 FILLCELL_X32 FILLER_205_1936 ();
 FILLCELL_X32 FILLER_205_1968 ();
 FILLCELL_X32 FILLER_205_2000 ();
 FILLCELL_X32 FILLER_205_2032 ();
 FILLCELL_X32 FILLER_205_2064 ();
 FILLCELL_X32 FILLER_205_2096 ();
 FILLCELL_X32 FILLER_205_2128 ();
 FILLCELL_X32 FILLER_205_2160 ();
 FILLCELL_X32 FILLER_205_2192 ();
 FILLCELL_X32 FILLER_205_2224 ();
 FILLCELL_X32 FILLER_205_2256 ();
 FILLCELL_X32 FILLER_205_2288 ();
 FILLCELL_X32 FILLER_205_2320 ();
 FILLCELL_X32 FILLER_205_2352 ();
 FILLCELL_X32 FILLER_205_2384 ();
 FILLCELL_X32 FILLER_205_2416 ();
 FILLCELL_X32 FILLER_205_2448 ();
 FILLCELL_X32 FILLER_205_2480 ();
 FILLCELL_X8 FILLER_205_2512 ();
 FILLCELL_X4 FILLER_205_2520 ();
 FILLCELL_X2 FILLER_205_2524 ();
 FILLCELL_X32 FILLER_205_2527 ();
 FILLCELL_X32 FILLER_205_2559 ();
 FILLCELL_X8 FILLER_205_2591 ();
 FILLCELL_X2 FILLER_205_2599 ();
 FILLCELL_X1 FILLER_205_2601 ();
 FILLCELL_X32 FILLER_206_1 ();
 FILLCELL_X32 FILLER_206_33 ();
 FILLCELL_X32 FILLER_206_65 ();
 FILLCELL_X32 FILLER_206_97 ();
 FILLCELL_X32 FILLER_206_129 ();
 FILLCELL_X32 FILLER_206_161 ();
 FILLCELL_X32 FILLER_206_193 ();
 FILLCELL_X32 FILLER_206_225 ();
 FILLCELL_X32 FILLER_206_257 ();
 FILLCELL_X32 FILLER_206_289 ();
 FILLCELL_X32 FILLER_206_321 ();
 FILLCELL_X32 FILLER_206_353 ();
 FILLCELL_X32 FILLER_206_385 ();
 FILLCELL_X32 FILLER_206_417 ();
 FILLCELL_X32 FILLER_206_449 ();
 FILLCELL_X32 FILLER_206_481 ();
 FILLCELL_X32 FILLER_206_513 ();
 FILLCELL_X32 FILLER_206_545 ();
 FILLCELL_X32 FILLER_206_577 ();
 FILLCELL_X16 FILLER_206_609 ();
 FILLCELL_X4 FILLER_206_625 ();
 FILLCELL_X2 FILLER_206_629 ();
 FILLCELL_X32 FILLER_206_632 ();
 FILLCELL_X32 FILLER_206_664 ();
 FILLCELL_X32 FILLER_206_696 ();
 FILLCELL_X32 FILLER_206_728 ();
 FILLCELL_X32 FILLER_206_760 ();
 FILLCELL_X32 FILLER_206_792 ();
 FILLCELL_X32 FILLER_206_824 ();
 FILLCELL_X32 FILLER_206_856 ();
 FILLCELL_X32 FILLER_206_888 ();
 FILLCELL_X32 FILLER_206_920 ();
 FILLCELL_X32 FILLER_206_952 ();
 FILLCELL_X32 FILLER_206_984 ();
 FILLCELL_X32 FILLER_206_1016 ();
 FILLCELL_X32 FILLER_206_1048 ();
 FILLCELL_X32 FILLER_206_1080 ();
 FILLCELL_X32 FILLER_206_1112 ();
 FILLCELL_X32 FILLER_206_1144 ();
 FILLCELL_X32 FILLER_206_1176 ();
 FILLCELL_X32 FILLER_206_1208 ();
 FILLCELL_X32 FILLER_206_1240 ();
 FILLCELL_X32 FILLER_206_1272 ();
 FILLCELL_X32 FILLER_206_1304 ();
 FILLCELL_X32 FILLER_206_1336 ();
 FILLCELL_X32 FILLER_206_1368 ();
 FILLCELL_X32 FILLER_206_1400 ();
 FILLCELL_X32 FILLER_206_1432 ();
 FILLCELL_X32 FILLER_206_1464 ();
 FILLCELL_X32 FILLER_206_1496 ();
 FILLCELL_X32 FILLER_206_1528 ();
 FILLCELL_X32 FILLER_206_1560 ();
 FILLCELL_X32 FILLER_206_1592 ();
 FILLCELL_X32 FILLER_206_1624 ();
 FILLCELL_X32 FILLER_206_1656 ();
 FILLCELL_X32 FILLER_206_1688 ();
 FILLCELL_X32 FILLER_206_1720 ();
 FILLCELL_X32 FILLER_206_1752 ();
 FILLCELL_X32 FILLER_206_1784 ();
 FILLCELL_X32 FILLER_206_1816 ();
 FILLCELL_X32 FILLER_206_1848 ();
 FILLCELL_X8 FILLER_206_1880 ();
 FILLCELL_X4 FILLER_206_1888 ();
 FILLCELL_X2 FILLER_206_1892 ();
 FILLCELL_X32 FILLER_206_1895 ();
 FILLCELL_X32 FILLER_206_1927 ();
 FILLCELL_X32 FILLER_206_1959 ();
 FILLCELL_X32 FILLER_206_1991 ();
 FILLCELL_X32 FILLER_206_2023 ();
 FILLCELL_X32 FILLER_206_2055 ();
 FILLCELL_X32 FILLER_206_2087 ();
 FILLCELL_X32 FILLER_206_2119 ();
 FILLCELL_X32 FILLER_206_2151 ();
 FILLCELL_X32 FILLER_206_2183 ();
 FILLCELL_X32 FILLER_206_2215 ();
 FILLCELL_X32 FILLER_206_2247 ();
 FILLCELL_X32 FILLER_206_2279 ();
 FILLCELL_X32 FILLER_206_2311 ();
 FILLCELL_X32 FILLER_206_2343 ();
 FILLCELL_X32 FILLER_206_2375 ();
 FILLCELL_X32 FILLER_206_2407 ();
 FILLCELL_X32 FILLER_206_2439 ();
 FILLCELL_X32 FILLER_206_2471 ();
 FILLCELL_X32 FILLER_206_2503 ();
 FILLCELL_X32 FILLER_206_2535 ();
 FILLCELL_X32 FILLER_206_2567 ();
 FILLCELL_X2 FILLER_206_2599 ();
 FILLCELL_X1 FILLER_206_2601 ();
 FILLCELL_X32 FILLER_207_1 ();
 FILLCELL_X32 FILLER_207_33 ();
 FILLCELL_X32 FILLER_207_65 ();
 FILLCELL_X32 FILLER_207_97 ();
 FILLCELL_X32 FILLER_207_129 ();
 FILLCELL_X32 FILLER_207_161 ();
 FILLCELL_X32 FILLER_207_193 ();
 FILLCELL_X32 FILLER_207_225 ();
 FILLCELL_X32 FILLER_207_257 ();
 FILLCELL_X32 FILLER_207_289 ();
 FILLCELL_X32 FILLER_207_321 ();
 FILLCELL_X32 FILLER_207_353 ();
 FILLCELL_X32 FILLER_207_385 ();
 FILLCELL_X32 FILLER_207_417 ();
 FILLCELL_X32 FILLER_207_449 ();
 FILLCELL_X32 FILLER_207_481 ();
 FILLCELL_X32 FILLER_207_513 ();
 FILLCELL_X32 FILLER_207_545 ();
 FILLCELL_X32 FILLER_207_577 ();
 FILLCELL_X32 FILLER_207_609 ();
 FILLCELL_X32 FILLER_207_641 ();
 FILLCELL_X32 FILLER_207_673 ();
 FILLCELL_X32 FILLER_207_705 ();
 FILLCELL_X32 FILLER_207_737 ();
 FILLCELL_X32 FILLER_207_769 ();
 FILLCELL_X32 FILLER_207_801 ();
 FILLCELL_X32 FILLER_207_833 ();
 FILLCELL_X32 FILLER_207_865 ();
 FILLCELL_X32 FILLER_207_897 ();
 FILLCELL_X32 FILLER_207_929 ();
 FILLCELL_X32 FILLER_207_961 ();
 FILLCELL_X32 FILLER_207_993 ();
 FILLCELL_X32 FILLER_207_1025 ();
 FILLCELL_X32 FILLER_207_1057 ();
 FILLCELL_X32 FILLER_207_1089 ();
 FILLCELL_X32 FILLER_207_1121 ();
 FILLCELL_X32 FILLER_207_1153 ();
 FILLCELL_X32 FILLER_207_1185 ();
 FILLCELL_X32 FILLER_207_1217 ();
 FILLCELL_X8 FILLER_207_1249 ();
 FILLCELL_X4 FILLER_207_1257 ();
 FILLCELL_X2 FILLER_207_1261 ();
 FILLCELL_X32 FILLER_207_1264 ();
 FILLCELL_X32 FILLER_207_1296 ();
 FILLCELL_X32 FILLER_207_1328 ();
 FILLCELL_X32 FILLER_207_1360 ();
 FILLCELL_X32 FILLER_207_1392 ();
 FILLCELL_X32 FILLER_207_1424 ();
 FILLCELL_X32 FILLER_207_1456 ();
 FILLCELL_X32 FILLER_207_1488 ();
 FILLCELL_X32 FILLER_207_1520 ();
 FILLCELL_X32 FILLER_207_1552 ();
 FILLCELL_X32 FILLER_207_1584 ();
 FILLCELL_X32 FILLER_207_1616 ();
 FILLCELL_X32 FILLER_207_1648 ();
 FILLCELL_X32 FILLER_207_1680 ();
 FILLCELL_X32 FILLER_207_1712 ();
 FILLCELL_X32 FILLER_207_1744 ();
 FILLCELL_X32 FILLER_207_1776 ();
 FILLCELL_X32 FILLER_207_1808 ();
 FILLCELL_X32 FILLER_207_1840 ();
 FILLCELL_X32 FILLER_207_1872 ();
 FILLCELL_X32 FILLER_207_1904 ();
 FILLCELL_X32 FILLER_207_1936 ();
 FILLCELL_X32 FILLER_207_1968 ();
 FILLCELL_X32 FILLER_207_2000 ();
 FILLCELL_X32 FILLER_207_2032 ();
 FILLCELL_X32 FILLER_207_2064 ();
 FILLCELL_X32 FILLER_207_2096 ();
 FILLCELL_X32 FILLER_207_2128 ();
 FILLCELL_X32 FILLER_207_2160 ();
 FILLCELL_X32 FILLER_207_2192 ();
 FILLCELL_X32 FILLER_207_2224 ();
 FILLCELL_X32 FILLER_207_2256 ();
 FILLCELL_X32 FILLER_207_2288 ();
 FILLCELL_X32 FILLER_207_2320 ();
 FILLCELL_X32 FILLER_207_2352 ();
 FILLCELL_X32 FILLER_207_2384 ();
 FILLCELL_X32 FILLER_207_2416 ();
 FILLCELL_X32 FILLER_207_2448 ();
 FILLCELL_X32 FILLER_207_2480 ();
 FILLCELL_X8 FILLER_207_2512 ();
 FILLCELL_X4 FILLER_207_2520 ();
 FILLCELL_X2 FILLER_207_2524 ();
 FILLCELL_X32 FILLER_207_2527 ();
 FILLCELL_X32 FILLER_207_2559 ();
 FILLCELL_X8 FILLER_207_2591 ();
 FILLCELL_X2 FILLER_207_2599 ();
 FILLCELL_X1 FILLER_207_2601 ();
 FILLCELL_X32 FILLER_208_1 ();
 FILLCELL_X32 FILLER_208_33 ();
 FILLCELL_X32 FILLER_208_65 ();
 FILLCELL_X32 FILLER_208_97 ();
 FILLCELL_X32 FILLER_208_129 ();
 FILLCELL_X32 FILLER_208_161 ();
 FILLCELL_X32 FILLER_208_193 ();
 FILLCELL_X32 FILLER_208_225 ();
 FILLCELL_X32 FILLER_208_257 ();
 FILLCELL_X32 FILLER_208_289 ();
 FILLCELL_X32 FILLER_208_321 ();
 FILLCELL_X32 FILLER_208_353 ();
 FILLCELL_X32 FILLER_208_385 ();
 FILLCELL_X32 FILLER_208_417 ();
 FILLCELL_X32 FILLER_208_449 ();
 FILLCELL_X32 FILLER_208_481 ();
 FILLCELL_X32 FILLER_208_513 ();
 FILLCELL_X32 FILLER_208_545 ();
 FILLCELL_X32 FILLER_208_577 ();
 FILLCELL_X16 FILLER_208_609 ();
 FILLCELL_X4 FILLER_208_625 ();
 FILLCELL_X2 FILLER_208_629 ();
 FILLCELL_X32 FILLER_208_632 ();
 FILLCELL_X32 FILLER_208_664 ();
 FILLCELL_X32 FILLER_208_696 ();
 FILLCELL_X32 FILLER_208_728 ();
 FILLCELL_X32 FILLER_208_760 ();
 FILLCELL_X32 FILLER_208_792 ();
 FILLCELL_X32 FILLER_208_824 ();
 FILLCELL_X32 FILLER_208_856 ();
 FILLCELL_X32 FILLER_208_888 ();
 FILLCELL_X32 FILLER_208_920 ();
 FILLCELL_X32 FILLER_208_952 ();
 FILLCELL_X32 FILLER_208_984 ();
 FILLCELL_X32 FILLER_208_1016 ();
 FILLCELL_X32 FILLER_208_1048 ();
 FILLCELL_X32 FILLER_208_1080 ();
 FILLCELL_X32 FILLER_208_1112 ();
 FILLCELL_X32 FILLER_208_1144 ();
 FILLCELL_X32 FILLER_208_1176 ();
 FILLCELL_X32 FILLER_208_1208 ();
 FILLCELL_X32 FILLER_208_1240 ();
 FILLCELL_X32 FILLER_208_1272 ();
 FILLCELL_X32 FILLER_208_1304 ();
 FILLCELL_X32 FILLER_208_1336 ();
 FILLCELL_X32 FILLER_208_1368 ();
 FILLCELL_X32 FILLER_208_1400 ();
 FILLCELL_X32 FILLER_208_1432 ();
 FILLCELL_X32 FILLER_208_1464 ();
 FILLCELL_X32 FILLER_208_1496 ();
 FILLCELL_X32 FILLER_208_1528 ();
 FILLCELL_X32 FILLER_208_1560 ();
 FILLCELL_X32 FILLER_208_1592 ();
 FILLCELL_X32 FILLER_208_1624 ();
 FILLCELL_X32 FILLER_208_1656 ();
 FILLCELL_X32 FILLER_208_1688 ();
 FILLCELL_X32 FILLER_208_1720 ();
 FILLCELL_X32 FILLER_208_1752 ();
 FILLCELL_X32 FILLER_208_1784 ();
 FILLCELL_X32 FILLER_208_1816 ();
 FILLCELL_X32 FILLER_208_1848 ();
 FILLCELL_X8 FILLER_208_1880 ();
 FILLCELL_X4 FILLER_208_1888 ();
 FILLCELL_X2 FILLER_208_1892 ();
 FILLCELL_X32 FILLER_208_1895 ();
 FILLCELL_X32 FILLER_208_1927 ();
 FILLCELL_X32 FILLER_208_1959 ();
 FILLCELL_X32 FILLER_208_1991 ();
 FILLCELL_X32 FILLER_208_2023 ();
 FILLCELL_X32 FILLER_208_2055 ();
 FILLCELL_X32 FILLER_208_2087 ();
 FILLCELL_X32 FILLER_208_2119 ();
 FILLCELL_X32 FILLER_208_2151 ();
 FILLCELL_X32 FILLER_208_2183 ();
 FILLCELL_X32 FILLER_208_2215 ();
 FILLCELL_X32 FILLER_208_2247 ();
 FILLCELL_X32 FILLER_208_2279 ();
 FILLCELL_X32 FILLER_208_2311 ();
 FILLCELL_X32 FILLER_208_2343 ();
 FILLCELL_X32 FILLER_208_2375 ();
 FILLCELL_X32 FILLER_208_2407 ();
 FILLCELL_X32 FILLER_208_2439 ();
 FILLCELL_X32 FILLER_208_2471 ();
 FILLCELL_X32 FILLER_208_2503 ();
 FILLCELL_X32 FILLER_208_2535 ();
 FILLCELL_X32 FILLER_208_2567 ();
 FILLCELL_X2 FILLER_208_2599 ();
 FILLCELL_X1 FILLER_208_2601 ();
 FILLCELL_X32 FILLER_209_1 ();
 FILLCELL_X32 FILLER_209_33 ();
 FILLCELL_X32 FILLER_209_65 ();
 FILLCELL_X32 FILLER_209_97 ();
 FILLCELL_X32 FILLER_209_129 ();
 FILLCELL_X32 FILLER_209_161 ();
 FILLCELL_X32 FILLER_209_193 ();
 FILLCELL_X32 FILLER_209_225 ();
 FILLCELL_X32 FILLER_209_257 ();
 FILLCELL_X32 FILLER_209_289 ();
 FILLCELL_X32 FILLER_209_321 ();
 FILLCELL_X32 FILLER_209_353 ();
 FILLCELL_X32 FILLER_209_385 ();
 FILLCELL_X32 FILLER_209_417 ();
 FILLCELL_X32 FILLER_209_449 ();
 FILLCELL_X32 FILLER_209_481 ();
 FILLCELL_X32 FILLER_209_513 ();
 FILLCELL_X32 FILLER_209_545 ();
 FILLCELL_X32 FILLER_209_577 ();
 FILLCELL_X32 FILLER_209_609 ();
 FILLCELL_X32 FILLER_209_641 ();
 FILLCELL_X32 FILLER_209_673 ();
 FILLCELL_X32 FILLER_209_705 ();
 FILLCELL_X32 FILLER_209_737 ();
 FILLCELL_X32 FILLER_209_769 ();
 FILLCELL_X32 FILLER_209_801 ();
 FILLCELL_X32 FILLER_209_833 ();
 FILLCELL_X32 FILLER_209_865 ();
 FILLCELL_X32 FILLER_209_897 ();
 FILLCELL_X32 FILLER_209_929 ();
 FILLCELL_X32 FILLER_209_961 ();
 FILLCELL_X32 FILLER_209_993 ();
 FILLCELL_X32 FILLER_209_1025 ();
 FILLCELL_X32 FILLER_209_1057 ();
 FILLCELL_X32 FILLER_209_1089 ();
 FILLCELL_X32 FILLER_209_1121 ();
 FILLCELL_X32 FILLER_209_1153 ();
 FILLCELL_X32 FILLER_209_1185 ();
 FILLCELL_X32 FILLER_209_1217 ();
 FILLCELL_X8 FILLER_209_1249 ();
 FILLCELL_X4 FILLER_209_1257 ();
 FILLCELL_X2 FILLER_209_1261 ();
 FILLCELL_X32 FILLER_209_1264 ();
 FILLCELL_X32 FILLER_209_1296 ();
 FILLCELL_X32 FILLER_209_1328 ();
 FILLCELL_X32 FILLER_209_1360 ();
 FILLCELL_X32 FILLER_209_1392 ();
 FILLCELL_X32 FILLER_209_1424 ();
 FILLCELL_X32 FILLER_209_1456 ();
 FILLCELL_X32 FILLER_209_1488 ();
 FILLCELL_X32 FILLER_209_1520 ();
 FILLCELL_X32 FILLER_209_1552 ();
 FILLCELL_X32 FILLER_209_1584 ();
 FILLCELL_X32 FILLER_209_1616 ();
 FILLCELL_X32 FILLER_209_1648 ();
 FILLCELL_X32 FILLER_209_1680 ();
 FILLCELL_X32 FILLER_209_1712 ();
 FILLCELL_X32 FILLER_209_1744 ();
 FILLCELL_X32 FILLER_209_1776 ();
 FILLCELL_X32 FILLER_209_1808 ();
 FILLCELL_X32 FILLER_209_1840 ();
 FILLCELL_X32 FILLER_209_1872 ();
 FILLCELL_X32 FILLER_209_1904 ();
 FILLCELL_X32 FILLER_209_1936 ();
 FILLCELL_X32 FILLER_209_1968 ();
 FILLCELL_X32 FILLER_209_2000 ();
 FILLCELL_X32 FILLER_209_2032 ();
 FILLCELL_X32 FILLER_209_2064 ();
 FILLCELL_X32 FILLER_209_2096 ();
 FILLCELL_X32 FILLER_209_2128 ();
 FILLCELL_X32 FILLER_209_2160 ();
 FILLCELL_X32 FILLER_209_2192 ();
 FILLCELL_X32 FILLER_209_2224 ();
 FILLCELL_X32 FILLER_209_2256 ();
 FILLCELL_X32 FILLER_209_2288 ();
 FILLCELL_X32 FILLER_209_2320 ();
 FILLCELL_X32 FILLER_209_2352 ();
 FILLCELL_X32 FILLER_209_2384 ();
 FILLCELL_X32 FILLER_209_2416 ();
 FILLCELL_X32 FILLER_209_2448 ();
 FILLCELL_X32 FILLER_209_2480 ();
 FILLCELL_X8 FILLER_209_2512 ();
 FILLCELL_X4 FILLER_209_2520 ();
 FILLCELL_X2 FILLER_209_2524 ();
 FILLCELL_X32 FILLER_209_2527 ();
 FILLCELL_X32 FILLER_209_2559 ();
 FILLCELL_X8 FILLER_209_2591 ();
 FILLCELL_X2 FILLER_209_2599 ();
 FILLCELL_X1 FILLER_209_2601 ();
 FILLCELL_X32 FILLER_210_1 ();
 FILLCELL_X32 FILLER_210_33 ();
 FILLCELL_X32 FILLER_210_65 ();
 FILLCELL_X32 FILLER_210_97 ();
 FILLCELL_X32 FILLER_210_129 ();
 FILLCELL_X32 FILLER_210_161 ();
 FILLCELL_X32 FILLER_210_193 ();
 FILLCELL_X32 FILLER_210_225 ();
 FILLCELL_X32 FILLER_210_257 ();
 FILLCELL_X32 FILLER_210_289 ();
 FILLCELL_X32 FILLER_210_321 ();
 FILLCELL_X32 FILLER_210_353 ();
 FILLCELL_X32 FILLER_210_385 ();
 FILLCELL_X32 FILLER_210_417 ();
 FILLCELL_X32 FILLER_210_449 ();
 FILLCELL_X32 FILLER_210_481 ();
 FILLCELL_X32 FILLER_210_513 ();
 FILLCELL_X32 FILLER_210_545 ();
 FILLCELL_X32 FILLER_210_577 ();
 FILLCELL_X16 FILLER_210_609 ();
 FILLCELL_X4 FILLER_210_625 ();
 FILLCELL_X2 FILLER_210_629 ();
 FILLCELL_X32 FILLER_210_632 ();
 FILLCELL_X32 FILLER_210_664 ();
 FILLCELL_X32 FILLER_210_696 ();
 FILLCELL_X32 FILLER_210_728 ();
 FILLCELL_X32 FILLER_210_760 ();
 FILLCELL_X32 FILLER_210_792 ();
 FILLCELL_X32 FILLER_210_824 ();
 FILLCELL_X32 FILLER_210_856 ();
 FILLCELL_X32 FILLER_210_888 ();
 FILLCELL_X32 FILLER_210_920 ();
 FILLCELL_X32 FILLER_210_952 ();
 FILLCELL_X32 FILLER_210_984 ();
 FILLCELL_X32 FILLER_210_1016 ();
 FILLCELL_X32 FILLER_210_1048 ();
 FILLCELL_X32 FILLER_210_1080 ();
 FILLCELL_X32 FILLER_210_1112 ();
 FILLCELL_X32 FILLER_210_1144 ();
 FILLCELL_X32 FILLER_210_1176 ();
 FILLCELL_X32 FILLER_210_1208 ();
 FILLCELL_X32 FILLER_210_1240 ();
 FILLCELL_X32 FILLER_210_1272 ();
 FILLCELL_X32 FILLER_210_1304 ();
 FILLCELL_X32 FILLER_210_1336 ();
 FILLCELL_X32 FILLER_210_1368 ();
 FILLCELL_X32 FILLER_210_1400 ();
 FILLCELL_X32 FILLER_210_1432 ();
 FILLCELL_X32 FILLER_210_1464 ();
 FILLCELL_X32 FILLER_210_1496 ();
 FILLCELL_X32 FILLER_210_1528 ();
 FILLCELL_X32 FILLER_210_1560 ();
 FILLCELL_X32 FILLER_210_1592 ();
 FILLCELL_X32 FILLER_210_1624 ();
 FILLCELL_X32 FILLER_210_1656 ();
 FILLCELL_X32 FILLER_210_1688 ();
 FILLCELL_X32 FILLER_210_1720 ();
 FILLCELL_X32 FILLER_210_1752 ();
 FILLCELL_X32 FILLER_210_1784 ();
 FILLCELL_X32 FILLER_210_1816 ();
 FILLCELL_X32 FILLER_210_1848 ();
 FILLCELL_X8 FILLER_210_1880 ();
 FILLCELL_X4 FILLER_210_1888 ();
 FILLCELL_X2 FILLER_210_1892 ();
 FILLCELL_X32 FILLER_210_1895 ();
 FILLCELL_X32 FILLER_210_1927 ();
 FILLCELL_X32 FILLER_210_1959 ();
 FILLCELL_X32 FILLER_210_1991 ();
 FILLCELL_X32 FILLER_210_2023 ();
 FILLCELL_X32 FILLER_210_2055 ();
 FILLCELL_X32 FILLER_210_2087 ();
 FILLCELL_X32 FILLER_210_2119 ();
 FILLCELL_X32 FILLER_210_2151 ();
 FILLCELL_X32 FILLER_210_2183 ();
 FILLCELL_X32 FILLER_210_2215 ();
 FILLCELL_X32 FILLER_210_2247 ();
 FILLCELL_X32 FILLER_210_2279 ();
 FILLCELL_X32 FILLER_210_2311 ();
 FILLCELL_X32 FILLER_210_2343 ();
 FILLCELL_X32 FILLER_210_2375 ();
 FILLCELL_X32 FILLER_210_2407 ();
 FILLCELL_X32 FILLER_210_2439 ();
 FILLCELL_X32 FILLER_210_2471 ();
 FILLCELL_X32 FILLER_210_2503 ();
 FILLCELL_X32 FILLER_210_2535 ();
 FILLCELL_X32 FILLER_210_2567 ();
 FILLCELL_X2 FILLER_210_2599 ();
 FILLCELL_X1 FILLER_210_2601 ();
 FILLCELL_X32 FILLER_211_1 ();
 FILLCELL_X32 FILLER_211_33 ();
 FILLCELL_X32 FILLER_211_65 ();
 FILLCELL_X32 FILLER_211_97 ();
 FILLCELL_X32 FILLER_211_129 ();
 FILLCELL_X32 FILLER_211_161 ();
 FILLCELL_X32 FILLER_211_193 ();
 FILLCELL_X32 FILLER_211_225 ();
 FILLCELL_X32 FILLER_211_257 ();
 FILLCELL_X32 FILLER_211_289 ();
 FILLCELL_X32 FILLER_211_321 ();
 FILLCELL_X32 FILLER_211_353 ();
 FILLCELL_X32 FILLER_211_385 ();
 FILLCELL_X32 FILLER_211_417 ();
 FILLCELL_X32 FILLER_211_449 ();
 FILLCELL_X32 FILLER_211_481 ();
 FILLCELL_X32 FILLER_211_513 ();
 FILLCELL_X32 FILLER_211_545 ();
 FILLCELL_X32 FILLER_211_577 ();
 FILLCELL_X32 FILLER_211_609 ();
 FILLCELL_X32 FILLER_211_641 ();
 FILLCELL_X32 FILLER_211_673 ();
 FILLCELL_X32 FILLER_211_705 ();
 FILLCELL_X32 FILLER_211_737 ();
 FILLCELL_X32 FILLER_211_769 ();
 FILLCELL_X32 FILLER_211_801 ();
 FILLCELL_X32 FILLER_211_833 ();
 FILLCELL_X32 FILLER_211_865 ();
 FILLCELL_X32 FILLER_211_897 ();
 FILLCELL_X32 FILLER_211_929 ();
 FILLCELL_X32 FILLER_211_961 ();
 FILLCELL_X32 FILLER_211_993 ();
 FILLCELL_X32 FILLER_211_1025 ();
 FILLCELL_X32 FILLER_211_1057 ();
 FILLCELL_X32 FILLER_211_1089 ();
 FILLCELL_X32 FILLER_211_1121 ();
 FILLCELL_X32 FILLER_211_1153 ();
 FILLCELL_X32 FILLER_211_1185 ();
 FILLCELL_X32 FILLER_211_1217 ();
 FILLCELL_X8 FILLER_211_1249 ();
 FILLCELL_X4 FILLER_211_1257 ();
 FILLCELL_X2 FILLER_211_1261 ();
 FILLCELL_X32 FILLER_211_1264 ();
 FILLCELL_X32 FILLER_211_1296 ();
 FILLCELL_X32 FILLER_211_1328 ();
 FILLCELL_X32 FILLER_211_1360 ();
 FILLCELL_X32 FILLER_211_1392 ();
 FILLCELL_X32 FILLER_211_1424 ();
 FILLCELL_X32 FILLER_211_1456 ();
 FILLCELL_X32 FILLER_211_1488 ();
 FILLCELL_X32 FILLER_211_1520 ();
 FILLCELL_X32 FILLER_211_1552 ();
 FILLCELL_X32 FILLER_211_1584 ();
 FILLCELL_X32 FILLER_211_1616 ();
 FILLCELL_X32 FILLER_211_1648 ();
 FILLCELL_X32 FILLER_211_1680 ();
 FILLCELL_X32 FILLER_211_1712 ();
 FILLCELL_X32 FILLER_211_1744 ();
 FILLCELL_X32 FILLER_211_1776 ();
 FILLCELL_X32 FILLER_211_1808 ();
 FILLCELL_X32 FILLER_211_1840 ();
 FILLCELL_X32 FILLER_211_1872 ();
 FILLCELL_X32 FILLER_211_1904 ();
 FILLCELL_X32 FILLER_211_1936 ();
 FILLCELL_X32 FILLER_211_1968 ();
 FILLCELL_X32 FILLER_211_2000 ();
 FILLCELL_X32 FILLER_211_2032 ();
 FILLCELL_X32 FILLER_211_2064 ();
 FILLCELL_X32 FILLER_211_2096 ();
 FILLCELL_X32 FILLER_211_2128 ();
 FILLCELL_X32 FILLER_211_2160 ();
 FILLCELL_X32 FILLER_211_2192 ();
 FILLCELL_X32 FILLER_211_2224 ();
 FILLCELL_X32 FILLER_211_2256 ();
 FILLCELL_X32 FILLER_211_2288 ();
 FILLCELL_X32 FILLER_211_2320 ();
 FILLCELL_X32 FILLER_211_2352 ();
 FILLCELL_X32 FILLER_211_2384 ();
 FILLCELL_X32 FILLER_211_2416 ();
 FILLCELL_X32 FILLER_211_2448 ();
 FILLCELL_X32 FILLER_211_2480 ();
 FILLCELL_X8 FILLER_211_2512 ();
 FILLCELL_X4 FILLER_211_2520 ();
 FILLCELL_X2 FILLER_211_2524 ();
 FILLCELL_X32 FILLER_211_2527 ();
 FILLCELL_X32 FILLER_211_2559 ();
 FILLCELL_X8 FILLER_211_2591 ();
 FILLCELL_X2 FILLER_211_2599 ();
 FILLCELL_X1 FILLER_211_2601 ();
 FILLCELL_X32 FILLER_212_1 ();
 FILLCELL_X32 FILLER_212_33 ();
 FILLCELL_X32 FILLER_212_65 ();
 FILLCELL_X32 FILLER_212_97 ();
 FILLCELL_X32 FILLER_212_129 ();
 FILLCELL_X32 FILLER_212_161 ();
 FILLCELL_X32 FILLER_212_193 ();
 FILLCELL_X32 FILLER_212_225 ();
 FILLCELL_X32 FILLER_212_257 ();
 FILLCELL_X32 FILLER_212_289 ();
 FILLCELL_X32 FILLER_212_321 ();
 FILLCELL_X32 FILLER_212_353 ();
 FILLCELL_X32 FILLER_212_385 ();
 FILLCELL_X32 FILLER_212_417 ();
 FILLCELL_X32 FILLER_212_449 ();
 FILLCELL_X32 FILLER_212_481 ();
 FILLCELL_X32 FILLER_212_513 ();
 FILLCELL_X32 FILLER_212_545 ();
 FILLCELL_X32 FILLER_212_577 ();
 FILLCELL_X16 FILLER_212_609 ();
 FILLCELL_X4 FILLER_212_625 ();
 FILLCELL_X2 FILLER_212_629 ();
 FILLCELL_X32 FILLER_212_632 ();
 FILLCELL_X32 FILLER_212_664 ();
 FILLCELL_X32 FILLER_212_696 ();
 FILLCELL_X32 FILLER_212_728 ();
 FILLCELL_X32 FILLER_212_760 ();
 FILLCELL_X32 FILLER_212_792 ();
 FILLCELL_X32 FILLER_212_824 ();
 FILLCELL_X32 FILLER_212_856 ();
 FILLCELL_X32 FILLER_212_888 ();
 FILLCELL_X32 FILLER_212_920 ();
 FILLCELL_X32 FILLER_212_952 ();
 FILLCELL_X32 FILLER_212_984 ();
 FILLCELL_X32 FILLER_212_1016 ();
 FILLCELL_X32 FILLER_212_1048 ();
 FILLCELL_X32 FILLER_212_1080 ();
 FILLCELL_X32 FILLER_212_1112 ();
 FILLCELL_X32 FILLER_212_1144 ();
 FILLCELL_X32 FILLER_212_1176 ();
 FILLCELL_X32 FILLER_212_1208 ();
 FILLCELL_X32 FILLER_212_1240 ();
 FILLCELL_X32 FILLER_212_1272 ();
 FILLCELL_X32 FILLER_212_1304 ();
 FILLCELL_X32 FILLER_212_1336 ();
 FILLCELL_X32 FILLER_212_1368 ();
 FILLCELL_X32 FILLER_212_1400 ();
 FILLCELL_X32 FILLER_212_1432 ();
 FILLCELL_X32 FILLER_212_1464 ();
 FILLCELL_X32 FILLER_212_1496 ();
 FILLCELL_X32 FILLER_212_1528 ();
 FILLCELL_X32 FILLER_212_1560 ();
 FILLCELL_X32 FILLER_212_1592 ();
 FILLCELL_X32 FILLER_212_1624 ();
 FILLCELL_X32 FILLER_212_1656 ();
 FILLCELL_X32 FILLER_212_1688 ();
 FILLCELL_X32 FILLER_212_1720 ();
 FILLCELL_X32 FILLER_212_1752 ();
 FILLCELL_X32 FILLER_212_1784 ();
 FILLCELL_X32 FILLER_212_1816 ();
 FILLCELL_X32 FILLER_212_1848 ();
 FILLCELL_X8 FILLER_212_1880 ();
 FILLCELL_X4 FILLER_212_1888 ();
 FILLCELL_X2 FILLER_212_1892 ();
 FILLCELL_X32 FILLER_212_1895 ();
 FILLCELL_X32 FILLER_212_1927 ();
 FILLCELL_X32 FILLER_212_1959 ();
 FILLCELL_X32 FILLER_212_1991 ();
 FILLCELL_X32 FILLER_212_2023 ();
 FILLCELL_X32 FILLER_212_2055 ();
 FILLCELL_X32 FILLER_212_2087 ();
 FILLCELL_X32 FILLER_212_2119 ();
 FILLCELL_X32 FILLER_212_2151 ();
 FILLCELL_X32 FILLER_212_2183 ();
 FILLCELL_X32 FILLER_212_2215 ();
 FILLCELL_X32 FILLER_212_2247 ();
 FILLCELL_X32 FILLER_212_2279 ();
 FILLCELL_X32 FILLER_212_2311 ();
 FILLCELL_X32 FILLER_212_2343 ();
 FILLCELL_X32 FILLER_212_2375 ();
 FILLCELL_X32 FILLER_212_2407 ();
 FILLCELL_X32 FILLER_212_2439 ();
 FILLCELL_X32 FILLER_212_2471 ();
 FILLCELL_X32 FILLER_212_2503 ();
 FILLCELL_X32 FILLER_212_2535 ();
 FILLCELL_X32 FILLER_212_2567 ();
 FILLCELL_X2 FILLER_212_2599 ();
 FILLCELL_X1 FILLER_212_2601 ();
 FILLCELL_X32 FILLER_213_1 ();
 FILLCELL_X32 FILLER_213_33 ();
 FILLCELL_X32 FILLER_213_65 ();
 FILLCELL_X32 FILLER_213_97 ();
 FILLCELL_X32 FILLER_213_129 ();
 FILLCELL_X32 FILLER_213_161 ();
 FILLCELL_X32 FILLER_213_193 ();
 FILLCELL_X32 FILLER_213_225 ();
 FILLCELL_X32 FILLER_213_257 ();
 FILLCELL_X32 FILLER_213_289 ();
 FILLCELL_X32 FILLER_213_321 ();
 FILLCELL_X32 FILLER_213_353 ();
 FILLCELL_X32 FILLER_213_385 ();
 FILLCELL_X32 FILLER_213_417 ();
 FILLCELL_X32 FILLER_213_449 ();
 FILLCELL_X32 FILLER_213_481 ();
 FILLCELL_X32 FILLER_213_513 ();
 FILLCELL_X32 FILLER_213_545 ();
 FILLCELL_X32 FILLER_213_577 ();
 FILLCELL_X32 FILLER_213_609 ();
 FILLCELL_X32 FILLER_213_641 ();
 FILLCELL_X32 FILLER_213_673 ();
 FILLCELL_X32 FILLER_213_705 ();
 FILLCELL_X32 FILLER_213_737 ();
 FILLCELL_X32 FILLER_213_769 ();
 FILLCELL_X32 FILLER_213_801 ();
 FILLCELL_X32 FILLER_213_833 ();
 FILLCELL_X32 FILLER_213_865 ();
 FILLCELL_X32 FILLER_213_897 ();
 FILLCELL_X32 FILLER_213_929 ();
 FILLCELL_X32 FILLER_213_961 ();
 FILLCELL_X32 FILLER_213_993 ();
 FILLCELL_X32 FILLER_213_1025 ();
 FILLCELL_X32 FILLER_213_1057 ();
 FILLCELL_X32 FILLER_213_1089 ();
 FILLCELL_X32 FILLER_213_1121 ();
 FILLCELL_X32 FILLER_213_1153 ();
 FILLCELL_X32 FILLER_213_1185 ();
 FILLCELL_X32 FILLER_213_1217 ();
 FILLCELL_X8 FILLER_213_1249 ();
 FILLCELL_X4 FILLER_213_1257 ();
 FILLCELL_X2 FILLER_213_1261 ();
 FILLCELL_X32 FILLER_213_1264 ();
 FILLCELL_X32 FILLER_213_1296 ();
 FILLCELL_X32 FILLER_213_1328 ();
 FILLCELL_X32 FILLER_213_1360 ();
 FILLCELL_X32 FILLER_213_1392 ();
 FILLCELL_X32 FILLER_213_1424 ();
 FILLCELL_X32 FILLER_213_1456 ();
 FILLCELL_X32 FILLER_213_1488 ();
 FILLCELL_X32 FILLER_213_1520 ();
 FILLCELL_X32 FILLER_213_1552 ();
 FILLCELL_X32 FILLER_213_1584 ();
 FILLCELL_X32 FILLER_213_1616 ();
 FILLCELL_X32 FILLER_213_1648 ();
 FILLCELL_X32 FILLER_213_1680 ();
 FILLCELL_X32 FILLER_213_1712 ();
 FILLCELL_X32 FILLER_213_1744 ();
 FILLCELL_X32 FILLER_213_1776 ();
 FILLCELL_X32 FILLER_213_1808 ();
 FILLCELL_X32 FILLER_213_1840 ();
 FILLCELL_X32 FILLER_213_1872 ();
 FILLCELL_X32 FILLER_213_1904 ();
 FILLCELL_X32 FILLER_213_1936 ();
 FILLCELL_X32 FILLER_213_1968 ();
 FILLCELL_X32 FILLER_213_2000 ();
 FILLCELL_X32 FILLER_213_2032 ();
 FILLCELL_X32 FILLER_213_2064 ();
 FILLCELL_X32 FILLER_213_2096 ();
 FILLCELL_X32 FILLER_213_2128 ();
 FILLCELL_X32 FILLER_213_2160 ();
 FILLCELL_X32 FILLER_213_2192 ();
 FILLCELL_X32 FILLER_213_2224 ();
 FILLCELL_X32 FILLER_213_2256 ();
 FILLCELL_X32 FILLER_213_2288 ();
 FILLCELL_X32 FILLER_213_2320 ();
 FILLCELL_X32 FILLER_213_2352 ();
 FILLCELL_X32 FILLER_213_2384 ();
 FILLCELL_X32 FILLER_213_2416 ();
 FILLCELL_X32 FILLER_213_2448 ();
 FILLCELL_X32 FILLER_213_2480 ();
 FILLCELL_X8 FILLER_213_2512 ();
 FILLCELL_X4 FILLER_213_2520 ();
 FILLCELL_X2 FILLER_213_2524 ();
 FILLCELL_X32 FILLER_213_2527 ();
 FILLCELL_X32 FILLER_213_2559 ();
 FILLCELL_X8 FILLER_213_2591 ();
 FILLCELL_X2 FILLER_213_2599 ();
 FILLCELL_X1 FILLER_213_2601 ();
 FILLCELL_X32 FILLER_214_1 ();
 FILLCELL_X32 FILLER_214_33 ();
 FILLCELL_X32 FILLER_214_65 ();
 FILLCELL_X32 FILLER_214_97 ();
 FILLCELL_X32 FILLER_214_129 ();
 FILLCELL_X32 FILLER_214_161 ();
 FILLCELL_X32 FILLER_214_193 ();
 FILLCELL_X32 FILLER_214_225 ();
 FILLCELL_X32 FILLER_214_257 ();
 FILLCELL_X32 FILLER_214_289 ();
 FILLCELL_X32 FILLER_214_321 ();
 FILLCELL_X32 FILLER_214_353 ();
 FILLCELL_X32 FILLER_214_385 ();
 FILLCELL_X32 FILLER_214_417 ();
 FILLCELL_X32 FILLER_214_449 ();
 FILLCELL_X32 FILLER_214_481 ();
 FILLCELL_X32 FILLER_214_513 ();
 FILLCELL_X32 FILLER_214_545 ();
 FILLCELL_X32 FILLER_214_577 ();
 FILLCELL_X16 FILLER_214_609 ();
 FILLCELL_X4 FILLER_214_625 ();
 FILLCELL_X2 FILLER_214_629 ();
 FILLCELL_X32 FILLER_214_632 ();
 FILLCELL_X32 FILLER_214_664 ();
 FILLCELL_X32 FILLER_214_696 ();
 FILLCELL_X32 FILLER_214_728 ();
 FILLCELL_X32 FILLER_214_760 ();
 FILLCELL_X32 FILLER_214_792 ();
 FILLCELL_X32 FILLER_214_824 ();
 FILLCELL_X32 FILLER_214_856 ();
 FILLCELL_X32 FILLER_214_888 ();
 FILLCELL_X32 FILLER_214_920 ();
 FILLCELL_X32 FILLER_214_952 ();
 FILLCELL_X32 FILLER_214_984 ();
 FILLCELL_X32 FILLER_214_1016 ();
 FILLCELL_X32 FILLER_214_1048 ();
 FILLCELL_X32 FILLER_214_1080 ();
 FILLCELL_X32 FILLER_214_1112 ();
 FILLCELL_X32 FILLER_214_1144 ();
 FILLCELL_X32 FILLER_214_1176 ();
 FILLCELL_X32 FILLER_214_1208 ();
 FILLCELL_X32 FILLER_214_1240 ();
 FILLCELL_X32 FILLER_214_1272 ();
 FILLCELL_X32 FILLER_214_1304 ();
 FILLCELL_X32 FILLER_214_1336 ();
 FILLCELL_X32 FILLER_214_1368 ();
 FILLCELL_X32 FILLER_214_1400 ();
 FILLCELL_X32 FILLER_214_1432 ();
 FILLCELL_X32 FILLER_214_1464 ();
 FILLCELL_X32 FILLER_214_1496 ();
 FILLCELL_X32 FILLER_214_1528 ();
 FILLCELL_X32 FILLER_214_1560 ();
 FILLCELL_X32 FILLER_214_1592 ();
 FILLCELL_X32 FILLER_214_1624 ();
 FILLCELL_X32 FILLER_214_1656 ();
 FILLCELL_X32 FILLER_214_1688 ();
 FILLCELL_X32 FILLER_214_1720 ();
 FILLCELL_X32 FILLER_214_1752 ();
 FILLCELL_X32 FILLER_214_1784 ();
 FILLCELL_X32 FILLER_214_1816 ();
 FILLCELL_X32 FILLER_214_1848 ();
 FILLCELL_X8 FILLER_214_1880 ();
 FILLCELL_X4 FILLER_214_1888 ();
 FILLCELL_X2 FILLER_214_1892 ();
 FILLCELL_X32 FILLER_214_1895 ();
 FILLCELL_X32 FILLER_214_1927 ();
 FILLCELL_X32 FILLER_214_1959 ();
 FILLCELL_X32 FILLER_214_1991 ();
 FILLCELL_X32 FILLER_214_2023 ();
 FILLCELL_X32 FILLER_214_2055 ();
 FILLCELL_X32 FILLER_214_2087 ();
 FILLCELL_X32 FILLER_214_2119 ();
 FILLCELL_X32 FILLER_214_2151 ();
 FILLCELL_X32 FILLER_214_2183 ();
 FILLCELL_X32 FILLER_214_2215 ();
 FILLCELL_X32 FILLER_214_2247 ();
 FILLCELL_X32 FILLER_214_2279 ();
 FILLCELL_X32 FILLER_214_2311 ();
 FILLCELL_X32 FILLER_214_2343 ();
 FILLCELL_X32 FILLER_214_2375 ();
 FILLCELL_X32 FILLER_214_2407 ();
 FILLCELL_X32 FILLER_214_2439 ();
 FILLCELL_X32 FILLER_214_2471 ();
 FILLCELL_X32 FILLER_214_2503 ();
 FILLCELL_X32 FILLER_214_2535 ();
 FILLCELL_X32 FILLER_214_2567 ();
 FILLCELL_X2 FILLER_214_2599 ();
 FILLCELL_X1 FILLER_214_2601 ();
 FILLCELL_X32 FILLER_215_1 ();
 FILLCELL_X32 FILLER_215_33 ();
 FILLCELL_X32 FILLER_215_65 ();
 FILLCELL_X32 FILLER_215_97 ();
 FILLCELL_X32 FILLER_215_129 ();
 FILLCELL_X32 FILLER_215_161 ();
 FILLCELL_X32 FILLER_215_193 ();
 FILLCELL_X32 FILLER_215_225 ();
 FILLCELL_X32 FILLER_215_257 ();
 FILLCELL_X32 FILLER_215_289 ();
 FILLCELL_X32 FILLER_215_321 ();
 FILLCELL_X32 FILLER_215_353 ();
 FILLCELL_X32 FILLER_215_385 ();
 FILLCELL_X32 FILLER_215_417 ();
 FILLCELL_X32 FILLER_215_449 ();
 FILLCELL_X32 FILLER_215_481 ();
 FILLCELL_X32 FILLER_215_513 ();
 FILLCELL_X32 FILLER_215_545 ();
 FILLCELL_X32 FILLER_215_577 ();
 FILLCELL_X32 FILLER_215_609 ();
 FILLCELL_X32 FILLER_215_641 ();
 FILLCELL_X32 FILLER_215_673 ();
 FILLCELL_X32 FILLER_215_705 ();
 FILLCELL_X32 FILLER_215_737 ();
 FILLCELL_X32 FILLER_215_769 ();
 FILLCELL_X32 FILLER_215_801 ();
 FILLCELL_X32 FILLER_215_833 ();
 FILLCELL_X32 FILLER_215_865 ();
 FILLCELL_X32 FILLER_215_897 ();
 FILLCELL_X32 FILLER_215_929 ();
 FILLCELL_X32 FILLER_215_961 ();
 FILLCELL_X32 FILLER_215_993 ();
 FILLCELL_X32 FILLER_215_1025 ();
 FILLCELL_X32 FILLER_215_1057 ();
 FILLCELL_X32 FILLER_215_1089 ();
 FILLCELL_X32 FILLER_215_1121 ();
 FILLCELL_X32 FILLER_215_1153 ();
 FILLCELL_X32 FILLER_215_1185 ();
 FILLCELL_X32 FILLER_215_1217 ();
 FILLCELL_X8 FILLER_215_1249 ();
 FILLCELL_X4 FILLER_215_1257 ();
 FILLCELL_X2 FILLER_215_1261 ();
 FILLCELL_X32 FILLER_215_1264 ();
 FILLCELL_X32 FILLER_215_1296 ();
 FILLCELL_X32 FILLER_215_1328 ();
 FILLCELL_X32 FILLER_215_1360 ();
 FILLCELL_X32 FILLER_215_1392 ();
 FILLCELL_X32 FILLER_215_1424 ();
 FILLCELL_X32 FILLER_215_1456 ();
 FILLCELL_X32 FILLER_215_1488 ();
 FILLCELL_X32 FILLER_215_1520 ();
 FILLCELL_X32 FILLER_215_1552 ();
 FILLCELL_X32 FILLER_215_1584 ();
 FILLCELL_X32 FILLER_215_1616 ();
 FILLCELL_X32 FILLER_215_1648 ();
 FILLCELL_X32 FILLER_215_1680 ();
 FILLCELL_X32 FILLER_215_1712 ();
 FILLCELL_X32 FILLER_215_1744 ();
 FILLCELL_X32 FILLER_215_1776 ();
 FILLCELL_X32 FILLER_215_1808 ();
 FILLCELL_X32 FILLER_215_1840 ();
 FILLCELL_X32 FILLER_215_1872 ();
 FILLCELL_X32 FILLER_215_1904 ();
 FILLCELL_X32 FILLER_215_1936 ();
 FILLCELL_X32 FILLER_215_1968 ();
 FILLCELL_X32 FILLER_215_2000 ();
 FILLCELL_X32 FILLER_215_2032 ();
 FILLCELL_X32 FILLER_215_2064 ();
 FILLCELL_X32 FILLER_215_2096 ();
 FILLCELL_X32 FILLER_215_2128 ();
 FILLCELL_X32 FILLER_215_2160 ();
 FILLCELL_X32 FILLER_215_2192 ();
 FILLCELL_X32 FILLER_215_2224 ();
 FILLCELL_X32 FILLER_215_2256 ();
 FILLCELL_X32 FILLER_215_2288 ();
 FILLCELL_X32 FILLER_215_2320 ();
 FILLCELL_X32 FILLER_215_2352 ();
 FILLCELL_X32 FILLER_215_2384 ();
 FILLCELL_X32 FILLER_215_2416 ();
 FILLCELL_X32 FILLER_215_2448 ();
 FILLCELL_X32 FILLER_215_2480 ();
 FILLCELL_X8 FILLER_215_2512 ();
 FILLCELL_X4 FILLER_215_2520 ();
 FILLCELL_X2 FILLER_215_2524 ();
 FILLCELL_X32 FILLER_215_2527 ();
 FILLCELL_X32 FILLER_215_2559 ();
 FILLCELL_X8 FILLER_215_2591 ();
 FILLCELL_X2 FILLER_215_2599 ();
 FILLCELL_X1 FILLER_215_2601 ();
 FILLCELL_X32 FILLER_216_1 ();
 FILLCELL_X32 FILLER_216_33 ();
 FILLCELL_X32 FILLER_216_65 ();
 FILLCELL_X32 FILLER_216_97 ();
 FILLCELL_X32 FILLER_216_129 ();
 FILLCELL_X32 FILLER_216_161 ();
 FILLCELL_X32 FILLER_216_193 ();
 FILLCELL_X32 FILLER_216_225 ();
 FILLCELL_X32 FILLER_216_257 ();
 FILLCELL_X32 FILLER_216_289 ();
 FILLCELL_X32 FILLER_216_321 ();
 FILLCELL_X32 FILLER_216_353 ();
 FILLCELL_X32 FILLER_216_385 ();
 FILLCELL_X32 FILLER_216_417 ();
 FILLCELL_X32 FILLER_216_449 ();
 FILLCELL_X32 FILLER_216_481 ();
 FILLCELL_X32 FILLER_216_513 ();
 FILLCELL_X32 FILLER_216_545 ();
 FILLCELL_X32 FILLER_216_577 ();
 FILLCELL_X16 FILLER_216_609 ();
 FILLCELL_X4 FILLER_216_625 ();
 FILLCELL_X2 FILLER_216_629 ();
 FILLCELL_X32 FILLER_216_632 ();
 FILLCELL_X32 FILLER_216_664 ();
 FILLCELL_X32 FILLER_216_696 ();
 FILLCELL_X32 FILLER_216_728 ();
 FILLCELL_X32 FILLER_216_760 ();
 FILLCELL_X32 FILLER_216_792 ();
 FILLCELL_X32 FILLER_216_824 ();
 FILLCELL_X32 FILLER_216_856 ();
 FILLCELL_X32 FILLER_216_888 ();
 FILLCELL_X32 FILLER_216_920 ();
 FILLCELL_X32 FILLER_216_952 ();
 FILLCELL_X32 FILLER_216_984 ();
 FILLCELL_X32 FILLER_216_1016 ();
 FILLCELL_X32 FILLER_216_1048 ();
 FILLCELL_X32 FILLER_216_1080 ();
 FILLCELL_X32 FILLER_216_1112 ();
 FILLCELL_X32 FILLER_216_1144 ();
 FILLCELL_X32 FILLER_216_1176 ();
 FILLCELL_X32 FILLER_216_1208 ();
 FILLCELL_X32 FILLER_216_1240 ();
 FILLCELL_X32 FILLER_216_1272 ();
 FILLCELL_X32 FILLER_216_1304 ();
 FILLCELL_X32 FILLER_216_1336 ();
 FILLCELL_X32 FILLER_216_1368 ();
 FILLCELL_X32 FILLER_216_1400 ();
 FILLCELL_X32 FILLER_216_1432 ();
 FILLCELL_X32 FILLER_216_1464 ();
 FILLCELL_X32 FILLER_216_1496 ();
 FILLCELL_X32 FILLER_216_1528 ();
 FILLCELL_X32 FILLER_216_1560 ();
 FILLCELL_X32 FILLER_216_1592 ();
 FILLCELL_X32 FILLER_216_1624 ();
 FILLCELL_X32 FILLER_216_1656 ();
 FILLCELL_X32 FILLER_216_1688 ();
 FILLCELL_X32 FILLER_216_1720 ();
 FILLCELL_X32 FILLER_216_1752 ();
 FILLCELL_X32 FILLER_216_1784 ();
 FILLCELL_X32 FILLER_216_1816 ();
 FILLCELL_X32 FILLER_216_1848 ();
 FILLCELL_X8 FILLER_216_1880 ();
 FILLCELL_X4 FILLER_216_1888 ();
 FILLCELL_X2 FILLER_216_1892 ();
 FILLCELL_X32 FILLER_216_1895 ();
 FILLCELL_X32 FILLER_216_1927 ();
 FILLCELL_X32 FILLER_216_1959 ();
 FILLCELL_X32 FILLER_216_1991 ();
 FILLCELL_X32 FILLER_216_2023 ();
 FILLCELL_X32 FILLER_216_2055 ();
 FILLCELL_X32 FILLER_216_2087 ();
 FILLCELL_X32 FILLER_216_2119 ();
 FILLCELL_X32 FILLER_216_2151 ();
 FILLCELL_X32 FILLER_216_2183 ();
 FILLCELL_X32 FILLER_216_2215 ();
 FILLCELL_X32 FILLER_216_2247 ();
 FILLCELL_X32 FILLER_216_2279 ();
 FILLCELL_X32 FILLER_216_2311 ();
 FILLCELL_X32 FILLER_216_2343 ();
 FILLCELL_X32 FILLER_216_2375 ();
 FILLCELL_X32 FILLER_216_2407 ();
 FILLCELL_X32 FILLER_216_2439 ();
 FILLCELL_X32 FILLER_216_2471 ();
 FILLCELL_X32 FILLER_216_2503 ();
 FILLCELL_X32 FILLER_216_2535 ();
 FILLCELL_X32 FILLER_216_2567 ();
 FILLCELL_X2 FILLER_216_2599 ();
 FILLCELL_X1 FILLER_216_2601 ();
 FILLCELL_X32 FILLER_217_1 ();
 FILLCELL_X32 FILLER_217_33 ();
 FILLCELL_X32 FILLER_217_65 ();
 FILLCELL_X32 FILLER_217_97 ();
 FILLCELL_X32 FILLER_217_129 ();
 FILLCELL_X32 FILLER_217_161 ();
 FILLCELL_X32 FILLER_217_193 ();
 FILLCELL_X32 FILLER_217_225 ();
 FILLCELL_X32 FILLER_217_257 ();
 FILLCELL_X32 FILLER_217_289 ();
 FILLCELL_X32 FILLER_217_321 ();
 FILLCELL_X32 FILLER_217_353 ();
 FILLCELL_X32 FILLER_217_385 ();
 FILLCELL_X32 FILLER_217_417 ();
 FILLCELL_X32 FILLER_217_449 ();
 FILLCELL_X32 FILLER_217_481 ();
 FILLCELL_X32 FILLER_217_513 ();
 FILLCELL_X32 FILLER_217_545 ();
 FILLCELL_X32 FILLER_217_577 ();
 FILLCELL_X32 FILLER_217_609 ();
 FILLCELL_X32 FILLER_217_641 ();
 FILLCELL_X32 FILLER_217_673 ();
 FILLCELL_X32 FILLER_217_705 ();
 FILLCELL_X32 FILLER_217_737 ();
 FILLCELL_X32 FILLER_217_769 ();
 FILLCELL_X32 FILLER_217_801 ();
 FILLCELL_X32 FILLER_217_833 ();
 FILLCELL_X32 FILLER_217_865 ();
 FILLCELL_X32 FILLER_217_897 ();
 FILLCELL_X32 FILLER_217_929 ();
 FILLCELL_X32 FILLER_217_961 ();
 FILLCELL_X32 FILLER_217_993 ();
 FILLCELL_X32 FILLER_217_1025 ();
 FILLCELL_X32 FILLER_217_1057 ();
 FILLCELL_X32 FILLER_217_1089 ();
 FILLCELL_X32 FILLER_217_1121 ();
 FILLCELL_X32 FILLER_217_1153 ();
 FILLCELL_X32 FILLER_217_1185 ();
 FILLCELL_X32 FILLER_217_1217 ();
 FILLCELL_X8 FILLER_217_1249 ();
 FILLCELL_X4 FILLER_217_1257 ();
 FILLCELL_X2 FILLER_217_1261 ();
 FILLCELL_X32 FILLER_217_1264 ();
 FILLCELL_X32 FILLER_217_1296 ();
 FILLCELL_X32 FILLER_217_1328 ();
 FILLCELL_X32 FILLER_217_1360 ();
 FILLCELL_X32 FILLER_217_1392 ();
 FILLCELL_X32 FILLER_217_1424 ();
 FILLCELL_X32 FILLER_217_1456 ();
 FILLCELL_X32 FILLER_217_1488 ();
 FILLCELL_X32 FILLER_217_1520 ();
 FILLCELL_X32 FILLER_217_1552 ();
 FILLCELL_X32 FILLER_217_1584 ();
 FILLCELL_X32 FILLER_217_1616 ();
 FILLCELL_X32 FILLER_217_1648 ();
 FILLCELL_X32 FILLER_217_1680 ();
 FILLCELL_X32 FILLER_217_1712 ();
 FILLCELL_X32 FILLER_217_1744 ();
 FILLCELL_X32 FILLER_217_1776 ();
 FILLCELL_X32 FILLER_217_1808 ();
 FILLCELL_X32 FILLER_217_1840 ();
 FILLCELL_X32 FILLER_217_1872 ();
 FILLCELL_X32 FILLER_217_1904 ();
 FILLCELL_X32 FILLER_217_1936 ();
 FILLCELL_X32 FILLER_217_1968 ();
 FILLCELL_X32 FILLER_217_2000 ();
 FILLCELL_X32 FILLER_217_2032 ();
 FILLCELL_X32 FILLER_217_2064 ();
 FILLCELL_X32 FILLER_217_2096 ();
 FILLCELL_X32 FILLER_217_2128 ();
 FILLCELL_X32 FILLER_217_2160 ();
 FILLCELL_X32 FILLER_217_2192 ();
 FILLCELL_X32 FILLER_217_2224 ();
 FILLCELL_X32 FILLER_217_2256 ();
 FILLCELL_X32 FILLER_217_2288 ();
 FILLCELL_X32 FILLER_217_2320 ();
 FILLCELL_X32 FILLER_217_2352 ();
 FILLCELL_X32 FILLER_217_2384 ();
 FILLCELL_X32 FILLER_217_2416 ();
 FILLCELL_X32 FILLER_217_2448 ();
 FILLCELL_X32 FILLER_217_2480 ();
 FILLCELL_X8 FILLER_217_2512 ();
 FILLCELL_X4 FILLER_217_2520 ();
 FILLCELL_X2 FILLER_217_2524 ();
 FILLCELL_X32 FILLER_217_2527 ();
 FILLCELL_X32 FILLER_217_2559 ();
 FILLCELL_X8 FILLER_217_2591 ();
 FILLCELL_X2 FILLER_217_2599 ();
 FILLCELL_X1 FILLER_217_2601 ();
 FILLCELL_X32 FILLER_218_1 ();
 FILLCELL_X32 FILLER_218_33 ();
 FILLCELL_X32 FILLER_218_65 ();
 FILLCELL_X32 FILLER_218_97 ();
 FILLCELL_X32 FILLER_218_129 ();
 FILLCELL_X32 FILLER_218_161 ();
 FILLCELL_X32 FILLER_218_193 ();
 FILLCELL_X32 FILLER_218_225 ();
 FILLCELL_X32 FILLER_218_257 ();
 FILLCELL_X32 FILLER_218_289 ();
 FILLCELL_X32 FILLER_218_321 ();
 FILLCELL_X32 FILLER_218_353 ();
 FILLCELL_X32 FILLER_218_385 ();
 FILLCELL_X32 FILLER_218_417 ();
 FILLCELL_X32 FILLER_218_449 ();
 FILLCELL_X32 FILLER_218_481 ();
 FILLCELL_X32 FILLER_218_513 ();
 FILLCELL_X32 FILLER_218_545 ();
 FILLCELL_X32 FILLER_218_577 ();
 FILLCELL_X16 FILLER_218_609 ();
 FILLCELL_X4 FILLER_218_625 ();
 FILLCELL_X2 FILLER_218_629 ();
 FILLCELL_X32 FILLER_218_632 ();
 FILLCELL_X32 FILLER_218_664 ();
 FILLCELL_X32 FILLER_218_696 ();
 FILLCELL_X32 FILLER_218_728 ();
 FILLCELL_X32 FILLER_218_760 ();
 FILLCELL_X32 FILLER_218_792 ();
 FILLCELL_X32 FILLER_218_824 ();
 FILLCELL_X32 FILLER_218_856 ();
 FILLCELL_X32 FILLER_218_888 ();
 FILLCELL_X32 FILLER_218_920 ();
 FILLCELL_X32 FILLER_218_952 ();
 FILLCELL_X32 FILLER_218_984 ();
 FILLCELL_X32 FILLER_218_1016 ();
 FILLCELL_X32 FILLER_218_1048 ();
 FILLCELL_X32 FILLER_218_1080 ();
 FILLCELL_X32 FILLER_218_1112 ();
 FILLCELL_X32 FILLER_218_1144 ();
 FILLCELL_X32 FILLER_218_1176 ();
 FILLCELL_X32 FILLER_218_1208 ();
 FILLCELL_X32 FILLER_218_1240 ();
 FILLCELL_X32 FILLER_218_1272 ();
 FILLCELL_X32 FILLER_218_1304 ();
 FILLCELL_X32 FILLER_218_1336 ();
 FILLCELL_X32 FILLER_218_1368 ();
 FILLCELL_X32 FILLER_218_1400 ();
 FILLCELL_X32 FILLER_218_1432 ();
 FILLCELL_X32 FILLER_218_1464 ();
 FILLCELL_X32 FILLER_218_1496 ();
 FILLCELL_X32 FILLER_218_1528 ();
 FILLCELL_X32 FILLER_218_1560 ();
 FILLCELL_X32 FILLER_218_1592 ();
 FILLCELL_X32 FILLER_218_1624 ();
 FILLCELL_X32 FILLER_218_1656 ();
 FILLCELL_X32 FILLER_218_1688 ();
 FILLCELL_X32 FILLER_218_1720 ();
 FILLCELL_X32 FILLER_218_1752 ();
 FILLCELL_X32 FILLER_218_1784 ();
 FILLCELL_X32 FILLER_218_1816 ();
 FILLCELL_X32 FILLER_218_1848 ();
 FILLCELL_X8 FILLER_218_1880 ();
 FILLCELL_X4 FILLER_218_1888 ();
 FILLCELL_X2 FILLER_218_1892 ();
 FILLCELL_X32 FILLER_218_1895 ();
 FILLCELL_X32 FILLER_218_1927 ();
 FILLCELL_X32 FILLER_218_1959 ();
 FILLCELL_X32 FILLER_218_1991 ();
 FILLCELL_X32 FILLER_218_2023 ();
 FILLCELL_X32 FILLER_218_2055 ();
 FILLCELL_X32 FILLER_218_2087 ();
 FILLCELL_X32 FILLER_218_2119 ();
 FILLCELL_X32 FILLER_218_2151 ();
 FILLCELL_X32 FILLER_218_2183 ();
 FILLCELL_X32 FILLER_218_2215 ();
 FILLCELL_X32 FILLER_218_2247 ();
 FILLCELL_X32 FILLER_218_2279 ();
 FILLCELL_X32 FILLER_218_2311 ();
 FILLCELL_X32 FILLER_218_2343 ();
 FILLCELL_X32 FILLER_218_2375 ();
 FILLCELL_X32 FILLER_218_2407 ();
 FILLCELL_X32 FILLER_218_2439 ();
 FILLCELL_X32 FILLER_218_2471 ();
 FILLCELL_X32 FILLER_218_2503 ();
 FILLCELL_X32 FILLER_218_2535 ();
 FILLCELL_X32 FILLER_218_2567 ();
 FILLCELL_X2 FILLER_218_2599 ();
 FILLCELL_X1 FILLER_218_2601 ();
 FILLCELL_X32 FILLER_219_1 ();
 FILLCELL_X32 FILLER_219_33 ();
 FILLCELL_X32 FILLER_219_65 ();
 FILLCELL_X32 FILLER_219_97 ();
 FILLCELL_X32 FILLER_219_129 ();
 FILLCELL_X32 FILLER_219_161 ();
 FILLCELL_X32 FILLER_219_193 ();
 FILLCELL_X32 FILLER_219_225 ();
 FILLCELL_X32 FILLER_219_257 ();
 FILLCELL_X32 FILLER_219_289 ();
 FILLCELL_X32 FILLER_219_321 ();
 FILLCELL_X32 FILLER_219_353 ();
 FILLCELL_X32 FILLER_219_385 ();
 FILLCELL_X32 FILLER_219_417 ();
 FILLCELL_X32 FILLER_219_449 ();
 FILLCELL_X32 FILLER_219_481 ();
 FILLCELL_X32 FILLER_219_513 ();
 FILLCELL_X32 FILLER_219_545 ();
 FILLCELL_X32 FILLER_219_577 ();
 FILLCELL_X32 FILLER_219_609 ();
 FILLCELL_X32 FILLER_219_641 ();
 FILLCELL_X32 FILLER_219_673 ();
 FILLCELL_X32 FILLER_219_705 ();
 FILLCELL_X32 FILLER_219_737 ();
 FILLCELL_X32 FILLER_219_769 ();
 FILLCELL_X32 FILLER_219_801 ();
 FILLCELL_X32 FILLER_219_833 ();
 FILLCELL_X32 FILLER_219_865 ();
 FILLCELL_X32 FILLER_219_897 ();
 FILLCELL_X32 FILLER_219_929 ();
 FILLCELL_X32 FILLER_219_961 ();
 FILLCELL_X32 FILLER_219_993 ();
 FILLCELL_X32 FILLER_219_1025 ();
 FILLCELL_X32 FILLER_219_1057 ();
 FILLCELL_X32 FILLER_219_1089 ();
 FILLCELL_X32 FILLER_219_1121 ();
 FILLCELL_X32 FILLER_219_1153 ();
 FILLCELL_X32 FILLER_219_1185 ();
 FILLCELL_X32 FILLER_219_1217 ();
 FILLCELL_X8 FILLER_219_1249 ();
 FILLCELL_X4 FILLER_219_1257 ();
 FILLCELL_X2 FILLER_219_1261 ();
 FILLCELL_X32 FILLER_219_1264 ();
 FILLCELL_X32 FILLER_219_1296 ();
 FILLCELL_X32 FILLER_219_1328 ();
 FILLCELL_X32 FILLER_219_1360 ();
 FILLCELL_X32 FILLER_219_1392 ();
 FILLCELL_X32 FILLER_219_1424 ();
 FILLCELL_X32 FILLER_219_1456 ();
 FILLCELL_X32 FILLER_219_1488 ();
 FILLCELL_X32 FILLER_219_1520 ();
 FILLCELL_X32 FILLER_219_1552 ();
 FILLCELL_X32 FILLER_219_1584 ();
 FILLCELL_X32 FILLER_219_1616 ();
 FILLCELL_X32 FILLER_219_1648 ();
 FILLCELL_X32 FILLER_219_1680 ();
 FILLCELL_X32 FILLER_219_1712 ();
 FILLCELL_X32 FILLER_219_1744 ();
 FILLCELL_X32 FILLER_219_1776 ();
 FILLCELL_X32 FILLER_219_1808 ();
 FILLCELL_X32 FILLER_219_1840 ();
 FILLCELL_X32 FILLER_219_1872 ();
 FILLCELL_X32 FILLER_219_1904 ();
 FILLCELL_X32 FILLER_219_1936 ();
 FILLCELL_X32 FILLER_219_1968 ();
 FILLCELL_X32 FILLER_219_2000 ();
 FILLCELL_X32 FILLER_219_2032 ();
 FILLCELL_X32 FILLER_219_2064 ();
 FILLCELL_X32 FILLER_219_2096 ();
 FILLCELL_X32 FILLER_219_2128 ();
 FILLCELL_X32 FILLER_219_2160 ();
 FILLCELL_X32 FILLER_219_2192 ();
 FILLCELL_X32 FILLER_219_2224 ();
 FILLCELL_X32 FILLER_219_2256 ();
 FILLCELL_X32 FILLER_219_2288 ();
 FILLCELL_X32 FILLER_219_2320 ();
 FILLCELL_X32 FILLER_219_2352 ();
 FILLCELL_X32 FILLER_219_2384 ();
 FILLCELL_X32 FILLER_219_2416 ();
 FILLCELL_X32 FILLER_219_2448 ();
 FILLCELL_X32 FILLER_219_2480 ();
 FILLCELL_X8 FILLER_219_2512 ();
 FILLCELL_X4 FILLER_219_2520 ();
 FILLCELL_X2 FILLER_219_2524 ();
 FILLCELL_X32 FILLER_219_2527 ();
 FILLCELL_X32 FILLER_219_2559 ();
 FILLCELL_X8 FILLER_219_2591 ();
 FILLCELL_X2 FILLER_219_2599 ();
 FILLCELL_X1 FILLER_219_2601 ();
 FILLCELL_X32 FILLER_220_1 ();
 FILLCELL_X32 FILLER_220_33 ();
 FILLCELL_X32 FILLER_220_65 ();
 FILLCELL_X32 FILLER_220_97 ();
 FILLCELL_X32 FILLER_220_129 ();
 FILLCELL_X32 FILLER_220_161 ();
 FILLCELL_X32 FILLER_220_193 ();
 FILLCELL_X32 FILLER_220_225 ();
 FILLCELL_X32 FILLER_220_257 ();
 FILLCELL_X32 FILLER_220_289 ();
 FILLCELL_X32 FILLER_220_321 ();
 FILLCELL_X32 FILLER_220_353 ();
 FILLCELL_X32 FILLER_220_385 ();
 FILLCELL_X32 FILLER_220_417 ();
 FILLCELL_X32 FILLER_220_449 ();
 FILLCELL_X32 FILLER_220_481 ();
 FILLCELL_X32 FILLER_220_513 ();
 FILLCELL_X32 FILLER_220_545 ();
 FILLCELL_X32 FILLER_220_577 ();
 FILLCELL_X16 FILLER_220_609 ();
 FILLCELL_X4 FILLER_220_625 ();
 FILLCELL_X2 FILLER_220_629 ();
 FILLCELL_X32 FILLER_220_632 ();
 FILLCELL_X32 FILLER_220_664 ();
 FILLCELL_X32 FILLER_220_696 ();
 FILLCELL_X32 FILLER_220_728 ();
 FILLCELL_X32 FILLER_220_760 ();
 FILLCELL_X32 FILLER_220_792 ();
 FILLCELL_X32 FILLER_220_824 ();
 FILLCELL_X32 FILLER_220_856 ();
 FILLCELL_X32 FILLER_220_888 ();
 FILLCELL_X32 FILLER_220_920 ();
 FILLCELL_X32 FILLER_220_952 ();
 FILLCELL_X32 FILLER_220_984 ();
 FILLCELL_X32 FILLER_220_1016 ();
 FILLCELL_X32 FILLER_220_1048 ();
 FILLCELL_X32 FILLER_220_1080 ();
 FILLCELL_X32 FILLER_220_1112 ();
 FILLCELL_X32 FILLER_220_1144 ();
 FILLCELL_X32 FILLER_220_1176 ();
 FILLCELL_X32 FILLER_220_1208 ();
 FILLCELL_X32 FILLER_220_1240 ();
 FILLCELL_X32 FILLER_220_1272 ();
 FILLCELL_X32 FILLER_220_1304 ();
 FILLCELL_X32 FILLER_220_1336 ();
 FILLCELL_X32 FILLER_220_1368 ();
 FILLCELL_X32 FILLER_220_1400 ();
 FILLCELL_X32 FILLER_220_1432 ();
 FILLCELL_X32 FILLER_220_1464 ();
 FILLCELL_X32 FILLER_220_1496 ();
 FILLCELL_X32 FILLER_220_1528 ();
 FILLCELL_X32 FILLER_220_1560 ();
 FILLCELL_X32 FILLER_220_1592 ();
 FILLCELL_X32 FILLER_220_1624 ();
 FILLCELL_X32 FILLER_220_1656 ();
 FILLCELL_X32 FILLER_220_1688 ();
 FILLCELL_X32 FILLER_220_1720 ();
 FILLCELL_X32 FILLER_220_1752 ();
 FILLCELL_X32 FILLER_220_1784 ();
 FILLCELL_X32 FILLER_220_1816 ();
 FILLCELL_X32 FILLER_220_1848 ();
 FILLCELL_X8 FILLER_220_1880 ();
 FILLCELL_X4 FILLER_220_1888 ();
 FILLCELL_X2 FILLER_220_1892 ();
 FILLCELL_X32 FILLER_220_1895 ();
 FILLCELL_X32 FILLER_220_1927 ();
 FILLCELL_X32 FILLER_220_1959 ();
 FILLCELL_X32 FILLER_220_1991 ();
 FILLCELL_X32 FILLER_220_2023 ();
 FILLCELL_X32 FILLER_220_2055 ();
 FILLCELL_X32 FILLER_220_2087 ();
 FILLCELL_X32 FILLER_220_2119 ();
 FILLCELL_X32 FILLER_220_2151 ();
 FILLCELL_X32 FILLER_220_2183 ();
 FILLCELL_X32 FILLER_220_2215 ();
 FILLCELL_X32 FILLER_220_2247 ();
 FILLCELL_X32 FILLER_220_2279 ();
 FILLCELL_X32 FILLER_220_2311 ();
 FILLCELL_X32 FILLER_220_2343 ();
 FILLCELL_X32 FILLER_220_2375 ();
 FILLCELL_X32 FILLER_220_2407 ();
 FILLCELL_X32 FILLER_220_2439 ();
 FILLCELL_X32 FILLER_220_2471 ();
 FILLCELL_X32 FILLER_220_2503 ();
 FILLCELL_X32 FILLER_220_2535 ();
 FILLCELL_X32 FILLER_220_2567 ();
 FILLCELL_X2 FILLER_220_2599 ();
 FILLCELL_X1 FILLER_220_2601 ();
 FILLCELL_X32 FILLER_221_1 ();
 FILLCELL_X32 FILLER_221_33 ();
 FILLCELL_X32 FILLER_221_65 ();
 FILLCELL_X32 FILLER_221_97 ();
 FILLCELL_X32 FILLER_221_129 ();
 FILLCELL_X32 FILLER_221_161 ();
 FILLCELL_X32 FILLER_221_193 ();
 FILLCELL_X32 FILLER_221_225 ();
 FILLCELL_X32 FILLER_221_257 ();
 FILLCELL_X32 FILLER_221_289 ();
 FILLCELL_X32 FILLER_221_321 ();
 FILLCELL_X32 FILLER_221_353 ();
 FILLCELL_X32 FILLER_221_385 ();
 FILLCELL_X32 FILLER_221_417 ();
 FILLCELL_X32 FILLER_221_449 ();
 FILLCELL_X32 FILLER_221_481 ();
 FILLCELL_X32 FILLER_221_513 ();
 FILLCELL_X32 FILLER_221_545 ();
 FILLCELL_X32 FILLER_221_577 ();
 FILLCELL_X32 FILLER_221_609 ();
 FILLCELL_X32 FILLER_221_641 ();
 FILLCELL_X32 FILLER_221_673 ();
 FILLCELL_X32 FILLER_221_705 ();
 FILLCELL_X32 FILLER_221_737 ();
 FILLCELL_X32 FILLER_221_769 ();
 FILLCELL_X32 FILLER_221_801 ();
 FILLCELL_X32 FILLER_221_833 ();
 FILLCELL_X32 FILLER_221_865 ();
 FILLCELL_X32 FILLER_221_897 ();
 FILLCELL_X32 FILLER_221_929 ();
 FILLCELL_X32 FILLER_221_961 ();
 FILLCELL_X32 FILLER_221_993 ();
 FILLCELL_X32 FILLER_221_1025 ();
 FILLCELL_X32 FILLER_221_1057 ();
 FILLCELL_X32 FILLER_221_1089 ();
 FILLCELL_X32 FILLER_221_1121 ();
 FILLCELL_X32 FILLER_221_1153 ();
 FILLCELL_X32 FILLER_221_1185 ();
 FILLCELL_X32 FILLER_221_1217 ();
 FILLCELL_X8 FILLER_221_1249 ();
 FILLCELL_X4 FILLER_221_1257 ();
 FILLCELL_X2 FILLER_221_1261 ();
 FILLCELL_X32 FILLER_221_1264 ();
 FILLCELL_X32 FILLER_221_1296 ();
 FILLCELL_X32 FILLER_221_1328 ();
 FILLCELL_X32 FILLER_221_1360 ();
 FILLCELL_X32 FILLER_221_1392 ();
 FILLCELL_X32 FILLER_221_1424 ();
 FILLCELL_X32 FILLER_221_1456 ();
 FILLCELL_X32 FILLER_221_1488 ();
 FILLCELL_X32 FILLER_221_1520 ();
 FILLCELL_X32 FILLER_221_1552 ();
 FILLCELL_X32 FILLER_221_1584 ();
 FILLCELL_X32 FILLER_221_1616 ();
 FILLCELL_X32 FILLER_221_1648 ();
 FILLCELL_X32 FILLER_221_1680 ();
 FILLCELL_X32 FILLER_221_1712 ();
 FILLCELL_X32 FILLER_221_1744 ();
 FILLCELL_X32 FILLER_221_1776 ();
 FILLCELL_X32 FILLER_221_1808 ();
 FILLCELL_X32 FILLER_221_1840 ();
 FILLCELL_X32 FILLER_221_1872 ();
 FILLCELL_X32 FILLER_221_1904 ();
 FILLCELL_X32 FILLER_221_1936 ();
 FILLCELL_X32 FILLER_221_1968 ();
 FILLCELL_X32 FILLER_221_2000 ();
 FILLCELL_X32 FILLER_221_2032 ();
 FILLCELL_X32 FILLER_221_2064 ();
 FILLCELL_X32 FILLER_221_2096 ();
 FILLCELL_X32 FILLER_221_2128 ();
 FILLCELL_X32 FILLER_221_2160 ();
 FILLCELL_X32 FILLER_221_2192 ();
 FILLCELL_X32 FILLER_221_2224 ();
 FILLCELL_X32 FILLER_221_2256 ();
 FILLCELL_X32 FILLER_221_2288 ();
 FILLCELL_X32 FILLER_221_2320 ();
 FILLCELL_X32 FILLER_221_2352 ();
 FILLCELL_X32 FILLER_221_2384 ();
 FILLCELL_X32 FILLER_221_2416 ();
 FILLCELL_X32 FILLER_221_2448 ();
 FILLCELL_X32 FILLER_221_2480 ();
 FILLCELL_X8 FILLER_221_2512 ();
 FILLCELL_X4 FILLER_221_2520 ();
 FILLCELL_X2 FILLER_221_2524 ();
 FILLCELL_X32 FILLER_221_2527 ();
 FILLCELL_X32 FILLER_221_2559 ();
 FILLCELL_X8 FILLER_221_2591 ();
 FILLCELL_X2 FILLER_221_2599 ();
 FILLCELL_X1 FILLER_221_2601 ();
 FILLCELL_X32 FILLER_222_1 ();
 FILLCELL_X32 FILLER_222_33 ();
 FILLCELL_X32 FILLER_222_65 ();
 FILLCELL_X32 FILLER_222_97 ();
 FILLCELL_X32 FILLER_222_129 ();
 FILLCELL_X32 FILLER_222_161 ();
 FILLCELL_X32 FILLER_222_193 ();
 FILLCELL_X32 FILLER_222_225 ();
 FILLCELL_X32 FILLER_222_257 ();
 FILLCELL_X32 FILLER_222_289 ();
 FILLCELL_X32 FILLER_222_321 ();
 FILLCELL_X32 FILLER_222_353 ();
 FILLCELL_X32 FILLER_222_385 ();
 FILLCELL_X32 FILLER_222_417 ();
 FILLCELL_X32 FILLER_222_449 ();
 FILLCELL_X32 FILLER_222_481 ();
 FILLCELL_X32 FILLER_222_513 ();
 FILLCELL_X32 FILLER_222_545 ();
 FILLCELL_X32 FILLER_222_577 ();
 FILLCELL_X16 FILLER_222_609 ();
 FILLCELL_X4 FILLER_222_625 ();
 FILLCELL_X2 FILLER_222_629 ();
 FILLCELL_X32 FILLER_222_632 ();
 FILLCELL_X32 FILLER_222_664 ();
 FILLCELL_X32 FILLER_222_696 ();
 FILLCELL_X32 FILLER_222_728 ();
 FILLCELL_X32 FILLER_222_760 ();
 FILLCELL_X32 FILLER_222_792 ();
 FILLCELL_X32 FILLER_222_824 ();
 FILLCELL_X32 FILLER_222_856 ();
 FILLCELL_X32 FILLER_222_888 ();
 FILLCELL_X32 FILLER_222_920 ();
 FILLCELL_X32 FILLER_222_952 ();
 FILLCELL_X32 FILLER_222_984 ();
 FILLCELL_X32 FILLER_222_1016 ();
 FILLCELL_X32 FILLER_222_1048 ();
 FILLCELL_X32 FILLER_222_1080 ();
 FILLCELL_X32 FILLER_222_1112 ();
 FILLCELL_X32 FILLER_222_1144 ();
 FILLCELL_X32 FILLER_222_1176 ();
 FILLCELL_X32 FILLER_222_1208 ();
 FILLCELL_X32 FILLER_222_1240 ();
 FILLCELL_X32 FILLER_222_1272 ();
 FILLCELL_X32 FILLER_222_1304 ();
 FILLCELL_X32 FILLER_222_1336 ();
 FILLCELL_X32 FILLER_222_1368 ();
 FILLCELL_X32 FILLER_222_1400 ();
 FILLCELL_X32 FILLER_222_1432 ();
 FILLCELL_X32 FILLER_222_1464 ();
 FILLCELL_X32 FILLER_222_1496 ();
 FILLCELL_X32 FILLER_222_1528 ();
 FILLCELL_X32 FILLER_222_1560 ();
 FILLCELL_X32 FILLER_222_1592 ();
 FILLCELL_X32 FILLER_222_1624 ();
 FILLCELL_X32 FILLER_222_1656 ();
 FILLCELL_X32 FILLER_222_1688 ();
 FILLCELL_X32 FILLER_222_1720 ();
 FILLCELL_X32 FILLER_222_1752 ();
 FILLCELL_X32 FILLER_222_1784 ();
 FILLCELL_X32 FILLER_222_1816 ();
 FILLCELL_X32 FILLER_222_1848 ();
 FILLCELL_X8 FILLER_222_1880 ();
 FILLCELL_X4 FILLER_222_1888 ();
 FILLCELL_X2 FILLER_222_1892 ();
 FILLCELL_X32 FILLER_222_1895 ();
 FILLCELL_X32 FILLER_222_1927 ();
 FILLCELL_X32 FILLER_222_1959 ();
 FILLCELL_X32 FILLER_222_1991 ();
 FILLCELL_X32 FILLER_222_2023 ();
 FILLCELL_X32 FILLER_222_2055 ();
 FILLCELL_X32 FILLER_222_2087 ();
 FILLCELL_X32 FILLER_222_2119 ();
 FILLCELL_X32 FILLER_222_2151 ();
 FILLCELL_X32 FILLER_222_2183 ();
 FILLCELL_X32 FILLER_222_2215 ();
 FILLCELL_X32 FILLER_222_2247 ();
 FILLCELL_X32 FILLER_222_2279 ();
 FILLCELL_X32 FILLER_222_2311 ();
 FILLCELL_X32 FILLER_222_2343 ();
 FILLCELL_X32 FILLER_222_2375 ();
 FILLCELL_X32 FILLER_222_2407 ();
 FILLCELL_X32 FILLER_222_2439 ();
 FILLCELL_X32 FILLER_222_2471 ();
 FILLCELL_X32 FILLER_222_2503 ();
 FILLCELL_X32 FILLER_222_2535 ();
 FILLCELL_X32 FILLER_222_2567 ();
 FILLCELL_X2 FILLER_222_2599 ();
 FILLCELL_X1 FILLER_222_2601 ();
 FILLCELL_X32 FILLER_223_1 ();
 FILLCELL_X32 FILLER_223_33 ();
 FILLCELL_X32 FILLER_223_65 ();
 FILLCELL_X32 FILLER_223_97 ();
 FILLCELL_X32 FILLER_223_129 ();
 FILLCELL_X32 FILLER_223_161 ();
 FILLCELL_X32 FILLER_223_193 ();
 FILLCELL_X32 FILLER_223_225 ();
 FILLCELL_X32 FILLER_223_257 ();
 FILLCELL_X32 FILLER_223_289 ();
 FILLCELL_X32 FILLER_223_321 ();
 FILLCELL_X32 FILLER_223_353 ();
 FILLCELL_X32 FILLER_223_385 ();
 FILLCELL_X32 FILLER_223_417 ();
 FILLCELL_X32 FILLER_223_449 ();
 FILLCELL_X32 FILLER_223_481 ();
 FILLCELL_X32 FILLER_223_513 ();
 FILLCELL_X32 FILLER_223_545 ();
 FILLCELL_X32 FILLER_223_577 ();
 FILLCELL_X32 FILLER_223_609 ();
 FILLCELL_X32 FILLER_223_641 ();
 FILLCELL_X32 FILLER_223_673 ();
 FILLCELL_X32 FILLER_223_705 ();
 FILLCELL_X32 FILLER_223_737 ();
 FILLCELL_X32 FILLER_223_769 ();
 FILLCELL_X32 FILLER_223_801 ();
 FILLCELL_X32 FILLER_223_833 ();
 FILLCELL_X32 FILLER_223_865 ();
 FILLCELL_X32 FILLER_223_897 ();
 FILLCELL_X32 FILLER_223_929 ();
 FILLCELL_X32 FILLER_223_961 ();
 FILLCELL_X32 FILLER_223_993 ();
 FILLCELL_X32 FILLER_223_1025 ();
 FILLCELL_X32 FILLER_223_1057 ();
 FILLCELL_X32 FILLER_223_1089 ();
 FILLCELL_X32 FILLER_223_1121 ();
 FILLCELL_X32 FILLER_223_1153 ();
 FILLCELL_X32 FILLER_223_1185 ();
 FILLCELL_X32 FILLER_223_1217 ();
 FILLCELL_X8 FILLER_223_1249 ();
 FILLCELL_X4 FILLER_223_1257 ();
 FILLCELL_X2 FILLER_223_1261 ();
 FILLCELL_X32 FILLER_223_1264 ();
 FILLCELL_X32 FILLER_223_1296 ();
 FILLCELL_X32 FILLER_223_1328 ();
 FILLCELL_X32 FILLER_223_1360 ();
 FILLCELL_X32 FILLER_223_1392 ();
 FILLCELL_X32 FILLER_223_1424 ();
 FILLCELL_X32 FILLER_223_1456 ();
 FILLCELL_X32 FILLER_223_1488 ();
 FILLCELL_X32 FILLER_223_1520 ();
 FILLCELL_X32 FILLER_223_1552 ();
 FILLCELL_X32 FILLER_223_1584 ();
 FILLCELL_X32 FILLER_223_1616 ();
 FILLCELL_X32 FILLER_223_1648 ();
 FILLCELL_X32 FILLER_223_1680 ();
 FILLCELL_X32 FILLER_223_1712 ();
 FILLCELL_X32 FILLER_223_1744 ();
 FILLCELL_X32 FILLER_223_1776 ();
 FILLCELL_X32 FILLER_223_1808 ();
 FILLCELL_X32 FILLER_223_1840 ();
 FILLCELL_X32 FILLER_223_1872 ();
 FILLCELL_X32 FILLER_223_1904 ();
 FILLCELL_X32 FILLER_223_1936 ();
 FILLCELL_X32 FILLER_223_1968 ();
 FILLCELL_X32 FILLER_223_2000 ();
 FILLCELL_X32 FILLER_223_2032 ();
 FILLCELL_X32 FILLER_223_2064 ();
 FILLCELL_X32 FILLER_223_2096 ();
 FILLCELL_X32 FILLER_223_2128 ();
 FILLCELL_X32 FILLER_223_2160 ();
 FILLCELL_X32 FILLER_223_2192 ();
 FILLCELL_X32 FILLER_223_2224 ();
 FILLCELL_X32 FILLER_223_2256 ();
 FILLCELL_X32 FILLER_223_2288 ();
 FILLCELL_X32 FILLER_223_2320 ();
 FILLCELL_X32 FILLER_223_2352 ();
 FILLCELL_X32 FILLER_223_2384 ();
 FILLCELL_X32 FILLER_223_2416 ();
 FILLCELL_X32 FILLER_223_2448 ();
 FILLCELL_X32 FILLER_223_2480 ();
 FILLCELL_X8 FILLER_223_2512 ();
 FILLCELL_X4 FILLER_223_2520 ();
 FILLCELL_X2 FILLER_223_2524 ();
 FILLCELL_X32 FILLER_223_2527 ();
 FILLCELL_X32 FILLER_223_2559 ();
 FILLCELL_X8 FILLER_223_2591 ();
 FILLCELL_X2 FILLER_223_2599 ();
 FILLCELL_X1 FILLER_223_2601 ();
 FILLCELL_X32 FILLER_224_1 ();
 FILLCELL_X32 FILLER_224_33 ();
 FILLCELL_X32 FILLER_224_65 ();
 FILLCELL_X32 FILLER_224_97 ();
 FILLCELL_X32 FILLER_224_129 ();
 FILLCELL_X32 FILLER_224_161 ();
 FILLCELL_X32 FILLER_224_193 ();
 FILLCELL_X32 FILLER_224_225 ();
 FILLCELL_X32 FILLER_224_257 ();
 FILLCELL_X32 FILLER_224_289 ();
 FILLCELL_X32 FILLER_224_321 ();
 FILLCELL_X32 FILLER_224_353 ();
 FILLCELL_X32 FILLER_224_385 ();
 FILLCELL_X32 FILLER_224_417 ();
 FILLCELL_X32 FILLER_224_449 ();
 FILLCELL_X32 FILLER_224_481 ();
 FILLCELL_X32 FILLER_224_513 ();
 FILLCELL_X32 FILLER_224_545 ();
 FILLCELL_X32 FILLER_224_577 ();
 FILLCELL_X16 FILLER_224_609 ();
 FILLCELL_X4 FILLER_224_625 ();
 FILLCELL_X2 FILLER_224_629 ();
 FILLCELL_X32 FILLER_224_632 ();
 FILLCELL_X32 FILLER_224_664 ();
 FILLCELL_X32 FILLER_224_696 ();
 FILLCELL_X32 FILLER_224_728 ();
 FILLCELL_X32 FILLER_224_760 ();
 FILLCELL_X32 FILLER_224_792 ();
 FILLCELL_X32 FILLER_224_824 ();
 FILLCELL_X32 FILLER_224_856 ();
 FILLCELL_X32 FILLER_224_888 ();
 FILLCELL_X32 FILLER_224_920 ();
 FILLCELL_X32 FILLER_224_952 ();
 FILLCELL_X32 FILLER_224_984 ();
 FILLCELL_X32 FILLER_224_1016 ();
 FILLCELL_X32 FILLER_224_1048 ();
 FILLCELL_X32 FILLER_224_1080 ();
 FILLCELL_X32 FILLER_224_1112 ();
 FILLCELL_X32 FILLER_224_1144 ();
 FILLCELL_X32 FILLER_224_1176 ();
 FILLCELL_X32 FILLER_224_1208 ();
 FILLCELL_X32 FILLER_224_1240 ();
 FILLCELL_X32 FILLER_224_1272 ();
 FILLCELL_X32 FILLER_224_1304 ();
 FILLCELL_X32 FILLER_224_1336 ();
 FILLCELL_X32 FILLER_224_1368 ();
 FILLCELL_X32 FILLER_224_1400 ();
 FILLCELL_X32 FILLER_224_1432 ();
 FILLCELL_X32 FILLER_224_1464 ();
 FILLCELL_X32 FILLER_224_1496 ();
 FILLCELL_X32 FILLER_224_1528 ();
 FILLCELL_X32 FILLER_224_1560 ();
 FILLCELL_X32 FILLER_224_1592 ();
 FILLCELL_X32 FILLER_224_1624 ();
 FILLCELL_X32 FILLER_224_1656 ();
 FILLCELL_X32 FILLER_224_1688 ();
 FILLCELL_X32 FILLER_224_1720 ();
 FILLCELL_X32 FILLER_224_1752 ();
 FILLCELL_X32 FILLER_224_1784 ();
 FILLCELL_X32 FILLER_224_1816 ();
 FILLCELL_X32 FILLER_224_1848 ();
 FILLCELL_X8 FILLER_224_1880 ();
 FILLCELL_X4 FILLER_224_1888 ();
 FILLCELL_X2 FILLER_224_1892 ();
 FILLCELL_X32 FILLER_224_1895 ();
 FILLCELL_X32 FILLER_224_1927 ();
 FILLCELL_X32 FILLER_224_1959 ();
 FILLCELL_X32 FILLER_224_1991 ();
 FILLCELL_X32 FILLER_224_2023 ();
 FILLCELL_X32 FILLER_224_2055 ();
 FILLCELL_X32 FILLER_224_2087 ();
 FILLCELL_X32 FILLER_224_2119 ();
 FILLCELL_X32 FILLER_224_2151 ();
 FILLCELL_X32 FILLER_224_2183 ();
 FILLCELL_X32 FILLER_224_2215 ();
 FILLCELL_X32 FILLER_224_2247 ();
 FILLCELL_X32 FILLER_224_2279 ();
 FILLCELL_X32 FILLER_224_2311 ();
 FILLCELL_X32 FILLER_224_2343 ();
 FILLCELL_X32 FILLER_224_2375 ();
 FILLCELL_X32 FILLER_224_2407 ();
 FILLCELL_X32 FILLER_224_2439 ();
 FILLCELL_X32 FILLER_224_2471 ();
 FILLCELL_X32 FILLER_224_2503 ();
 FILLCELL_X32 FILLER_224_2535 ();
 FILLCELL_X32 FILLER_224_2567 ();
 FILLCELL_X2 FILLER_224_2599 ();
 FILLCELL_X1 FILLER_224_2601 ();
 FILLCELL_X32 FILLER_225_1 ();
 FILLCELL_X32 FILLER_225_33 ();
 FILLCELL_X32 FILLER_225_65 ();
 FILLCELL_X32 FILLER_225_97 ();
 FILLCELL_X32 FILLER_225_129 ();
 FILLCELL_X32 FILLER_225_161 ();
 FILLCELL_X32 FILLER_225_193 ();
 FILLCELL_X32 FILLER_225_225 ();
 FILLCELL_X32 FILLER_225_257 ();
 FILLCELL_X32 FILLER_225_289 ();
 FILLCELL_X32 FILLER_225_321 ();
 FILLCELL_X32 FILLER_225_353 ();
 FILLCELL_X32 FILLER_225_385 ();
 FILLCELL_X32 FILLER_225_417 ();
 FILLCELL_X32 FILLER_225_449 ();
 FILLCELL_X32 FILLER_225_481 ();
 FILLCELL_X32 FILLER_225_513 ();
 FILLCELL_X32 FILLER_225_545 ();
 FILLCELL_X32 FILLER_225_577 ();
 FILLCELL_X32 FILLER_225_609 ();
 FILLCELL_X32 FILLER_225_641 ();
 FILLCELL_X32 FILLER_225_673 ();
 FILLCELL_X32 FILLER_225_705 ();
 FILLCELL_X32 FILLER_225_737 ();
 FILLCELL_X32 FILLER_225_769 ();
 FILLCELL_X32 FILLER_225_801 ();
 FILLCELL_X32 FILLER_225_833 ();
 FILLCELL_X32 FILLER_225_865 ();
 FILLCELL_X32 FILLER_225_897 ();
 FILLCELL_X32 FILLER_225_929 ();
 FILLCELL_X32 FILLER_225_961 ();
 FILLCELL_X32 FILLER_225_993 ();
 FILLCELL_X32 FILLER_225_1025 ();
 FILLCELL_X32 FILLER_225_1057 ();
 FILLCELL_X32 FILLER_225_1089 ();
 FILLCELL_X32 FILLER_225_1121 ();
 FILLCELL_X32 FILLER_225_1153 ();
 FILLCELL_X32 FILLER_225_1185 ();
 FILLCELL_X32 FILLER_225_1217 ();
 FILLCELL_X8 FILLER_225_1249 ();
 FILLCELL_X4 FILLER_225_1257 ();
 FILLCELL_X2 FILLER_225_1261 ();
 FILLCELL_X32 FILLER_225_1264 ();
 FILLCELL_X32 FILLER_225_1296 ();
 FILLCELL_X32 FILLER_225_1328 ();
 FILLCELL_X32 FILLER_225_1360 ();
 FILLCELL_X32 FILLER_225_1392 ();
 FILLCELL_X32 FILLER_225_1424 ();
 FILLCELL_X32 FILLER_225_1456 ();
 FILLCELL_X32 FILLER_225_1488 ();
 FILLCELL_X32 FILLER_225_1520 ();
 FILLCELL_X32 FILLER_225_1552 ();
 FILLCELL_X32 FILLER_225_1584 ();
 FILLCELL_X32 FILLER_225_1616 ();
 FILLCELL_X32 FILLER_225_1648 ();
 FILLCELL_X32 FILLER_225_1680 ();
 FILLCELL_X32 FILLER_225_1712 ();
 FILLCELL_X32 FILLER_225_1744 ();
 FILLCELL_X32 FILLER_225_1776 ();
 FILLCELL_X32 FILLER_225_1808 ();
 FILLCELL_X32 FILLER_225_1840 ();
 FILLCELL_X32 FILLER_225_1872 ();
 FILLCELL_X32 FILLER_225_1904 ();
 FILLCELL_X32 FILLER_225_1936 ();
 FILLCELL_X32 FILLER_225_1968 ();
 FILLCELL_X32 FILLER_225_2000 ();
 FILLCELL_X32 FILLER_225_2032 ();
 FILLCELL_X32 FILLER_225_2064 ();
 FILLCELL_X32 FILLER_225_2096 ();
 FILLCELL_X32 FILLER_225_2128 ();
 FILLCELL_X32 FILLER_225_2160 ();
 FILLCELL_X32 FILLER_225_2192 ();
 FILLCELL_X32 FILLER_225_2224 ();
 FILLCELL_X32 FILLER_225_2256 ();
 FILLCELL_X32 FILLER_225_2288 ();
 FILLCELL_X32 FILLER_225_2320 ();
 FILLCELL_X32 FILLER_225_2352 ();
 FILLCELL_X32 FILLER_225_2384 ();
 FILLCELL_X32 FILLER_225_2416 ();
 FILLCELL_X32 FILLER_225_2448 ();
 FILLCELL_X32 FILLER_225_2480 ();
 FILLCELL_X8 FILLER_225_2512 ();
 FILLCELL_X4 FILLER_225_2520 ();
 FILLCELL_X2 FILLER_225_2524 ();
 FILLCELL_X32 FILLER_225_2527 ();
 FILLCELL_X32 FILLER_225_2559 ();
 FILLCELL_X8 FILLER_225_2591 ();
 FILLCELL_X2 FILLER_225_2599 ();
 FILLCELL_X1 FILLER_225_2601 ();
 FILLCELL_X32 FILLER_226_1 ();
 FILLCELL_X32 FILLER_226_33 ();
 FILLCELL_X32 FILLER_226_65 ();
 FILLCELL_X32 FILLER_226_97 ();
 FILLCELL_X32 FILLER_226_129 ();
 FILLCELL_X32 FILLER_226_161 ();
 FILLCELL_X32 FILLER_226_193 ();
 FILLCELL_X32 FILLER_226_225 ();
 FILLCELL_X32 FILLER_226_257 ();
 FILLCELL_X32 FILLER_226_289 ();
 FILLCELL_X32 FILLER_226_321 ();
 FILLCELL_X32 FILLER_226_353 ();
 FILLCELL_X32 FILLER_226_385 ();
 FILLCELL_X32 FILLER_226_417 ();
 FILLCELL_X32 FILLER_226_449 ();
 FILLCELL_X32 FILLER_226_481 ();
 FILLCELL_X32 FILLER_226_513 ();
 FILLCELL_X32 FILLER_226_545 ();
 FILLCELL_X32 FILLER_226_577 ();
 FILLCELL_X16 FILLER_226_609 ();
 FILLCELL_X4 FILLER_226_625 ();
 FILLCELL_X2 FILLER_226_629 ();
 FILLCELL_X32 FILLER_226_632 ();
 FILLCELL_X32 FILLER_226_664 ();
 FILLCELL_X32 FILLER_226_696 ();
 FILLCELL_X32 FILLER_226_728 ();
 FILLCELL_X32 FILLER_226_760 ();
 FILLCELL_X32 FILLER_226_792 ();
 FILLCELL_X32 FILLER_226_824 ();
 FILLCELL_X32 FILLER_226_856 ();
 FILLCELL_X32 FILLER_226_888 ();
 FILLCELL_X32 FILLER_226_920 ();
 FILLCELL_X32 FILLER_226_952 ();
 FILLCELL_X32 FILLER_226_984 ();
 FILLCELL_X32 FILLER_226_1016 ();
 FILLCELL_X32 FILLER_226_1048 ();
 FILLCELL_X32 FILLER_226_1080 ();
 FILLCELL_X32 FILLER_226_1112 ();
 FILLCELL_X32 FILLER_226_1144 ();
 FILLCELL_X32 FILLER_226_1176 ();
 FILLCELL_X32 FILLER_226_1208 ();
 FILLCELL_X32 FILLER_226_1240 ();
 FILLCELL_X32 FILLER_226_1272 ();
 FILLCELL_X32 FILLER_226_1304 ();
 FILLCELL_X32 FILLER_226_1336 ();
 FILLCELL_X32 FILLER_226_1368 ();
 FILLCELL_X32 FILLER_226_1400 ();
 FILLCELL_X32 FILLER_226_1432 ();
 FILLCELL_X32 FILLER_226_1464 ();
 FILLCELL_X32 FILLER_226_1496 ();
 FILLCELL_X32 FILLER_226_1528 ();
 FILLCELL_X32 FILLER_226_1560 ();
 FILLCELL_X32 FILLER_226_1592 ();
 FILLCELL_X32 FILLER_226_1624 ();
 FILLCELL_X32 FILLER_226_1656 ();
 FILLCELL_X32 FILLER_226_1688 ();
 FILLCELL_X32 FILLER_226_1720 ();
 FILLCELL_X32 FILLER_226_1752 ();
 FILLCELL_X32 FILLER_226_1784 ();
 FILLCELL_X32 FILLER_226_1816 ();
 FILLCELL_X32 FILLER_226_1848 ();
 FILLCELL_X8 FILLER_226_1880 ();
 FILLCELL_X4 FILLER_226_1888 ();
 FILLCELL_X2 FILLER_226_1892 ();
 FILLCELL_X32 FILLER_226_1895 ();
 FILLCELL_X32 FILLER_226_1927 ();
 FILLCELL_X32 FILLER_226_1959 ();
 FILLCELL_X32 FILLER_226_1991 ();
 FILLCELL_X32 FILLER_226_2023 ();
 FILLCELL_X32 FILLER_226_2055 ();
 FILLCELL_X32 FILLER_226_2087 ();
 FILLCELL_X32 FILLER_226_2119 ();
 FILLCELL_X32 FILLER_226_2151 ();
 FILLCELL_X32 FILLER_226_2183 ();
 FILLCELL_X32 FILLER_226_2215 ();
 FILLCELL_X32 FILLER_226_2247 ();
 FILLCELL_X32 FILLER_226_2279 ();
 FILLCELL_X32 FILLER_226_2311 ();
 FILLCELL_X32 FILLER_226_2343 ();
 FILLCELL_X32 FILLER_226_2375 ();
 FILLCELL_X32 FILLER_226_2407 ();
 FILLCELL_X32 FILLER_226_2439 ();
 FILLCELL_X32 FILLER_226_2471 ();
 FILLCELL_X32 FILLER_226_2503 ();
 FILLCELL_X32 FILLER_226_2535 ();
 FILLCELL_X32 FILLER_226_2567 ();
 FILLCELL_X2 FILLER_226_2599 ();
 FILLCELL_X1 FILLER_226_2601 ();
 FILLCELL_X32 FILLER_227_1 ();
 FILLCELL_X32 FILLER_227_33 ();
 FILLCELL_X32 FILLER_227_65 ();
 FILLCELL_X32 FILLER_227_97 ();
 FILLCELL_X32 FILLER_227_129 ();
 FILLCELL_X32 FILLER_227_161 ();
 FILLCELL_X32 FILLER_227_193 ();
 FILLCELL_X32 FILLER_227_225 ();
 FILLCELL_X32 FILLER_227_257 ();
 FILLCELL_X32 FILLER_227_289 ();
 FILLCELL_X32 FILLER_227_321 ();
 FILLCELL_X32 FILLER_227_353 ();
 FILLCELL_X32 FILLER_227_385 ();
 FILLCELL_X32 FILLER_227_417 ();
 FILLCELL_X32 FILLER_227_449 ();
 FILLCELL_X32 FILLER_227_481 ();
 FILLCELL_X32 FILLER_227_513 ();
 FILLCELL_X32 FILLER_227_545 ();
 FILLCELL_X32 FILLER_227_577 ();
 FILLCELL_X32 FILLER_227_609 ();
 FILLCELL_X32 FILLER_227_641 ();
 FILLCELL_X32 FILLER_227_673 ();
 FILLCELL_X32 FILLER_227_705 ();
 FILLCELL_X32 FILLER_227_737 ();
 FILLCELL_X32 FILLER_227_769 ();
 FILLCELL_X32 FILLER_227_801 ();
 FILLCELL_X32 FILLER_227_833 ();
 FILLCELL_X32 FILLER_227_865 ();
 FILLCELL_X32 FILLER_227_897 ();
 FILLCELL_X32 FILLER_227_929 ();
 FILLCELL_X32 FILLER_227_961 ();
 FILLCELL_X32 FILLER_227_993 ();
 FILLCELL_X32 FILLER_227_1025 ();
 FILLCELL_X32 FILLER_227_1057 ();
 FILLCELL_X32 FILLER_227_1089 ();
 FILLCELL_X32 FILLER_227_1121 ();
 FILLCELL_X32 FILLER_227_1153 ();
 FILLCELL_X32 FILLER_227_1185 ();
 FILLCELL_X32 FILLER_227_1217 ();
 FILLCELL_X8 FILLER_227_1249 ();
 FILLCELL_X4 FILLER_227_1257 ();
 FILLCELL_X2 FILLER_227_1261 ();
 FILLCELL_X32 FILLER_227_1264 ();
 FILLCELL_X32 FILLER_227_1296 ();
 FILLCELL_X32 FILLER_227_1328 ();
 FILLCELL_X32 FILLER_227_1360 ();
 FILLCELL_X32 FILLER_227_1392 ();
 FILLCELL_X32 FILLER_227_1424 ();
 FILLCELL_X32 FILLER_227_1456 ();
 FILLCELL_X32 FILLER_227_1488 ();
 FILLCELL_X32 FILLER_227_1520 ();
 FILLCELL_X32 FILLER_227_1552 ();
 FILLCELL_X32 FILLER_227_1584 ();
 FILLCELL_X32 FILLER_227_1616 ();
 FILLCELL_X32 FILLER_227_1648 ();
 FILLCELL_X32 FILLER_227_1680 ();
 FILLCELL_X32 FILLER_227_1712 ();
 FILLCELL_X32 FILLER_227_1744 ();
 FILLCELL_X32 FILLER_227_1776 ();
 FILLCELL_X32 FILLER_227_1808 ();
 FILLCELL_X32 FILLER_227_1840 ();
 FILLCELL_X32 FILLER_227_1872 ();
 FILLCELL_X32 FILLER_227_1904 ();
 FILLCELL_X32 FILLER_227_1936 ();
 FILLCELL_X32 FILLER_227_1968 ();
 FILLCELL_X32 FILLER_227_2000 ();
 FILLCELL_X32 FILLER_227_2032 ();
 FILLCELL_X32 FILLER_227_2064 ();
 FILLCELL_X32 FILLER_227_2096 ();
 FILLCELL_X32 FILLER_227_2128 ();
 FILLCELL_X32 FILLER_227_2160 ();
 FILLCELL_X32 FILLER_227_2192 ();
 FILLCELL_X32 FILLER_227_2224 ();
 FILLCELL_X32 FILLER_227_2256 ();
 FILLCELL_X32 FILLER_227_2288 ();
 FILLCELL_X32 FILLER_227_2320 ();
 FILLCELL_X32 FILLER_227_2352 ();
 FILLCELL_X32 FILLER_227_2384 ();
 FILLCELL_X32 FILLER_227_2416 ();
 FILLCELL_X32 FILLER_227_2448 ();
 FILLCELL_X32 FILLER_227_2480 ();
 FILLCELL_X8 FILLER_227_2512 ();
 FILLCELL_X4 FILLER_227_2520 ();
 FILLCELL_X2 FILLER_227_2524 ();
 FILLCELL_X32 FILLER_227_2527 ();
 FILLCELL_X32 FILLER_227_2559 ();
 FILLCELL_X8 FILLER_227_2591 ();
 FILLCELL_X2 FILLER_227_2599 ();
 FILLCELL_X1 FILLER_227_2601 ();
 FILLCELL_X32 FILLER_228_1 ();
 FILLCELL_X32 FILLER_228_33 ();
 FILLCELL_X32 FILLER_228_65 ();
 FILLCELL_X32 FILLER_228_97 ();
 FILLCELL_X32 FILLER_228_129 ();
 FILLCELL_X32 FILLER_228_161 ();
 FILLCELL_X32 FILLER_228_193 ();
 FILLCELL_X32 FILLER_228_225 ();
 FILLCELL_X32 FILLER_228_257 ();
 FILLCELL_X32 FILLER_228_289 ();
 FILLCELL_X32 FILLER_228_321 ();
 FILLCELL_X32 FILLER_228_353 ();
 FILLCELL_X32 FILLER_228_385 ();
 FILLCELL_X32 FILLER_228_417 ();
 FILLCELL_X32 FILLER_228_449 ();
 FILLCELL_X32 FILLER_228_481 ();
 FILLCELL_X32 FILLER_228_513 ();
 FILLCELL_X32 FILLER_228_545 ();
 FILLCELL_X32 FILLER_228_577 ();
 FILLCELL_X16 FILLER_228_609 ();
 FILLCELL_X4 FILLER_228_625 ();
 FILLCELL_X2 FILLER_228_629 ();
 FILLCELL_X32 FILLER_228_632 ();
 FILLCELL_X32 FILLER_228_664 ();
 FILLCELL_X32 FILLER_228_696 ();
 FILLCELL_X32 FILLER_228_728 ();
 FILLCELL_X32 FILLER_228_760 ();
 FILLCELL_X32 FILLER_228_792 ();
 FILLCELL_X32 FILLER_228_824 ();
 FILLCELL_X32 FILLER_228_856 ();
 FILLCELL_X32 FILLER_228_888 ();
 FILLCELL_X32 FILLER_228_920 ();
 FILLCELL_X32 FILLER_228_952 ();
 FILLCELL_X32 FILLER_228_984 ();
 FILLCELL_X32 FILLER_228_1016 ();
 FILLCELL_X32 FILLER_228_1048 ();
 FILLCELL_X32 FILLER_228_1080 ();
 FILLCELL_X32 FILLER_228_1112 ();
 FILLCELL_X32 FILLER_228_1144 ();
 FILLCELL_X32 FILLER_228_1176 ();
 FILLCELL_X32 FILLER_228_1208 ();
 FILLCELL_X32 FILLER_228_1240 ();
 FILLCELL_X32 FILLER_228_1272 ();
 FILLCELL_X32 FILLER_228_1304 ();
 FILLCELL_X32 FILLER_228_1336 ();
 FILLCELL_X32 FILLER_228_1368 ();
 FILLCELL_X32 FILLER_228_1400 ();
 FILLCELL_X32 FILLER_228_1432 ();
 FILLCELL_X32 FILLER_228_1464 ();
 FILLCELL_X32 FILLER_228_1496 ();
 FILLCELL_X32 FILLER_228_1528 ();
 FILLCELL_X32 FILLER_228_1560 ();
 FILLCELL_X32 FILLER_228_1592 ();
 FILLCELL_X32 FILLER_228_1624 ();
 FILLCELL_X32 FILLER_228_1656 ();
 FILLCELL_X32 FILLER_228_1688 ();
 FILLCELL_X32 FILLER_228_1720 ();
 FILLCELL_X32 FILLER_228_1752 ();
 FILLCELL_X32 FILLER_228_1784 ();
 FILLCELL_X32 FILLER_228_1816 ();
 FILLCELL_X32 FILLER_228_1848 ();
 FILLCELL_X8 FILLER_228_1880 ();
 FILLCELL_X4 FILLER_228_1888 ();
 FILLCELL_X2 FILLER_228_1892 ();
 FILLCELL_X32 FILLER_228_1895 ();
 FILLCELL_X32 FILLER_228_1927 ();
 FILLCELL_X32 FILLER_228_1959 ();
 FILLCELL_X32 FILLER_228_1991 ();
 FILLCELL_X32 FILLER_228_2023 ();
 FILLCELL_X32 FILLER_228_2055 ();
 FILLCELL_X32 FILLER_228_2087 ();
 FILLCELL_X32 FILLER_228_2119 ();
 FILLCELL_X32 FILLER_228_2151 ();
 FILLCELL_X32 FILLER_228_2183 ();
 FILLCELL_X32 FILLER_228_2215 ();
 FILLCELL_X32 FILLER_228_2247 ();
 FILLCELL_X32 FILLER_228_2279 ();
 FILLCELL_X32 FILLER_228_2311 ();
 FILLCELL_X32 FILLER_228_2343 ();
 FILLCELL_X32 FILLER_228_2375 ();
 FILLCELL_X32 FILLER_228_2407 ();
 FILLCELL_X32 FILLER_228_2439 ();
 FILLCELL_X32 FILLER_228_2471 ();
 FILLCELL_X32 FILLER_228_2503 ();
 FILLCELL_X32 FILLER_228_2535 ();
 FILLCELL_X32 FILLER_228_2567 ();
 FILLCELL_X2 FILLER_228_2599 ();
 FILLCELL_X1 FILLER_228_2601 ();
 FILLCELL_X32 FILLER_229_1 ();
 FILLCELL_X32 FILLER_229_33 ();
 FILLCELL_X32 FILLER_229_65 ();
 FILLCELL_X32 FILLER_229_97 ();
 FILLCELL_X32 FILLER_229_129 ();
 FILLCELL_X32 FILLER_229_161 ();
 FILLCELL_X32 FILLER_229_193 ();
 FILLCELL_X32 FILLER_229_225 ();
 FILLCELL_X32 FILLER_229_257 ();
 FILLCELL_X32 FILLER_229_289 ();
 FILLCELL_X32 FILLER_229_321 ();
 FILLCELL_X32 FILLER_229_353 ();
 FILLCELL_X32 FILLER_229_385 ();
 FILLCELL_X32 FILLER_229_417 ();
 FILLCELL_X32 FILLER_229_449 ();
 FILLCELL_X32 FILLER_229_481 ();
 FILLCELL_X32 FILLER_229_513 ();
 FILLCELL_X32 FILLER_229_545 ();
 FILLCELL_X32 FILLER_229_577 ();
 FILLCELL_X32 FILLER_229_609 ();
 FILLCELL_X32 FILLER_229_641 ();
 FILLCELL_X32 FILLER_229_673 ();
 FILLCELL_X32 FILLER_229_705 ();
 FILLCELL_X32 FILLER_229_737 ();
 FILLCELL_X32 FILLER_229_769 ();
 FILLCELL_X32 FILLER_229_801 ();
 FILLCELL_X32 FILLER_229_833 ();
 FILLCELL_X32 FILLER_229_865 ();
 FILLCELL_X32 FILLER_229_897 ();
 FILLCELL_X32 FILLER_229_929 ();
 FILLCELL_X32 FILLER_229_961 ();
 FILLCELL_X32 FILLER_229_993 ();
 FILLCELL_X32 FILLER_229_1025 ();
 FILLCELL_X32 FILLER_229_1057 ();
 FILLCELL_X32 FILLER_229_1089 ();
 FILLCELL_X32 FILLER_229_1121 ();
 FILLCELL_X32 FILLER_229_1153 ();
 FILLCELL_X32 FILLER_229_1185 ();
 FILLCELL_X32 FILLER_229_1217 ();
 FILLCELL_X8 FILLER_229_1249 ();
 FILLCELL_X4 FILLER_229_1257 ();
 FILLCELL_X2 FILLER_229_1261 ();
 FILLCELL_X32 FILLER_229_1264 ();
 FILLCELL_X32 FILLER_229_1296 ();
 FILLCELL_X32 FILLER_229_1328 ();
 FILLCELL_X32 FILLER_229_1360 ();
 FILLCELL_X32 FILLER_229_1392 ();
 FILLCELL_X32 FILLER_229_1424 ();
 FILLCELL_X32 FILLER_229_1456 ();
 FILLCELL_X32 FILLER_229_1488 ();
 FILLCELL_X32 FILLER_229_1520 ();
 FILLCELL_X32 FILLER_229_1552 ();
 FILLCELL_X32 FILLER_229_1584 ();
 FILLCELL_X32 FILLER_229_1616 ();
 FILLCELL_X32 FILLER_229_1648 ();
 FILLCELL_X32 FILLER_229_1680 ();
 FILLCELL_X32 FILLER_229_1712 ();
 FILLCELL_X32 FILLER_229_1744 ();
 FILLCELL_X32 FILLER_229_1776 ();
 FILLCELL_X32 FILLER_229_1808 ();
 FILLCELL_X32 FILLER_229_1840 ();
 FILLCELL_X32 FILLER_229_1872 ();
 FILLCELL_X32 FILLER_229_1904 ();
 FILLCELL_X32 FILLER_229_1936 ();
 FILLCELL_X32 FILLER_229_1968 ();
 FILLCELL_X32 FILLER_229_2000 ();
 FILLCELL_X32 FILLER_229_2032 ();
 FILLCELL_X32 FILLER_229_2064 ();
 FILLCELL_X32 FILLER_229_2096 ();
 FILLCELL_X32 FILLER_229_2128 ();
 FILLCELL_X32 FILLER_229_2160 ();
 FILLCELL_X32 FILLER_229_2192 ();
 FILLCELL_X32 FILLER_229_2224 ();
 FILLCELL_X32 FILLER_229_2256 ();
 FILLCELL_X32 FILLER_229_2288 ();
 FILLCELL_X32 FILLER_229_2320 ();
 FILLCELL_X32 FILLER_229_2352 ();
 FILLCELL_X32 FILLER_229_2384 ();
 FILLCELL_X32 FILLER_229_2416 ();
 FILLCELL_X32 FILLER_229_2448 ();
 FILLCELL_X32 FILLER_229_2480 ();
 FILLCELL_X8 FILLER_229_2512 ();
 FILLCELL_X4 FILLER_229_2520 ();
 FILLCELL_X2 FILLER_229_2524 ();
 FILLCELL_X32 FILLER_229_2527 ();
 FILLCELL_X32 FILLER_229_2559 ();
 FILLCELL_X8 FILLER_229_2591 ();
 FILLCELL_X2 FILLER_229_2599 ();
 FILLCELL_X1 FILLER_229_2601 ();
 FILLCELL_X32 FILLER_230_1 ();
 FILLCELL_X32 FILLER_230_33 ();
 FILLCELL_X32 FILLER_230_65 ();
 FILLCELL_X32 FILLER_230_97 ();
 FILLCELL_X32 FILLER_230_129 ();
 FILLCELL_X32 FILLER_230_161 ();
 FILLCELL_X32 FILLER_230_193 ();
 FILLCELL_X32 FILLER_230_225 ();
 FILLCELL_X32 FILLER_230_257 ();
 FILLCELL_X32 FILLER_230_289 ();
 FILLCELL_X32 FILLER_230_321 ();
 FILLCELL_X32 FILLER_230_353 ();
 FILLCELL_X32 FILLER_230_385 ();
 FILLCELL_X32 FILLER_230_417 ();
 FILLCELL_X32 FILLER_230_449 ();
 FILLCELL_X32 FILLER_230_481 ();
 FILLCELL_X32 FILLER_230_513 ();
 FILLCELL_X32 FILLER_230_545 ();
 FILLCELL_X32 FILLER_230_577 ();
 FILLCELL_X16 FILLER_230_609 ();
 FILLCELL_X4 FILLER_230_625 ();
 FILLCELL_X2 FILLER_230_629 ();
 FILLCELL_X32 FILLER_230_632 ();
 FILLCELL_X32 FILLER_230_664 ();
 FILLCELL_X32 FILLER_230_696 ();
 FILLCELL_X32 FILLER_230_728 ();
 FILLCELL_X32 FILLER_230_760 ();
 FILLCELL_X32 FILLER_230_792 ();
 FILLCELL_X32 FILLER_230_824 ();
 FILLCELL_X32 FILLER_230_856 ();
 FILLCELL_X32 FILLER_230_888 ();
 FILLCELL_X32 FILLER_230_920 ();
 FILLCELL_X32 FILLER_230_952 ();
 FILLCELL_X32 FILLER_230_984 ();
 FILLCELL_X32 FILLER_230_1016 ();
 FILLCELL_X32 FILLER_230_1048 ();
 FILLCELL_X32 FILLER_230_1080 ();
 FILLCELL_X32 FILLER_230_1112 ();
 FILLCELL_X32 FILLER_230_1144 ();
 FILLCELL_X32 FILLER_230_1176 ();
 FILLCELL_X32 FILLER_230_1208 ();
 FILLCELL_X32 FILLER_230_1240 ();
 FILLCELL_X32 FILLER_230_1272 ();
 FILLCELL_X32 FILLER_230_1304 ();
 FILLCELL_X32 FILLER_230_1336 ();
 FILLCELL_X32 FILLER_230_1368 ();
 FILLCELL_X32 FILLER_230_1400 ();
 FILLCELL_X32 FILLER_230_1432 ();
 FILLCELL_X32 FILLER_230_1464 ();
 FILLCELL_X32 FILLER_230_1496 ();
 FILLCELL_X32 FILLER_230_1528 ();
 FILLCELL_X32 FILLER_230_1560 ();
 FILLCELL_X32 FILLER_230_1592 ();
 FILLCELL_X32 FILLER_230_1624 ();
 FILLCELL_X32 FILLER_230_1656 ();
 FILLCELL_X32 FILLER_230_1688 ();
 FILLCELL_X32 FILLER_230_1720 ();
 FILLCELL_X32 FILLER_230_1752 ();
 FILLCELL_X32 FILLER_230_1784 ();
 FILLCELL_X32 FILLER_230_1816 ();
 FILLCELL_X32 FILLER_230_1848 ();
 FILLCELL_X8 FILLER_230_1880 ();
 FILLCELL_X4 FILLER_230_1888 ();
 FILLCELL_X2 FILLER_230_1892 ();
 FILLCELL_X32 FILLER_230_1895 ();
 FILLCELL_X32 FILLER_230_1927 ();
 FILLCELL_X32 FILLER_230_1959 ();
 FILLCELL_X32 FILLER_230_1991 ();
 FILLCELL_X32 FILLER_230_2023 ();
 FILLCELL_X32 FILLER_230_2055 ();
 FILLCELL_X32 FILLER_230_2087 ();
 FILLCELL_X32 FILLER_230_2119 ();
 FILLCELL_X32 FILLER_230_2151 ();
 FILLCELL_X32 FILLER_230_2183 ();
 FILLCELL_X32 FILLER_230_2215 ();
 FILLCELL_X32 FILLER_230_2247 ();
 FILLCELL_X32 FILLER_230_2279 ();
 FILLCELL_X32 FILLER_230_2311 ();
 FILLCELL_X32 FILLER_230_2343 ();
 FILLCELL_X32 FILLER_230_2375 ();
 FILLCELL_X32 FILLER_230_2407 ();
 FILLCELL_X32 FILLER_230_2439 ();
 FILLCELL_X32 FILLER_230_2471 ();
 FILLCELL_X32 FILLER_230_2503 ();
 FILLCELL_X32 FILLER_230_2535 ();
 FILLCELL_X32 FILLER_230_2567 ();
 FILLCELL_X2 FILLER_230_2599 ();
 FILLCELL_X1 FILLER_230_2601 ();
 FILLCELL_X32 FILLER_231_1 ();
 FILLCELL_X32 FILLER_231_33 ();
 FILLCELL_X32 FILLER_231_65 ();
 FILLCELL_X32 FILLER_231_97 ();
 FILLCELL_X32 FILLER_231_129 ();
 FILLCELL_X32 FILLER_231_161 ();
 FILLCELL_X32 FILLER_231_193 ();
 FILLCELL_X32 FILLER_231_225 ();
 FILLCELL_X32 FILLER_231_257 ();
 FILLCELL_X32 FILLER_231_289 ();
 FILLCELL_X32 FILLER_231_321 ();
 FILLCELL_X32 FILLER_231_353 ();
 FILLCELL_X32 FILLER_231_385 ();
 FILLCELL_X32 FILLER_231_417 ();
 FILLCELL_X32 FILLER_231_449 ();
 FILLCELL_X32 FILLER_231_481 ();
 FILLCELL_X32 FILLER_231_513 ();
 FILLCELL_X32 FILLER_231_545 ();
 FILLCELL_X32 FILLER_231_577 ();
 FILLCELL_X32 FILLER_231_609 ();
 FILLCELL_X32 FILLER_231_641 ();
 FILLCELL_X32 FILLER_231_673 ();
 FILLCELL_X32 FILLER_231_705 ();
 FILLCELL_X32 FILLER_231_737 ();
 FILLCELL_X32 FILLER_231_769 ();
 FILLCELL_X32 FILLER_231_801 ();
 FILLCELL_X32 FILLER_231_833 ();
 FILLCELL_X32 FILLER_231_865 ();
 FILLCELL_X32 FILLER_231_897 ();
 FILLCELL_X32 FILLER_231_929 ();
 FILLCELL_X32 FILLER_231_961 ();
 FILLCELL_X32 FILLER_231_993 ();
 FILLCELL_X32 FILLER_231_1025 ();
 FILLCELL_X32 FILLER_231_1057 ();
 FILLCELL_X32 FILLER_231_1089 ();
 FILLCELL_X32 FILLER_231_1121 ();
 FILLCELL_X32 FILLER_231_1153 ();
 FILLCELL_X32 FILLER_231_1185 ();
 FILLCELL_X32 FILLER_231_1217 ();
 FILLCELL_X8 FILLER_231_1249 ();
 FILLCELL_X4 FILLER_231_1257 ();
 FILLCELL_X2 FILLER_231_1261 ();
 FILLCELL_X32 FILLER_231_1264 ();
 FILLCELL_X32 FILLER_231_1296 ();
 FILLCELL_X32 FILLER_231_1328 ();
 FILLCELL_X32 FILLER_231_1360 ();
 FILLCELL_X32 FILLER_231_1392 ();
 FILLCELL_X32 FILLER_231_1424 ();
 FILLCELL_X32 FILLER_231_1456 ();
 FILLCELL_X32 FILLER_231_1488 ();
 FILLCELL_X32 FILLER_231_1520 ();
 FILLCELL_X32 FILLER_231_1552 ();
 FILLCELL_X32 FILLER_231_1584 ();
 FILLCELL_X32 FILLER_231_1616 ();
 FILLCELL_X32 FILLER_231_1648 ();
 FILLCELL_X32 FILLER_231_1680 ();
 FILLCELL_X32 FILLER_231_1712 ();
 FILLCELL_X32 FILLER_231_1744 ();
 FILLCELL_X32 FILLER_231_1776 ();
 FILLCELL_X32 FILLER_231_1808 ();
 FILLCELL_X32 FILLER_231_1840 ();
 FILLCELL_X32 FILLER_231_1872 ();
 FILLCELL_X32 FILLER_231_1904 ();
 FILLCELL_X32 FILLER_231_1936 ();
 FILLCELL_X32 FILLER_231_1968 ();
 FILLCELL_X32 FILLER_231_2000 ();
 FILLCELL_X32 FILLER_231_2032 ();
 FILLCELL_X32 FILLER_231_2064 ();
 FILLCELL_X32 FILLER_231_2096 ();
 FILLCELL_X32 FILLER_231_2128 ();
 FILLCELL_X32 FILLER_231_2160 ();
 FILLCELL_X32 FILLER_231_2192 ();
 FILLCELL_X32 FILLER_231_2224 ();
 FILLCELL_X32 FILLER_231_2256 ();
 FILLCELL_X32 FILLER_231_2288 ();
 FILLCELL_X32 FILLER_231_2320 ();
 FILLCELL_X32 FILLER_231_2352 ();
 FILLCELL_X32 FILLER_231_2384 ();
 FILLCELL_X32 FILLER_231_2416 ();
 FILLCELL_X32 FILLER_231_2448 ();
 FILLCELL_X32 FILLER_231_2480 ();
 FILLCELL_X8 FILLER_231_2512 ();
 FILLCELL_X4 FILLER_231_2520 ();
 FILLCELL_X2 FILLER_231_2524 ();
 FILLCELL_X32 FILLER_231_2527 ();
 FILLCELL_X32 FILLER_231_2559 ();
 FILLCELL_X8 FILLER_231_2591 ();
 FILLCELL_X2 FILLER_231_2599 ();
 FILLCELL_X1 FILLER_231_2601 ();
 FILLCELL_X32 FILLER_232_1 ();
 FILLCELL_X32 FILLER_232_33 ();
 FILLCELL_X32 FILLER_232_65 ();
 FILLCELL_X32 FILLER_232_97 ();
 FILLCELL_X32 FILLER_232_129 ();
 FILLCELL_X32 FILLER_232_161 ();
 FILLCELL_X32 FILLER_232_193 ();
 FILLCELL_X32 FILLER_232_225 ();
 FILLCELL_X32 FILLER_232_257 ();
 FILLCELL_X32 FILLER_232_289 ();
 FILLCELL_X32 FILLER_232_321 ();
 FILLCELL_X32 FILLER_232_353 ();
 FILLCELL_X32 FILLER_232_385 ();
 FILLCELL_X32 FILLER_232_417 ();
 FILLCELL_X32 FILLER_232_449 ();
 FILLCELL_X32 FILLER_232_481 ();
 FILLCELL_X32 FILLER_232_513 ();
 FILLCELL_X32 FILLER_232_545 ();
 FILLCELL_X32 FILLER_232_577 ();
 FILLCELL_X16 FILLER_232_609 ();
 FILLCELL_X4 FILLER_232_625 ();
 FILLCELL_X2 FILLER_232_629 ();
 FILLCELL_X32 FILLER_232_632 ();
 FILLCELL_X32 FILLER_232_664 ();
 FILLCELL_X32 FILLER_232_696 ();
 FILLCELL_X32 FILLER_232_728 ();
 FILLCELL_X32 FILLER_232_760 ();
 FILLCELL_X32 FILLER_232_792 ();
 FILLCELL_X32 FILLER_232_824 ();
 FILLCELL_X32 FILLER_232_856 ();
 FILLCELL_X32 FILLER_232_888 ();
 FILLCELL_X32 FILLER_232_920 ();
 FILLCELL_X32 FILLER_232_952 ();
 FILLCELL_X32 FILLER_232_984 ();
 FILLCELL_X32 FILLER_232_1016 ();
 FILLCELL_X32 FILLER_232_1048 ();
 FILLCELL_X32 FILLER_232_1080 ();
 FILLCELL_X32 FILLER_232_1112 ();
 FILLCELL_X32 FILLER_232_1144 ();
 FILLCELL_X32 FILLER_232_1176 ();
 FILLCELL_X32 FILLER_232_1208 ();
 FILLCELL_X32 FILLER_232_1240 ();
 FILLCELL_X32 FILLER_232_1272 ();
 FILLCELL_X32 FILLER_232_1304 ();
 FILLCELL_X32 FILLER_232_1336 ();
 FILLCELL_X32 FILLER_232_1368 ();
 FILLCELL_X32 FILLER_232_1400 ();
 FILLCELL_X32 FILLER_232_1432 ();
 FILLCELL_X32 FILLER_232_1464 ();
 FILLCELL_X32 FILLER_232_1496 ();
 FILLCELL_X32 FILLER_232_1528 ();
 FILLCELL_X32 FILLER_232_1560 ();
 FILLCELL_X32 FILLER_232_1592 ();
 FILLCELL_X32 FILLER_232_1624 ();
 FILLCELL_X32 FILLER_232_1656 ();
 FILLCELL_X32 FILLER_232_1688 ();
 FILLCELL_X32 FILLER_232_1720 ();
 FILLCELL_X32 FILLER_232_1752 ();
 FILLCELL_X32 FILLER_232_1784 ();
 FILLCELL_X32 FILLER_232_1816 ();
 FILLCELL_X32 FILLER_232_1848 ();
 FILLCELL_X8 FILLER_232_1880 ();
 FILLCELL_X4 FILLER_232_1888 ();
 FILLCELL_X2 FILLER_232_1892 ();
 FILLCELL_X32 FILLER_232_1895 ();
 FILLCELL_X32 FILLER_232_1927 ();
 FILLCELL_X32 FILLER_232_1959 ();
 FILLCELL_X32 FILLER_232_1991 ();
 FILLCELL_X32 FILLER_232_2023 ();
 FILLCELL_X32 FILLER_232_2055 ();
 FILLCELL_X32 FILLER_232_2087 ();
 FILLCELL_X32 FILLER_232_2119 ();
 FILLCELL_X32 FILLER_232_2151 ();
 FILLCELL_X32 FILLER_232_2183 ();
 FILLCELL_X32 FILLER_232_2215 ();
 FILLCELL_X32 FILLER_232_2247 ();
 FILLCELL_X32 FILLER_232_2279 ();
 FILLCELL_X32 FILLER_232_2311 ();
 FILLCELL_X32 FILLER_232_2343 ();
 FILLCELL_X32 FILLER_232_2375 ();
 FILLCELL_X32 FILLER_232_2407 ();
 FILLCELL_X32 FILLER_232_2439 ();
 FILLCELL_X32 FILLER_232_2471 ();
 FILLCELL_X32 FILLER_232_2503 ();
 FILLCELL_X32 FILLER_232_2535 ();
 FILLCELL_X32 FILLER_232_2567 ();
 FILLCELL_X2 FILLER_232_2599 ();
 FILLCELL_X1 FILLER_232_2601 ();
 FILLCELL_X32 FILLER_233_1 ();
 FILLCELL_X32 FILLER_233_33 ();
 FILLCELL_X32 FILLER_233_65 ();
 FILLCELL_X32 FILLER_233_97 ();
 FILLCELL_X32 FILLER_233_129 ();
 FILLCELL_X32 FILLER_233_161 ();
 FILLCELL_X32 FILLER_233_193 ();
 FILLCELL_X32 FILLER_233_225 ();
 FILLCELL_X32 FILLER_233_257 ();
 FILLCELL_X32 FILLER_233_289 ();
 FILLCELL_X32 FILLER_233_321 ();
 FILLCELL_X32 FILLER_233_353 ();
 FILLCELL_X32 FILLER_233_385 ();
 FILLCELL_X32 FILLER_233_417 ();
 FILLCELL_X32 FILLER_233_449 ();
 FILLCELL_X32 FILLER_233_481 ();
 FILLCELL_X32 FILLER_233_513 ();
 FILLCELL_X32 FILLER_233_545 ();
 FILLCELL_X32 FILLER_233_577 ();
 FILLCELL_X32 FILLER_233_609 ();
 FILLCELL_X32 FILLER_233_641 ();
 FILLCELL_X32 FILLER_233_673 ();
 FILLCELL_X32 FILLER_233_705 ();
 FILLCELL_X32 FILLER_233_737 ();
 FILLCELL_X32 FILLER_233_769 ();
 FILLCELL_X32 FILLER_233_801 ();
 FILLCELL_X32 FILLER_233_833 ();
 FILLCELL_X32 FILLER_233_865 ();
 FILLCELL_X32 FILLER_233_897 ();
 FILLCELL_X32 FILLER_233_929 ();
 FILLCELL_X32 FILLER_233_961 ();
 FILLCELL_X32 FILLER_233_993 ();
 FILLCELL_X32 FILLER_233_1025 ();
 FILLCELL_X32 FILLER_233_1057 ();
 FILLCELL_X32 FILLER_233_1089 ();
 FILLCELL_X32 FILLER_233_1121 ();
 FILLCELL_X32 FILLER_233_1153 ();
 FILLCELL_X32 FILLER_233_1185 ();
 FILLCELL_X32 FILLER_233_1217 ();
 FILLCELL_X8 FILLER_233_1249 ();
 FILLCELL_X4 FILLER_233_1257 ();
 FILLCELL_X2 FILLER_233_1261 ();
 FILLCELL_X32 FILLER_233_1264 ();
 FILLCELL_X32 FILLER_233_1296 ();
 FILLCELL_X32 FILLER_233_1328 ();
 FILLCELL_X32 FILLER_233_1360 ();
 FILLCELL_X32 FILLER_233_1392 ();
 FILLCELL_X32 FILLER_233_1424 ();
 FILLCELL_X32 FILLER_233_1456 ();
 FILLCELL_X32 FILLER_233_1488 ();
 FILLCELL_X32 FILLER_233_1520 ();
 FILLCELL_X32 FILLER_233_1552 ();
 FILLCELL_X32 FILLER_233_1584 ();
 FILLCELL_X32 FILLER_233_1616 ();
 FILLCELL_X32 FILLER_233_1648 ();
 FILLCELL_X32 FILLER_233_1680 ();
 FILLCELL_X32 FILLER_233_1712 ();
 FILLCELL_X32 FILLER_233_1744 ();
 FILLCELL_X32 FILLER_233_1776 ();
 FILLCELL_X32 FILLER_233_1808 ();
 FILLCELL_X32 FILLER_233_1840 ();
 FILLCELL_X32 FILLER_233_1872 ();
 FILLCELL_X32 FILLER_233_1904 ();
 FILLCELL_X32 FILLER_233_1936 ();
 FILLCELL_X32 FILLER_233_1968 ();
 FILLCELL_X32 FILLER_233_2000 ();
 FILLCELL_X32 FILLER_233_2032 ();
 FILLCELL_X32 FILLER_233_2064 ();
 FILLCELL_X32 FILLER_233_2096 ();
 FILLCELL_X32 FILLER_233_2128 ();
 FILLCELL_X32 FILLER_233_2160 ();
 FILLCELL_X32 FILLER_233_2192 ();
 FILLCELL_X32 FILLER_233_2224 ();
 FILLCELL_X32 FILLER_233_2256 ();
 FILLCELL_X32 FILLER_233_2288 ();
 FILLCELL_X32 FILLER_233_2320 ();
 FILLCELL_X32 FILLER_233_2352 ();
 FILLCELL_X32 FILLER_233_2384 ();
 FILLCELL_X32 FILLER_233_2416 ();
 FILLCELL_X32 FILLER_233_2448 ();
 FILLCELL_X32 FILLER_233_2480 ();
 FILLCELL_X8 FILLER_233_2512 ();
 FILLCELL_X4 FILLER_233_2520 ();
 FILLCELL_X2 FILLER_233_2524 ();
 FILLCELL_X32 FILLER_233_2527 ();
 FILLCELL_X32 FILLER_233_2559 ();
 FILLCELL_X8 FILLER_233_2591 ();
 FILLCELL_X2 FILLER_233_2599 ();
 FILLCELL_X1 FILLER_233_2601 ();
 FILLCELL_X32 FILLER_234_1 ();
 FILLCELL_X32 FILLER_234_33 ();
 FILLCELL_X32 FILLER_234_65 ();
 FILLCELL_X32 FILLER_234_97 ();
 FILLCELL_X32 FILLER_234_129 ();
 FILLCELL_X32 FILLER_234_161 ();
 FILLCELL_X32 FILLER_234_193 ();
 FILLCELL_X32 FILLER_234_225 ();
 FILLCELL_X32 FILLER_234_257 ();
 FILLCELL_X32 FILLER_234_289 ();
 FILLCELL_X32 FILLER_234_321 ();
 FILLCELL_X32 FILLER_234_353 ();
 FILLCELL_X32 FILLER_234_385 ();
 FILLCELL_X32 FILLER_234_417 ();
 FILLCELL_X32 FILLER_234_449 ();
 FILLCELL_X32 FILLER_234_481 ();
 FILLCELL_X32 FILLER_234_513 ();
 FILLCELL_X32 FILLER_234_545 ();
 FILLCELL_X32 FILLER_234_577 ();
 FILLCELL_X16 FILLER_234_609 ();
 FILLCELL_X4 FILLER_234_625 ();
 FILLCELL_X2 FILLER_234_629 ();
 FILLCELL_X32 FILLER_234_632 ();
 FILLCELL_X32 FILLER_234_664 ();
 FILLCELL_X32 FILLER_234_696 ();
 FILLCELL_X32 FILLER_234_728 ();
 FILLCELL_X32 FILLER_234_760 ();
 FILLCELL_X32 FILLER_234_792 ();
 FILLCELL_X32 FILLER_234_824 ();
 FILLCELL_X32 FILLER_234_856 ();
 FILLCELL_X32 FILLER_234_888 ();
 FILLCELL_X32 FILLER_234_920 ();
 FILLCELL_X32 FILLER_234_952 ();
 FILLCELL_X32 FILLER_234_984 ();
 FILLCELL_X32 FILLER_234_1016 ();
 FILLCELL_X32 FILLER_234_1048 ();
 FILLCELL_X32 FILLER_234_1080 ();
 FILLCELL_X32 FILLER_234_1112 ();
 FILLCELL_X32 FILLER_234_1144 ();
 FILLCELL_X32 FILLER_234_1176 ();
 FILLCELL_X32 FILLER_234_1208 ();
 FILLCELL_X32 FILLER_234_1240 ();
 FILLCELL_X32 FILLER_234_1272 ();
 FILLCELL_X32 FILLER_234_1304 ();
 FILLCELL_X32 FILLER_234_1336 ();
 FILLCELL_X32 FILLER_234_1368 ();
 FILLCELL_X32 FILLER_234_1400 ();
 FILLCELL_X32 FILLER_234_1432 ();
 FILLCELL_X32 FILLER_234_1464 ();
 FILLCELL_X32 FILLER_234_1496 ();
 FILLCELL_X32 FILLER_234_1528 ();
 FILLCELL_X32 FILLER_234_1560 ();
 FILLCELL_X32 FILLER_234_1592 ();
 FILLCELL_X32 FILLER_234_1624 ();
 FILLCELL_X32 FILLER_234_1656 ();
 FILLCELL_X32 FILLER_234_1688 ();
 FILLCELL_X32 FILLER_234_1720 ();
 FILLCELL_X32 FILLER_234_1752 ();
 FILLCELL_X32 FILLER_234_1784 ();
 FILLCELL_X32 FILLER_234_1816 ();
 FILLCELL_X32 FILLER_234_1848 ();
 FILLCELL_X8 FILLER_234_1880 ();
 FILLCELL_X4 FILLER_234_1888 ();
 FILLCELL_X2 FILLER_234_1892 ();
 FILLCELL_X32 FILLER_234_1895 ();
 FILLCELL_X32 FILLER_234_1927 ();
 FILLCELL_X32 FILLER_234_1959 ();
 FILLCELL_X32 FILLER_234_1991 ();
 FILLCELL_X32 FILLER_234_2023 ();
 FILLCELL_X32 FILLER_234_2055 ();
 FILLCELL_X32 FILLER_234_2087 ();
 FILLCELL_X32 FILLER_234_2119 ();
 FILLCELL_X32 FILLER_234_2151 ();
 FILLCELL_X32 FILLER_234_2183 ();
 FILLCELL_X32 FILLER_234_2215 ();
 FILLCELL_X32 FILLER_234_2247 ();
 FILLCELL_X32 FILLER_234_2279 ();
 FILLCELL_X32 FILLER_234_2311 ();
 FILLCELL_X32 FILLER_234_2343 ();
 FILLCELL_X32 FILLER_234_2375 ();
 FILLCELL_X32 FILLER_234_2407 ();
 FILLCELL_X32 FILLER_234_2439 ();
 FILLCELL_X32 FILLER_234_2471 ();
 FILLCELL_X32 FILLER_234_2503 ();
 FILLCELL_X32 FILLER_234_2535 ();
 FILLCELL_X32 FILLER_234_2567 ();
 FILLCELL_X2 FILLER_234_2599 ();
 FILLCELL_X1 FILLER_234_2601 ();
 FILLCELL_X32 FILLER_235_1 ();
 FILLCELL_X32 FILLER_235_33 ();
 FILLCELL_X32 FILLER_235_65 ();
 FILLCELL_X32 FILLER_235_97 ();
 FILLCELL_X32 FILLER_235_129 ();
 FILLCELL_X32 FILLER_235_161 ();
 FILLCELL_X32 FILLER_235_193 ();
 FILLCELL_X32 FILLER_235_225 ();
 FILLCELL_X32 FILLER_235_257 ();
 FILLCELL_X32 FILLER_235_289 ();
 FILLCELL_X32 FILLER_235_321 ();
 FILLCELL_X32 FILLER_235_353 ();
 FILLCELL_X32 FILLER_235_385 ();
 FILLCELL_X32 FILLER_235_417 ();
 FILLCELL_X32 FILLER_235_449 ();
 FILLCELL_X32 FILLER_235_481 ();
 FILLCELL_X32 FILLER_235_513 ();
 FILLCELL_X32 FILLER_235_545 ();
 FILLCELL_X32 FILLER_235_577 ();
 FILLCELL_X32 FILLER_235_609 ();
 FILLCELL_X32 FILLER_235_641 ();
 FILLCELL_X32 FILLER_235_673 ();
 FILLCELL_X32 FILLER_235_705 ();
 FILLCELL_X32 FILLER_235_737 ();
 FILLCELL_X32 FILLER_235_769 ();
 FILLCELL_X32 FILLER_235_801 ();
 FILLCELL_X32 FILLER_235_833 ();
 FILLCELL_X32 FILLER_235_865 ();
 FILLCELL_X32 FILLER_235_897 ();
 FILLCELL_X32 FILLER_235_929 ();
 FILLCELL_X32 FILLER_235_961 ();
 FILLCELL_X32 FILLER_235_993 ();
 FILLCELL_X32 FILLER_235_1025 ();
 FILLCELL_X32 FILLER_235_1057 ();
 FILLCELL_X32 FILLER_235_1089 ();
 FILLCELL_X32 FILLER_235_1121 ();
 FILLCELL_X32 FILLER_235_1153 ();
 FILLCELL_X32 FILLER_235_1185 ();
 FILLCELL_X32 FILLER_235_1217 ();
 FILLCELL_X8 FILLER_235_1249 ();
 FILLCELL_X4 FILLER_235_1257 ();
 FILLCELL_X2 FILLER_235_1261 ();
 FILLCELL_X32 FILLER_235_1264 ();
 FILLCELL_X32 FILLER_235_1296 ();
 FILLCELL_X32 FILLER_235_1328 ();
 FILLCELL_X32 FILLER_235_1360 ();
 FILLCELL_X32 FILLER_235_1392 ();
 FILLCELL_X32 FILLER_235_1424 ();
 FILLCELL_X32 FILLER_235_1456 ();
 FILLCELL_X32 FILLER_235_1488 ();
 FILLCELL_X32 FILLER_235_1520 ();
 FILLCELL_X32 FILLER_235_1552 ();
 FILLCELL_X32 FILLER_235_1584 ();
 FILLCELL_X32 FILLER_235_1616 ();
 FILLCELL_X32 FILLER_235_1648 ();
 FILLCELL_X32 FILLER_235_1680 ();
 FILLCELL_X32 FILLER_235_1712 ();
 FILLCELL_X32 FILLER_235_1744 ();
 FILLCELL_X32 FILLER_235_1776 ();
 FILLCELL_X32 FILLER_235_1808 ();
 FILLCELL_X32 FILLER_235_1840 ();
 FILLCELL_X32 FILLER_235_1872 ();
 FILLCELL_X32 FILLER_235_1904 ();
 FILLCELL_X32 FILLER_235_1936 ();
 FILLCELL_X32 FILLER_235_1968 ();
 FILLCELL_X32 FILLER_235_2000 ();
 FILLCELL_X32 FILLER_235_2032 ();
 FILLCELL_X32 FILLER_235_2064 ();
 FILLCELL_X32 FILLER_235_2096 ();
 FILLCELL_X32 FILLER_235_2128 ();
 FILLCELL_X32 FILLER_235_2160 ();
 FILLCELL_X32 FILLER_235_2192 ();
 FILLCELL_X32 FILLER_235_2224 ();
 FILLCELL_X32 FILLER_235_2256 ();
 FILLCELL_X32 FILLER_235_2288 ();
 FILLCELL_X32 FILLER_235_2320 ();
 FILLCELL_X32 FILLER_235_2352 ();
 FILLCELL_X32 FILLER_235_2384 ();
 FILLCELL_X32 FILLER_235_2416 ();
 FILLCELL_X32 FILLER_235_2448 ();
 FILLCELL_X32 FILLER_235_2480 ();
 FILLCELL_X8 FILLER_235_2512 ();
 FILLCELL_X4 FILLER_235_2520 ();
 FILLCELL_X2 FILLER_235_2524 ();
 FILLCELL_X32 FILLER_235_2527 ();
 FILLCELL_X32 FILLER_235_2559 ();
 FILLCELL_X8 FILLER_235_2591 ();
 FILLCELL_X2 FILLER_235_2599 ();
 FILLCELL_X1 FILLER_235_2601 ();
 FILLCELL_X32 FILLER_236_1 ();
 FILLCELL_X32 FILLER_236_33 ();
 FILLCELL_X32 FILLER_236_65 ();
 FILLCELL_X32 FILLER_236_97 ();
 FILLCELL_X32 FILLER_236_129 ();
 FILLCELL_X32 FILLER_236_161 ();
 FILLCELL_X32 FILLER_236_193 ();
 FILLCELL_X32 FILLER_236_225 ();
 FILLCELL_X32 FILLER_236_257 ();
 FILLCELL_X32 FILLER_236_289 ();
 FILLCELL_X32 FILLER_236_321 ();
 FILLCELL_X32 FILLER_236_353 ();
 FILLCELL_X32 FILLER_236_385 ();
 FILLCELL_X32 FILLER_236_417 ();
 FILLCELL_X32 FILLER_236_449 ();
 FILLCELL_X32 FILLER_236_481 ();
 FILLCELL_X32 FILLER_236_513 ();
 FILLCELL_X32 FILLER_236_545 ();
 FILLCELL_X32 FILLER_236_577 ();
 FILLCELL_X16 FILLER_236_609 ();
 FILLCELL_X4 FILLER_236_625 ();
 FILLCELL_X2 FILLER_236_629 ();
 FILLCELL_X32 FILLER_236_632 ();
 FILLCELL_X32 FILLER_236_664 ();
 FILLCELL_X32 FILLER_236_696 ();
 FILLCELL_X32 FILLER_236_728 ();
 FILLCELL_X32 FILLER_236_760 ();
 FILLCELL_X32 FILLER_236_792 ();
 FILLCELL_X32 FILLER_236_824 ();
 FILLCELL_X32 FILLER_236_856 ();
 FILLCELL_X32 FILLER_236_888 ();
 FILLCELL_X32 FILLER_236_920 ();
 FILLCELL_X32 FILLER_236_952 ();
 FILLCELL_X32 FILLER_236_984 ();
 FILLCELL_X32 FILLER_236_1016 ();
 FILLCELL_X32 FILLER_236_1048 ();
 FILLCELL_X32 FILLER_236_1080 ();
 FILLCELL_X32 FILLER_236_1112 ();
 FILLCELL_X32 FILLER_236_1144 ();
 FILLCELL_X32 FILLER_236_1176 ();
 FILLCELL_X32 FILLER_236_1208 ();
 FILLCELL_X32 FILLER_236_1240 ();
 FILLCELL_X32 FILLER_236_1272 ();
 FILLCELL_X32 FILLER_236_1304 ();
 FILLCELL_X32 FILLER_236_1336 ();
 FILLCELL_X32 FILLER_236_1368 ();
 FILLCELL_X32 FILLER_236_1400 ();
 FILLCELL_X32 FILLER_236_1432 ();
 FILLCELL_X32 FILLER_236_1464 ();
 FILLCELL_X32 FILLER_236_1496 ();
 FILLCELL_X32 FILLER_236_1528 ();
 FILLCELL_X32 FILLER_236_1560 ();
 FILLCELL_X32 FILLER_236_1592 ();
 FILLCELL_X32 FILLER_236_1624 ();
 FILLCELL_X32 FILLER_236_1656 ();
 FILLCELL_X32 FILLER_236_1688 ();
 FILLCELL_X32 FILLER_236_1720 ();
 FILLCELL_X32 FILLER_236_1752 ();
 FILLCELL_X32 FILLER_236_1784 ();
 FILLCELL_X32 FILLER_236_1816 ();
 FILLCELL_X32 FILLER_236_1848 ();
 FILLCELL_X8 FILLER_236_1880 ();
 FILLCELL_X4 FILLER_236_1888 ();
 FILLCELL_X2 FILLER_236_1892 ();
 FILLCELL_X32 FILLER_236_1895 ();
 FILLCELL_X32 FILLER_236_1927 ();
 FILLCELL_X32 FILLER_236_1959 ();
 FILLCELL_X32 FILLER_236_1991 ();
 FILLCELL_X32 FILLER_236_2023 ();
 FILLCELL_X32 FILLER_236_2055 ();
 FILLCELL_X32 FILLER_236_2087 ();
 FILLCELL_X32 FILLER_236_2119 ();
 FILLCELL_X32 FILLER_236_2151 ();
 FILLCELL_X32 FILLER_236_2183 ();
 FILLCELL_X32 FILLER_236_2215 ();
 FILLCELL_X32 FILLER_236_2247 ();
 FILLCELL_X32 FILLER_236_2279 ();
 FILLCELL_X32 FILLER_236_2311 ();
 FILLCELL_X32 FILLER_236_2343 ();
 FILLCELL_X32 FILLER_236_2375 ();
 FILLCELL_X32 FILLER_236_2407 ();
 FILLCELL_X32 FILLER_236_2439 ();
 FILLCELL_X32 FILLER_236_2471 ();
 FILLCELL_X32 FILLER_236_2503 ();
 FILLCELL_X32 FILLER_236_2535 ();
 FILLCELL_X32 FILLER_236_2567 ();
 FILLCELL_X2 FILLER_236_2599 ();
 FILLCELL_X1 FILLER_236_2601 ();
 FILLCELL_X32 FILLER_237_1 ();
 FILLCELL_X32 FILLER_237_33 ();
 FILLCELL_X32 FILLER_237_65 ();
 FILLCELL_X32 FILLER_237_97 ();
 FILLCELL_X32 FILLER_237_129 ();
 FILLCELL_X32 FILLER_237_161 ();
 FILLCELL_X32 FILLER_237_193 ();
 FILLCELL_X32 FILLER_237_225 ();
 FILLCELL_X32 FILLER_237_257 ();
 FILLCELL_X32 FILLER_237_289 ();
 FILLCELL_X32 FILLER_237_321 ();
 FILLCELL_X32 FILLER_237_353 ();
 FILLCELL_X32 FILLER_237_385 ();
 FILLCELL_X32 FILLER_237_417 ();
 FILLCELL_X32 FILLER_237_449 ();
 FILLCELL_X32 FILLER_237_481 ();
 FILLCELL_X32 FILLER_237_513 ();
 FILLCELL_X32 FILLER_237_545 ();
 FILLCELL_X32 FILLER_237_577 ();
 FILLCELL_X32 FILLER_237_609 ();
 FILLCELL_X32 FILLER_237_641 ();
 FILLCELL_X32 FILLER_237_673 ();
 FILLCELL_X32 FILLER_237_705 ();
 FILLCELL_X32 FILLER_237_737 ();
 FILLCELL_X32 FILLER_237_769 ();
 FILLCELL_X32 FILLER_237_801 ();
 FILLCELL_X32 FILLER_237_833 ();
 FILLCELL_X32 FILLER_237_865 ();
 FILLCELL_X32 FILLER_237_897 ();
 FILLCELL_X32 FILLER_237_929 ();
 FILLCELL_X32 FILLER_237_961 ();
 FILLCELL_X32 FILLER_237_993 ();
 FILLCELL_X32 FILLER_237_1025 ();
 FILLCELL_X32 FILLER_237_1057 ();
 FILLCELL_X32 FILLER_237_1089 ();
 FILLCELL_X32 FILLER_237_1121 ();
 FILLCELL_X32 FILLER_237_1153 ();
 FILLCELL_X32 FILLER_237_1185 ();
 FILLCELL_X32 FILLER_237_1217 ();
 FILLCELL_X8 FILLER_237_1249 ();
 FILLCELL_X4 FILLER_237_1257 ();
 FILLCELL_X2 FILLER_237_1261 ();
 FILLCELL_X32 FILLER_237_1264 ();
 FILLCELL_X32 FILLER_237_1296 ();
 FILLCELL_X32 FILLER_237_1328 ();
 FILLCELL_X32 FILLER_237_1360 ();
 FILLCELL_X32 FILLER_237_1392 ();
 FILLCELL_X32 FILLER_237_1424 ();
 FILLCELL_X32 FILLER_237_1456 ();
 FILLCELL_X32 FILLER_237_1488 ();
 FILLCELL_X32 FILLER_237_1520 ();
 FILLCELL_X32 FILLER_237_1552 ();
 FILLCELL_X32 FILLER_237_1584 ();
 FILLCELL_X32 FILLER_237_1616 ();
 FILLCELL_X32 FILLER_237_1648 ();
 FILLCELL_X32 FILLER_237_1680 ();
 FILLCELL_X32 FILLER_237_1712 ();
 FILLCELL_X32 FILLER_237_1744 ();
 FILLCELL_X32 FILLER_237_1776 ();
 FILLCELL_X32 FILLER_237_1808 ();
 FILLCELL_X32 FILLER_237_1840 ();
 FILLCELL_X32 FILLER_237_1872 ();
 FILLCELL_X32 FILLER_237_1904 ();
 FILLCELL_X32 FILLER_237_1936 ();
 FILLCELL_X32 FILLER_237_1968 ();
 FILLCELL_X32 FILLER_237_2000 ();
 FILLCELL_X32 FILLER_237_2032 ();
 FILLCELL_X32 FILLER_237_2064 ();
 FILLCELL_X32 FILLER_237_2096 ();
 FILLCELL_X32 FILLER_237_2128 ();
 FILLCELL_X32 FILLER_237_2160 ();
 FILLCELL_X32 FILLER_237_2192 ();
 FILLCELL_X32 FILLER_237_2224 ();
 FILLCELL_X32 FILLER_237_2256 ();
 FILLCELL_X32 FILLER_237_2288 ();
 FILLCELL_X32 FILLER_237_2320 ();
 FILLCELL_X32 FILLER_237_2352 ();
 FILLCELL_X32 FILLER_237_2384 ();
 FILLCELL_X32 FILLER_237_2416 ();
 FILLCELL_X32 FILLER_237_2448 ();
 FILLCELL_X32 FILLER_237_2480 ();
 FILLCELL_X8 FILLER_237_2512 ();
 FILLCELL_X4 FILLER_237_2520 ();
 FILLCELL_X2 FILLER_237_2524 ();
 FILLCELL_X32 FILLER_237_2527 ();
 FILLCELL_X32 FILLER_237_2559 ();
 FILLCELL_X8 FILLER_237_2591 ();
 FILLCELL_X2 FILLER_237_2599 ();
 FILLCELL_X1 FILLER_237_2601 ();
 FILLCELL_X32 FILLER_238_1 ();
 FILLCELL_X32 FILLER_238_33 ();
 FILLCELL_X32 FILLER_238_65 ();
 FILLCELL_X32 FILLER_238_97 ();
 FILLCELL_X32 FILLER_238_129 ();
 FILLCELL_X32 FILLER_238_161 ();
 FILLCELL_X32 FILLER_238_193 ();
 FILLCELL_X32 FILLER_238_225 ();
 FILLCELL_X32 FILLER_238_257 ();
 FILLCELL_X32 FILLER_238_289 ();
 FILLCELL_X32 FILLER_238_321 ();
 FILLCELL_X32 FILLER_238_353 ();
 FILLCELL_X32 FILLER_238_385 ();
 FILLCELL_X32 FILLER_238_417 ();
 FILLCELL_X32 FILLER_238_449 ();
 FILLCELL_X32 FILLER_238_481 ();
 FILLCELL_X32 FILLER_238_513 ();
 FILLCELL_X32 FILLER_238_545 ();
 FILLCELL_X32 FILLER_238_577 ();
 FILLCELL_X16 FILLER_238_609 ();
 FILLCELL_X4 FILLER_238_625 ();
 FILLCELL_X2 FILLER_238_629 ();
 FILLCELL_X32 FILLER_238_632 ();
 FILLCELL_X32 FILLER_238_664 ();
 FILLCELL_X32 FILLER_238_696 ();
 FILLCELL_X32 FILLER_238_728 ();
 FILLCELL_X32 FILLER_238_760 ();
 FILLCELL_X32 FILLER_238_792 ();
 FILLCELL_X32 FILLER_238_824 ();
 FILLCELL_X32 FILLER_238_856 ();
 FILLCELL_X32 FILLER_238_888 ();
 FILLCELL_X32 FILLER_238_920 ();
 FILLCELL_X32 FILLER_238_952 ();
 FILLCELL_X32 FILLER_238_984 ();
 FILLCELL_X32 FILLER_238_1016 ();
 FILLCELL_X32 FILLER_238_1048 ();
 FILLCELL_X32 FILLER_238_1080 ();
 FILLCELL_X32 FILLER_238_1112 ();
 FILLCELL_X32 FILLER_238_1144 ();
 FILLCELL_X32 FILLER_238_1176 ();
 FILLCELL_X32 FILLER_238_1208 ();
 FILLCELL_X32 FILLER_238_1240 ();
 FILLCELL_X32 FILLER_238_1272 ();
 FILLCELL_X32 FILLER_238_1304 ();
 FILLCELL_X32 FILLER_238_1336 ();
 FILLCELL_X32 FILLER_238_1368 ();
 FILLCELL_X32 FILLER_238_1400 ();
 FILLCELL_X32 FILLER_238_1432 ();
 FILLCELL_X32 FILLER_238_1464 ();
 FILLCELL_X32 FILLER_238_1496 ();
 FILLCELL_X32 FILLER_238_1528 ();
 FILLCELL_X32 FILLER_238_1560 ();
 FILLCELL_X32 FILLER_238_1592 ();
 FILLCELL_X32 FILLER_238_1624 ();
 FILLCELL_X32 FILLER_238_1656 ();
 FILLCELL_X32 FILLER_238_1688 ();
 FILLCELL_X32 FILLER_238_1720 ();
 FILLCELL_X32 FILLER_238_1752 ();
 FILLCELL_X32 FILLER_238_1784 ();
 FILLCELL_X32 FILLER_238_1816 ();
 FILLCELL_X32 FILLER_238_1848 ();
 FILLCELL_X8 FILLER_238_1880 ();
 FILLCELL_X4 FILLER_238_1888 ();
 FILLCELL_X2 FILLER_238_1892 ();
 FILLCELL_X32 FILLER_238_1895 ();
 FILLCELL_X32 FILLER_238_1927 ();
 FILLCELL_X32 FILLER_238_1959 ();
 FILLCELL_X32 FILLER_238_1991 ();
 FILLCELL_X32 FILLER_238_2023 ();
 FILLCELL_X32 FILLER_238_2055 ();
 FILLCELL_X32 FILLER_238_2087 ();
 FILLCELL_X32 FILLER_238_2119 ();
 FILLCELL_X32 FILLER_238_2151 ();
 FILLCELL_X32 FILLER_238_2183 ();
 FILLCELL_X32 FILLER_238_2215 ();
 FILLCELL_X32 FILLER_238_2247 ();
 FILLCELL_X32 FILLER_238_2279 ();
 FILLCELL_X32 FILLER_238_2311 ();
 FILLCELL_X32 FILLER_238_2343 ();
 FILLCELL_X32 FILLER_238_2375 ();
 FILLCELL_X32 FILLER_238_2407 ();
 FILLCELL_X32 FILLER_238_2439 ();
 FILLCELL_X32 FILLER_238_2471 ();
 FILLCELL_X32 FILLER_238_2503 ();
 FILLCELL_X32 FILLER_238_2535 ();
 FILLCELL_X32 FILLER_238_2567 ();
 FILLCELL_X2 FILLER_238_2599 ();
 FILLCELL_X1 FILLER_238_2601 ();
 FILLCELL_X32 FILLER_239_1 ();
 FILLCELL_X32 FILLER_239_33 ();
 FILLCELL_X32 FILLER_239_65 ();
 FILLCELL_X32 FILLER_239_97 ();
 FILLCELL_X32 FILLER_239_129 ();
 FILLCELL_X32 FILLER_239_161 ();
 FILLCELL_X32 FILLER_239_193 ();
 FILLCELL_X32 FILLER_239_225 ();
 FILLCELL_X32 FILLER_239_257 ();
 FILLCELL_X32 FILLER_239_289 ();
 FILLCELL_X32 FILLER_239_321 ();
 FILLCELL_X32 FILLER_239_353 ();
 FILLCELL_X32 FILLER_239_385 ();
 FILLCELL_X32 FILLER_239_417 ();
 FILLCELL_X32 FILLER_239_449 ();
 FILLCELL_X32 FILLER_239_481 ();
 FILLCELL_X32 FILLER_239_513 ();
 FILLCELL_X32 FILLER_239_545 ();
 FILLCELL_X32 FILLER_239_577 ();
 FILLCELL_X32 FILLER_239_609 ();
 FILLCELL_X32 FILLER_239_641 ();
 FILLCELL_X32 FILLER_239_673 ();
 FILLCELL_X32 FILLER_239_705 ();
 FILLCELL_X32 FILLER_239_737 ();
 FILLCELL_X32 FILLER_239_769 ();
 FILLCELL_X32 FILLER_239_801 ();
 FILLCELL_X32 FILLER_239_833 ();
 FILLCELL_X32 FILLER_239_865 ();
 FILLCELL_X32 FILLER_239_897 ();
 FILLCELL_X32 FILLER_239_929 ();
 FILLCELL_X32 FILLER_239_961 ();
 FILLCELL_X32 FILLER_239_993 ();
 FILLCELL_X32 FILLER_239_1025 ();
 FILLCELL_X32 FILLER_239_1057 ();
 FILLCELL_X32 FILLER_239_1089 ();
 FILLCELL_X32 FILLER_239_1121 ();
 FILLCELL_X32 FILLER_239_1153 ();
 FILLCELL_X32 FILLER_239_1185 ();
 FILLCELL_X32 FILLER_239_1217 ();
 FILLCELL_X8 FILLER_239_1249 ();
 FILLCELL_X4 FILLER_239_1257 ();
 FILLCELL_X2 FILLER_239_1261 ();
 FILLCELL_X32 FILLER_239_1264 ();
 FILLCELL_X32 FILLER_239_1296 ();
 FILLCELL_X32 FILLER_239_1328 ();
 FILLCELL_X32 FILLER_239_1360 ();
 FILLCELL_X32 FILLER_239_1392 ();
 FILLCELL_X32 FILLER_239_1424 ();
 FILLCELL_X32 FILLER_239_1456 ();
 FILLCELL_X32 FILLER_239_1488 ();
 FILLCELL_X32 FILLER_239_1520 ();
 FILLCELL_X32 FILLER_239_1552 ();
 FILLCELL_X32 FILLER_239_1584 ();
 FILLCELL_X32 FILLER_239_1616 ();
 FILLCELL_X32 FILLER_239_1648 ();
 FILLCELL_X32 FILLER_239_1680 ();
 FILLCELL_X32 FILLER_239_1712 ();
 FILLCELL_X32 FILLER_239_1744 ();
 FILLCELL_X32 FILLER_239_1776 ();
 FILLCELL_X32 FILLER_239_1808 ();
 FILLCELL_X32 FILLER_239_1840 ();
 FILLCELL_X32 FILLER_239_1872 ();
 FILLCELL_X32 FILLER_239_1904 ();
 FILLCELL_X32 FILLER_239_1936 ();
 FILLCELL_X32 FILLER_239_1968 ();
 FILLCELL_X32 FILLER_239_2000 ();
 FILLCELL_X32 FILLER_239_2032 ();
 FILLCELL_X32 FILLER_239_2064 ();
 FILLCELL_X32 FILLER_239_2096 ();
 FILLCELL_X32 FILLER_239_2128 ();
 FILLCELL_X32 FILLER_239_2160 ();
 FILLCELL_X32 FILLER_239_2192 ();
 FILLCELL_X32 FILLER_239_2224 ();
 FILLCELL_X32 FILLER_239_2256 ();
 FILLCELL_X32 FILLER_239_2288 ();
 FILLCELL_X32 FILLER_239_2320 ();
 FILLCELL_X32 FILLER_239_2352 ();
 FILLCELL_X32 FILLER_239_2384 ();
 FILLCELL_X32 FILLER_239_2416 ();
 FILLCELL_X32 FILLER_239_2448 ();
 FILLCELL_X32 FILLER_239_2480 ();
 FILLCELL_X8 FILLER_239_2512 ();
 FILLCELL_X4 FILLER_239_2520 ();
 FILLCELL_X2 FILLER_239_2524 ();
 FILLCELL_X32 FILLER_239_2527 ();
 FILLCELL_X32 FILLER_239_2559 ();
 FILLCELL_X8 FILLER_239_2591 ();
 FILLCELL_X2 FILLER_239_2599 ();
 FILLCELL_X1 FILLER_239_2601 ();
 FILLCELL_X32 FILLER_240_1 ();
 FILLCELL_X32 FILLER_240_33 ();
 FILLCELL_X32 FILLER_240_65 ();
 FILLCELL_X32 FILLER_240_97 ();
 FILLCELL_X32 FILLER_240_129 ();
 FILLCELL_X32 FILLER_240_161 ();
 FILLCELL_X32 FILLER_240_193 ();
 FILLCELL_X32 FILLER_240_225 ();
 FILLCELL_X32 FILLER_240_257 ();
 FILLCELL_X32 FILLER_240_289 ();
 FILLCELL_X32 FILLER_240_321 ();
 FILLCELL_X32 FILLER_240_353 ();
 FILLCELL_X32 FILLER_240_385 ();
 FILLCELL_X32 FILLER_240_417 ();
 FILLCELL_X32 FILLER_240_449 ();
 FILLCELL_X32 FILLER_240_481 ();
 FILLCELL_X32 FILLER_240_513 ();
 FILLCELL_X32 FILLER_240_545 ();
 FILLCELL_X32 FILLER_240_577 ();
 FILLCELL_X16 FILLER_240_609 ();
 FILLCELL_X4 FILLER_240_625 ();
 FILLCELL_X2 FILLER_240_629 ();
 FILLCELL_X32 FILLER_240_632 ();
 FILLCELL_X32 FILLER_240_664 ();
 FILLCELL_X32 FILLER_240_696 ();
 FILLCELL_X32 FILLER_240_728 ();
 FILLCELL_X32 FILLER_240_760 ();
 FILLCELL_X32 FILLER_240_792 ();
 FILLCELL_X32 FILLER_240_824 ();
 FILLCELL_X32 FILLER_240_856 ();
 FILLCELL_X32 FILLER_240_888 ();
 FILLCELL_X32 FILLER_240_920 ();
 FILLCELL_X32 FILLER_240_952 ();
 FILLCELL_X32 FILLER_240_984 ();
 FILLCELL_X32 FILLER_240_1016 ();
 FILLCELL_X32 FILLER_240_1048 ();
 FILLCELL_X32 FILLER_240_1080 ();
 FILLCELL_X32 FILLER_240_1112 ();
 FILLCELL_X32 FILLER_240_1144 ();
 FILLCELL_X32 FILLER_240_1176 ();
 FILLCELL_X32 FILLER_240_1208 ();
 FILLCELL_X32 FILLER_240_1240 ();
 FILLCELL_X32 FILLER_240_1272 ();
 FILLCELL_X32 FILLER_240_1304 ();
 FILLCELL_X32 FILLER_240_1336 ();
 FILLCELL_X32 FILLER_240_1368 ();
 FILLCELL_X32 FILLER_240_1400 ();
 FILLCELL_X32 FILLER_240_1432 ();
 FILLCELL_X32 FILLER_240_1464 ();
 FILLCELL_X32 FILLER_240_1496 ();
 FILLCELL_X32 FILLER_240_1528 ();
 FILLCELL_X32 FILLER_240_1560 ();
 FILLCELL_X32 FILLER_240_1592 ();
 FILLCELL_X32 FILLER_240_1624 ();
 FILLCELL_X32 FILLER_240_1656 ();
 FILLCELL_X32 FILLER_240_1688 ();
 FILLCELL_X32 FILLER_240_1720 ();
 FILLCELL_X32 FILLER_240_1752 ();
 FILLCELL_X32 FILLER_240_1784 ();
 FILLCELL_X32 FILLER_240_1816 ();
 FILLCELL_X32 FILLER_240_1848 ();
 FILLCELL_X8 FILLER_240_1880 ();
 FILLCELL_X4 FILLER_240_1888 ();
 FILLCELL_X2 FILLER_240_1892 ();
 FILLCELL_X32 FILLER_240_1895 ();
 FILLCELL_X32 FILLER_240_1927 ();
 FILLCELL_X32 FILLER_240_1959 ();
 FILLCELL_X32 FILLER_240_1991 ();
 FILLCELL_X32 FILLER_240_2023 ();
 FILLCELL_X32 FILLER_240_2055 ();
 FILLCELL_X32 FILLER_240_2087 ();
 FILLCELL_X32 FILLER_240_2119 ();
 FILLCELL_X32 FILLER_240_2151 ();
 FILLCELL_X32 FILLER_240_2183 ();
 FILLCELL_X32 FILLER_240_2215 ();
 FILLCELL_X32 FILLER_240_2247 ();
 FILLCELL_X32 FILLER_240_2279 ();
 FILLCELL_X32 FILLER_240_2311 ();
 FILLCELL_X32 FILLER_240_2343 ();
 FILLCELL_X32 FILLER_240_2375 ();
 FILLCELL_X32 FILLER_240_2407 ();
 FILLCELL_X32 FILLER_240_2439 ();
 FILLCELL_X32 FILLER_240_2471 ();
 FILLCELL_X32 FILLER_240_2503 ();
 FILLCELL_X32 FILLER_240_2535 ();
 FILLCELL_X32 FILLER_240_2567 ();
 FILLCELL_X2 FILLER_240_2599 ();
 FILLCELL_X1 FILLER_240_2601 ();
 FILLCELL_X32 FILLER_241_1 ();
 FILLCELL_X32 FILLER_241_33 ();
 FILLCELL_X32 FILLER_241_65 ();
 FILLCELL_X32 FILLER_241_97 ();
 FILLCELL_X32 FILLER_241_129 ();
 FILLCELL_X32 FILLER_241_161 ();
 FILLCELL_X32 FILLER_241_193 ();
 FILLCELL_X32 FILLER_241_225 ();
 FILLCELL_X32 FILLER_241_257 ();
 FILLCELL_X32 FILLER_241_289 ();
 FILLCELL_X32 FILLER_241_321 ();
 FILLCELL_X32 FILLER_241_353 ();
 FILLCELL_X32 FILLER_241_385 ();
 FILLCELL_X32 FILLER_241_417 ();
 FILLCELL_X32 FILLER_241_449 ();
 FILLCELL_X32 FILLER_241_481 ();
 FILLCELL_X32 FILLER_241_513 ();
 FILLCELL_X32 FILLER_241_545 ();
 FILLCELL_X32 FILLER_241_577 ();
 FILLCELL_X32 FILLER_241_609 ();
 FILLCELL_X32 FILLER_241_641 ();
 FILLCELL_X32 FILLER_241_673 ();
 FILLCELL_X32 FILLER_241_705 ();
 FILLCELL_X32 FILLER_241_737 ();
 FILLCELL_X32 FILLER_241_769 ();
 FILLCELL_X32 FILLER_241_801 ();
 FILLCELL_X32 FILLER_241_833 ();
 FILLCELL_X32 FILLER_241_865 ();
 FILLCELL_X32 FILLER_241_897 ();
 FILLCELL_X32 FILLER_241_929 ();
 FILLCELL_X32 FILLER_241_961 ();
 FILLCELL_X32 FILLER_241_993 ();
 FILLCELL_X32 FILLER_241_1025 ();
 FILLCELL_X32 FILLER_241_1057 ();
 FILLCELL_X32 FILLER_241_1089 ();
 FILLCELL_X32 FILLER_241_1121 ();
 FILLCELL_X32 FILLER_241_1153 ();
 FILLCELL_X32 FILLER_241_1185 ();
 FILLCELL_X32 FILLER_241_1217 ();
 FILLCELL_X8 FILLER_241_1249 ();
 FILLCELL_X4 FILLER_241_1257 ();
 FILLCELL_X2 FILLER_241_1261 ();
 FILLCELL_X32 FILLER_241_1264 ();
 FILLCELL_X32 FILLER_241_1296 ();
 FILLCELL_X32 FILLER_241_1328 ();
 FILLCELL_X32 FILLER_241_1360 ();
 FILLCELL_X32 FILLER_241_1392 ();
 FILLCELL_X32 FILLER_241_1424 ();
 FILLCELL_X32 FILLER_241_1456 ();
 FILLCELL_X32 FILLER_241_1488 ();
 FILLCELL_X32 FILLER_241_1520 ();
 FILLCELL_X32 FILLER_241_1552 ();
 FILLCELL_X32 FILLER_241_1584 ();
 FILLCELL_X32 FILLER_241_1616 ();
 FILLCELL_X32 FILLER_241_1648 ();
 FILLCELL_X32 FILLER_241_1680 ();
 FILLCELL_X32 FILLER_241_1712 ();
 FILLCELL_X32 FILLER_241_1744 ();
 FILLCELL_X32 FILLER_241_1776 ();
 FILLCELL_X32 FILLER_241_1808 ();
 FILLCELL_X32 FILLER_241_1840 ();
 FILLCELL_X32 FILLER_241_1872 ();
 FILLCELL_X32 FILLER_241_1904 ();
 FILLCELL_X32 FILLER_241_1936 ();
 FILLCELL_X32 FILLER_241_1968 ();
 FILLCELL_X32 FILLER_241_2000 ();
 FILLCELL_X32 FILLER_241_2032 ();
 FILLCELL_X32 FILLER_241_2064 ();
 FILLCELL_X32 FILLER_241_2096 ();
 FILLCELL_X32 FILLER_241_2128 ();
 FILLCELL_X32 FILLER_241_2160 ();
 FILLCELL_X32 FILLER_241_2192 ();
 FILLCELL_X32 FILLER_241_2224 ();
 FILLCELL_X32 FILLER_241_2256 ();
 FILLCELL_X32 FILLER_241_2288 ();
 FILLCELL_X32 FILLER_241_2320 ();
 FILLCELL_X32 FILLER_241_2352 ();
 FILLCELL_X32 FILLER_241_2384 ();
 FILLCELL_X32 FILLER_241_2416 ();
 FILLCELL_X32 FILLER_241_2448 ();
 FILLCELL_X32 FILLER_241_2480 ();
 FILLCELL_X8 FILLER_241_2512 ();
 FILLCELL_X4 FILLER_241_2520 ();
 FILLCELL_X2 FILLER_241_2524 ();
 FILLCELL_X32 FILLER_241_2527 ();
 FILLCELL_X32 FILLER_241_2559 ();
 FILLCELL_X8 FILLER_241_2591 ();
 FILLCELL_X2 FILLER_241_2599 ();
 FILLCELL_X1 FILLER_241_2601 ();
 FILLCELL_X32 FILLER_242_1 ();
 FILLCELL_X32 FILLER_242_33 ();
 FILLCELL_X32 FILLER_242_65 ();
 FILLCELL_X32 FILLER_242_97 ();
 FILLCELL_X32 FILLER_242_129 ();
 FILLCELL_X32 FILLER_242_161 ();
 FILLCELL_X32 FILLER_242_193 ();
 FILLCELL_X32 FILLER_242_225 ();
 FILLCELL_X32 FILLER_242_257 ();
 FILLCELL_X32 FILLER_242_289 ();
 FILLCELL_X32 FILLER_242_321 ();
 FILLCELL_X32 FILLER_242_353 ();
 FILLCELL_X32 FILLER_242_385 ();
 FILLCELL_X32 FILLER_242_417 ();
 FILLCELL_X32 FILLER_242_449 ();
 FILLCELL_X32 FILLER_242_481 ();
 FILLCELL_X32 FILLER_242_513 ();
 FILLCELL_X32 FILLER_242_545 ();
 FILLCELL_X32 FILLER_242_577 ();
 FILLCELL_X16 FILLER_242_609 ();
 FILLCELL_X4 FILLER_242_625 ();
 FILLCELL_X2 FILLER_242_629 ();
 FILLCELL_X32 FILLER_242_632 ();
 FILLCELL_X32 FILLER_242_664 ();
 FILLCELL_X32 FILLER_242_696 ();
 FILLCELL_X32 FILLER_242_728 ();
 FILLCELL_X32 FILLER_242_760 ();
 FILLCELL_X32 FILLER_242_792 ();
 FILLCELL_X32 FILLER_242_824 ();
 FILLCELL_X32 FILLER_242_856 ();
 FILLCELL_X32 FILLER_242_888 ();
 FILLCELL_X32 FILLER_242_920 ();
 FILLCELL_X32 FILLER_242_952 ();
 FILLCELL_X32 FILLER_242_984 ();
 FILLCELL_X32 FILLER_242_1016 ();
 FILLCELL_X32 FILLER_242_1048 ();
 FILLCELL_X32 FILLER_242_1080 ();
 FILLCELL_X32 FILLER_242_1112 ();
 FILLCELL_X32 FILLER_242_1144 ();
 FILLCELL_X32 FILLER_242_1176 ();
 FILLCELL_X32 FILLER_242_1208 ();
 FILLCELL_X32 FILLER_242_1240 ();
 FILLCELL_X32 FILLER_242_1272 ();
 FILLCELL_X32 FILLER_242_1304 ();
 FILLCELL_X32 FILLER_242_1336 ();
 FILLCELL_X32 FILLER_242_1368 ();
 FILLCELL_X32 FILLER_242_1400 ();
 FILLCELL_X32 FILLER_242_1432 ();
 FILLCELL_X32 FILLER_242_1464 ();
 FILLCELL_X32 FILLER_242_1496 ();
 FILLCELL_X32 FILLER_242_1528 ();
 FILLCELL_X32 FILLER_242_1560 ();
 FILLCELL_X32 FILLER_242_1592 ();
 FILLCELL_X32 FILLER_242_1624 ();
 FILLCELL_X32 FILLER_242_1656 ();
 FILLCELL_X32 FILLER_242_1688 ();
 FILLCELL_X32 FILLER_242_1720 ();
 FILLCELL_X32 FILLER_242_1752 ();
 FILLCELL_X32 FILLER_242_1784 ();
 FILLCELL_X32 FILLER_242_1816 ();
 FILLCELL_X32 FILLER_242_1848 ();
 FILLCELL_X8 FILLER_242_1880 ();
 FILLCELL_X4 FILLER_242_1888 ();
 FILLCELL_X2 FILLER_242_1892 ();
 FILLCELL_X32 FILLER_242_1895 ();
 FILLCELL_X32 FILLER_242_1927 ();
 FILLCELL_X32 FILLER_242_1959 ();
 FILLCELL_X32 FILLER_242_1991 ();
 FILLCELL_X32 FILLER_242_2023 ();
 FILLCELL_X32 FILLER_242_2055 ();
 FILLCELL_X32 FILLER_242_2087 ();
 FILLCELL_X32 FILLER_242_2119 ();
 FILLCELL_X32 FILLER_242_2151 ();
 FILLCELL_X32 FILLER_242_2183 ();
 FILLCELL_X32 FILLER_242_2215 ();
 FILLCELL_X32 FILLER_242_2247 ();
 FILLCELL_X32 FILLER_242_2279 ();
 FILLCELL_X32 FILLER_242_2311 ();
 FILLCELL_X32 FILLER_242_2343 ();
 FILLCELL_X32 FILLER_242_2375 ();
 FILLCELL_X32 FILLER_242_2407 ();
 FILLCELL_X32 FILLER_242_2439 ();
 FILLCELL_X32 FILLER_242_2471 ();
 FILLCELL_X32 FILLER_242_2503 ();
 FILLCELL_X32 FILLER_242_2535 ();
 FILLCELL_X32 FILLER_242_2567 ();
 FILLCELL_X2 FILLER_242_2599 ();
 FILLCELL_X1 FILLER_242_2601 ();
 FILLCELL_X32 FILLER_243_1 ();
 FILLCELL_X32 FILLER_243_33 ();
 FILLCELL_X32 FILLER_243_65 ();
 FILLCELL_X32 FILLER_243_97 ();
 FILLCELL_X32 FILLER_243_129 ();
 FILLCELL_X32 FILLER_243_161 ();
 FILLCELL_X32 FILLER_243_193 ();
 FILLCELL_X32 FILLER_243_225 ();
 FILLCELL_X32 FILLER_243_257 ();
 FILLCELL_X32 FILLER_243_289 ();
 FILLCELL_X32 FILLER_243_321 ();
 FILLCELL_X32 FILLER_243_353 ();
 FILLCELL_X32 FILLER_243_385 ();
 FILLCELL_X32 FILLER_243_417 ();
 FILLCELL_X32 FILLER_243_449 ();
 FILLCELL_X32 FILLER_243_481 ();
 FILLCELL_X32 FILLER_243_513 ();
 FILLCELL_X32 FILLER_243_545 ();
 FILLCELL_X32 FILLER_243_577 ();
 FILLCELL_X32 FILLER_243_609 ();
 FILLCELL_X32 FILLER_243_641 ();
 FILLCELL_X32 FILLER_243_673 ();
 FILLCELL_X32 FILLER_243_705 ();
 FILLCELL_X32 FILLER_243_737 ();
 FILLCELL_X32 FILLER_243_769 ();
 FILLCELL_X32 FILLER_243_801 ();
 FILLCELL_X32 FILLER_243_833 ();
 FILLCELL_X32 FILLER_243_865 ();
 FILLCELL_X32 FILLER_243_897 ();
 FILLCELL_X32 FILLER_243_929 ();
 FILLCELL_X32 FILLER_243_961 ();
 FILLCELL_X32 FILLER_243_993 ();
 FILLCELL_X32 FILLER_243_1025 ();
 FILLCELL_X32 FILLER_243_1057 ();
 FILLCELL_X32 FILLER_243_1089 ();
 FILLCELL_X32 FILLER_243_1121 ();
 FILLCELL_X32 FILLER_243_1153 ();
 FILLCELL_X32 FILLER_243_1185 ();
 FILLCELL_X32 FILLER_243_1217 ();
 FILLCELL_X8 FILLER_243_1249 ();
 FILLCELL_X4 FILLER_243_1257 ();
 FILLCELL_X2 FILLER_243_1261 ();
 FILLCELL_X32 FILLER_243_1264 ();
 FILLCELL_X32 FILLER_243_1296 ();
 FILLCELL_X32 FILLER_243_1328 ();
 FILLCELL_X32 FILLER_243_1360 ();
 FILLCELL_X32 FILLER_243_1392 ();
 FILLCELL_X32 FILLER_243_1424 ();
 FILLCELL_X32 FILLER_243_1456 ();
 FILLCELL_X32 FILLER_243_1488 ();
 FILLCELL_X32 FILLER_243_1520 ();
 FILLCELL_X32 FILLER_243_1552 ();
 FILLCELL_X32 FILLER_243_1584 ();
 FILLCELL_X32 FILLER_243_1616 ();
 FILLCELL_X32 FILLER_243_1648 ();
 FILLCELL_X32 FILLER_243_1680 ();
 FILLCELL_X32 FILLER_243_1712 ();
 FILLCELL_X32 FILLER_243_1744 ();
 FILLCELL_X32 FILLER_243_1776 ();
 FILLCELL_X32 FILLER_243_1808 ();
 FILLCELL_X32 FILLER_243_1840 ();
 FILLCELL_X32 FILLER_243_1872 ();
 FILLCELL_X32 FILLER_243_1904 ();
 FILLCELL_X32 FILLER_243_1936 ();
 FILLCELL_X32 FILLER_243_1968 ();
 FILLCELL_X32 FILLER_243_2000 ();
 FILLCELL_X32 FILLER_243_2032 ();
 FILLCELL_X32 FILLER_243_2064 ();
 FILLCELL_X32 FILLER_243_2096 ();
 FILLCELL_X32 FILLER_243_2128 ();
 FILLCELL_X32 FILLER_243_2160 ();
 FILLCELL_X32 FILLER_243_2192 ();
 FILLCELL_X32 FILLER_243_2224 ();
 FILLCELL_X32 FILLER_243_2256 ();
 FILLCELL_X32 FILLER_243_2288 ();
 FILLCELL_X32 FILLER_243_2320 ();
 FILLCELL_X32 FILLER_243_2352 ();
 FILLCELL_X32 FILLER_243_2384 ();
 FILLCELL_X32 FILLER_243_2416 ();
 FILLCELL_X32 FILLER_243_2448 ();
 FILLCELL_X32 FILLER_243_2480 ();
 FILLCELL_X8 FILLER_243_2512 ();
 FILLCELL_X4 FILLER_243_2520 ();
 FILLCELL_X2 FILLER_243_2524 ();
 FILLCELL_X32 FILLER_243_2527 ();
 FILLCELL_X32 FILLER_243_2559 ();
 FILLCELL_X8 FILLER_243_2591 ();
 FILLCELL_X2 FILLER_243_2599 ();
 FILLCELL_X1 FILLER_243_2601 ();
 FILLCELL_X32 FILLER_244_1 ();
 FILLCELL_X32 FILLER_244_33 ();
 FILLCELL_X32 FILLER_244_65 ();
 FILLCELL_X32 FILLER_244_97 ();
 FILLCELL_X32 FILLER_244_129 ();
 FILLCELL_X32 FILLER_244_161 ();
 FILLCELL_X32 FILLER_244_193 ();
 FILLCELL_X32 FILLER_244_225 ();
 FILLCELL_X32 FILLER_244_257 ();
 FILLCELL_X32 FILLER_244_289 ();
 FILLCELL_X32 FILLER_244_321 ();
 FILLCELL_X32 FILLER_244_353 ();
 FILLCELL_X32 FILLER_244_385 ();
 FILLCELL_X32 FILLER_244_417 ();
 FILLCELL_X32 FILLER_244_449 ();
 FILLCELL_X32 FILLER_244_481 ();
 FILLCELL_X32 FILLER_244_513 ();
 FILLCELL_X32 FILLER_244_545 ();
 FILLCELL_X32 FILLER_244_577 ();
 FILLCELL_X16 FILLER_244_609 ();
 FILLCELL_X4 FILLER_244_625 ();
 FILLCELL_X2 FILLER_244_629 ();
 FILLCELL_X32 FILLER_244_632 ();
 FILLCELL_X32 FILLER_244_664 ();
 FILLCELL_X32 FILLER_244_696 ();
 FILLCELL_X32 FILLER_244_728 ();
 FILLCELL_X32 FILLER_244_760 ();
 FILLCELL_X32 FILLER_244_792 ();
 FILLCELL_X32 FILLER_244_824 ();
 FILLCELL_X32 FILLER_244_856 ();
 FILLCELL_X32 FILLER_244_888 ();
 FILLCELL_X32 FILLER_244_920 ();
 FILLCELL_X32 FILLER_244_952 ();
 FILLCELL_X32 FILLER_244_984 ();
 FILLCELL_X32 FILLER_244_1016 ();
 FILLCELL_X32 FILLER_244_1048 ();
 FILLCELL_X32 FILLER_244_1080 ();
 FILLCELL_X32 FILLER_244_1112 ();
 FILLCELL_X32 FILLER_244_1144 ();
 FILLCELL_X32 FILLER_244_1176 ();
 FILLCELL_X32 FILLER_244_1208 ();
 FILLCELL_X32 FILLER_244_1240 ();
 FILLCELL_X32 FILLER_244_1272 ();
 FILLCELL_X32 FILLER_244_1304 ();
 FILLCELL_X32 FILLER_244_1336 ();
 FILLCELL_X32 FILLER_244_1368 ();
 FILLCELL_X32 FILLER_244_1400 ();
 FILLCELL_X32 FILLER_244_1432 ();
 FILLCELL_X32 FILLER_244_1464 ();
 FILLCELL_X32 FILLER_244_1496 ();
 FILLCELL_X32 FILLER_244_1528 ();
 FILLCELL_X32 FILLER_244_1560 ();
 FILLCELL_X32 FILLER_244_1592 ();
 FILLCELL_X32 FILLER_244_1624 ();
 FILLCELL_X32 FILLER_244_1656 ();
 FILLCELL_X32 FILLER_244_1688 ();
 FILLCELL_X32 FILLER_244_1720 ();
 FILLCELL_X32 FILLER_244_1752 ();
 FILLCELL_X32 FILLER_244_1784 ();
 FILLCELL_X32 FILLER_244_1816 ();
 FILLCELL_X32 FILLER_244_1848 ();
 FILLCELL_X8 FILLER_244_1880 ();
 FILLCELL_X4 FILLER_244_1888 ();
 FILLCELL_X2 FILLER_244_1892 ();
 FILLCELL_X32 FILLER_244_1895 ();
 FILLCELL_X32 FILLER_244_1927 ();
 FILLCELL_X32 FILLER_244_1959 ();
 FILLCELL_X32 FILLER_244_1991 ();
 FILLCELL_X32 FILLER_244_2023 ();
 FILLCELL_X32 FILLER_244_2055 ();
 FILLCELL_X32 FILLER_244_2087 ();
 FILLCELL_X32 FILLER_244_2119 ();
 FILLCELL_X32 FILLER_244_2151 ();
 FILLCELL_X32 FILLER_244_2183 ();
 FILLCELL_X32 FILLER_244_2215 ();
 FILLCELL_X32 FILLER_244_2247 ();
 FILLCELL_X32 FILLER_244_2279 ();
 FILLCELL_X32 FILLER_244_2311 ();
 FILLCELL_X32 FILLER_244_2343 ();
 FILLCELL_X32 FILLER_244_2375 ();
 FILLCELL_X32 FILLER_244_2407 ();
 FILLCELL_X32 FILLER_244_2439 ();
 FILLCELL_X32 FILLER_244_2471 ();
 FILLCELL_X32 FILLER_244_2503 ();
 FILLCELL_X32 FILLER_244_2535 ();
 FILLCELL_X32 FILLER_244_2567 ();
 FILLCELL_X2 FILLER_244_2599 ();
 FILLCELL_X1 FILLER_244_2601 ();
 FILLCELL_X32 FILLER_245_1 ();
 FILLCELL_X32 FILLER_245_33 ();
 FILLCELL_X32 FILLER_245_65 ();
 FILLCELL_X32 FILLER_245_97 ();
 FILLCELL_X32 FILLER_245_129 ();
 FILLCELL_X32 FILLER_245_161 ();
 FILLCELL_X32 FILLER_245_193 ();
 FILLCELL_X32 FILLER_245_225 ();
 FILLCELL_X32 FILLER_245_257 ();
 FILLCELL_X32 FILLER_245_289 ();
 FILLCELL_X32 FILLER_245_321 ();
 FILLCELL_X32 FILLER_245_353 ();
 FILLCELL_X32 FILLER_245_385 ();
 FILLCELL_X32 FILLER_245_417 ();
 FILLCELL_X32 FILLER_245_449 ();
 FILLCELL_X32 FILLER_245_481 ();
 FILLCELL_X32 FILLER_245_513 ();
 FILLCELL_X32 FILLER_245_545 ();
 FILLCELL_X32 FILLER_245_577 ();
 FILLCELL_X32 FILLER_245_609 ();
 FILLCELL_X32 FILLER_245_641 ();
 FILLCELL_X32 FILLER_245_673 ();
 FILLCELL_X32 FILLER_245_705 ();
 FILLCELL_X32 FILLER_245_737 ();
 FILLCELL_X32 FILLER_245_769 ();
 FILLCELL_X32 FILLER_245_801 ();
 FILLCELL_X32 FILLER_245_833 ();
 FILLCELL_X32 FILLER_245_865 ();
 FILLCELL_X32 FILLER_245_897 ();
 FILLCELL_X32 FILLER_245_929 ();
 FILLCELL_X32 FILLER_245_961 ();
 FILLCELL_X32 FILLER_245_993 ();
 FILLCELL_X32 FILLER_245_1025 ();
 FILLCELL_X32 FILLER_245_1057 ();
 FILLCELL_X32 FILLER_245_1089 ();
 FILLCELL_X32 FILLER_245_1121 ();
 FILLCELL_X32 FILLER_245_1153 ();
 FILLCELL_X32 FILLER_245_1185 ();
 FILLCELL_X32 FILLER_245_1217 ();
 FILLCELL_X8 FILLER_245_1249 ();
 FILLCELL_X4 FILLER_245_1257 ();
 FILLCELL_X2 FILLER_245_1261 ();
 FILLCELL_X32 FILLER_245_1264 ();
 FILLCELL_X32 FILLER_245_1296 ();
 FILLCELL_X32 FILLER_245_1328 ();
 FILLCELL_X32 FILLER_245_1360 ();
 FILLCELL_X32 FILLER_245_1392 ();
 FILLCELL_X32 FILLER_245_1424 ();
 FILLCELL_X32 FILLER_245_1456 ();
 FILLCELL_X32 FILLER_245_1488 ();
 FILLCELL_X32 FILLER_245_1520 ();
 FILLCELL_X32 FILLER_245_1552 ();
 FILLCELL_X32 FILLER_245_1584 ();
 FILLCELL_X32 FILLER_245_1616 ();
 FILLCELL_X32 FILLER_245_1648 ();
 FILLCELL_X32 FILLER_245_1680 ();
 FILLCELL_X32 FILLER_245_1712 ();
 FILLCELL_X32 FILLER_245_1744 ();
 FILLCELL_X32 FILLER_245_1776 ();
 FILLCELL_X32 FILLER_245_1808 ();
 FILLCELL_X32 FILLER_245_1840 ();
 FILLCELL_X32 FILLER_245_1872 ();
 FILLCELL_X32 FILLER_245_1904 ();
 FILLCELL_X32 FILLER_245_1936 ();
 FILLCELL_X32 FILLER_245_1968 ();
 FILLCELL_X32 FILLER_245_2000 ();
 FILLCELL_X32 FILLER_245_2032 ();
 FILLCELL_X32 FILLER_245_2064 ();
 FILLCELL_X32 FILLER_245_2096 ();
 FILLCELL_X32 FILLER_245_2128 ();
 FILLCELL_X32 FILLER_245_2160 ();
 FILLCELL_X32 FILLER_245_2192 ();
 FILLCELL_X32 FILLER_245_2224 ();
 FILLCELL_X32 FILLER_245_2256 ();
 FILLCELL_X32 FILLER_245_2288 ();
 FILLCELL_X32 FILLER_245_2320 ();
 FILLCELL_X32 FILLER_245_2352 ();
 FILLCELL_X32 FILLER_245_2384 ();
 FILLCELL_X32 FILLER_245_2416 ();
 FILLCELL_X32 FILLER_245_2448 ();
 FILLCELL_X32 FILLER_245_2480 ();
 FILLCELL_X8 FILLER_245_2512 ();
 FILLCELL_X4 FILLER_245_2520 ();
 FILLCELL_X2 FILLER_245_2524 ();
 FILLCELL_X32 FILLER_245_2527 ();
 FILLCELL_X32 FILLER_245_2559 ();
 FILLCELL_X8 FILLER_245_2591 ();
 FILLCELL_X2 FILLER_245_2599 ();
 FILLCELL_X1 FILLER_245_2601 ();
 FILLCELL_X32 FILLER_246_1 ();
 FILLCELL_X32 FILLER_246_33 ();
 FILLCELL_X32 FILLER_246_65 ();
 FILLCELL_X32 FILLER_246_97 ();
 FILLCELL_X32 FILLER_246_129 ();
 FILLCELL_X32 FILLER_246_161 ();
 FILLCELL_X32 FILLER_246_193 ();
 FILLCELL_X32 FILLER_246_225 ();
 FILLCELL_X32 FILLER_246_257 ();
 FILLCELL_X32 FILLER_246_289 ();
 FILLCELL_X32 FILLER_246_321 ();
 FILLCELL_X32 FILLER_246_353 ();
 FILLCELL_X32 FILLER_246_385 ();
 FILLCELL_X32 FILLER_246_417 ();
 FILLCELL_X32 FILLER_246_449 ();
 FILLCELL_X32 FILLER_246_481 ();
 FILLCELL_X32 FILLER_246_513 ();
 FILLCELL_X32 FILLER_246_545 ();
 FILLCELL_X32 FILLER_246_577 ();
 FILLCELL_X16 FILLER_246_609 ();
 FILLCELL_X4 FILLER_246_625 ();
 FILLCELL_X2 FILLER_246_629 ();
 FILLCELL_X32 FILLER_246_632 ();
 FILLCELL_X32 FILLER_246_664 ();
 FILLCELL_X32 FILLER_246_696 ();
 FILLCELL_X32 FILLER_246_728 ();
 FILLCELL_X32 FILLER_246_760 ();
 FILLCELL_X32 FILLER_246_792 ();
 FILLCELL_X32 FILLER_246_824 ();
 FILLCELL_X32 FILLER_246_856 ();
 FILLCELL_X32 FILLER_246_888 ();
 FILLCELL_X32 FILLER_246_920 ();
 FILLCELL_X32 FILLER_246_952 ();
 FILLCELL_X32 FILLER_246_984 ();
 FILLCELL_X32 FILLER_246_1016 ();
 FILLCELL_X32 FILLER_246_1048 ();
 FILLCELL_X32 FILLER_246_1080 ();
 FILLCELL_X32 FILLER_246_1112 ();
 FILLCELL_X32 FILLER_246_1144 ();
 FILLCELL_X32 FILLER_246_1176 ();
 FILLCELL_X32 FILLER_246_1208 ();
 FILLCELL_X32 FILLER_246_1240 ();
 FILLCELL_X32 FILLER_246_1272 ();
 FILLCELL_X32 FILLER_246_1304 ();
 FILLCELL_X32 FILLER_246_1336 ();
 FILLCELL_X32 FILLER_246_1368 ();
 FILLCELL_X32 FILLER_246_1400 ();
 FILLCELL_X32 FILLER_246_1432 ();
 FILLCELL_X32 FILLER_246_1464 ();
 FILLCELL_X32 FILLER_246_1496 ();
 FILLCELL_X32 FILLER_246_1528 ();
 FILLCELL_X32 FILLER_246_1560 ();
 FILLCELL_X32 FILLER_246_1592 ();
 FILLCELL_X32 FILLER_246_1624 ();
 FILLCELL_X32 FILLER_246_1656 ();
 FILLCELL_X32 FILLER_246_1688 ();
 FILLCELL_X32 FILLER_246_1720 ();
 FILLCELL_X32 FILLER_246_1752 ();
 FILLCELL_X32 FILLER_246_1784 ();
 FILLCELL_X32 FILLER_246_1816 ();
 FILLCELL_X32 FILLER_246_1848 ();
 FILLCELL_X8 FILLER_246_1880 ();
 FILLCELL_X4 FILLER_246_1888 ();
 FILLCELL_X2 FILLER_246_1892 ();
 FILLCELL_X32 FILLER_246_1895 ();
 FILLCELL_X32 FILLER_246_1927 ();
 FILLCELL_X32 FILLER_246_1959 ();
 FILLCELL_X32 FILLER_246_1991 ();
 FILLCELL_X32 FILLER_246_2023 ();
 FILLCELL_X32 FILLER_246_2055 ();
 FILLCELL_X32 FILLER_246_2087 ();
 FILLCELL_X32 FILLER_246_2119 ();
 FILLCELL_X32 FILLER_246_2151 ();
 FILLCELL_X32 FILLER_246_2183 ();
 FILLCELL_X32 FILLER_246_2215 ();
 FILLCELL_X32 FILLER_246_2247 ();
 FILLCELL_X32 FILLER_246_2279 ();
 FILLCELL_X32 FILLER_246_2311 ();
 FILLCELL_X32 FILLER_246_2343 ();
 FILLCELL_X32 FILLER_246_2375 ();
 FILLCELL_X32 FILLER_246_2407 ();
 FILLCELL_X32 FILLER_246_2439 ();
 FILLCELL_X32 FILLER_246_2471 ();
 FILLCELL_X32 FILLER_246_2503 ();
 FILLCELL_X32 FILLER_246_2535 ();
 FILLCELL_X32 FILLER_246_2567 ();
 FILLCELL_X2 FILLER_246_2599 ();
 FILLCELL_X1 FILLER_246_2601 ();
 FILLCELL_X32 FILLER_247_1 ();
 FILLCELL_X32 FILLER_247_33 ();
 FILLCELL_X32 FILLER_247_65 ();
 FILLCELL_X32 FILLER_247_97 ();
 FILLCELL_X32 FILLER_247_129 ();
 FILLCELL_X32 FILLER_247_161 ();
 FILLCELL_X32 FILLER_247_193 ();
 FILLCELL_X32 FILLER_247_225 ();
 FILLCELL_X32 FILLER_247_257 ();
 FILLCELL_X32 FILLER_247_289 ();
 FILLCELL_X32 FILLER_247_321 ();
 FILLCELL_X32 FILLER_247_353 ();
 FILLCELL_X32 FILLER_247_385 ();
 FILLCELL_X32 FILLER_247_417 ();
 FILLCELL_X32 FILLER_247_449 ();
 FILLCELL_X32 FILLER_247_481 ();
 FILLCELL_X32 FILLER_247_513 ();
 FILLCELL_X32 FILLER_247_545 ();
 FILLCELL_X32 FILLER_247_577 ();
 FILLCELL_X32 FILLER_247_609 ();
 FILLCELL_X32 FILLER_247_641 ();
 FILLCELL_X32 FILLER_247_673 ();
 FILLCELL_X32 FILLER_247_705 ();
 FILLCELL_X32 FILLER_247_737 ();
 FILLCELL_X32 FILLER_247_769 ();
 FILLCELL_X32 FILLER_247_801 ();
 FILLCELL_X32 FILLER_247_833 ();
 FILLCELL_X32 FILLER_247_865 ();
 FILLCELL_X32 FILLER_247_897 ();
 FILLCELL_X32 FILLER_247_929 ();
 FILLCELL_X32 FILLER_247_961 ();
 FILLCELL_X32 FILLER_247_993 ();
 FILLCELL_X32 FILLER_247_1025 ();
 FILLCELL_X32 FILLER_247_1057 ();
 FILLCELL_X32 FILLER_247_1089 ();
 FILLCELL_X32 FILLER_247_1121 ();
 FILLCELL_X32 FILLER_247_1153 ();
 FILLCELL_X32 FILLER_247_1185 ();
 FILLCELL_X32 FILLER_247_1217 ();
 FILLCELL_X8 FILLER_247_1249 ();
 FILLCELL_X4 FILLER_247_1257 ();
 FILLCELL_X2 FILLER_247_1261 ();
 FILLCELL_X32 FILLER_247_1264 ();
 FILLCELL_X32 FILLER_247_1296 ();
 FILLCELL_X32 FILLER_247_1328 ();
 FILLCELL_X32 FILLER_247_1360 ();
 FILLCELL_X32 FILLER_247_1392 ();
 FILLCELL_X32 FILLER_247_1424 ();
 FILLCELL_X32 FILLER_247_1456 ();
 FILLCELL_X32 FILLER_247_1488 ();
 FILLCELL_X32 FILLER_247_1520 ();
 FILLCELL_X32 FILLER_247_1552 ();
 FILLCELL_X32 FILLER_247_1584 ();
 FILLCELL_X32 FILLER_247_1616 ();
 FILLCELL_X32 FILLER_247_1648 ();
 FILLCELL_X32 FILLER_247_1680 ();
 FILLCELL_X32 FILLER_247_1712 ();
 FILLCELL_X32 FILLER_247_1744 ();
 FILLCELL_X32 FILLER_247_1776 ();
 FILLCELL_X32 FILLER_247_1808 ();
 FILLCELL_X32 FILLER_247_1840 ();
 FILLCELL_X32 FILLER_247_1872 ();
 FILLCELL_X32 FILLER_247_1904 ();
 FILLCELL_X32 FILLER_247_1936 ();
 FILLCELL_X32 FILLER_247_1968 ();
 FILLCELL_X32 FILLER_247_2000 ();
 FILLCELL_X32 FILLER_247_2032 ();
 FILLCELL_X32 FILLER_247_2064 ();
 FILLCELL_X32 FILLER_247_2096 ();
 FILLCELL_X32 FILLER_247_2128 ();
 FILLCELL_X32 FILLER_247_2160 ();
 FILLCELL_X32 FILLER_247_2192 ();
 FILLCELL_X32 FILLER_247_2224 ();
 FILLCELL_X32 FILLER_247_2256 ();
 FILLCELL_X32 FILLER_247_2288 ();
 FILLCELL_X32 FILLER_247_2320 ();
 FILLCELL_X32 FILLER_247_2352 ();
 FILLCELL_X32 FILLER_247_2384 ();
 FILLCELL_X32 FILLER_247_2416 ();
 FILLCELL_X32 FILLER_247_2448 ();
 FILLCELL_X32 FILLER_247_2480 ();
 FILLCELL_X8 FILLER_247_2512 ();
 FILLCELL_X4 FILLER_247_2520 ();
 FILLCELL_X2 FILLER_247_2524 ();
 FILLCELL_X32 FILLER_247_2527 ();
 FILLCELL_X32 FILLER_247_2559 ();
 FILLCELL_X8 FILLER_247_2591 ();
 FILLCELL_X2 FILLER_247_2599 ();
 FILLCELL_X1 FILLER_247_2601 ();
 FILLCELL_X32 FILLER_248_1 ();
 FILLCELL_X32 FILLER_248_33 ();
 FILLCELL_X32 FILLER_248_65 ();
 FILLCELL_X32 FILLER_248_97 ();
 FILLCELL_X32 FILLER_248_129 ();
 FILLCELL_X32 FILLER_248_161 ();
 FILLCELL_X32 FILLER_248_193 ();
 FILLCELL_X32 FILLER_248_225 ();
 FILLCELL_X32 FILLER_248_257 ();
 FILLCELL_X32 FILLER_248_289 ();
 FILLCELL_X32 FILLER_248_321 ();
 FILLCELL_X32 FILLER_248_353 ();
 FILLCELL_X32 FILLER_248_385 ();
 FILLCELL_X32 FILLER_248_417 ();
 FILLCELL_X32 FILLER_248_449 ();
 FILLCELL_X32 FILLER_248_481 ();
 FILLCELL_X32 FILLER_248_513 ();
 FILLCELL_X32 FILLER_248_545 ();
 FILLCELL_X32 FILLER_248_577 ();
 FILLCELL_X16 FILLER_248_609 ();
 FILLCELL_X4 FILLER_248_625 ();
 FILLCELL_X2 FILLER_248_629 ();
 FILLCELL_X32 FILLER_248_632 ();
 FILLCELL_X32 FILLER_248_664 ();
 FILLCELL_X32 FILLER_248_696 ();
 FILLCELL_X32 FILLER_248_728 ();
 FILLCELL_X32 FILLER_248_760 ();
 FILLCELL_X32 FILLER_248_792 ();
 FILLCELL_X32 FILLER_248_824 ();
 FILLCELL_X32 FILLER_248_856 ();
 FILLCELL_X32 FILLER_248_888 ();
 FILLCELL_X32 FILLER_248_920 ();
 FILLCELL_X32 FILLER_248_952 ();
 FILLCELL_X32 FILLER_248_984 ();
 FILLCELL_X32 FILLER_248_1016 ();
 FILLCELL_X32 FILLER_248_1048 ();
 FILLCELL_X32 FILLER_248_1080 ();
 FILLCELL_X32 FILLER_248_1112 ();
 FILLCELL_X32 FILLER_248_1144 ();
 FILLCELL_X32 FILLER_248_1176 ();
 FILLCELL_X32 FILLER_248_1208 ();
 FILLCELL_X32 FILLER_248_1240 ();
 FILLCELL_X32 FILLER_248_1272 ();
 FILLCELL_X32 FILLER_248_1304 ();
 FILLCELL_X32 FILLER_248_1336 ();
 FILLCELL_X32 FILLER_248_1368 ();
 FILLCELL_X32 FILLER_248_1400 ();
 FILLCELL_X32 FILLER_248_1432 ();
 FILLCELL_X32 FILLER_248_1464 ();
 FILLCELL_X32 FILLER_248_1496 ();
 FILLCELL_X32 FILLER_248_1528 ();
 FILLCELL_X32 FILLER_248_1560 ();
 FILLCELL_X32 FILLER_248_1592 ();
 FILLCELL_X32 FILLER_248_1624 ();
 FILLCELL_X32 FILLER_248_1656 ();
 FILLCELL_X32 FILLER_248_1688 ();
 FILLCELL_X32 FILLER_248_1720 ();
 FILLCELL_X32 FILLER_248_1752 ();
 FILLCELL_X32 FILLER_248_1784 ();
 FILLCELL_X32 FILLER_248_1816 ();
 FILLCELL_X32 FILLER_248_1848 ();
 FILLCELL_X8 FILLER_248_1880 ();
 FILLCELL_X4 FILLER_248_1888 ();
 FILLCELL_X2 FILLER_248_1892 ();
 FILLCELL_X32 FILLER_248_1895 ();
 FILLCELL_X32 FILLER_248_1927 ();
 FILLCELL_X32 FILLER_248_1959 ();
 FILLCELL_X32 FILLER_248_1991 ();
 FILLCELL_X32 FILLER_248_2023 ();
 FILLCELL_X32 FILLER_248_2055 ();
 FILLCELL_X32 FILLER_248_2087 ();
 FILLCELL_X32 FILLER_248_2119 ();
 FILLCELL_X32 FILLER_248_2151 ();
 FILLCELL_X32 FILLER_248_2183 ();
 FILLCELL_X32 FILLER_248_2215 ();
 FILLCELL_X32 FILLER_248_2247 ();
 FILLCELL_X32 FILLER_248_2279 ();
 FILLCELL_X32 FILLER_248_2311 ();
 FILLCELL_X32 FILLER_248_2343 ();
 FILLCELL_X32 FILLER_248_2375 ();
 FILLCELL_X32 FILLER_248_2407 ();
 FILLCELL_X32 FILLER_248_2439 ();
 FILLCELL_X32 FILLER_248_2471 ();
 FILLCELL_X32 FILLER_248_2503 ();
 FILLCELL_X32 FILLER_248_2535 ();
 FILLCELL_X32 FILLER_248_2567 ();
 FILLCELL_X2 FILLER_248_2599 ();
 FILLCELL_X1 FILLER_248_2601 ();
 FILLCELL_X32 FILLER_249_1 ();
 FILLCELL_X32 FILLER_249_33 ();
 FILLCELL_X32 FILLER_249_65 ();
 FILLCELL_X32 FILLER_249_97 ();
 FILLCELL_X32 FILLER_249_129 ();
 FILLCELL_X32 FILLER_249_161 ();
 FILLCELL_X32 FILLER_249_193 ();
 FILLCELL_X32 FILLER_249_225 ();
 FILLCELL_X32 FILLER_249_257 ();
 FILLCELL_X32 FILLER_249_289 ();
 FILLCELL_X32 FILLER_249_321 ();
 FILLCELL_X32 FILLER_249_353 ();
 FILLCELL_X32 FILLER_249_385 ();
 FILLCELL_X32 FILLER_249_417 ();
 FILLCELL_X32 FILLER_249_449 ();
 FILLCELL_X32 FILLER_249_481 ();
 FILLCELL_X32 FILLER_249_513 ();
 FILLCELL_X32 FILLER_249_545 ();
 FILLCELL_X32 FILLER_249_577 ();
 FILLCELL_X32 FILLER_249_609 ();
 FILLCELL_X32 FILLER_249_641 ();
 FILLCELL_X32 FILLER_249_673 ();
 FILLCELL_X32 FILLER_249_705 ();
 FILLCELL_X32 FILLER_249_737 ();
 FILLCELL_X32 FILLER_249_769 ();
 FILLCELL_X32 FILLER_249_801 ();
 FILLCELL_X32 FILLER_249_833 ();
 FILLCELL_X32 FILLER_249_865 ();
 FILLCELL_X32 FILLER_249_897 ();
 FILLCELL_X32 FILLER_249_929 ();
 FILLCELL_X32 FILLER_249_961 ();
 FILLCELL_X32 FILLER_249_993 ();
 FILLCELL_X32 FILLER_249_1025 ();
 FILLCELL_X32 FILLER_249_1057 ();
 FILLCELL_X32 FILLER_249_1089 ();
 FILLCELL_X32 FILLER_249_1121 ();
 FILLCELL_X32 FILLER_249_1153 ();
 FILLCELL_X32 FILLER_249_1185 ();
 FILLCELL_X32 FILLER_249_1217 ();
 FILLCELL_X8 FILLER_249_1249 ();
 FILLCELL_X4 FILLER_249_1257 ();
 FILLCELL_X2 FILLER_249_1261 ();
 FILLCELL_X32 FILLER_249_1264 ();
 FILLCELL_X32 FILLER_249_1296 ();
 FILLCELL_X32 FILLER_249_1328 ();
 FILLCELL_X32 FILLER_249_1360 ();
 FILLCELL_X32 FILLER_249_1392 ();
 FILLCELL_X32 FILLER_249_1424 ();
 FILLCELL_X32 FILLER_249_1456 ();
 FILLCELL_X32 FILLER_249_1488 ();
 FILLCELL_X32 FILLER_249_1520 ();
 FILLCELL_X32 FILLER_249_1552 ();
 FILLCELL_X32 FILLER_249_1584 ();
 FILLCELL_X32 FILLER_249_1616 ();
 FILLCELL_X32 FILLER_249_1648 ();
 FILLCELL_X32 FILLER_249_1680 ();
 FILLCELL_X32 FILLER_249_1712 ();
 FILLCELL_X32 FILLER_249_1744 ();
 FILLCELL_X32 FILLER_249_1776 ();
 FILLCELL_X32 FILLER_249_1808 ();
 FILLCELL_X32 FILLER_249_1840 ();
 FILLCELL_X32 FILLER_249_1872 ();
 FILLCELL_X32 FILLER_249_1904 ();
 FILLCELL_X32 FILLER_249_1936 ();
 FILLCELL_X32 FILLER_249_1968 ();
 FILLCELL_X32 FILLER_249_2000 ();
 FILLCELL_X32 FILLER_249_2032 ();
 FILLCELL_X32 FILLER_249_2064 ();
 FILLCELL_X32 FILLER_249_2096 ();
 FILLCELL_X32 FILLER_249_2128 ();
 FILLCELL_X32 FILLER_249_2160 ();
 FILLCELL_X32 FILLER_249_2192 ();
 FILLCELL_X32 FILLER_249_2224 ();
 FILLCELL_X32 FILLER_249_2256 ();
 FILLCELL_X32 FILLER_249_2288 ();
 FILLCELL_X32 FILLER_249_2320 ();
 FILLCELL_X32 FILLER_249_2352 ();
 FILLCELL_X32 FILLER_249_2384 ();
 FILLCELL_X32 FILLER_249_2416 ();
 FILLCELL_X32 FILLER_249_2448 ();
 FILLCELL_X32 FILLER_249_2480 ();
 FILLCELL_X8 FILLER_249_2512 ();
 FILLCELL_X4 FILLER_249_2520 ();
 FILLCELL_X2 FILLER_249_2524 ();
 FILLCELL_X32 FILLER_249_2527 ();
 FILLCELL_X32 FILLER_249_2559 ();
 FILLCELL_X8 FILLER_249_2591 ();
 FILLCELL_X2 FILLER_249_2599 ();
 FILLCELL_X1 FILLER_249_2601 ();
 FILLCELL_X32 FILLER_250_1 ();
 FILLCELL_X32 FILLER_250_33 ();
 FILLCELL_X32 FILLER_250_65 ();
 FILLCELL_X32 FILLER_250_97 ();
 FILLCELL_X32 FILLER_250_129 ();
 FILLCELL_X32 FILLER_250_161 ();
 FILLCELL_X32 FILLER_250_193 ();
 FILLCELL_X32 FILLER_250_225 ();
 FILLCELL_X32 FILLER_250_257 ();
 FILLCELL_X32 FILLER_250_289 ();
 FILLCELL_X32 FILLER_250_321 ();
 FILLCELL_X32 FILLER_250_353 ();
 FILLCELL_X32 FILLER_250_385 ();
 FILLCELL_X32 FILLER_250_417 ();
 FILLCELL_X32 FILLER_250_449 ();
 FILLCELL_X32 FILLER_250_481 ();
 FILLCELL_X32 FILLER_250_513 ();
 FILLCELL_X32 FILLER_250_545 ();
 FILLCELL_X32 FILLER_250_577 ();
 FILLCELL_X16 FILLER_250_609 ();
 FILLCELL_X4 FILLER_250_625 ();
 FILLCELL_X2 FILLER_250_629 ();
 FILLCELL_X32 FILLER_250_632 ();
 FILLCELL_X32 FILLER_250_664 ();
 FILLCELL_X32 FILLER_250_696 ();
 FILLCELL_X32 FILLER_250_728 ();
 FILLCELL_X32 FILLER_250_760 ();
 FILLCELL_X32 FILLER_250_792 ();
 FILLCELL_X32 FILLER_250_824 ();
 FILLCELL_X32 FILLER_250_856 ();
 FILLCELL_X32 FILLER_250_888 ();
 FILLCELL_X32 FILLER_250_920 ();
 FILLCELL_X32 FILLER_250_952 ();
 FILLCELL_X32 FILLER_250_984 ();
 FILLCELL_X32 FILLER_250_1016 ();
 FILLCELL_X32 FILLER_250_1048 ();
 FILLCELL_X32 FILLER_250_1080 ();
 FILLCELL_X32 FILLER_250_1112 ();
 FILLCELL_X32 FILLER_250_1144 ();
 FILLCELL_X32 FILLER_250_1176 ();
 FILLCELL_X32 FILLER_250_1208 ();
 FILLCELL_X32 FILLER_250_1240 ();
 FILLCELL_X32 FILLER_250_1272 ();
 FILLCELL_X32 FILLER_250_1304 ();
 FILLCELL_X32 FILLER_250_1336 ();
 FILLCELL_X32 FILLER_250_1368 ();
 FILLCELL_X32 FILLER_250_1400 ();
 FILLCELL_X32 FILLER_250_1432 ();
 FILLCELL_X32 FILLER_250_1464 ();
 FILLCELL_X32 FILLER_250_1496 ();
 FILLCELL_X32 FILLER_250_1528 ();
 FILLCELL_X32 FILLER_250_1560 ();
 FILLCELL_X32 FILLER_250_1592 ();
 FILLCELL_X32 FILLER_250_1624 ();
 FILLCELL_X32 FILLER_250_1656 ();
 FILLCELL_X32 FILLER_250_1688 ();
 FILLCELL_X32 FILLER_250_1720 ();
 FILLCELL_X32 FILLER_250_1752 ();
 FILLCELL_X32 FILLER_250_1784 ();
 FILLCELL_X32 FILLER_250_1816 ();
 FILLCELL_X32 FILLER_250_1848 ();
 FILLCELL_X8 FILLER_250_1880 ();
 FILLCELL_X4 FILLER_250_1888 ();
 FILLCELL_X2 FILLER_250_1892 ();
 FILLCELL_X32 FILLER_250_1895 ();
 FILLCELL_X32 FILLER_250_1927 ();
 FILLCELL_X32 FILLER_250_1959 ();
 FILLCELL_X32 FILLER_250_1991 ();
 FILLCELL_X32 FILLER_250_2023 ();
 FILLCELL_X32 FILLER_250_2055 ();
 FILLCELL_X32 FILLER_250_2087 ();
 FILLCELL_X32 FILLER_250_2119 ();
 FILLCELL_X32 FILLER_250_2151 ();
 FILLCELL_X32 FILLER_250_2183 ();
 FILLCELL_X32 FILLER_250_2215 ();
 FILLCELL_X32 FILLER_250_2247 ();
 FILLCELL_X32 FILLER_250_2279 ();
 FILLCELL_X32 FILLER_250_2311 ();
 FILLCELL_X32 FILLER_250_2343 ();
 FILLCELL_X32 FILLER_250_2375 ();
 FILLCELL_X32 FILLER_250_2407 ();
 FILLCELL_X32 FILLER_250_2439 ();
 FILLCELL_X32 FILLER_250_2471 ();
 FILLCELL_X32 FILLER_250_2503 ();
 FILLCELL_X32 FILLER_250_2535 ();
 FILLCELL_X32 FILLER_250_2567 ();
 FILLCELL_X2 FILLER_250_2599 ();
 FILLCELL_X1 FILLER_250_2601 ();
 FILLCELL_X32 FILLER_251_1 ();
 FILLCELL_X32 FILLER_251_33 ();
 FILLCELL_X32 FILLER_251_65 ();
 FILLCELL_X32 FILLER_251_97 ();
 FILLCELL_X32 FILLER_251_129 ();
 FILLCELL_X32 FILLER_251_161 ();
 FILLCELL_X32 FILLER_251_193 ();
 FILLCELL_X32 FILLER_251_225 ();
 FILLCELL_X32 FILLER_251_257 ();
 FILLCELL_X32 FILLER_251_289 ();
 FILLCELL_X32 FILLER_251_321 ();
 FILLCELL_X32 FILLER_251_353 ();
 FILLCELL_X32 FILLER_251_385 ();
 FILLCELL_X32 FILLER_251_417 ();
 FILLCELL_X32 FILLER_251_449 ();
 FILLCELL_X32 FILLER_251_481 ();
 FILLCELL_X32 FILLER_251_513 ();
 FILLCELL_X32 FILLER_251_545 ();
 FILLCELL_X32 FILLER_251_577 ();
 FILLCELL_X32 FILLER_251_609 ();
 FILLCELL_X32 FILLER_251_641 ();
 FILLCELL_X32 FILLER_251_673 ();
 FILLCELL_X32 FILLER_251_705 ();
 FILLCELL_X32 FILLER_251_737 ();
 FILLCELL_X32 FILLER_251_769 ();
 FILLCELL_X32 FILLER_251_801 ();
 FILLCELL_X32 FILLER_251_833 ();
 FILLCELL_X32 FILLER_251_865 ();
 FILLCELL_X32 FILLER_251_897 ();
 FILLCELL_X32 FILLER_251_929 ();
 FILLCELL_X32 FILLER_251_961 ();
 FILLCELL_X32 FILLER_251_993 ();
 FILLCELL_X32 FILLER_251_1025 ();
 FILLCELL_X32 FILLER_251_1057 ();
 FILLCELL_X32 FILLER_251_1089 ();
 FILLCELL_X32 FILLER_251_1121 ();
 FILLCELL_X32 FILLER_251_1153 ();
 FILLCELL_X32 FILLER_251_1185 ();
 FILLCELL_X32 FILLER_251_1217 ();
 FILLCELL_X8 FILLER_251_1249 ();
 FILLCELL_X4 FILLER_251_1257 ();
 FILLCELL_X2 FILLER_251_1261 ();
 FILLCELL_X32 FILLER_251_1264 ();
 FILLCELL_X32 FILLER_251_1296 ();
 FILLCELL_X32 FILLER_251_1328 ();
 FILLCELL_X32 FILLER_251_1360 ();
 FILLCELL_X32 FILLER_251_1392 ();
 FILLCELL_X32 FILLER_251_1424 ();
 FILLCELL_X32 FILLER_251_1456 ();
 FILLCELL_X32 FILLER_251_1488 ();
 FILLCELL_X32 FILLER_251_1520 ();
 FILLCELL_X32 FILLER_251_1552 ();
 FILLCELL_X32 FILLER_251_1584 ();
 FILLCELL_X32 FILLER_251_1616 ();
 FILLCELL_X32 FILLER_251_1648 ();
 FILLCELL_X32 FILLER_251_1680 ();
 FILLCELL_X32 FILLER_251_1712 ();
 FILLCELL_X32 FILLER_251_1744 ();
 FILLCELL_X32 FILLER_251_1776 ();
 FILLCELL_X32 FILLER_251_1808 ();
 FILLCELL_X32 FILLER_251_1840 ();
 FILLCELL_X32 FILLER_251_1872 ();
 FILLCELL_X32 FILLER_251_1904 ();
 FILLCELL_X32 FILLER_251_1936 ();
 FILLCELL_X32 FILLER_251_1968 ();
 FILLCELL_X32 FILLER_251_2000 ();
 FILLCELL_X32 FILLER_251_2032 ();
 FILLCELL_X32 FILLER_251_2064 ();
 FILLCELL_X32 FILLER_251_2096 ();
 FILLCELL_X32 FILLER_251_2128 ();
 FILLCELL_X32 FILLER_251_2160 ();
 FILLCELL_X32 FILLER_251_2192 ();
 FILLCELL_X32 FILLER_251_2224 ();
 FILLCELL_X32 FILLER_251_2256 ();
 FILLCELL_X32 FILLER_251_2288 ();
 FILLCELL_X32 FILLER_251_2320 ();
 FILLCELL_X32 FILLER_251_2352 ();
 FILLCELL_X32 FILLER_251_2384 ();
 FILLCELL_X32 FILLER_251_2416 ();
 FILLCELL_X32 FILLER_251_2448 ();
 FILLCELL_X32 FILLER_251_2480 ();
 FILLCELL_X8 FILLER_251_2512 ();
 FILLCELL_X4 FILLER_251_2520 ();
 FILLCELL_X2 FILLER_251_2524 ();
 FILLCELL_X32 FILLER_251_2527 ();
 FILLCELL_X32 FILLER_251_2559 ();
 FILLCELL_X8 FILLER_251_2591 ();
 FILLCELL_X2 FILLER_251_2599 ();
 FILLCELL_X1 FILLER_251_2601 ();
 FILLCELL_X32 FILLER_252_1 ();
 FILLCELL_X32 FILLER_252_33 ();
 FILLCELL_X32 FILLER_252_65 ();
 FILLCELL_X32 FILLER_252_97 ();
 FILLCELL_X32 FILLER_252_129 ();
 FILLCELL_X32 FILLER_252_161 ();
 FILLCELL_X32 FILLER_252_193 ();
 FILLCELL_X32 FILLER_252_225 ();
 FILLCELL_X32 FILLER_252_257 ();
 FILLCELL_X32 FILLER_252_289 ();
 FILLCELL_X32 FILLER_252_321 ();
 FILLCELL_X32 FILLER_252_353 ();
 FILLCELL_X32 FILLER_252_385 ();
 FILLCELL_X32 FILLER_252_417 ();
 FILLCELL_X32 FILLER_252_449 ();
 FILLCELL_X32 FILLER_252_481 ();
 FILLCELL_X32 FILLER_252_513 ();
 FILLCELL_X32 FILLER_252_545 ();
 FILLCELL_X32 FILLER_252_577 ();
 FILLCELL_X16 FILLER_252_609 ();
 FILLCELL_X4 FILLER_252_625 ();
 FILLCELL_X2 FILLER_252_629 ();
 FILLCELL_X32 FILLER_252_632 ();
 FILLCELL_X32 FILLER_252_664 ();
 FILLCELL_X32 FILLER_252_696 ();
 FILLCELL_X32 FILLER_252_728 ();
 FILLCELL_X32 FILLER_252_760 ();
 FILLCELL_X32 FILLER_252_792 ();
 FILLCELL_X32 FILLER_252_824 ();
 FILLCELL_X32 FILLER_252_856 ();
 FILLCELL_X32 FILLER_252_888 ();
 FILLCELL_X32 FILLER_252_920 ();
 FILLCELL_X32 FILLER_252_952 ();
 FILLCELL_X32 FILLER_252_984 ();
 FILLCELL_X32 FILLER_252_1016 ();
 FILLCELL_X32 FILLER_252_1048 ();
 FILLCELL_X32 FILLER_252_1080 ();
 FILLCELL_X32 FILLER_252_1112 ();
 FILLCELL_X32 FILLER_252_1144 ();
 FILLCELL_X32 FILLER_252_1176 ();
 FILLCELL_X32 FILLER_252_1208 ();
 FILLCELL_X32 FILLER_252_1240 ();
 FILLCELL_X32 FILLER_252_1272 ();
 FILLCELL_X32 FILLER_252_1304 ();
 FILLCELL_X32 FILLER_252_1336 ();
 FILLCELL_X32 FILLER_252_1368 ();
 FILLCELL_X32 FILLER_252_1400 ();
 FILLCELL_X32 FILLER_252_1432 ();
 FILLCELL_X32 FILLER_252_1464 ();
 FILLCELL_X32 FILLER_252_1496 ();
 FILLCELL_X32 FILLER_252_1528 ();
 FILLCELL_X32 FILLER_252_1560 ();
 FILLCELL_X32 FILLER_252_1592 ();
 FILLCELL_X32 FILLER_252_1624 ();
 FILLCELL_X32 FILLER_252_1656 ();
 FILLCELL_X32 FILLER_252_1688 ();
 FILLCELL_X32 FILLER_252_1720 ();
 FILLCELL_X32 FILLER_252_1752 ();
 FILLCELL_X32 FILLER_252_1784 ();
 FILLCELL_X32 FILLER_252_1816 ();
 FILLCELL_X32 FILLER_252_1848 ();
 FILLCELL_X8 FILLER_252_1880 ();
 FILLCELL_X4 FILLER_252_1888 ();
 FILLCELL_X2 FILLER_252_1892 ();
 FILLCELL_X32 FILLER_252_1895 ();
 FILLCELL_X32 FILLER_252_1927 ();
 FILLCELL_X32 FILLER_252_1959 ();
 FILLCELL_X32 FILLER_252_1991 ();
 FILLCELL_X32 FILLER_252_2023 ();
 FILLCELL_X32 FILLER_252_2055 ();
 FILLCELL_X32 FILLER_252_2087 ();
 FILLCELL_X32 FILLER_252_2119 ();
 FILLCELL_X32 FILLER_252_2151 ();
 FILLCELL_X32 FILLER_252_2183 ();
 FILLCELL_X32 FILLER_252_2215 ();
 FILLCELL_X32 FILLER_252_2247 ();
 FILLCELL_X32 FILLER_252_2279 ();
 FILLCELL_X32 FILLER_252_2311 ();
 FILLCELL_X32 FILLER_252_2343 ();
 FILLCELL_X32 FILLER_252_2375 ();
 FILLCELL_X32 FILLER_252_2407 ();
 FILLCELL_X32 FILLER_252_2439 ();
 FILLCELL_X32 FILLER_252_2471 ();
 FILLCELL_X32 FILLER_252_2503 ();
 FILLCELL_X32 FILLER_252_2535 ();
 FILLCELL_X32 FILLER_252_2567 ();
 FILLCELL_X2 FILLER_252_2599 ();
 FILLCELL_X1 FILLER_252_2601 ();
 FILLCELL_X32 FILLER_253_1 ();
 FILLCELL_X32 FILLER_253_33 ();
 FILLCELL_X32 FILLER_253_65 ();
 FILLCELL_X32 FILLER_253_97 ();
 FILLCELL_X32 FILLER_253_129 ();
 FILLCELL_X32 FILLER_253_161 ();
 FILLCELL_X32 FILLER_253_193 ();
 FILLCELL_X32 FILLER_253_225 ();
 FILLCELL_X32 FILLER_253_257 ();
 FILLCELL_X32 FILLER_253_289 ();
 FILLCELL_X32 FILLER_253_321 ();
 FILLCELL_X32 FILLER_253_353 ();
 FILLCELL_X32 FILLER_253_385 ();
 FILLCELL_X32 FILLER_253_417 ();
 FILLCELL_X32 FILLER_253_449 ();
 FILLCELL_X32 FILLER_253_481 ();
 FILLCELL_X32 FILLER_253_513 ();
 FILLCELL_X32 FILLER_253_545 ();
 FILLCELL_X32 FILLER_253_577 ();
 FILLCELL_X32 FILLER_253_609 ();
 FILLCELL_X32 FILLER_253_641 ();
 FILLCELL_X32 FILLER_253_673 ();
 FILLCELL_X32 FILLER_253_705 ();
 FILLCELL_X32 FILLER_253_737 ();
 FILLCELL_X32 FILLER_253_769 ();
 FILLCELL_X32 FILLER_253_801 ();
 FILLCELL_X32 FILLER_253_833 ();
 FILLCELL_X32 FILLER_253_865 ();
 FILLCELL_X32 FILLER_253_897 ();
 FILLCELL_X32 FILLER_253_929 ();
 FILLCELL_X32 FILLER_253_961 ();
 FILLCELL_X32 FILLER_253_993 ();
 FILLCELL_X32 FILLER_253_1025 ();
 FILLCELL_X32 FILLER_253_1057 ();
 FILLCELL_X32 FILLER_253_1089 ();
 FILLCELL_X32 FILLER_253_1121 ();
 FILLCELL_X32 FILLER_253_1153 ();
 FILLCELL_X32 FILLER_253_1185 ();
 FILLCELL_X32 FILLER_253_1217 ();
 FILLCELL_X8 FILLER_253_1249 ();
 FILLCELL_X4 FILLER_253_1257 ();
 FILLCELL_X2 FILLER_253_1261 ();
 FILLCELL_X32 FILLER_253_1264 ();
 FILLCELL_X32 FILLER_253_1296 ();
 FILLCELL_X32 FILLER_253_1328 ();
 FILLCELL_X32 FILLER_253_1360 ();
 FILLCELL_X32 FILLER_253_1392 ();
 FILLCELL_X32 FILLER_253_1424 ();
 FILLCELL_X32 FILLER_253_1456 ();
 FILLCELL_X32 FILLER_253_1488 ();
 FILLCELL_X32 FILLER_253_1520 ();
 FILLCELL_X32 FILLER_253_1552 ();
 FILLCELL_X32 FILLER_253_1584 ();
 FILLCELL_X32 FILLER_253_1616 ();
 FILLCELL_X32 FILLER_253_1648 ();
 FILLCELL_X32 FILLER_253_1680 ();
 FILLCELL_X32 FILLER_253_1712 ();
 FILLCELL_X32 FILLER_253_1744 ();
 FILLCELL_X32 FILLER_253_1776 ();
 FILLCELL_X32 FILLER_253_1808 ();
 FILLCELL_X32 FILLER_253_1840 ();
 FILLCELL_X32 FILLER_253_1872 ();
 FILLCELL_X32 FILLER_253_1904 ();
 FILLCELL_X32 FILLER_253_1936 ();
 FILLCELL_X32 FILLER_253_1968 ();
 FILLCELL_X32 FILLER_253_2000 ();
 FILLCELL_X32 FILLER_253_2032 ();
 FILLCELL_X32 FILLER_253_2064 ();
 FILLCELL_X32 FILLER_253_2096 ();
 FILLCELL_X32 FILLER_253_2128 ();
 FILLCELL_X32 FILLER_253_2160 ();
 FILLCELL_X32 FILLER_253_2192 ();
 FILLCELL_X32 FILLER_253_2224 ();
 FILLCELL_X32 FILLER_253_2256 ();
 FILLCELL_X32 FILLER_253_2288 ();
 FILLCELL_X32 FILLER_253_2320 ();
 FILLCELL_X32 FILLER_253_2352 ();
 FILLCELL_X32 FILLER_253_2384 ();
 FILLCELL_X32 FILLER_253_2416 ();
 FILLCELL_X32 FILLER_253_2448 ();
 FILLCELL_X32 FILLER_253_2480 ();
 FILLCELL_X8 FILLER_253_2512 ();
 FILLCELL_X4 FILLER_253_2520 ();
 FILLCELL_X2 FILLER_253_2524 ();
 FILLCELL_X32 FILLER_253_2527 ();
 FILLCELL_X32 FILLER_253_2559 ();
 FILLCELL_X8 FILLER_253_2591 ();
 FILLCELL_X2 FILLER_253_2599 ();
 FILLCELL_X1 FILLER_253_2601 ();
 FILLCELL_X32 FILLER_254_1 ();
 FILLCELL_X32 FILLER_254_33 ();
 FILLCELL_X32 FILLER_254_65 ();
 FILLCELL_X32 FILLER_254_97 ();
 FILLCELL_X32 FILLER_254_129 ();
 FILLCELL_X32 FILLER_254_161 ();
 FILLCELL_X32 FILLER_254_193 ();
 FILLCELL_X32 FILLER_254_225 ();
 FILLCELL_X32 FILLER_254_257 ();
 FILLCELL_X32 FILLER_254_289 ();
 FILLCELL_X32 FILLER_254_321 ();
 FILLCELL_X32 FILLER_254_353 ();
 FILLCELL_X32 FILLER_254_385 ();
 FILLCELL_X32 FILLER_254_417 ();
 FILLCELL_X32 FILLER_254_449 ();
 FILLCELL_X32 FILLER_254_481 ();
 FILLCELL_X32 FILLER_254_513 ();
 FILLCELL_X32 FILLER_254_545 ();
 FILLCELL_X32 FILLER_254_577 ();
 FILLCELL_X16 FILLER_254_609 ();
 FILLCELL_X4 FILLER_254_625 ();
 FILLCELL_X2 FILLER_254_629 ();
 FILLCELL_X32 FILLER_254_632 ();
 FILLCELL_X32 FILLER_254_664 ();
 FILLCELL_X32 FILLER_254_696 ();
 FILLCELL_X32 FILLER_254_728 ();
 FILLCELL_X32 FILLER_254_760 ();
 FILLCELL_X32 FILLER_254_792 ();
 FILLCELL_X32 FILLER_254_824 ();
 FILLCELL_X32 FILLER_254_856 ();
 FILLCELL_X32 FILLER_254_888 ();
 FILLCELL_X32 FILLER_254_920 ();
 FILLCELL_X32 FILLER_254_952 ();
 FILLCELL_X32 FILLER_254_984 ();
 FILLCELL_X32 FILLER_254_1016 ();
 FILLCELL_X32 FILLER_254_1048 ();
 FILLCELL_X32 FILLER_254_1080 ();
 FILLCELL_X32 FILLER_254_1112 ();
 FILLCELL_X32 FILLER_254_1144 ();
 FILLCELL_X32 FILLER_254_1176 ();
 FILLCELL_X32 FILLER_254_1208 ();
 FILLCELL_X32 FILLER_254_1240 ();
 FILLCELL_X32 FILLER_254_1272 ();
 FILLCELL_X32 FILLER_254_1304 ();
 FILLCELL_X32 FILLER_254_1336 ();
 FILLCELL_X32 FILLER_254_1368 ();
 FILLCELL_X32 FILLER_254_1400 ();
 FILLCELL_X32 FILLER_254_1432 ();
 FILLCELL_X32 FILLER_254_1464 ();
 FILLCELL_X32 FILLER_254_1496 ();
 FILLCELL_X32 FILLER_254_1528 ();
 FILLCELL_X32 FILLER_254_1560 ();
 FILLCELL_X32 FILLER_254_1592 ();
 FILLCELL_X32 FILLER_254_1624 ();
 FILLCELL_X32 FILLER_254_1656 ();
 FILLCELL_X32 FILLER_254_1688 ();
 FILLCELL_X32 FILLER_254_1720 ();
 FILLCELL_X32 FILLER_254_1752 ();
 FILLCELL_X32 FILLER_254_1784 ();
 FILLCELL_X32 FILLER_254_1816 ();
 FILLCELL_X32 FILLER_254_1848 ();
 FILLCELL_X8 FILLER_254_1880 ();
 FILLCELL_X4 FILLER_254_1888 ();
 FILLCELL_X2 FILLER_254_1892 ();
 FILLCELL_X32 FILLER_254_1895 ();
 FILLCELL_X32 FILLER_254_1927 ();
 FILLCELL_X32 FILLER_254_1959 ();
 FILLCELL_X32 FILLER_254_1991 ();
 FILLCELL_X32 FILLER_254_2023 ();
 FILLCELL_X32 FILLER_254_2055 ();
 FILLCELL_X32 FILLER_254_2087 ();
 FILLCELL_X32 FILLER_254_2119 ();
 FILLCELL_X32 FILLER_254_2151 ();
 FILLCELL_X32 FILLER_254_2183 ();
 FILLCELL_X32 FILLER_254_2215 ();
 FILLCELL_X32 FILLER_254_2247 ();
 FILLCELL_X32 FILLER_254_2279 ();
 FILLCELL_X32 FILLER_254_2311 ();
 FILLCELL_X32 FILLER_254_2343 ();
 FILLCELL_X32 FILLER_254_2375 ();
 FILLCELL_X32 FILLER_254_2407 ();
 FILLCELL_X32 FILLER_254_2439 ();
 FILLCELL_X32 FILLER_254_2471 ();
 FILLCELL_X32 FILLER_254_2503 ();
 FILLCELL_X32 FILLER_254_2535 ();
 FILLCELL_X32 FILLER_254_2567 ();
 FILLCELL_X2 FILLER_254_2599 ();
 FILLCELL_X1 FILLER_254_2601 ();
 FILLCELL_X32 FILLER_255_1 ();
 FILLCELL_X32 FILLER_255_33 ();
 FILLCELL_X32 FILLER_255_65 ();
 FILLCELL_X32 FILLER_255_97 ();
 FILLCELL_X32 FILLER_255_129 ();
 FILLCELL_X32 FILLER_255_161 ();
 FILLCELL_X32 FILLER_255_193 ();
 FILLCELL_X32 FILLER_255_225 ();
 FILLCELL_X32 FILLER_255_257 ();
 FILLCELL_X32 FILLER_255_289 ();
 FILLCELL_X32 FILLER_255_321 ();
 FILLCELL_X32 FILLER_255_353 ();
 FILLCELL_X32 FILLER_255_385 ();
 FILLCELL_X32 FILLER_255_417 ();
 FILLCELL_X32 FILLER_255_449 ();
 FILLCELL_X32 FILLER_255_481 ();
 FILLCELL_X32 FILLER_255_513 ();
 FILLCELL_X32 FILLER_255_545 ();
 FILLCELL_X32 FILLER_255_577 ();
 FILLCELL_X32 FILLER_255_609 ();
 FILLCELL_X32 FILLER_255_641 ();
 FILLCELL_X32 FILLER_255_673 ();
 FILLCELL_X32 FILLER_255_705 ();
 FILLCELL_X32 FILLER_255_737 ();
 FILLCELL_X32 FILLER_255_769 ();
 FILLCELL_X32 FILLER_255_801 ();
 FILLCELL_X32 FILLER_255_833 ();
 FILLCELL_X32 FILLER_255_865 ();
 FILLCELL_X32 FILLER_255_897 ();
 FILLCELL_X32 FILLER_255_929 ();
 FILLCELL_X32 FILLER_255_961 ();
 FILLCELL_X32 FILLER_255_993 ();
 FILLCELL_X32 FILLER_255_1025 ();
 FILLCELL_X32 FILLER_255_1057 ();
 FILLCELL_X32 FILLER_255_1089 ();
 FILLCELL_X32 FILLER_255_1121 ();
 FILLCELL_X32 FILLER_255_1153 ();
 FILLCELL_X32 FILLER_255_1185 ();
 FILLCELL_X32 FILLER_255_1217 ();
 FILLCELL_X8 FILLER_255_1249 ();
 FILLCELL_X4 FILLER_255_1257 ();
 FILLCELL_X2 FILLER_255_1261 ();
 FILLCELL_X32 FILLER_255_1264 ();
 FILLCELL_X32 FILLER_255_1296 ();
 FILLCELL_X32 FILLER_255_1328 ();
 FILLCELL_X32 FILLER_255_1360 ();
 FILLCELL_X32 FILLER_255_1392 ();
 FILLCELL_X32 FILLER_255_1424 ();
 FILLCELL_X32 FILLER_255_1456 ();
 FILLCELL_X32 FILLER_255_1488 ();
 FILLCELL_X32 FILLER_255_1520 ();
 FILLCELL_X32 FILLER_255_1552 ();
 FILLCELL_X32 FILLER_255_1584 ();
 FILLCELL_X32 FILLER_255_1616 ();
 FILLCELL_X32 FILLER_255_1648 ();
 FILLCELL_X32 FILLER_255_1680 ();
 FILLCELL_X32 FILLER_255_1712 ();
 FILLCELL_X32 FILLER_255_1744 ();
 FILLCELL_X32 FILLER_255_1776 ();
 FILLCELL_X32 FILLER_255_1808 ();
 FILLCELL_X32 FILLER_255_1840 ();
 FILLCELL_X32 FILLER_255_1872 ();
 FILLCELL_X32 FILLER_255_1904 ();
 FILLCELL_X32 FILLER_255_1936 ();
 FILLCELL_X32 FILLER_255_1968 ();
 FILLCELL_X32 FILLER_255_2000 ();
 FILLCELL_X32 FILLER_255_2032 ();
 FILLCELL_X32 FILLER_255_2064 ();
 FILLCELL_X32 FILLER_255_2096 ();
 FILLCELL_X32 FILLER_255_2128 ();
 FILLCELL_X32 FILLER_255_2160 ();
 FILLCELL_X32 FILLER_255_2192 ();
 FILLCELL_X32 FILLER_255_2224 ();
 FILLCELL_X32 FILLER_255_2256 ();
 FILLCELL_X32 FILLER_255_2288 ();
 FILLCELL_X32 FILLER_255_2320 ();
 FILLCELL_X32 FILLER_255_2352 ();
 FILLCELL_X32 FILLER_255_2384 ();
 FILLCELL_X32 FILLER_255_2416 ();
 FILLCELL_X32 FILLER_255_2448 ();
 FILLCELL_X32 FILLER_255_2480 ();
 FILLCELL_X8 FILLER_255_2512 ();
 FILLCELL_X4 FILLER_255_2520 ();
 FILLCELL_X2 FILLER_255_2524 ();
 FILLCELL_X32 FILLER_255_2527 ();
 FILLCELL_X32 FILLER_255_2559 ();
 FILLCELL_X8 FILLER_255_2591 ();
 FILLCELL_X2 FILLER_255_2599 ();
 FILLCELL_X1 FILLER_255_2601 ();
 FILLCELL_X32 FILLER_256_1 ();
 FILLCELL_X32 FILLER_256_33 ();
 FILLCELL_X32 FILLER_256_65 ();
 FILLCELL_X32 FILLER_256_97 ();
 FILLCELL_X32 FILLER_256_129 ();
 FILLCELL_X32 FILLER_256_161 ();
 FILLCELL_X32 FILLER_256_193 ();
 FILLCELL_X32 FILLER_256_225 ();
 FILLCELL_X32 FILLER_256_257 ();
 FILLCELL_X32 FILLER_256_289 ();
 FILLCELL_X32 FILLER_256_321 ();
 FILLCELL_X32 FILLER_256_353 ();
 FILLCELL_X32 FILLER_256_385 ();
 FILLCELL_X32 FILLER_256_417 ();
 FILLCELL_X32 FILLER_256_449 ();
 FILLCELL_X32 FILLER_256_481 ();
 FILLCELL_X32 FILLER_256_513 ();
 FILLCELL_X32 FILLER_256_545 ();
 FILLCELL_X32 FILLER_256_577 ();
 FILLCELL_X16 FILLER_256_609 ();
 FILLCELL_X4 FILLER_256_625 ();
 FILLCELL_X2 FILLER_256_629 ();
 FILLCELL_X32 FILLER_256_632 ();
 FILLCELL_X32 FILLER_256_664 ();
 FILLCELL_X32 FILLER_256_696 ();
 FILLCELL_X32 FILLER_256_728 ();
 FILLCELL_X32 FILLER_256_760 ();
 FILLCELL_X32 FILLER_256_792 ();
 FILLCELL_X32 FILLER_256_824 ();
 FILLCELL_X32 FILLER_256_856 ();
 FILLCELL_X32 FILLER_256_888 ();
 FILLCELL_X32 FILLER_256_920 ();
 FILLCELL_X32 FILLER_256_952 ();
 FILLCELL_X32 FILLER_256_984 ();
 FILLCELL_X32 FILLER_256_1016 ();
 FILLCELL_X32 FILLER_256_1048 ();
 FILLCELL_X32 FILLER_256_1080 ();
 FILLCELL_X32 FILLER_256_1112 ();
 FILLCELL_X32 FILLER_256_1144 ();
 FILLCELL_X32 FILLER_256_1176 ();
 FILLCELL_X32 FILLER_256_1208 ();
 FILLCELL_X32 FILLER_256_1240 ();
 FILLCELL_X32 FILLER_256_1272 ();
 FILLCELL_X32 FILLER_256_1304 ();
 FILLCELL_X32 FILLER_256_1336 ();
 FILLCELL_X32 FILLER_256_1368 ();
 FILLCELL_X32 FILLER_256_1400 ();
 FILLCELL_X32 FILLER_256_1432 ();
 FILLCELL_X32 FILLER_256_1464 ();
 FILLCELL_X32 FILLER_256_1496 ();
 FILLCELL_X32 FILLER_256_1528 ();
 FILLCELL_X32 FILLER_256_1560 ();
 FILLCELL_X32 FILLER_256_1592 ();
 FILLCELL_X32 FILLER_256_1624 ();
 FILLCELL_X32 FILLER_256_1656 ();
 FILLCELL_X32 FILLER_256_1688 ();
 FILLCELL_X32 FILLER_256_1720 ();
 FILLCELL_X32 FILLER_256_1752 ();
 FILLCELL_X32 FILLER_256_1784 ();
 FILLCELL_X32 FILLER_256_1816 ();
 FILLCELL_X32 FILLER_256_1848 ();
 FILLCELL_X8 FILLER_256_1880 ();
 FILLCELL_X4 FILLER_256_1888 ();
 FILLCELL_X2 FILLER_256_1892 ();
 FILLCELL_X32 FILLER_256_1895 ();
 FILLCELL_X32 FILLER_256_1927 ();
 FILLCELL_X32 FILLER_256_1959 ();
 FILLCELL_X32 FILLER_256_1991 ();
 FILLCELL_X32 FILLER_256_2023 ();
 FILLCELL_X32 FILLER_256_2055 ();
 FILLCELL_X32 FILLER_256_2087 ();
 FILLCELL_X32 FILLER_256_2119 ();
 FILLCELL_X32 FILLER_256_2151 ();
 FILLCELL_X32 FILLER_256_2183 ();
 FILLCELL_X32 FILLER_256_2215 ();
 FILLCELL_X32 FILLER_256_2247 ();
 FILLCELL_X32 FILLER_256_2279 ();
 FILLCELL_X32 FILLER_256_2311 ();
 FILLCELL_X32 FILLER_256_2343 ();
 FILLCELL_X32 FILLER_256_2375 ();
 FILLCELL_X32 FILLER_256_2407 ();
 FILLCELL_X32 FILLER_256_2439 ();
 FILLCELL_X32 FILLER_256_2471 ();
 FILLCELL_X32 FILLER_256_2503 ();
 FILLCELL_X32 FILLER_256_2535 ();
 FILLCELL_X32 FILLER_256_2567 ();
 FILLCELL_X2 FILLER_256_2599 ();
 FILLCELL_X1 FILLER_256_2601 ();
 FILLCELL_X32 FILLER_257_1 ();
 FILLCELL_X32 FILLER_257_33 ();
 FILLCELL_X32 FILLER_257_65 ();
 FILLCELL_X32 FILLER_257_97 ();
 FILLCELL_X32 FILLER_257_129 ();
 FILLCELL_X32 FILLER_257_161 ();
 FILLCELL_X32 FILLER_257_193 ();
 FILLCELL_X32 FILLER_257_225 ();
 FILLCELL_X32 FILLER_257_257 ();
 FILLCELL_X32 FILLER_257_289 ();
 FILLCELL_X32 FILLER_257_321 ();
 FILLCELL_X32 FILLER_257_353 ();
 FILLCELL_X32 FILLER_257_385 ();
 FILLCELL_X32 FILLER_257_417 ();
 FILLCELL_X32 FILLER_257_449 ();
 FILLCELL_X32 FILLER_257_481 ();
 FILLCELL_X32 FILLER_257_513 ();
 FILLCELL_X32 FILLER_257_545 ();
 FILLCELL_X32 FILLER_257_577 ();
 FILLCELL_X32 FILLER_257_609 ();
 FILLCELL_X32 FILLER_257_641 ();
 FILLCELL_X32 FILLER_257_673 ();
 FILLCELL_X32 FILLER_257_705 ();
 FILLCELL_X32 FILLER_257_737 ();
 FILLCELL_X32 FILLER_257_769 ();
 FILLCELL_X32 FILLER_257_801 ();
 FILLCELL_X32 FILLER_257_833 ();
 FILLCELL_X32 FILLER_257_865 ();
 FILLCELL_X32 FILLER_257_897 ();
 FILLCELL_X32 FILLER_257_929 ();
 FILLCELL_X32 FILLER_257_961 ();
 FILLCELL_X32 FILLER_257_993 ();
 FILLCELL_X32 FILLER_257_1025 ();
 FILLCELL_X32 FILLER_257_1057 ();
 FILLCELL_X32 FILLER_257_1089 ();
 FILLCELL_X32 FILLER_257_1121 ();
 FILLCELL_X32 FILLER_257_1153 ();
 FILLCELL_X32 FILLER_257_1185 ();
 FILLCELL_X32 FILLER_257_1217 ();
 FILLCELL_X8 FILLER_257_1249 ();
 FILLCELL_X4 FILLER_257_1257 ();
 FILLCELL_X2 FILLER_257_1261 ();
 FILLCELL_X32 FILLER_257_1264 ();
 FILLCELL_X32 FILLER_257_1296 ();
 FILLCELL_X32 FILLER_257_1328 ();
 FILLCELL_X32 FILLER_257_1360 ();
 FILLCELL_X32 FILLER_257_1392 ();
 FILLCELL_X32 FILLER_257_1424 ();
 FILLCELL_X32 FILLER_257_1456 ();
 FILLCELL_X32 FILLER_257_1488 ();
 FILLCELL_X32 FILLER_257_1520 ();
 FILLCELL_X32 FILLER_257_1552 ();
 FILLCELL_X32 FILLER_257_1584 ();
 FILLCELL_X32 FILLER_257_1616 ();
 FILLCELL_X32 FILLER_257_1648 ();
 FILLCELL_X32 FILLER_257_1680 ();
 FILLCELL_X32 FILLER_257_1712 ();
 FILLCELL_X32 FILLER_257_1744 ();
 FILLCELL_X32 FILLER_257_1776 ();
 FILLCELL_X32 FILLER_257_1808 ();
 FILLCELL_X32 FILLER_257_1840 ();
 FILLCELL_X32 FILLER_257_1872 ();
 FILLCELL_X32 FILLER_257_1904 ();
 FILLCELL_X32 FILLER_257_1936 ();
 FILLCELL_X32 FILLER_257_1968 ();
 FILLCELL_X32 FILLER_257_2000 ();
 FILLCELL_X32 FILLER_257_2032 ();
 FILLCELL_X32 FILLER_257_2064 ();
 FILLCELL_X32 FILLER_257_2096 ();
 FILLCELL_X32 FILLER_257_2128 ();
 FILLCELL_X32 FILLER_257_2160 ();
 FILLCELL_X32 FILLER_257_2192 ();
 FILLCELL_X32 FILLER_257_2224 ();
 FILLCELL_X32 FILLER_257_2256 ();
 FILLCELL_X32 FILLER_257_2288 ();
 FILLCELL_X32 FILLER_257_2320 ();
 FILLCELL_X32 FILLER_257_2352 ();
 FILLCELL_X32 FILLER_257_2384 ();
 FILLCELL_X32 FILLER_257_2416 ();
 FILLCELL_X32 FILLER_257_2448 ();
 FILLCELL_X32 FILLER_257_2480 ();
 FILLCELL_X8 FILLER_257_2512 ();
 FILLCELL_X4 FILLER_257_2520 ();
 FILLCELL_X2 FILLER_257_2524 ();
 FILLCELL_X32 FILLER_257_2527 ();
 FILLCELL_X32 FILLER_257_2559 ();
 FILLCELL_X8 FILLER_257_2591 ();
 FILLCELL_X2 FILLER_257_2599 ();
 FILLCELL_X1 FILLER_257_2601 ();
 FILLCELL_X32 FILLER_258_1 ();
 FILLCELL_X32 FILLER_258_33 ();
 FILLCELL_X32 FILLER_258_65 ();
 FILLCELL_X32 FILLER_258_97 ();
 FILLCELL_X32 FILLER_258_129 ();
 FILLCELL_X32 FILLER_258_161 ();
 FILLCELL_X32 FILLER_258_193 ();
 FILLCELL_X32 FILLER_258_225 ();
 FILLCELL_X32 FILLER_258_257 ();
 FILLCELL_X32 FILLER_258_289 ();
 FILLCELL_X32 FILLER_258_321 ();
 FILLCELL_X32 FILLER_258_353 ();
 FILLCELL_X32 FILLER_258_385 ();
 FILLCELL_X32 FILLER_258_417 ();
 FILLCELL_X32 FILLER_258_449 ();
 FILLCELL_X32 FILLER_258_481 ();
 FILLCELL_X32 FILLER_258_513 ();
 FILLCELL_X32 FILLER_258_545 ();
 FILLCELL_X32 FILLER_258_577 ();
 FILLCELL_X16 FILLER_258_609 ();
 FILLCELL_X4 FILLER_258_625 ();
 FILLCELL_X2 FILLER_258_629 ();
 FILLCELL_X32 FILLER_258_632 ();
 FILLCELL_X32 FILLER_258_664 ();
 FILLCELL_X32 FILLER_258_696 ();
 FILLCELL_X32 FILLER_258_728 ();
 FILLCELL_X32 FILLER_258_760 ();
 FILLCELL_X32 FILLER_258_792 ();
 FILLCELL_X32 FILLER_258_824 ();
 FILLCELL_X32 FILLER_258_856 ();
 FILLCELL_X32 FILLER_258_888 ();
 FILLCELL_X32 FILLER_258_920 ();
 FILLCELL_X32 FILLER_258_952 ();
 FILLCELL_X32 FILLER_258_984 ();
 FILLCELL_X32 FILLER_258_1016 ();
 FILLCELL_X32 FILLER_258_1048 ();
 FILLCELL_X32 FILLER_258_1080 ();
 FILLCELL_X32 FILLER_258_1112 ();
 FILLCELL_X32 FILLER_258_1144 ();
 FILLCELL_X32 FILLER_258_1176 ();
 FILLCELL_X32 FILLER_258_1208 ();
 FILLCELL_X32 FILLER_258_1240 ();
 FILLCELL_X32 FILLER_258_1272 ();
 FILLCELL_X32 FILLER_258_1304 ();
 FILLCELL_X32 FILLER_258_1336 ();
 FILLCELL_X32 FILLER_258_1368 ();
 FILLCELL_X32 FILLER_258_1400 ();
 FILLCELL_X32 FILLER_258_1432 ();
 FILLCELL_X32 FILLER_258_1464 ();
 FILLCELL_X32 FILLER_258_1496 ();
 FILLCELL_X32 FILLER_258_1528 ();
 FILLCELL_X32 FILLER_258_1560 ();
 FILLCELL_X32 FILLER_258_1592 ();
 FILLCELL_X32 FILLER_258_1624 ();
 FILLCELL_X32 FILLER_258_1656 ();
 FILLCELL_X32 FILLER_258_1688 ();
 FILLCELL_X32 FILLER_258_1720 ();
 FILLCELL_X32 FILLER_258_1752 ();
 FILLCELL_X32 FILLER_258_1784 ();
 FILLCELL_X32 FILLER_258_1816 ();
 FILLCELL_X32 FILLER_258_1848 ();
 FILLCELL_X8 FILLER_258_1880 ();
 FILLCELL_X4 FILLER_258_1888 ();
 FILLCELL_X2 FILLER_258_1892 ();
 FILLCELL_X32 FILLER_258_1895 ();
 FILLCELL_X32 FILLER_258_1927 ();
 FILLCELL_X32 FILLER_258_1959 ();
 FILLCELL_X32 FILLER_258_1991 ();
 FILLCELL_X32 FILLER_258_2023 ();
 FILLCELL_X32 FILLER_258_2055 ();
 FILLCELL_X32 FILLER_258_2087 ();
 FILLCELL_X32 FILLER_258_2119 ();
 FILLCELL_X32 FILLER_258_2151 ();
 FILLCELL_X32 FILLER_258_2183 ();
 FILLCELL_X32 FILLER_258_2215 ();
 FILLCELL_X32 FILLER_258_2247 ();
 FILLCELL_X32 FILLER_258_2279 ();
 FILLCELL_X32 FILLER_258_2311 ();
 FILLCELL_X32 FILLER_258_2343 ();
 FILLCELL_X32 FILLER_258_2375 ();
 FILLCELL_X32 FILLER_258_2407 ();
 FILLCELL_X32 FILLER_258_2439 ();
 FILLCELL_X32 FILLER_258_2471 ();
 FILLCELL_X32 FILLER_258_2503 ();
 FILLCELL_X32 FILLER_258_2535 ();
 FILLCELL_X32 FILLER_258_2567 ();
 FILLCELL_X2 FILLER_258_2599 ();
 FILLCELL_X1 FILLER_258_2601 ();
 FILLCELL_X32 FILLER_259_1 ();
 FILLCELL_X32 FILLER_259_33 ();
 FILLCELL_X32 FILLER_259_65 ();
 FILLCELL_X32 FILLER_259_97 ();
 FILLCELL_X32 FILLER_259_129 ();
 FILLCELL_X32 FILLER_259_161 ();
 FILLCELL_X32 FILLER_259_193 ();
 FILLCELL_X32 FILLER_259_225 ();
 FILLCELL_X32 FILLER_259_257 ();
 FILLCELL_X32 FILLER_259_289 ();
 FILLCELL_X32 FILLER_259_321 ();
 FILLCELL_X32 FILLER_259_353 ();
 FILLCELL_X32 FILLER_259_385 ();
 FILLCELL_X32 FILLER_259_417 ();
 FILLCELL_X32 FILLER_259_449 ();
 FILLCELL_X32 FILLER_259_481 ();
 FILLCELL_X32 FILLER_259_513 ();
 FILLCELL_X32 FILLER_259_545 ();
 FILLCELL_X32 FILLER_259_577 ();
 FILLCELL_X32 FILLER_259_609 ();
 FILLCELL_X32 FILLER_259_641 ();
 FILLCELL_X32 FILLER_259_673 ();
 FILLCELL_X32 FILLER_259_705 ();
 FILLCELL_X32 FILLER_259_737 ();
 FILLCELL_X32 FILLER_259_769 ();
 FILLCELL_X32 FILLER_259_801 ();
 FILLCELL_X32 FILLER_259_833 ();
 FILLCELL_X32 FILLER_259_865 ();
 FILLCELL_X32 FILLER_259_897 ();
 FILLCELL_X32 FILLER_259_929 ();
 FILLCELL_X32 FILLER_259_961 ();
 FILLCELL_X32 FILLER_259_993 ();
 FILLCELL_X32 FILLER_259_1025 ();
 FILLCELL_X32 FILLER_259_1057 ();
 FILLCELL_X32 FILLER_259_1089 ();
 FILLCELL_X32 FILLER_259_1121 ();
 FILLCELL_X32 FILLER_259_1153 ();
 FILLCELL_X32 FILLER_259_1185 ();
 FILLCELL_X32 FILLER_259_1217 ();
 FILLCELL_X8 FILLER_259_1249 ();
 FILLCELL_X4 FILLER_259_1257 ();
 FILLCELL_X2 FILLER_259_1261 ();
 FILLCELL_X32 FILLER_259_1264 ();
 FILLCELL_X32 FILLER_259_1296 ();
 FILLCELL_X32 FILLER_259_1328 ();
 FILLCELL_X32 FILLER_259_1360 ();
 FILLCELL_X32 FILLER_259_1392 ();
 FILLCELL_X32 FILLER_259_1424 ();
 FILLCELL_X32 FILLER_259_1456 ();
 FILLCELL_X32 FILLER_259_1488 ();
 FILLCELL_X32 FILLER_259_1520 ();
 FILLCELL_X32 FILLER_259_1552 ();
 FILLCELL_X32 FILLER_259_1584 ();
 FILLCELL_X32 FILLER_259_1616 ();
 FILLCELL_X32 FILLER_259_1648 ();
 FILLCELL_X32 FILLER_259_1680 ();
 FILLCELL_X32 FILLER_259_1712 ();
 FILLCELL_X32 FILLER_259_1744 ();
 FILLCELL_X32 FILLER_259_1776 ();
 FILLCELL_X32 FILLER_259_1808 ();
 FILLCELL_X32 FILLER_259_1840 ();
 FILLCELL_X32 FILLER_259_1872 ();
 FILLCELL_X32 FILLER_259_1904 ();
 FILLCELL_X32 FILLER_259_1936 ();
 FILLCELL_X32 FILLER_259_1968 ();
 FILLCELL_X32 FILLER_259_2000 ();
 FILLCELL_X32 FILLER_259_2032 ();
 FILLCELL_X32 FILLER_259_2064 ();
 FILLCELL_X32 FILLER_259_2096 ();
 FILLCELL_X32 FILLER_259_2128 ();
 FILLCELL_X32 FILLER_259_2160 ();
 FILLCELL_X32 FILLER_259_2192 ();
 FILLCELL_X32 FILLER_259_2224 ();
 FILLCELL_X32 FILLER_259_2256 ();
 FILLCELL_X32 FILLER_259_2288 ();
 FILLCELL_X32 FILLER_259_2320 ();
 FILLCELL_X32 FILLER_259_2352 ();
 FILLCELL_X32 FILLER_259_2384 ();
 FILLCELL_X32 FILLER_259_2416 ();
 FILLCELL_X32 FILLER_259_2448 ();
 FILLCELL_X32 FILLER_259_2480 ();
 FILLCELL_X8 FILLER_259_2512 ();
 FILLCELL_X4 FILLER_259_2520 ();
 FILLCELL_X2 FILLER_259_2524 ();
 FILLCELL_X32 FILLER_259_2527 ();
 FILLCELL_X32 FILLER_259_2559 ();
 FILLCELL_X8 FILLER_259_2591 ();
 FILLCELL_X2 FILLER_259_2599 ();
 FILLCELL_X1 FILLER_259_2601 ();
 FILLCELL_X32 FILLER_260_1 ();
 FILLCELL_X32 FILLER_260_33 ();
 FILLCELL_X32 FILLER_260_65 ();
 FILLCELL_X32 FILLER_260_97 ();
 FILLCELL_X32 FILLER_260_129 ();
 FILLCELL_X32 FILLER_260_161 ();
 FILLCELL_X32 FILLER_260_193 ();
 FILLCELL_X32 FILLER_260_225 ();
 FILLCELL_X32 FILLER_260_257 ();
 FILLCELL_X32 FILLER_260_289 ();
 FILLCELL_X32 FILLER_260_321 ();
 FILLCELL_X32 FILLER_260_353 ();
 FILLCELL_X32 FILLER_260_385 ();
 FILLCELL_X32 FILLER_260_417 ();
 FILLCELL_X32 FILLER_260_449 ();
 FILLCELL_X32 FILLER_260_481 ();
 FILLCELL_X32 FILLER_260_513 ();
 FILLCELL_X32 FILLER_260_545 ();
 FILLCELL_X32 FILLER_260_577 ();
 FILLCELL_X16 FILLER_260_609 ();
 FILLCELL_X4 FILLER_260_625 ();
 FILLCELL_X2 FILLER_260_629 ();
 FILLCELL_X32 FILLER_260_632 ();
 FILLCELL_X32 FILLER_260_664 ();
 FILLCELL_X32 FILLER_260_696 ();
 FILLCELL_X32 FILLER_260_728 ();
 FILLCELL_X32 FILLER_260_760 ();
 FILLCELL_X32 FILLER_260_792 ();
 FILLCELL_X32 FILLER_260_824 ();
 FILLCELL_X32 FILLER_260_856 ();
 FILLCELL_X32 FILLER_260_888 ();
 FILLCELL_X32 FILLER_260_920 ();
 FILLCELL_X32 FILLER_260_952 ();
 FILLCELL_X32 FILLER_260_984 ();
 FILLCELL_X32 FILLER_260_1016 ();
 FILLCELL_X32 FILLER_260_1048 ();
 FILLCELL_X32 FILLER_260_1080 ();
 FILLCELL_X32 FILLER_260_1112 ();
 FILLCELL_X32 FILLER_260_1144 ();
 FILLCELL_X32 FILLER_260_1176 ();
 FILLCELL_X32 FILLER_260_1208 ();
 FILLCELL_X32 FILLER_260_1240 ();
 FILLCELL_X32 FILLER_260_1272 ();
 FILLCELL_X32 FILLER_260_1304 ();
 FILLCELL_X32 FILLER_260_1336 ();
 FILLCELL_X32 FILLER_260_1368 ();
 FILLCELL_X32 FILLER_260_1400 ();
 FILLCELL_X32 FILLER_260_1432 ();
 FILLCELL_X32 FILLER_260_1464 ();
 FILLCELL_X32 FILLER_260_1496 ();
 FILLCELL_X32 FILLER_260_1528 ();
 FILLCELL_X32 FILLER_260_1560 ();
 FILLCELL_X32 FILLER_260_1592 ();
 FILLCELL_X32 FILLER_260_1624 ();
 FILLCELL_X32 FILLER_260_1656 ();
 FILLCELL_X32 FILLER_260_1688 ();
 FILLCELL_X32 FILLER_260_1720 ();
 FILLCELL_X32 FILLER_260_1752 ();
 FILLCELL_X32 FILLER_260_1784 ();
 FILLCELL_X32 FILLER_260_1816 ();
 FILLCELL_X32 FILLER_260_1848 ();
 FILLCELL_X8 FILLER_260_1880 ();
 FILLCELL_X4 FILLER_260_1888 ();
 FILLCELL_X2 FILLER_260_1892 ();
 FILLCELL_X32 FILLER_260_1895 ();
 FILLCELL_X32 FILLER_260_1927 ();
 FILLCELL_X32 FILLER_260_1959 ();
 FILLCELL_X32 FILLER_260_1991 ();
 FILLCELL_X32 FILLER_260_2023 ();
 FILLCELL_X32 FILLER_260_2055 ();
 FILLCELL_X32 FILLER_260_2087 ();
 FILLCELL_X32 FILLER_260_2119 ();
 FILLCELL_X32 FILLER_260_2151 ();
 FILLCELL_X32 FILLER_260_2183 ();
 FILLCELL_X32 FILLER_260_2215 ();
 FILLCELL_X32 FILLER_260_2247 ();
 FILLCELL_X32 FILLER_260_2279 ();
 FILLCELL_X32 FILLER_260_2311 ();
 FILLCELL_X32 FILLER_260_2343 ();
 FILLCELL_X32 FILLER_260_2375 ();
 FILLCELL_X32 FILLER_260_2407 ();
 FILLCELL_X32 FILLER_260_2439 ();
 FILLCELL_X32 FILLER_260_2471 ();
 FILLCELL_X32 FILLER_260_2503 ();
 FILLCELL_X32 FILLER_260_2535 ();
 FILLCELL_X32 FILLER_260_2567 ();
 FILLCELL_X2 FILLER_260_2599 ();
 FILLCELL_X1 FILLER_260_2601 ();
 FILLCELL_X32 FILLER_261_1 ();
 FILLCELL_X32 FILLER_261_33 ();
 FILLCELL_X32 FILLER_261_65 ();
 FILLCELL_X32 FILLER_261_97 ();
 FILLCELL_X32 FILLER_261_129 ();
 FILLCELL_X32 FILLER_261_161 ();
 FILLCELL_X32 FILLER_261_193 ();
 FILLCELL_X32 FILLER_261_225 ();
 FILLCELL_X32 FILLER_261_257 ();
 FILLCELL_X32 FILLER_261_289 ();
 FILLCELL_X32 FILLER_261_321 ();
 FILLCELL_X32 FILLER_261_353 ();
 FILLCELL_X32 FILLER_261_385 ();
 FILLCELL_X32 FILLER_261_417 ();
 FILLCELL_X32 FILLER_261_449 ();
 FILLCELL_X32 FILLER_261_481 ();
 FILLCELL_X32 FILLER_261_513 ();
 FILLCELL_X32 FILLER_261_545 ();
 FILLCELL_X32 FILLER_261_577 ();
 FILLCELL_X32 FILLER_261_609 ();
 FILLCELL_X32 FILLER_261_641 ();
 FILLCELL_X32 FILLER_261_673 ();
 FILLCELL_X32 FILLER_261_705 ();
 FILLCELL_X32 FILLER_261_737 ();
 FILLCELL_X32 FILLER_261_769 ();
 FILLCELL_X32 FILLER_261_801 ();
 FILLCELL_X32 FILLER_261_833 ();
 FILLCELL_X32 FILLER_261_865 ();
 FILLCELL_X32 FILLER_261_897 ();
 FILLCELL_X32 FILLER_261_929 ();
 FILLCELL_X32 FILLER_261_961 ();
 FILLCELL_X32 FILLER_261_993 ();
 FILLCELL_X32 FILLER_261_1025 ();
 FILLCELL_X32 FILLER_261_1057 ();
 FILLCELL_X32 FILLER_261_1089 ();
 FILLCELL_X32 FILLER_261_1121 ();
 FILLCELL_X32 FILLER_261_1153 ();
 FILLCELL_X32 FILLER_261_1185 ();
 FILLCELL_X32 FILLER_261_1217 ();
 FILLCELL_X8 FILLER_261_1249 ();
 FILLCELL_X4 FILLER_261_1257 ();
 FILLCELL_X2 FILLER_261_1261 ();
 FILLCELL_X32 FILLER_261_1264 ();
 FILLCELL_X32 FILLER_261_1296 ();
 FILLCELL_X32 FILLER_261_1328 ();
 FILLCELL_X32 FILLER_261_1360 ();
 FILLCELL_X32 FILLER_261_1392 ();
 FILLCELL_X32 FILLER_261_1424 ();
 FILLCELL_X32 FILLER_261_1456 ();
 FILLCELL_X32 FILLER_261_1488 ();
 FILLCELL_X32 FILLER_261_1520 ();
 FILLCELL_X32 FILLER_261_1552 ();
 FILLCELL_X32 FILLER_261_1584 ();
 FILLCELL_X32 FILLER_261_1616 ();
 FILLCELL_X32 FILLER_261_1648 ();
 FILLCELL_X32 FILLER_261_1680 ();
 FILLCELL_X32 FILLER_261_1712 ();
 FILLCELL_X32 FILLER_261_1744 ();
 FILLCELL_X32 FILLER_261_1776 ();
 FILLCELL_X32 FILLER_261_1808 ();
 FILLCELL_X32 FILLER_261_1840 ();
 FILLCELL_X32 FILLER_261_1872 ();
 FILLCELL_X32 FILLER_261_1904 ();
 FILLCELL_X32 FILLER_261_1936 ();
 FILLCELL_X32 FILLER_261_1968 ();
 FILLCELL_X32 FILLER_261_2000 ();
 FILLCELL_X32 FILLER_261_2032 ();
 FILLCELL_X32 FILLER_261_2064 ();
 FILLCELL_X32 FILLER_261_2096 ();
 FILLCELL_X32 FILLER_261_2128 ();
 FILLCELL_X32 FILLER_261_2160 ();
 FILLCELL_X32 FILLER_261_2192 ();
 FILLCELL_X32 FILLER_261_2224 ();
 FILLCELL_X32 FILLER_261_2256 ();
 FILLCELL_X32 FILLER_261_2288 ();
 FILLCELL_X32 FILLER_261_2320 ();
 FILLCELL_X32 FILLER_261_2352 ();
 FILLCELL_X32 FILLER_261_2384 ();
 FILLCELL_X32 FILLER_261_2416 ();
 FILLCELL_X32 FILLER_261_2448 ();
 FILLCELL_X32 FILLER_261_2480 ();
 FILLCELL_X8 FILLER_261_2512 ();
 FILLCELL_X4 FILLER_261_2520 ();
 FILLCELL_X2 FILLER_261_2524 ();
 FILLCELL_X32 FILLER_261_2527 ();
 FILLCELL_X32 FILLER_261_2559 ();
 FILLCELL_X8 FILLER_261_2591 ();
 FILLCELL_X2 FILLER_261_2599 ();
 FILLCELL_X1 FILLER_261_2601 ();
 FILLCELL_X32 FILLER_262_1 ();
 FILLCELL_X32 FILLER_262_33 ();
 FILLCELL_X32 FILLER_262_65 ();
 FILLCELL_X32 FILLER_262_97 ();
 FILLCELL_X32 FILLER_262_129 ();
 FILLCELL_X32 FILLER_262_161 ();
 FILLCELL_X32 FILLER_262_193 ();
 FILLCELL_X32 FILLER_262_225 ();
 FILLCELL_X32 FILLER_262_257 ();
 FILLCELL_X32 FILLER_262_289 ();
 FILLCELL_X32 FILLER_262_321 ();
 FILLCELL_X32 FILLER_262_353 ();
 FILLCELL_X32 FILLER_262_385 ();
 FILLCELL_X32 FILLER_262_417 ();
 FILLCELL_X32 FILLER_262_449 ();
 FILLCELL_X32 FILLER_262_481 ();
 FILLCELL_X32 FILLER_262_513 ();
 FILLCELL_X32 FILLER_262_545 ();
 FILLCELL_X32 FILLER_262_577 ();
 FILLCELL_X16 FILLER_262_609 ();
 FILLCELL_X4 FILLER_262_625 ();
 FILLCELL_X2 FILLER_262_629 ();
 FILLCELL_X32 FILLER_262_632 ();
 FILLCELL_X32 FILLER_262_664 ();
 FILLCELL_X32 FILLER_262_696 ();
 FILLCELL_X32 FILLER_262_728 ();
 FILLCELL_X32 FILLER_262_760 ();
 FILLCELL_X32 FILLER_262_792 ();
 FILLCELL_X32 FILLER_262_824 ();
 FILLCELL_X32 FILLER_262_856 ();
 FILLCELL_X32 FILLER_262_888 ();
 FILLCELL_X32 FILLER_262_920 ();
 FILLCELL_X32 FILLER_262_952 ();
 FILLCELL_X32 FILLER_262_984 ();
 FILLCELL_X32 FILLER_262_1016 ();
 FILLCELL_X32 FILLER_262_1048 ();
 FILLCELL_X32 FILLER_262_1080 ();
 FILLCELL_X32 FILLER_262_1112 ();
 FILLCELL_X32 FILLER_262_1144 ();
 FILLCELL_X32 FILLER_262_1176 ();
 FILLCELL_X32 FILLER_262_1208 ();
 FILLCELL_X32 FILLER_262_1240 ();
 FILLCELL_X32 FILLER_262_1272 ();
 FILLCELL_X32 FILLER_262_1304 ();
 FILLCELL_X32 FILLER_262_1336 ();
 FILLCELL_X32 FILLER_262_1368 ();
 FILLCELL_X32 FILLER_262_1400 ();
 FILLCELL_X32 FILLER_262_1432 ();
 FILLCELL_X32 FILLER_262_1464 ();
 FILLCELL_X32 FILLER_262_1496 ();
 FILLCELL_X32 FILLER_262_1528 ();
 FILLCELL_X32 FILLER_262_1560 ();
 FILLCELL_X32 FILLER_262_1592 ();
 FILLCELL_X32 FILLER_262_1624 ();
 FILLCELL_X32 FILLER_262_1656 ();
 FILLCELL_X32 FILLER_262_1688 ();
 FILLCELL_X32 FILLER_262_1720 ();
 FILLCELL_X32 FILLER_262_1752 ();
 FILLCELL_X32 FILLER_262_1784 ();
 FILLCELL_X32 FILLER_262_1816 ();
 FILLCELL_X32 FILLER_262_1848 ();
 FILLCELL_X8 FILLER_262_1880 ();
 FILLCELL_X4 FILLER_262_1888 ();
 FILLCELL_X2 FILLER_262_1892 ();
 FILLCELL_X32 FILLER_262_1895 ();
 FILLCELL_X32 FILLER_262_1927 ();
 FILLCELL_X32 FILLER_262_1959 ();
 FILLCELL_X32 FILLER_262_1991 ();
 FILLCELL_X32 FILLER_262_2023 ();
 FILLCELL_X32 FILLER_262_2055 ();
 FILLCELL_X32 FILLER_262_2087 ();
 FILLCELL_X32 FILLER_262_2119 ();
 FILLCELL_X32 FILLER_262_2151 ();
 FILLCELL_X32 FILLER_262_2183 ();
 FILLCELL_X32 FILLER_262_2215 ();
 FILLCELL_X32 FILLER_262_2247 ();
 FILLCELL_X32 FILLER_262_2279 ();
 FILLCELL_X32 FILLER_262_2311 ();
 FILLCELL_X32 FILLER_262_2343 ();
 FILLCELL_X32 FILLER_262_2375 ();
 FILLCELL_X32 FILLER_262_2407 ();
 FILLCELL_X32 FILLER_262_2439 ();
 FILLCELL_X32 FILLER_262_2471 ();
 FILLCELL_X32 FILLER_262_2503 ();
 FILLCELL_X32 FILLER_262_2535 ();
 FILLCELL_X32 FILLER_262_2567 ();
 FILLCELL_X2 FILLER_262_2599 ();
 FILLCELL_X1 FILLER_262_2601 ();
 FILLCELL_X32 FILLER_263_1 ();
 FILLCELL_X32 FILLER_263_33 ();
 FILLCELL_X32 FILLER_263_65 ();
 FILLCELL_X32 FILLER_263_97 ();
 FILLCELL_X32 FILLER_263_129 ();
 FILLCELL_X32 FILLER_263_161 ();
 FILLCELL_X32 FILLER_263_193 ();
 FILLCELL_X32 FILLER_263_225 ();
 FILLCELL_X32 FILLER_263_257 ();
 FILLCELL_X32 FILLER_263_289 ();
 FILLCELL_X32 FILLER_263_321 ();
 FILLCELL_X32 FILLER_263_353 ();
 FILLCELL_X32 FILLER_263_385 ();
 FILLCELL_X32 FILLER_263_417 ();
 FILLCELL_X32 FILLER_263_449 ();
 FILLCELL_X32 FILLER_263_481 ();
 FILLCELL_X32 FILLER_263_513 ();
 FILLCELL_X32 FILLER_263_545 ();
 FILLCELL_X32 FILLER_263_577 ();
 FILLCELL_X32 FILLER_263_609 ();
 FILLCELL_X32 FILLER_263_641 ();
 FILLCELL_X32 FILLER_263_673 ();
 FILLCELL_X32 FILLER_263_705 ();
 FILLCELL_X32 FILLER_263_737 ();
 FILLCELL_X32 FILLER_263_769 ();
 FILLCELL_X32 FILLER_263_801 ();
 FILLCELL_X32 FILLER_263_833 ();
 FILLCELL_X32 FILLER_263_865 ();
 FILLCELL_X32 FILLER_263_897 ();
 FILLCELL_X32 FILLER_263_929 ();
 FILLCELL_X32 FILLER_263_961 ();
 FILLCELL_X32 FILLER_263_993 ();
 FILLCELL_X32 FILLER_263_1025 ();
 FILLCELL_X32 FILLER_263_1057 ();
 FILLCELL_X32 FILLER_263_1089 ();
 FILLCELL_X32 FILLER_263_1121 ();
 FILLCELL_X32 FILLER_263_1153 ();
 FILLCELL_X32 FILLER_263_1185 ();
 FILLCELL_X32 FILLER_263_1217 ();
 FILLCELL_X8 FILLER_263_1249 ();
 FILLCELL_X4 FILLER_263_1257 ();
 FILLCELL_X2 FILLER_263_1261 ();
 FILLCELL_X32 FILLER_263_1264 ();
 FILLCELL_X32 FILLER_263_1296 ();
 FILLCELL_X32 FILLER_263_1328 ();
 FILLCELL_X32 FILLER_263_1360 ();
 FILLCELL_X32 FILLER_263_1392 ();
 FILLCELL_X32 FILLER_263_1424 ();
 FILLCELL_X32 FILLER_263_1456 ();
 FILLCELL_X32 FILLER_263_1488 ();
 FILLCELL_X32 FILLER_263_1520 ();
 FILLCELL_X32 FILLER_263_1552 ();
 FILLCELL_X32 FILLER_263_1584 ();
 FILLCELL_X32 FILLER_263_1616 ();
 FILLCELL_X32 FILLER_263_1648 ();
 FILLCELL_X32 FILLER_263_1680 ();
 FILLCELL_X32 FILLER_263_1712 ();
 FILLCELL_X32 FILLER_263_1744 ();
 FILLCELL_X32 FILLER_263_1776 ();
 FILLCELL_X32 FILLER_263_1808 ();
 FILLCELL_X32 FILLER_263_1840 ();
 FILLCELL_X32 FILLER_263_1872 ();
 FILLCELL_X32 FILLER_263_1904 ();
 FILLCELL_X32 FILLER_263_1936 ();
 FILLCELL_X32 FILLER_263_1968 ();
 FILLCELL_X32 FILLER_263_2000 ();
 FILLCELL_X32 FILLER_263_2032 ();
 FILLCELL_X32 FILLER_263_2064 ();
 FILLCELL_X32 FILLER_263_2096 ();
 FILLCELL_X32 FILLER_263_2128 ();
 FILLCELL_X32 FILLER_263_2160 ();
 FILLCELL_X32 FILLER_263_2192 ();
 FILLCELL_X32 FILLER_263_2224 ();
 FILLCELL_X32 FILLER_263_2256 ();
 FILLCELL_X32 FILLER_263_2288 ();
 FILLCELL_X32 FILLER_263_2320 ();
 FILLCELL_X32 FILLER_263_2352 ();
 FILLCELL_X32 FILLER_263_2384 ();
 FILLCELL_X32 FILLER_263_2416 ();
 FILLCELL_X32 FILLER_263_2448 ();
 FILLCELL_X32 FILLER_263_2480 ();
 FILLCELL_X8 FILLER_263_2512 ();
 FILLCELL_X4 FILLER_263_2520 ();
 FILLCELL_X2 FILLER_263_2524 ();
 FILLCELL_X32 FILLER_263_2527 ();
 FILLCELL_X32 FILLER_263_2559 ();
 FILLCELL_X8 FILLER_263_2591 ();
 FILLCELL_X2 FILLER_263_2599 ();
 FILLCELL_X1 FILLER_263_2601 ();
 FILLCELL_X32 FILLER_264_1 ();
 FILLCELL_X32 FILLER_264_33 ();
 FILLCELL_X32 FILLER_264_65 ();
 FILLCELL_X32 FILLER_264_97 ();
 FILLCELL_X32 FILLER_264_129 ();
 FILLCELL_X32 FILLER_264_161 ();
 FILLCELL_X32 FILLER_264_193 ();
 FILLCELL_X32 FILLER_264_225 ();
 FILLCELL_X32 FILLER_264_257 ();
 FILLCELL_X32 FILLER_264_289 ();
 FILLCELL_X32 FILLER_264_321 ();
 FILLCELL_X32 FILLER_264_353 ();
 FILLCELL_X32 FILLER_264_385 ();
 FILLCELL_X32 FILLER_264_417 ();
 FILLCELL_X32 FILLER_264_449 ();
 FILLCELL_X32 FILLER_264_481 ();
 FILLCELL_X32 FILLER_264_513 ();
 FILLCELL_X32 FILLER_264_545 ();
 FILLCELL_X32 FILLER_264_577 ();
 FILLCELL_X16 FILLER_264_609 ();
 FILLCELL_X4 FILLER_264_625 ();
 FILLCELL_X2 FILLER_264_629 ();
 FILLCELL_X32 FILLER_264_632 ();
 FILLCELL_X32 FILLER_264_664 ();
 FILLCELL_X32 FILLER_264_696 ();
 FILLCELL_X32 FILLER_264_728 ();
 FILLCELL_X32 FILLER_264_760 ();
 FILLCELL_X32 FILLER_264_792 ();
 FILLCELL_X32 FILLER_264_824 ();
 FILLCELL_X32 FILLER_264_856 ();
 FILLCELL_X32 FILLER_264_888 ();
 FILLCELL_X32 FILLER_264_920 ();
 FILLCELL_X32 FILLER_264_952 ();
 FILLCELL_X32 FILLER_264_984 ();
 FILLCELL_X32 FILLER_264_1016 ();
 FILLCELL_X32 FILLER_264_1048 ();
 FILLCELL_X32 FILLER_264_1080 ();
 FILLCELL_X32 FILLER_264_1112 ();
 FILLCELL_X32 FILLER_264_1144 ();
 FILLCELL_X32 FILLER_264_1176 ();
 FILLCELL_X32 FILLER_264_1208 ();
 FILLCELL_X32 FILLER_264_1240 ();
 FILLCELL_X32 FILLER_264_1272 ();
 FILLCELL_X32 FILLER_264_1304 ();
 FILLCELL_X32 FILLER_264_1336 ();
 FILLCELL_X32 FILLER_264_1368 ();
 FILLCELL_X32 FILLER_264_1400 ();
 FILLCELL_X32 FILLER_264_1432 ();
 FILLCELL_X32 FILLER_264_1464 ();
 FILLCELL_X32 FILLER_264_1496 ();
 FILLCELL_X32 FILLER_264_1528 ();
 FILLCELL_X32 FILLER_264_1560 ();
 FILLCELL_X32 FILLER_264_1592 ();
 FILLCELL_X32 FILLER_264_1624 ();
 FILLCELL_X32 FILLER_264_1656 ();
 FILLCELL_X32 FILLER_264_1688 ();
 FILLCELL_X32 FILLER_264_1720 ();
 FILLCELL_X32 FILLER_264_1752 ();
 FILLCELL_X32 FILLER_264_1784 ();
 FILLCELL_X32 FILLER_264_1816 ();
 FILLCELL_X32 FILLER_264_1848 ();
 FILLCELL_X8 FILLER_264_1880 ();
 FILLCELL_X4 FILLER_264_1888 ();
 FILLCELL_X2 FILLER_264_1892 ();
 FILLCELL_X32 FILLER_264_1895 ();
 FILLCELL_X32 FILLER_264_1927 ();
 FILLCELL_X32 FILLER_264_1959 ();
 FILLCELL_X32 FILLER_264_1991 ();
 FILLCELL_X32 FILLER_264_2023 ();
 FILLCELL_X32 FILLER_264_2055 ();
 FILLCELL_X32 FILLER_264_2087 ();
 FILLCELL_X32 FILLER_264_2119 ();
 FILLCELL_X32 FILLER_264_2151 ();
 FILLCELL_X32 FILLER_264_2183 ();
 FILLCELL_X32 FILLER_264_2215 ();
 FILLCELL_X32 FILLER_264_2247 ();
 FILLCELL_X32 FILLER_264_2279 ();
 FILLCELL_X32 FILLER_264_2311 ();
 FILLCELL_X32 FILLER_264_2343 ();
 FILLCELL_X32 FILLER_264_2375 ();
 FILLCELL_X32 FILLER_264_2407 ();
 FILLCELL_X32 FILLER_264_2439 ();
 FILLCELL_X32 FILLER_264_2471 ();
 FILLCELL_X32 FILLER_264_2503 ();
 FILLCELL_X32 FILLER_264_2535 ();
 FILLCELL_X32 FILLER_264_2567 ();
 FILLCELL_X2 FILLER_264_2599 ();
 FILLCELL_X1 FILLER_264_2601 ();
 FILLCELL_X32 FILLER_265_1 ();
 FILLCELL_X32 FILLER_265_33 ();
 FILLCELL_X32 FILLER_265_65 ();
 FILLCELL_X32 FILLER_265_97 ();
 FILLCELL_X32 FILLER_265_129 ();
 FILLCELL_X32 FILLER_265_161 ();
 FILLCELL_X32 FILLER_265_193 ();
 FILLCELL_X32 FILLER_265_225 ();
 FILLCELL_X32 FILLER_265_257 ();
 FILLCELL_X32 FILLER_265_289 ();
 FILLCELL_X32 FILLER_265_321 ();
 FILLCELL_X32 FILLER_265_353 ();
 FILLCELL_X32 FILLER_265_385 ();
 FILLCELL_X32 FILLER_265_417 ();
 FILLCELL_X32 FILLER_265_449 ();
 FILLCELL_X32 FILLER_265_481 ();
 FILLCELL_X32 FILLER_265_513 ();
 FILLCELL_X32 FILLER_265_545 ();
 FILLCELL_X32 FILLER_265_577 ();
 FILLCELL_X32 FILLER_265_609 ();
 FILLCELL_X32 FILLER_265_641 ();
 FILLCELL_X32 FILLER_265_673 ();
 FILLCELL_X32 FILLER_265_705 ();
 FILLCELL_X32 FILLER_265_737 ();
 FILLCELL_X32 FILLER_265_769 ();
 FILLCELL_X32 FILLER_265_801 ();
 FILLCELL_X32 FILLER_265_833 ();
 FILLCELL_X32 FILLER_265_865 ();
 FILLCELL_X32 FILLER_265_897 ();
 FILLCELL_X32 FILLER_265_929 ();
 FILLCELL_X32 FILLER_265_961 ();
 FILLCELL_X32 FILLER_265_993 ();
 FILLCELL_X32 FILLER_265_1025 ();
 FILLCELL_X32 FILLER_265_1057 ();
 FILLCELL_X32 FILLER_265_1089 ();
 FILLCELL_X32 FILLER_265_1121 ();
 FILLCELL_X32 FILLER_265_1153 ();
 FILLCELL_X32 FILLER_265_1185 ();
 FILLCELL_X32 FILLER_265_1217 ();
 FILLCELL_X8 FILLER_265_1249 ();
 FILLCELL_X4 FILLER_265_1257 ();
 FILLCELL_X2 FILLER_265_1261 ();
 FILLCELL_X32 FILLER_265_1264 ();
 FILLCELL_X32 FILLER_265_1296 ();
 FILLCELL_X32 FILLER_265_1328 ();
 FILLCELL_X32 FILLER_265_1360 ();
 FILLCELL_X32 FILLER_265_1392 ();
 FILLCELL_X32 FILLER_265_1424 ();
 FILLCELL_X32 FILLER_265_1456 ();
 FILLCELL_X32 FILLER_265_1488 ();
 FILLCELL_X32 FILLER_265_1520 ();
 FILLCELL_X32 FILLER_265_1552 ();
 FILLCELL_X32 FILLER_265_1584 ();
 FILLCELL_X32 FILLER_265_1616 ();
 FILLCELL_X32 FILLER_265_1648 ();
 FILLCELL_X32 FILLER_265_1680 ();
 FILLCELL_X32 FILLER_265_1712 ();
 FILLCELL_X32 FILLER_265_1744 ();
 FILLCELL_X32 FILLER_265_1776 ();
 FILLCELL_X32 FILLER_265_1808 ();
 FILLCELL_X32 FILLER_265_1840 ();
 FILLCELL_X32 FILLER_265_1872 ();
 FILLCELL_X32 FILLER_265_1904 ();
 FILLCELL_X32 FILLER_265_1936 ();
 FILLCELL_X32 FILLER_265_1968 ();
 FILLCELL_X32 FILLER_265_2000 ();
 FILLCELL_X32 FILLER_265_2032 ();
 FILLCELL_X32 FILLER_265_2064 ();
 FILLCELL_X32 FILLER_265_2096 ();
 FILLCELL_X32 FILLER_265_2128 ();
 FILLCELL_X32 FILLER_265_2160 ();
 FILLCELL_X32 FILLER_265_2192 ();
 FILLCELL_X32 FILLER_265_2224 ();
 FILLCELL_X32 FILLER_265_2256 ();
 FILLCELL_X32 FILLER_265_2288 ();
 FILLCELL_X32 FILLER_265_2320 ();
 FILLCELL_X32 FILLER_265_2352 ();
 FILLCELL_X32 FILLER_265_2384 ();
 FILLCELL_X32 FILLER_265_2416 ();
 FILLCELL_X32 FILLER_265_2448 ();
 FILLCELL_X32 FILLER_265_2480 ();
 FILLCELL_X8 FILLER_265_2512 ();
 FILLCELL_X4 FILLER_265_2520 ();
 FILLCELL_X2 FILLER_265_2524 ();
 FILLCELL_X32 FILLER_265_2527 ();
 FILLCELL_X32 FILLER_265_2559 ();
 FILLCELL_X8 FILLER_265_2591 ();
 FILLCELL_X2 FILLER_265_2599 ();
 FILLCELL_X1 FILLER_265_2601 ();
 FILLCELL_X32 FILLER_266_1 ();
 FILLCELL_X32 FILLER_266_33 ();
 FILLCELL_X32 FILLER_266_65 ();
 FILLCELL_X32 FILLER_266_97 ();
 FILLCELL_X32 FILLER_266_129 ();
 FILLCELL_X32 FILLER_266_161 ();
 FILLCELL_X32 FILLER_266_193 ();
 FILLCELL_X32 FILLER_266_225 ();
 FILLCELL_X32 FILLER_266_257 ();
 FILLCELL_X32 FILLER_266_289 ();
 FILLCELL_X32 FILLER_266_321 ();
 FILLCELL_X32 FILLER_266_353 ();
 FILLCELL_X32 FILLER_266_385 ();
 FILLCELL_X32 FILLER_266_417 ();
 FILLCELL_X32 FILLER_266_449 ();
 FILLCELL_X32 FILLER_266_481 ();
 FILLCELL_X32 FILLER_266_513 ();
 FILLCELL_X32 FILLER_266_545 ();
 FILLCELL_X32 FILLER_266_577 ();
 FILLCELL_X16 FILLER_266_609 ();
 FILLCELL_X4 FILLER_266_625 ();
 FILLCELL_X2 FILLER_266_629 ();
 FILLCELL_X32 FILLER_266_632 ();
 FILLCELL_X32 FILLER_266_664 ();
 FILLCELL_X32 FILLER_266_696 ();
 FILLCELL_X32 FILLER_266_728 ();
 FILLCELL_X32 FILLER_266_760 ();
 FILLCELL_X32 FILLER_266_792 ();
 FILLCELL_X32 FILLER_266_824 ();
 FILLCELL_X32 FILLER_266_856 ();
 FILLCELL_X32 FILLER_266_888 ();
 FILLCELL_X32 FILLER_266_920 ();
 FILLCELL_X32 FILLER_266_952 ();
 FILLCELL_X32 FILLER_266_984 ();
 FILLCELL_X32 FILLER_266_1016 ();
 FILLCELL_X32 FILLER_266_1048 ();
 FILLCELL_X32 FILLER_266_1080 ();
 FILLCELL_X32 FILLER_266_1112 ();
 FILLCELL_X32 FILLER_266_1144 ();
 FILLCELL_X32 FILLER_266_1176 ();
 FILLCELL_X32 FILLER_266_1208 ();
 FILLCELL_X32 FILLER_266_1240 ();
 FILLCELL_X32 FILLER_266_1272 ();
 FILLCELL_X32 FILLER_266_1304 ();
 FILLCELL_X32 FILLER_266_1336 ();
 FILLCELL_X32 FILLER_266_1368 ();
 FILLCELL_X32 FILLER_266_1400 ();
 FILLCELL_X32 FILLER_266_1432 ();
 FILLCELL_X32 FILLER_266_1464 ();
 FILLCELL_X32 FILLER_266_1496 ();
 FILLCELL_X32 FILLER_266_1528 ();
 FILLCELL_X32 FILLER_266_1560 ();
 FILLCELL_X32 FILLER_266_1592 ();
 FILLCELL_X32 FILLER_266_1624 ();
 FILLCELL_X32 FILLER_266_1656 ();
 FILLCELL_X32 FILLER_266_1688 ();
 FILLCELL_X32 FILLER_266_1720 ();
 FILLCELL_X32 FILLER_266_1752 ();
 FILLCELL_X32 FILLER_266_1784 ();
 FILLCELL_X32 FILLER_266_1816 ();
 FILLCELL_X32 FILLER_266_1848 ();
 FILLCELL_X8 FILLER_266_1880 ();
 FILLCELL_X4 FILLER_266_1888 ();
 FILLCELL_X2 FILLER_266_1892 ();
 FILLCELL_X32 FILLER_266_1895 ();
 FILLCELL_X32 FILLER_266_1927 ();
 FILLCELL_X32 FILLER_266_1959 ();
 FILLCELL_X32 FILLER_266_1991 ();
 FILLCELL_X32 FILLER_266_2023 ();
 FILLCELL_X32 FILLER_266_2055 ();
 FILLCELL_X32 FILLER_266_2087 ();
 FILLCELL_X32 FILLER_266_2119 ();
 FILLCELL_X32 FILLER_266_2151 ();
 FILLCELL_X32 FILLER_266_2183 ();
 FILLCELL_X32 FILLER_266_2215 ();
 FILLCELL_X32 FILLER_266_2247 ();
 FILLCELL_X32 FILLER_266_2279 ();
 FILLCELL_X32 FILLER_266_2311 ();
 FILLCELL_X32 FILLER_266_2343 ();
 FILLCELL_X32 FILLER_266_2375 ();
 FILLCELL_X32 FILLER_266_2407 ();
 FILLCELL_X32 FILLER_266_2439 ();
 FILLCELL_X32 FILLER_266_2471 ();
 FILLCELL_X32 FILLER_266_2503 ();
 FILLCELL_X32 FILLER_266_2535 ();
 FILLCELL_X32 FILLER_266_2567 ();
 FILLCELL_X2 FILLER_266_2599 ();
 FILLCELL_X1 FILLER_266_2601 ();
 FILLCELL_X32 FILLER_267_1 ();
 FILLCELL_X32 FILLER_267_33 ();
 FILLCELL_X32 FILLER_267_65 ();
 FILLCELL_X32 FILLER_267_97 ();
 FILLCELL_X32 FILLER_267_129 ();
 FILLCELL_X32 FILLER_267_161 ();
 FILLCELL_X32 FILLER_267_193 ();
 FILLCELL_X32 FILLER_267_225 ();
 FILLCELL_X32 FILLER_267_257 ();
 FILLCELL_X32 FILLER_267_289 ();
 FILLCELL_X32 FILLER_267_321 ();
 FILLCELL_X32 FILLER_267_353 ();
 FILLCELL_X32 FILLER_267_385 ();
 FILLCELL_X32 FILLER_267_417 ();
 FILLCELL_X32 FILLER_267_449 ();
 FILLCELL_X32 FILLER_267_481 ();
 FILLCELL_X32 FILLER_267_513 ();
 FILLCELL_X32 FILLER_267_545 ();
 FILLCELL_X32 FILLER_267_577 ();
 FILLCELL_X32 FILLER_267_609 ();
 FILLCELL_X32 FILLER_267_641 ();
 FILLCELL_X32 FILLER_267_673 ();
 FILLCELL_X32 FILLER_267_705 ();
 FILLCELL_X32 FILLER_267_737 ();
 FILLCELL_X32 FILLER_267_769 ();
 FILLCELL_X32 FILLER_267_801 ();
 FILLCELL_X32 FILLER_267_833 ();
 FILLCELL_X32 FILLER_267_865 ();
 FILLCELL_X32 FILLER_267_897 ();
 FILLCELL_X32 FILLER_267_929 ();
 FILLCELL_X32 FILLER_267_961 ();
 FILLCELL_X32 FILLER_267_993 ();
 FILLCELL_X32 FILLER_267_1025 ();
 FILLCELL_X32 FILLER_267_1057 ();
 FILLCELL_X32 FILLER_267_1089 ();
 FILLCELL_X32 FILLER_267_1121 ();
 FILLCELL_X32 FILLER_267_1153 ();
 FILLCELL_X32 FILLER_267_1185 ();
 FILLCELL_X32 FILLER_267_1217 ();
 FILLCELL_X8 FILLER_267_1249 ();
 FILLCELL_X4 FILLER_267_1257 ();
 FILLCELL_X2 FILLER_267_1261 ();
 FILLCELL_X32 FILLER_267_1264 ();
 FILLCELL_X32 FILLER_267_1296 ();
 FILLCELL_X32 FILLER_267_1328 ();
 FILLCELL_X32 FILLER_267_1360 ();
 FILLCELL_X32 FILLER_267_1392 ();
 FILLCELL_X32 FILLER_267_1424 ();
 FILLCELL_X32 FILLER_267_1456 ();
 FILLCELL_X32 FILLER_267_1488 ();
 FILLCELL_X32 FILLER_267_1520 ();
 FILLCELL_X32 FILLER_267_1552 ();
 FILLCELL_X32 FILLER_267_1584 ();
 FILLCELL_X32 FILLER_267_1616 ();
 FILLCELL_X32 FILLER_267_1648 ();
 FILLCELL_X32 FILLER_267_1680 ();
 FILLCELL_X32 FILLER_267_1712 ();
 FILLCELL_X32 FILLER_267_1744 ();
 FILLCELL_X32 FILLER_267_1776 ();
 FILLCELL_X32 FILLER_267_1808 ();
 FILLCELL_X32 FILLER_267_1840 ();
 FILLCELL_X32 FILLER_267_1872 ();
 FILLCELL_X32 FILLER_267_1904 ();
 FILLCELL_X32 FILLER_267_1936 ();
 FILLCELL_X32 FILLER_267_1968 ();
 FILLCELL_X32 FILLER_267_2000 ();
 FILLCELL_X32 FILLER_267_2032 ();
 FILLCELL_X32 FILLER_267_2064 ();
 FILLCELL_X32 FILLER_267_2096 ();
 FILLCELL_X32 FILLER_267_2128 ();
 FILLCELL_X32 FILLER_267_2160 ();
 FILLCELL_X32 FILLER_267_2192 ();
 FILLCELL_X32 FILLER_267_2224 ();
 FILLCELL_X32 FILLER_267_2256 ();
 FILLCELL_X32 FILLER_267_2288 ();
 FILLCELL_X32 FILLER_267_2320 ();
 FILLCELL_X32 FILLER_267_2352 ();
 FILLCELL_X32 FILLER_267_2384 ();
 FILLCELL_X32 FILLER_267_2416 ();
 FILLCELL_X32 FILLER_267_2448 ();
 FILLCELL_X32 FILLER_267_2480 ();
 FILLCELL_X8 FILLER_267_2512 ();
 FILLCELL_X4 FILLER_267_2520 ();
 FILLCELL_X2 FILLER_267_2524 ();
 FILLCELL_X32 FILLER_267_2527 ();
 FILLCELL_X32 FILLER_267_2559 ();
 FILLCELL_X8 FILLER_267_2591 ();
 FILLCELL_X2 FILLER_267_2599 ();
 FILLCELL_X1 FILLER_267_2601 ();
 FILLCELL_X32 FILLER_268_1 ();
 FILLCELL_X32 FILLER_268_33 ();
 FILLCELL_X32 FILLER_268_65 ();
 FILLCELL_X32 FILLER_268_97 ();
 FILLCELL_X32 FILLER_268_129 ();
 FILLCELL_X32 FILLER_268_161 ();
 FILLCELL_X32 FILLER_268_193 ();
 FILLCELL_X32 FILLER_268_225 ();
 FILLCELL_X32 FILLER_268_257 ();
 FILLCELL_X32 FILLER_268_289 ();
 FILLCELL_X32 FILLER_268_321 ();
 FILLCELL_X32 FILLER_268_353 ();
 FILLCELL_X32 FILLER_268_385 ();
 FILLCELL_X32 FILLER_268_417 ();
 FILLCELL_X32 FILLER_268_449 ();
 FILLCELL_X32 FILLER_268_481 ();
 FILLCELL_X32 FILLER_268_513 ();
 FILLCELL_X32 FILLER_268_545 ();
 FILLCELL_X32 FILLER_268_577 ();
 FILLCELL_X16 FILLER_268_609 ();
 FILLCELL_X4 FILLER_268_625 ();
 FILLCELL_X2 FILLER_268_629 ();
 FILLCELL_X32 FILLER_268_632 ();
 FILLCELL_X32 FILLER_268_664 ();
 FILLCELL_X32 FILLER_268_696 ();
 FILLCELL_X32 FILLER_268_728 ();
 FILLCELL_X32 FILLER_268_760 ();
 FILLCELL_X32 FILLER_268_792 ();
 FILLCELL_X32 FILLER_268_824 ();
 FILLCELL_X32 FILLER_268_856 ();
 FILLCELL_X32 FILLER_268_888 ();
 FILLCELL_X32 FILLER_268_920 ();
 FILLCELL_X32 FILLER_268_952 ();
 FILLCELL_X32 FILLER_268_984 ();
 FILLCELL_X32 FILLER_268_1016 ();
 FILLCELL_X32 FILLER_268_1048 ();
 FILLCELL_X32 FILLER_268_1080 ();
 FILLCELL_X32 FILLER_268_1112 ();
 FILLCELL_X32 FILLER_268_1144 ();
 FILLCELL_X32 FILLER_268_1176 ();
 FILLCELL_X32 FILLER_268_1208 ();
 FILLCELL_X32 FILLER_268_1240 ();
 FILLCELL_X32 FILLER_268_1272 ();
 FILLCELL_X32 FILLER_268_1304 ();
 FILLCELL_X32 FILLER_268_1336 ();
 FILLCELL_X32 FILLER_268_1368 ();
 FILLCELL_X32 FILLER_268_1400 ();
 FILLCELL_X32 FILLER_268_1432 ();
 FILLCELL_X32 FILLER_268_1464 ();
 FILLCELL_X32 FILLER_268_1496 ();
 FILLCELL_X32 FILLER_268_1528 ();
 FILLCELL_X32 FILLER_268_1560 ();
 FILLCELL_X32 FILLER_268_1592 ();
 FILLCELL_X32 FILLER_268_1624 ();
 FILLCELL_X32 FILLER_268_1656 ();
 FILLCELL_X32 FILLER_268_1688 ();
 FILLCELL_X32 FILLER_268_1720 ();
 FILLCELL_X32 FILLER_268_1752 ();
 FILLCELL_X32 FILLER_268_1784 ();
 FILLCELL_X32 FILLER_268_1816 ();
 FILLCELL_X32 FILLER_268_1848 ();
 FILLCELL_X8 FILLER_268_1880 ();
 FILLCELL_X4 FILLER_268_1888 ();
 FILLCELL_X2 FILLER_268_1892 ();
 FILLCELL_X32 FILLER_268_1895 ();
 FILLCELL_X32 FILLER_268_1927 ();
 FILLCELL_X32 FILLER_268_1959 ();
 FILLCELL_X32 FILLER_268_1991 ();
 FILLCELL_X32 FILLER_268_2023 ();
 FILLCELL_X32 FILLER_268_2055 ();
 FILLCELL_X32 FILLER_268_2087 ();
 FILLCELL_X32 FILLER_268_2119 ();
 FILLCELL_X32 FILLER_268_2151 ();
 FILLCELL_X32 FILLER_268_2183 ();
 FILLCELL_X32 FILLER_268_2215 ();
 FILLCELL_X32 FILLER_268_2247 ();
 FILLCELL_X32 FILLER_268_2279 ();
 FILLCELL_X32 FILLER_268_2311 ();
 FILLCELL_X32 FILLER_268_2343 ();
 FILLCELL_X32 FILLER_268_2375 ();
 FILLCELL_X32 FILLER_268_2407 ();
 FILLCELL_X32 FILLER_268_2439 ();
 FILLCELL_X32 FILLER_268_2471 ();
 FILLCELL_X32 FILLER_268_2503 ();
 FILLCELL_X32 FILLER_268_2535 ();
 FILLCELL_X32 FILLER_268_2567 ();
 FILLCELL_X2 FILLER_268_2599 ();
 FILLCELL_X1 FILLER_268_2601 ();
 FILLCELL_X32 FILLER_269_1 ();
 FILLCELL_X32 FILLER_269_33 ();
 FILLCELL_X32 FILLER_269_65 ();
 FILLCELL_X32 FILLER_269_97 ();
 FILLCELL_X32 FILLER_269_129 ();
 FILLCELL_X32 FILLER_269_161 ();
 FILLCELL_X32 FILLER_269_193 ();
 FILLCELL_X32 FILLER_269_225 ();
 FILLCELL_X32 FILLER_269_257 ();
 FILLCELL_X32 FILLER_269_289 ();
 FILLCELL_X32 FILLER_269_321 ();
 FILLCELL_X32 FILLER_269_353 ();
 FILLCELL_X32 FILLER_269_385 ();
 FILLCELL_X32 FILLER_269_417 ();
 FILLCELL_X32 FILLER_269_449 ();
 FILLCELL_X32 FILLER_269_481 ();
 FILLCELL_X32 FILLER_269_513 ();
 FILLCELL_X32 FILLER_269_545 ();
 FILLCELL_X32 FILLER_269_577 ();
 FILLCELL_X32 FILLER_269_609 ();
 FILLCELL_X32 FILLER_269_641 ();
 FILLCELL_X32 FILLER_269_673 ();
 FILLCELL_X32 FILLER_269_705 ();
 FILLCELL_X32 FILLER_269_737 ();
 FILLCELL_X32 FILLER_269_769 ();
 FILLCELL_X32 FILLER_269_801 ();
 FILLCELL_X32 FILLER_269_833 ();
 FILLCELL_X32 FILLER_269_865 ();
 FILLCELL_X32 FILLER_269_897 ();
 FILLCELL_X32 FILLER_269_929 ();
 FILLCELL_X32 FILLER_269_961 ();
 FILLCELL_X32 FILLER_269_993 ();
 FILLCELL_X32 FILLER_269_1025 ();
 FILLCELL_X32 FILLER_269_1057 ();
 FILLCELL_X32 FILLER_269_1089 ();
 FILLCELL_X32 FILLER_269_1121 ();
 FILLCELL_X32 FILLER_269_1153 ();
 FILLCELL_X32 FILLER_269_1185 ();
 FILLCELL_X32 FILLER_269_1217 ();
 FILLCELL_X8 FILLER_269_1249 ();
 FILLCELL_X4 FILLER_269_1257 ();
 FILLCELL_X2 FILLER_269_1261 ();
 FILLCELL_X32 FILLER_269_1264 ();
 FILLCELL_X32 FILLER_269_1296 ();
 FILLCELL_X32 FILLER_269_1328 ();
 FILLCELL_X32 FILLER_269_1360 ();
 FILLCELL_X32 FILLER_269_1392 ();
 FILLCELL_X32 FILLER_269_1424 ();
 FILLCELL_X32 FILLER_269_1456 ();
 FILLCELL_X32 FILLER_269_1488 ();
 FILLCELL_X32 FILLER_269_1520 ();
 FILLCELL_X32 FILLER_269_1552 ();
 FILLCELL_X32 FILLER_269_1584 ();
 FILLCELL_X32 FILLER_269_1616 ();
 FILLCELL_X32 FILLER_269_1648 ();
 FILLCELL_X32 FILLER_269_1680 ();
 FILLCELL_X32 FILLER_269_1712 ();
 FILLCELL_X32 FILLER_269_1744 ();
 FILLCELL_X32 FILLER_269_1776 ();
 FILLCELL_X32 FILLER_269_1808 ();
 FILLCELL_X32 FILLER_269_1840 ();
 FILLCELL_X32 FILLER_269_1872 ();
 FILLCELL_X32 FILLER_269_1904 ();
 FILLCELL_X32 FILLER_269_1936 ();
 FILLCELL_X32 FILLER_269_1968 ();
 FILLCELL_X32 FILLER_269_2000 ();
 FILLCELL_X32 FILLER_269_2032 ();
 FILLCELL_X32 FILLER_269_2064 ();
 FILLCELL_X32 FILLER_269_2096 ();
 FILLCELL_X32 FILLER_269_2128 ();
 FILLCELL_X32 FILLER_269_2160 ();
 FILLCELL_X32 FILLER_269_2192 ();
 FILLCELL_X32 FILLER_269_2224 ();
 FILLCELL_X32 FILLER_269_2256 ();
 FILLCELL_X32 FILLER_269_2288 ();
 FILLCELL_X32 FILLER_269_2320 ();
 FILLCELL_X32 FILLER_269_2352 ();
 FILLCELL_X32 FILLER_269_2384 ();
 FILLCELL_X32 FILLER_269_2416 ();
 FILLCELL_X32 FILLER_269_2448 ();
 FILLCELL_X32 FILLER_269_2480 ();
 FILLCELL_X8 FILLER_269_2512 ();
 FILLCELL_X4 FILLER_269_2520 ();
 FILLCELL_X2 FILLER_269_2524 ();
 FILLCELL_X32 FILLER_269_2527 ();
 FILLCELL_X32 FILLER_269_2559 ();
 FILLCELL_X8 FILLER_269_2591 ();
 FILLCELL_X2 FILLER_269_2599 ();
 FILLCELL_X1 FILLER_269_2601 ();
 FILLCELL_X32 FILLER_270_1 ();
 FILLCELL_X32 FILLER_270_33 ();
 FILLCELL_X32 FILLER_270_65 ();
 FILLCELL_X32 FILLER_270_97 ();
 FILLCELL_X32 FILLER_270_129 ();
 FILLCELL_X32 FILLER_270_161 ();
 FILLCELL_X32 FILLER_270_193 ();
 FILLCELL_X32 FILLER_270_225 ();
 FILLCELL_X32 FILLER_270_257 ();
 FILLCELL_X32 FILLER_270_289 ();
 FILLCELL_X32 FILLER_270_321 ();
 FILLCELL_X32 FILLER_270_353 ();
 FILLCELL_X32 FILLER_270_385 ();
 FILLCELL_X32 FILLER_270_417 ();
 FILLCELL_X32 FILLER_270_449 ();
 FILLCELL_X32 FILLER_270_481 ();
 FILLCELL_X32 FILLER_270_513 ();
 FILLCELL_X32 FILLER_270_545 ();
 FILLCELL_X32 FILLER_270_577 ();
 FILLCELL_X16 FILLER_270_609 ();
 FILLCELL_X4 FILLER_270_625 ();
 FILLCELL_X2 FILLER_270_629 ();
 FILLCELL_X32 FILLER_270_632 ();
 FILLCELL_X32 FILLER_270_664 ();
 FILLCELL_X32 FILLER_270_696 ();
 FILLCELL_X32 FILLER_270_728 ();
 FILLCELL_X32 FILLER_270_760 ();
 FILLCELL_X32 FILLER_270_792 ();
 FILLCELL_X32 FILLER_270_824 ();
 FILLCELL_X32 FILLER_270_856 ();
 FILLCELL_X32 FILLER_270_888 ();
 FILLCELL_X32 FILLER_270_920 ();
 FILLCELL_X32 FILLER_270_952 ();
 FILLCELL_X32 FILLER_270_984 ();
 FILLCELL_X32 FILLER_270_1016 ();
 FILLCELL_X32 FILLER_270_1048 ();
 FILLCELL_X32 FILLER_270_1080 ();
 FILLCELL_X32 FILLER_270_1112 ();
 FILLCELL_X32 FILLER_270_1144 ();
 FILLCELL_X32 FILLER_270_1176 ();
 FILLCELL_X32 FILLER_270_1208 ();
 FILLCELL_X32 FILLER_270_1240 ();
 FILLCELL_X32 FILLER_270_1272 ();
 FILLCELL_X32 FILLER_270_1304 ();
 FILLCELL_X32 FILLER_270_1336 ();
 FILLCELL_X32 FILLER_270_1368 ();
 FILLCELL_X32 FILLER_270_1400 ();
 FILLCELL_X32 FILLER_270_1432 ();
 FILLCELL_X32 FILLER_270_1464 ();
 FILLCELL_X32 FILLER_270_1496 ();
 FILLCELL_X32 FILLER_270_1528 ();
 FILLCELL_X32 FILLER_270_1560 ();
 FILLCELL_X32 FILLER_270_1592 ();
 FILLCELL_X32 FILLER_270_1624 ();
 FILLCELL_X32 FILLER_270_1656 ();
 FILLCELL_X32 FILLER_270_1688 ();
 FILLCELL_X32 FILLER_270_1720 ();
 FILLCELL_X32 FILLER_270_1752 ();
 FILLCELL_X32 FILLER_270_1784 ();
 FILLCELL_X32 FILLER_270_1816 ();
 FILLCELL_X32 FILLER_270_1848 ();
 FILLCELL_X8 FILLER_270_1880 ();
 FILLCELL_X4 FILLER_270_1888 ();
 FILLCELL_X2 FILLER_270_1892 ();
 FILLCELL_X32 FILLER_270_1895 ();
 FILLCELL_X32 FILLER_270_1927 ();
 FILLCELL_X32 FILLER_270_1959 ();
 FILLCELL_X32 FILLER_270_1991 ();
 FILLCELL_X32 FILLER_270_2023 ();
 FILLCELL_X32 FILLER_270_2055 ();
 FILLCELL_X32 FILLER_270_2087 ();
 FILLCELL_X32 FILLER_270_2119 ();
 FILLCELL_X32 FILLER_270_2151 ();
 FILLCELL_X32 FILLER_270_2183 ();
 FILLCELL_X32 FILLER_270_2215 ();
 FILLCELL_X32 FILLER_270_2247 ();
 FILLCELL_X32 FILLER_270_2279 ();
 FILLCELL_X32 FILLER_270_2311 ();
 FILLCELL_X32 FILLER_270_2343 ();
 FILLCELL_X32 FILLER_270_2375 ();
 FILLCELL_X32 FILLER_270_2407 ();
 FILLCELL_X32 FILLER_270_2439 ();
 FILLCELL_X32 FILLER_270_2471 ();
 FILLCELL_X32 FILLER_270_2503 ();
 FILLCELL_X32 FILLER_270_2535 ();
 FILLCELL_X32 FILLER_270_2567 ();
 FILLCELL_X2 FILLER_270_2599 ();
 FILLCELL_X1 FILLER_270_2601 ();
 FILLCELL_X32 FILLER_271_1 ();
 FILLCELL_X32 FILLER_271_33 ();
 FILLCELL_X32 FILLER_271_65 ();
 FILLCELL_X32 FILLER_271_97 ();
 FILLCELL_X32 FILLER_271_129 ();
 FILLCELL_X32 FILLER_271_161 ();
 FILLCELL_X32 FILLER_271_193 ();
 FILLCELL_X32 FILLER_271_225 ();
 FILLCELL_X32 FILLER_271_257 ();
 FILLCELL_X32 FILLER_271_289 ();
 FILLCELL_X32 FILLER_271_321 ();
 FILLCELL_X32 FILLER_271_353 ();
 FILLCELL_X32 FILLER_271_385 ();
 FILLCELL_X32 FILLER_271_417 ();
 FILLCELL_X32 FILLER_271_449 ();
 FILLCELL_X32 FILLER_271_481 ();
 FILLCELL_X32 FILLER_271_513 ();
 FILLCELL_X32 FILLER_271_545 ();
 FILLCELL_X32 FILLER_271_577 ();
 FILLCELL_X32 FILLER_271_609 ();
 FILLCELL_X32 FILLER_271_641 ();
 FILLCELL_X32 FILLER_271_673 ();
 FILLCELL_X32 FILLER_271_705 ();
 FILLCELL_X32 FILLER_271_737 ();
 FILLCELL_X32 FILLER_271_769 ();
 FILLCELL_X32 FILLER_271_801 ();
 FILLCELL_X32 FILLER_271_833 ();
 FILLCELL_X32 FILLER_271_865 ();
 FILLCELL_X32 FILLER_271_897 ();
 FILLCELL_X32 FILLER_271_929 ();
 FILLCELL_X32 FILLER_271_961 ();
 FILLCELL_X32 FILLER_271_993 ();
 FILLCELL_X32 FILLER_271_1025 ();
 FILLCELL_X32 FILLER_271_1057 ();
 FILLCELL_X32 FILLER_271_1089 ();
 FILLCELL_X32 FILLER_271_1121 ();
 FILLCELL_X32 FILLER_271_1153 ();
 FILLCELL_X32 FILLER_271_1185 ();
 FILLCELL_X32 FILLER_271_1217 ();
 FILLCELL_X8 FILLER_271_1249 ();
 FILLCELL_X4 FILLER_271_1257 ();
 FILLCELL_X2 FILLER_271_1261 ();
 FILLCELL_X32 FILLER_271_1264 ();
 FILLCELL_X32 FILLER_271_1296 ();
 FILLCELL_X32 FILLER_271_1328 ();
 FILLCELL_X32 FILLER_271_1360 ();
 FILLCELL_X32 FILLER_271_1392 ();
 FILLCELL_X32 FILLER_271_1424 ();
 FILLCELL_X32 FILLER_271_1456 ();
 FILLCELL_X32 FILLER_271_1488 ();
 FILLCELL_X32 FILLER_271_1520 ();
 FILLCELL_X32 FILLER_271_1552 ();
 FILLCELL_X32 FILLER_271_1584 ();
 FILLCELL_X32 FILLER_271_1616 ();
 FILLCELL_X32 FILLER_271_1648 ();
 FILLCELL_X32 FILLER_271_1680 ();
 FILLCELL_X32 FILLER_271_1712 ();
 FILLCELL_X32 FILLER_271_1744 ();
 FILLCELL_X32 FILLER_271_1776 ();
 FILLCELL_X32 FILLER_271_1808 ();
 FILLCELL_X32 FILLER_271_1840 ();
 FILLCELL_X32 FILLER_271_1872 ();
 FILLCELL_X32 FILLER_271_1904 ();
 FILLCELL_X32 FILLER_271_1936 ();
 FILLCELL_X32 FILLER_271_1968 ();
 FILLCELL_X32 FILLER_271_2000 ();
 FILLCELL_X32 FILLER_271_2032 ();
 FILLCELL_X32 FILLER_271_2064 ();
 FILLCELL_X32 FILLER_271_2096 ();
 FILLCELL_X32 FILLER_271_2128 ();
 FILLCELL_X32 FILLER_271_2160 ();
 FILLCELL_X32 FILLER_271_2192 ();
 FILLCELL_X32 FILLER_271_2224 ();
 FILLCELL_X32 FILLER_271_2256 ();
 FILLCELL_X32 FILLER_271_2288 ();
 FILLCELL_X32 FILLER_271_2320 ();
 FILLCELL_X32 FILLER_271_2352 ();
 FILLCELL_X32 FILLER_271_2384 ();
 FILLCELL_X32 FILLER_271_2416 ();
 FILLCELL_X32 FILLER_271_2448 ();
 FILLCELL_X32 FILLER_271_2480 ();
 FILLCELL_X8 FILLER_271_2512 ();
 FILLCELL_X4 FILLER_271_2520 ();
 FILLCELL_X2 FILLER_271_2524 ();
 FILLCELL_X32 FILLER_271_2527 ();
 FILLCELL_X32 FILLER_271_2559 ();
 FILLCELL_X8 FILLER_271_2591 ();
 FILLCELL_X2 FILLER_271_2599 ();
 FILLCELL_X1 FILLER_271_2601 ();
 FILLCELL_X32 FILLER_272_1 ();
 FILLCELL_X32 FILLER_272_33 ();
 FILLCELL_X32 FILLER_272_65 ();
 FILLCELL_X32 FILLER_272_97 ();
 FILLCELL_X32 FILLER_272_129 ();
 FILLCELL_X32 FILLER_272_161 ();
 FILLCELL_X32 FILLER_272_193 ();
 FILLCELL_X32 FILLER_272_225 ();
 FILLCELL_X32 FILLER_272_257 ();
 FILLCELL_X32 FILLER_272_289 ();
 FILLCELL_X32 FILLER_272_321 ();
 FILLCELL_X32 FILLER_272_353 ();
 FILLCELL_X32 FILLER_272_385 ();
 FILLCELL_X32 FILLER_272_417 ();
 FILLCELL_X32 FILLER_272_449 ();
 FILLCELL_X32 FILLER_272_481 ();
 FILLCELL_X32 FILLER_272_513 ();
 FILLCELL_X32 FILLER_272_545 ();
 FILLCELL_X32 FILLER_272_577 ();
 FILLCELL_X16 FILLER_272_609 ();
 FILLCELL_X4 FILLER_272_625 ();
 FILLCELL_X2 FILLER_272_629 ();
 FILLCELL_X32 FILLER_272_632 ();
 FILLCELL_X32 FILLER_272_664 ();
 FILLCELL_X32 FILLER_272_696 ();
 FILLCELL_X32 FILLER_272_728 ();
 FILLCELL_X32 FILLER_272_760 ();
 FILLCELL_X32 FILLER_272_792 ();
 FILLCELL_X32 FILLER_272_824 ();
 FILLCELL_X32 FILLER_272_856 ();
 FILLCELL_X32 FILLER_272_888 ();
 FILLCELL_X32 FILLER_272_920 ();
 FILLCELL_X32 FILLER_272_952 ();
 FILLCELL_X32 FILLER_272_984 ();
 FILLCELL_X32 FILLER_272_1016 ();
 FILLCELL_X32 FILLER_272_1048 ();
 FILLCELL_X32 FILLER_272_1080 ();
 FILLCELL_X32 FILLER_272_1112 ();
 FILLCELL_X32 FILLER_272_1144 ();
 FILLCELL_X32 FILLER_272_1176 ();
 FILLCELL_X32 FILLER_272_1208 ();
 FILLCELL_X32 FILLER_272_1240 ();
 FILLCELL_X32 FILLER_272_1272 ();
 FILLCELL_X32 FILLER_272_1304 ();
 FILLCELL_X32 FILLER_272_1336 ();
 FILLCELL_X32 FILLER_272_1368 ();
 FILLCELL_X32 FILLER_272_1400 ();
 FILLCELL_X32 FILLER_272_1432 ();
 FILLCELL_X32 FILLER_272_1464 ();
 FILLCELL_X32 FILLER_272_1496 ();
 FILLCELL_X32 FILLER_272_1528 ();
 FILLCELL_X32 FILLER_272_1560 ();
 FILLCELL_X32 FILLER_272_1592 ();
 FILLCELL_X32 FILLER_272_1624 ();
 FILLCELL_X32 FILLER_272_1656 ();
 FILLCELL_X32 FILLER_272_1688 ();
 FILLCELL_X32 FILLER_272_1720 ();
 FILLCELL_X32 FILLER_272_1752 ();
 FILLCELL_X32 FILLER_272_1784 ();
 FILLCELL_X32 FILLER_272_1816 ();
 FILLCELL_X32 FILLER_272_1848 ();
 FILLCELL_X8 FILLER_272_1880 ();
 FILLCELL_X4 FILLER_272_1888 ();
 FILLCELL_X2 FILLER_272_1892 ();
 FILLCELL_X32 FILLER_272_1895 ();
 FILLCELL_X32 FILLER_272_1927 ();
 FILLCELL_X32 FILLER_272_1959 ();
 FILLCELL_X32 FILLER_272_1991 ();
 FILLCELL_X32 FILLER_272_2023 ();
 FILLCELL_X32 FILLER_272_2055 ();
 FILLCELL_X32 FILLER_272_2087 ();
 FILLCELL_X32 FILLER_272_2119 ();
 FILLCELL_X32 FILLER_272_2151 ();
 FILLCELL_X32 FILLER_272_2183 ();
 FILLCELL_X32 FILLER_272_2215 ();
 FILLCELL_X32 FILLER_272_2247 ();
 FILLCELL_X32 FILLER_272_2279 ();
 FILLCELL_X32 FILLER_272_2311 ();
 FILLCELL_X32 FILLER_272_2343 ();
 FILLCELL_X32 FILLER_272_2375 ();
 FILLCELL_X32 FILLER_272_2407 ();
 FILLCELL_X32 FILLER_272_2439 ();
 FILLCELL_X32 FILLER_272_2471 ();
 FILLCELL_X32 FILLER_272_2503 ();
 FILLCELL_X32 FILLER_272_2535 ();
 FILLCELL_X32 FILLER_272_2567 ();
 FILLCELL_X2 FILLER_272_2599 ();
 FILLCELL_X1 FILLER_272_2601 ();
 FILLCELL_X32 FILLER_273_1 ();
 FILLCELL_X32 FILLER_273_33 ();
 FILLCELL_X32 FILLER_273_65 ();
 FILLCELL_X32 FILLER_273_97 ();
 FILLCELL_X32 FILLER_273_129 ();
 FILLCELL_X32 FILLER_273_161 ();
 FILLCELL_X32 FILLER_273_193 ();
 FILLCELL_X32 FILLER_273_225 ();
 FILLCELL_X32 FILLER_273_257 ();
 FILLCELL_X32 FILLER_273_289 ();
 FILLCELL_X32 FILLER_273_321 ();
 FILLCELL_X32 FILLER_273_353 ();
 FILLCELL_X32 FILLER_273_385 ();
 FILLCELL_X32 FILLER_273_417 ();
 FILLCELL_X32 FILLER_273_449 ();
 FILLCELL_X32 FILLER_273_481 ();
 FILLCELL_X32 FILLER_273_513 ();
 FILLCELL_X32 FILLER_273_545 ();
 FILLCELL_X32 FILLER_273_577 ();
 FILLCELL_X32 FILLER_273_609 ();
 FILLCELL_X32 FILLER_273_641 ();
 FILLCELL_X32 FILLER_273_673 ();
 FILLCELL_X32 FILLER_273_705 ();
 FILLCELL_X32 FILLER_273_737 ();
 FILLCELL_X32 FILLER_273_769 ();
 FILLCELL_X32 FILLER_273_801 ();
 FILLCELL_X32 FILLER_273_833 ();
 FILLCELL_X32 FILLER_273_865 ();
 FILLCELL_X32 FILLER_273_897 ();
 FILLCELL_X32 FILLER_273_929 ();
 FILLCELL_X32 FILLER_273_961 ();
 FILLCELL_X32 FILLER_273_993 ();
 FILLCELL_X32 FILLER_273_1025 ();
 FILLCELL_X32 FILLER_273_1057 ();
 FILLCELL_X32 FILLER_273_1089 ();
 FILLCELL_X32 FILLER_273_1121 ();
 FILLCELL_X32 FILLER_273_1153 ();
 FILLCELL_X32 FILLER_273_1185 ();
 FILLCELL_X32 FILLER_273_1217 ();
 FILLCELL_X8 FILLER_273_1249 ();
 FILLCELL_X4 FILLER_273_1257 ();
 FILLCELL_X2 FILLER_273_1261 ();
 FILLCELL_X32 FILLER_273_1264 ();
 FILLCELL_X32 FILLER_273_1296 ();
 FILLCELL_X32 FILLER_273_1328 ();
 FILLCELL_X32 FILLER_273_1360 ();
 FILLCELL_X32 FILLER_273_1392 ();
 FILLCELL_X32 FILLER_273_1424 ();
 FILLCELL_X32 FILLER_273_1456 ();
 FILLCELL_X32 FILLER_273_1488 ();
 FILLCELL_X32 FILLER_273_1520 ();
 FILLCELL_X32 FILLER_273_1552 ();
 FILLCELL_X32 FILLER_273_1584 ();
 FILLCELL_X32 FILLER_273_1616 ();
 FILLCELL_X32 FILLER_273_1648 ();
 FILLCELL_X32 FILLER_273_1680 ();
 FILLCELL_X32 FILLER_273_1712 ();
 FILLCELL_X32 FILLER_273_1744 ();
 FILLCELL_X32 FILLER_273_1776 ();
 FILLCELL_X32 FILLER_273_1808 ();
 FILLCELL_X32 FILLER_273_1840 ();
 FILLCELL_X32 FILLER_273_1872 ();
 FILLCELL_X32 FILLER_273_1904 ();
 FILLCELL_X32 FILLER_273_1936 ();
 FILLCELL_X32 FILLER_273_1968 ();
 FILLCELL_X32 FILLER_273_2000 ();
 FILLCELL_X32 FILLER_273_2032 ();
 FILLCELL_X32 FILLER_273_2064 ();
 FILLCELL_X32 FILLER_273_2096 ();
 FILLCELL_X32 FILLER_273_2128 ();
 FILLCELL_X32 FILLER_273_2160 ();
 FILLCELL_X32 FILLER_273_2192 ();
 FILLCELL_X32 FILLER_273_2224 ();
 FILLCELL_X32 FILLER_273_2256 ();
 FILLCELL_X32 FILLER_273_2288 ();
 FILLCELL_X32 FILLER_273_2320 ();
 FILLCELL_X32 FILLER_273_2352 ();
 FILLCELL_X32 FILLER_273_2384 ();
 FILLCELL_X32 FILLER_273_2416 ();
 FILLCELL_X32 FILLER_273_2448 ();
 FILLCELL_X32 FILLER_273_2480 ();
 FILLCELL_X8 FILLER_273_2512 ();
 FILLCELL_X4 FILLER_273_2520 ();
 FILLCELL_X2 FILLER_273_2524 ();
 FILLCELL_X32 FILLER_273_2527 ();
 FILLCELL_X32 FILLER_273_2559 ();
 FILLCELL_X8 FILLER_273_2591 ();
 FILLCELL_X2 FILLER_273_2599 ();
 FILLCELL_X1 FILLER_273_2601 ();
 FILLCELL_X32 FILLER_274_1 ();
 FILLCELL_X32 FILLER_274_33 ();
 FILLCELL_X32 FILLER_274_65 ();
 FILLCELL_X32 FILLER_274_97 ();
 FILLCELL_X32 FILLER_274_129 ();
 FILLCELL_X32 FILLER_274_161 ();
 FILLCELL_X32 FILLER_274_193 ();
 FILLCELL_X32 FILLER_274_225 ();
 FILLCELL_X32 FILLER_274_257 ();
 FILLCELL_X32 FILLER_274_289 ();
 FILLCELL_X32 FILLER_274_321 ();
 FILLCELL_X32 FILLER_274_353 ();
 FILLCELL_X32 FILLER_274_385 ();
 FILLCELL_X32 FILLER_274_417 ();
 FILLCELL_X32 FILLER_274_449 ();
 FILLCELL_X32 FILLER_274_481 ();
 FILLCELL_X32 FILLER_274_513 ();
 FILLCELL_X32 FILLER_274_545 ();
 FILLCELL_X32 FILLER_274_577 ();
 FILLCELL_X16 FILLER_274_609 ();
 FILLCELL_X4 FILLER_274_625 ();
 FILLCELL_X2 FILLER_274_629 ();
 FILLCELL_X32 FILLER_274_632 ();
 FILLCELL_X32 FILLER_274_664 ();
 FILLCELL_X32 FILLER_274_696 ();
 FILLCELL_X32 FILLER_274_728 ();
 FILLCELL_X32 FILLER_274_760 ();
 FILLCELL_X32 FILLER_274_792 ();
 FILLCELL_X32 FILLER_274_824 ();
 FILLCELL_X32 FILLER_274_856 ();
 FILLCELL_X32 FILLER_274_888 ();
 FILLCELL_X32 FILLER_274_920 ();
 FILLCELL_X32 FILLER_274_952 ();
 FILLCELL_X32 FILLER_274_984 ();
 FILLCELL_X32 FILLER_274_1016 ();
 FILLCELL_X32 FILLER_274_1048 ();
 FILLCELL_X32 FILLER_274_1080 ();
 FILLCELL_X32 FILLER_274_1112 ();
 FILLCELL_X32 FILLER_274_1144 ();
 FILLCELL_X32 FILLER_274_1176 ();
 FILLCELL_X32 FILLER_274_1208 ();
 FILLCELL_X32 FILLER_274_1240 ();
 FILLCELL_X32 FILLER_274_1272 ();
 FILLCELL_X32 FILLER_274_1304 ();
 FILLCELL_X32 FILLER_274_1336 ();
 FILLCELL_X32 FILLER_274_1368 ();
 FILLCELL_X32 FILLER_274_1400 ();
 FILLCELL_X32 FILLER_274_1432 ();
 FILLCELL_X32 FILLER_274_1464 ();
 FILLCELL_X32 FILLER_274_1496 ();
 FILLCELL_X32 FILLER_274_1528 ();
 FILLCELL_X32 FILLER_274_1560 ();
 FILLCELL_X32 FILLER_274_1592 ();
 FILLCELL_X32 FILLER_274_1624 ();
 FILLCELL_X32 FILLER_274_1656 ();
 FILLCELL_X32 FILLER_274_1688 ();
 FILLCELL_X32 FILLER_274_1720 ();
 FILLCELL_X32 FILLER_274_1752 ();
 FILLCELL_X32 FILLER_274_1784 ();
 FILLCELL_X32 FILLER_274_1816 ();
 FILLCELL_X32 FILLER_274_1848 ();
 FILLCELL_X8 FILLER_274_1880 ();
 FILLCELL_X4 FILLER_274_1888 ();
 FILLCELL_X2 FILLER_274_1892 ();
 FILLCELL_X32 FILLER_274_1895 ();
 FILLCELL_X32 FILLER_274_1927 ();
 FILLCELL_X32 FILLER_274_1959 ();
 FILLCELL_X32 FILLER_274_1991 ();
 FILLCELL_X32 FILLER_274_2023 ();
 FILLCELL_X32 FILLER_274_2055 ();
 FILLCELL_X32 FILLER_274_2087 ();
 FILLCELL_X32 FILLER_274_2119 ();
 FILLCELL_X32 FILLER_274_2151 ();
 FILLCELL_X32 FILLER_274_2183 ();
 FILLCELL_X32 FILLER_274_2215 ();
 FILLCELL_X32 FILLER_274_2247 ();
 FILLCELL_X32 FILLER_274_2279 ();
 FILLCELL_X32 FILLER_274_2311 ();
 FILLCELL_X32 FILLER_274_2343 ();
 FILLCELL_X32 FILLER_274_2375 ();
 FILLCELL_X32 FILLER_274_2407 ();
 FILLCELL_X32 FILLER_274_2439 ();
 FILLCELL_X32 FILLER_274_2471 ();
 FILLCELL_X32 FILLER_274_2503 ();
 FILLCELL_X32 FILLER_274_2535 ();
 FILLCELL_X32 FILLER_274_2567 ();
 FILLCELL_X2 FILLER_274_2599 ();
 FILLCELL_X1 FILLER_274_2601 ();
 FILLCELL_X32 FILLER_275_1 ();
 FILLCELL_X32 FILLER_275_33 ();
 FILLCELL_X32 FILLER_275_65 ();
 FILLCELL_X32 FILLER_275_97 ();
 FILLCELL_X32 FILLER_275_129 ();
 FILLCELL_X32 FILLER_275_161 ();
 FILLCELL_X32 FILLER_275_193 ();
 FILLCELL_X32 FILLER_275_225 ();
 FILLCELL_X32 FILLER_275_257 ();
 FILLCELL_X32 FILLER_275_289 ();
 FILLCELL_X32 FILLER_275_321 ();
 FILLCELL_X32 FILLER_275_353 ();
 FILLCELL_X32 FILLER_275_385 ();
 FILLCELL_X32 FILLER_275_417 ();
 FILLCELL_X32 FILLER_275_449 ();
 FILLCELL_X32 FILLER_275_481 ();
 FILLCELL_X32 FILLER_275_513 ();
 FILLCELL_X32 FILLER_275_545 ();
 FILLCELL_X32 FILLER_275_577 ();
 FILLCELL_X32 FILLER_275_609 ();
 FILLCELL_X32 FILLER_275_641 ();
 FILLCELL_X32 FILLER_275_673 ();
 FILLCELL_X32 FILLER_275_705 ();
 FILLCELL_X32 FILLER_275_737 ();
 FILLCELL_X32 FILLER_275_769 ();
 FILLCELL_X32 FILLER_275_801 ();
 FILLCELL_X32 FILLER_275_833 ();
 FILLCELL_X32 FILLER_275_865 ();
 FILLCELL_X32 FILLER_275_897 ();
 FILLCELL_X32 FILLER_275_929 ();
 FILLCELL_X32 FILLER_275_961 ();
 FILLCELL_X32 FILLER_275_993 ();
 FILLCELL_X32 FILLER_275_1025 ();
 FILLCELL_X32 FILLER_275_1057 ();
 FILLCELL_X32 FILLER_275_1089 ();
 FILLCELL_X32 FILLER_275_1121 ();
 FILLCELL_X32 FILLER_275_1153 ();
 FILLCELL_X32 FILLER_275_1185 ();
 FILLCELL_X32 FILLER_275_1217 ();
 FILLCELL_X8 FILLER_275_1249 ();
 FILLCELL_X4 FILLER_275_1257 ();
 FILLCELL_X2 FILLER_275_1261 ();
 FILLCELL_X32 FILLER_275_1264 ();
 FILLCELL_X32 FILLER_275_1296 ();
 FILLCELL_X32 FILLER_275_1328 ();
 FILLCELL_X32 FILLER_275_1360 ();
 FILLCELL_X32 FILLER_275_1392 ();
 FILLCELL_X32 FILLER_275_1424 ();
 FILLCELL_X32 FILLER_275_1456 ();
 FILLCELL_X32 FILLER_275_1488 ();
 FILLCELL_X32 FILLER_275_1520 ();
 FILLCELL_X32 FILLER_275_1552 ();
 FILLCELL_X32 FILLER_275_1584 ();
 FILLCELL_X32 FILLER_275_1616 ();
 FILLCELL_X32 FILLER_275_1648 ();
 FILLCELL_X32 FILLER_275_1680 ();
 FILLCELL_X32 FILLER_275_1712 ();
 FILLCELL_X32 FILLER_275_1744 ();
 FILLCELL_X32 FILLER_275_1776 ();
 FILLCELL_X32 FILLER_275_1808 ();
 FILLCELL_X32 FILLER_275_1840 ();
 FILLCELL_X32 FILLER_275_1872 ();
 FILLCELL_X32 FILLER_275_1904 ();
 FILLCELL_X32 FILLER_275_1936 ();
 FILLCELL_X32 FILLER_275_1968 ();
 FILLCELL_X32 FILLER_275_2000 ();
 FILLCELL_X32 FILLER_275_2032 ();
 FILLCELL_X32 FILLER_275_2064 ();
 FILLCELL_X32 FILLER_275_2096 ();
 FILLCELL_X32 FILLER_275_2128 ();
 FILLCELL_X32 FILLER_275_2160 ();
 FILLCELL_X32 FILLER_275_2192 ();
 FILLCELL_X32 FILLER_275_2224 ();
 FILLCELL_X32 FILLER_275_2256 ();
 FILLCELL_X32 FILLER_275_2288 ();
 FILLCELL_X32 FILLER_275_2320 ();
 FILLCELL_X32 FILLER_275_2352 ();
 FILLCELL_X32 FILLER_275_2384 ();
 FILLCELL_X32 FILLER_275_2416 ();
 FILLCELL_X32 FILLER_275_2448 ();
 FILLCELL_X32 FILLER_275_2480 ();
 FILLCELL_X8 FILLER_275_2512 ();
 FILLCELL_X4 FILLER_275_2520 ();
 FILLCELL_X2 FILLER_275_2524 ();
 FILLCELL_X32 FILLER_275_2527 ();
 FILLCELL_X32 FILLER_275_2559 ();
 FILLCELL_X8 FILLER_275_2591 ();
 FILLCELL_X2 FILLER_275_2599 ();
 FILLCELL_X1 FILLER_275_2601 ();
 FILLCELL_X32 FILLER_276_1 ();
 FILLCELL_X32 FILLER_276_33 ();
 FILLCELL_X32 FILLER_276_65 ();
 FILLCELL_X32 FILLER_276_97 ();
 FILLCELL_X32 FILLER_276_129 ();
 FILLCELL_X32 FILLER_276_161 ();
 FILLCELL_X32 FILLER_276_193 ();
 FILLCELL_X32 FILLER_276_225 ();
 FILLCELL_X32 FILLER_276_257 ();
 FILLCELL_X32 FILLER_276_289 ();
 FILLCELL_X32 FILLER_276_321 ();
 FILLCELL_X32 FILLER_276_353 ();
 FILLCELL_X32 FILLER_276_385 ();
 FILLCELL_X32 FILLER_276_417 ();
 FILLCELL_X32 FILLER_276_449 ();
 FILLCELL_X32 FILLER_276_481 ();
 FILLCELL_X32 FILLER_276_513 ();
 FILLCELL_X32 FILLER_276_545 ();
 FILLCELL_X32 FILLER_276_577 ();
 FILLCELL_X16 FILLER_276_609 ();
 FILLCELL_X4 FILLER_276_625 ();
 FILLCELL_X2 FILLER_276_629 ();
 FILLCELL_X32 FILLER_276_632 ();
 FILLCELL_X32 FILLER_276_664 ();
 FILLCELL_X32 FILLER_276_696 ();
 FILLCELL_X32 FILLER_276_728 ();
 FILLCELL_X32 FILLER_276_760 ();
 FILLCELL_X32 FILLER_276_792 ();
 FILLCELL_X32 FILLER_276_824 ();
 FILLCELL_X32 FILLER_276_856 ();
 FILLCELL_X32 FILLER_276_888 ();
 FILLCELL_X32 FILLER_276_920 ();
 FILLCELL_X32 FILLER_276_952 ();
 FILLCELL_X32 FILLER_276_984 ();
 FILLCELL_X32 FILLER_276_1016 ();
 FILLCELL_X32 FILLER_276_1048 ();
 FILLCELL_X32 FILLER_276_1080 ();
 FILLCELL_X32 FILLER_276_1112 ();
 FILLCELL_X32 FILLER_276_1144 ();
 FILLCELL_X32 FILLER_276_1176 ();
 FILLCELL_X32 FILLER_276_1208 ();
 FILLCELL_X32 FILLER_276_1240 ();
 FILLCELL_X32 FILLER_276_1272 ();
 FILLCELL_X32 FILLER_276_1304 ();
 FILLCELL_X32 FILLER_276_1336 ();
 FILLCELL_X32 FILLER_276_1368 ();
 FILLCELL_X32 FILLER_276_1400 ();
 FILLCELL_X32 FILLER_276_1432 ();
 FILLCELL_X32 FILLER_276_1464 ();
 FILLCELL_X32 FILLER_276_1496 ();
 FILLCELL_X32 FILLER_276_1528 ();
 FILLCELL_X32 FILLER_276_1560 ();
 FILLCELL_X32 FILLER_276_1592 ();
 FILLCELL_X32 FILLER_276_1624 ();
 FILLCELL_X32 FILLER_276_1656 ();
 FILLCELL_X32 FILLER_276_1688 ();
 FILLCELL_X32 FILLER_276_1720 ();
 FILLCELL_X32 FILLER_276_1752 ();
 FILLCELL_X32 FILLER_276_1784 ();
 FILLCELL_X32 FILLER_276_1816 ();
 FILLCELL_X32 FILLER_276_1848 ();
 FILLCELL_X8 FILLER_276_1880 ();
 FILLCELL_X4 FILLER_276_1888 ();
 FILLCELL_X2 FILLER_276_1892 ();
 FILLCELL_X32 FILLER_276_1895 ();
 FILLCELL_X32 FILLER_276_1927 ();
 FILLCELL_X32 FILLER_276_1959 ();
 FILLCELL_X32 FILLER_276_1991 ();
 FILLCELL_X32 FILLER_276_2023 ();
 FILLCELL_X32 FILLER_276_2055 ();
 FILLCELL_X32 FILLER_276_2087 ();
 FILLCELL_X32 FILLER_276_2119 ();
 FILLCELL_X32 FILLER_276_2151 ();
 FILLCELL_X32 FILLER_276_2183 ();
 FILLCELL_X32 FILLER_276_2215 ();
 FILLCELL_X32 FILLER_276_2247 ();
 FILLCELL_X32 FILLER_276_2279 ();
 FILLCELL_X32 FILLER_276_2311 ();
 FILLCELL_X32 FILLER_276_2343 ();
 FILLCELL_X32 FILLER_276_2375 ();
 FILLCELL_X32 FILLER_276_2407 ();
 FILLCELL_X32 FILLER_276_2439 ();
 FILLCELL_X32 FILLER_276_2471 ();
 FILLCELL_X32 FILLER_276_2503 ();
 FILLCELL_X32 FILLER_276_2535 ();
 FILLCELL_X32 FILLER_276_2567 ();
 FILLCELL_X2 FILLER_276_2599 ();
 FILLCELL_X1 FILLER_276_2601 ();
 FILLCELL_X32 FILLER_277_1 ();
 FILLCELL_X32 FILLER_277_33 ();
 FILLCELL_X32 FILLER_277_65 ();
 FILLCELL_X32 FILLER_277_97 ();
 FILLCELL_X32 FILLER_277_129 ();
 FILLCELL_X32 FILLER_277_161 ();
 FILLCELL_X32 FILLER_277_193 ();
 FILLCELL_X32 FILLER_277_225 ();
 FILLCELL_X32 FILLER_277_257 ();
 FILLCELL_X32 FILLER_277_289 ();
 FILLCELL_X32 FILLER_277_321 ();
 FILLCELL_X32 FILLER_277_353 ();
 FILLCELL_X32 FILLER_277_385 ();
 FILLCELL_X32 FILLER_277_417 ();
 FILLCELL_X32 FILLER_277_449 ();
 FILLCELL_X32 FILLER_277_481 ();
 FILLCELL_X32 FILLER_277_513 ();
 FILLCELL_X32 FILLER_277_545 ();
 FILLCELL_X32 FILLER_277_577 ();
 FILLCELL_X32 FILLER_277_609 ();
 FILLCELL_X32 FILLER_277_641 ();
 FILLCELL_X32 FILLER_277_673 ();
 FILLCELL_X32 FILLER_277_705 ();
 FILLCELL_X32 FILLER_277_737 ();
 FILLCELL_X32 FILLER_277_769 ();
 FILLCELL_X32 FILLER_277_801 ();
 FILLCELL_X32 FILLER_277_833 ();
 FILLCELL_X32 FILLER_277_865 ();
 FILLCELL_X32 FILLER_277_897 ();
 FILLCELL_X32 FILLER_277_929 ();
 FILLCELL_X32 FILLER_277_961 ();
 FILLCELL_X32 FILLER_277_993 ();
 FILLCELL_X32 FILLER_277_1025 ();
 FILLCELL_X32 FILLER_277_1057 ();
 FILLCELL_X32 FILLER_277_1089 ();
 FILLCELL_X32 FILLER_277_1121 ();
 FILLCELL_X32 FILLER_277_1153 ();
 FILLCELL_X32 FILLER_277_1185 ();
 FILLCELL_X32 FILLER_277_1217 ();
 FILLCELL_X8 FILLER_277_1249 ();
 FILLCELL_X4 FILLER_277_1257 ();
 FILLCELL_X2 FILLER_277_1261 ();
 FILLCELL_X32 FILLER_277_1264 ();
 FILLCELL_X32 FILLER_277_1296 ();
 FILLCELL_X32 FILLER_277_1328 ();
 FILLCELL_X32 FILLER_277_1360 ();
 FILLCELL_X32 FILLER_277_1392 ();
 FILLCELL_X32 FILLER_277_1424 ();
 FILLCELL_X32 FILLER_277_1456 ();
 FILLCELL_X32 FILLER_277_1488 ();
 FILLCELL_X32 FILLER_277_1520 ();
 FILLCELL_X32 FILLER_277_1552 ();
 FILLCELL_X32 FILLER_277_1584 ();
 FILLCELL_X32 FILLER_277_1616 ();
 FILLCELL_X32 FILLER_277_1648 ();
 FILLCELL_X32 FILLER_277_1680 ();
 FILLCELL_X32 FILLER_277_1712 ();
 FILLCELL_X32 FILLER_277_1744 ();
 FILLCELL_X32 FILLER_277_1776 ();
 FILLCELL_X32 FILLER_277_1808 ();
 FILLCELL_X32 FILLER_277_1840 ();
 FILLCELL_X32 FILLER_277_1872 ();
 FILLCELL_X32 FILLER_277_1904 ();
 FILLCELL_X32 FILLER_277_1936 ();
 FILLCELL_X32 FILLER_277_1968 ();
 FILLCELL_X32 FILLER_277_2000 ();
 FILLCELL_X32 FILLER_277_2032 ();
 FILLCELL_X32 FILLER_277_2064 ();
 FILLCELL_X32 FILLER_277_2096 ();
 FILLCELL_X32 FILLER_277_2128 ();
 FILLCELL_X32 FILLER_277_2160 ();
 FILLCELL_X32 FILLER_277_2192 ();
 FILLCELL_X32 FILLER_277_2224 ();
 FILLCELL_X32 FILLER_277_2256 ();
 FILLCELL_X32 FILLER_277_2288 ();
 FILLCELL_X32 FILLER_277_2320 ();
 FILLCELL_X32 FILLER_277_2352 ();
 FILLCELL_X32 FILLER_277_2384 ();
 FILLCELL_X32 FILLER_277_2416 ();
 FILLCELL_X32 FILLER_277_2448 ();
 FILLCELL_X32 FILLER_277_2480 ();
 FILLCELL_X8 FILLER_277_2512 ();
 FILLCELL_X4 FILLER_277_2520 ();
 FILLCELL_X2 FILLER_277_2524 ();
 FILLCELL_X32 FILLER_277_2527 ();
 FILLCELL_X32 FILLER_277_2559 ();
 FILLCELL_X8 FILLER_277_2591 ();
 FILLCELL_X2 FILLER_277_2599 ();
 FILLCELL_X1 FILLER_277_2601 ();
 FILLCELL_X32 FILLER_278_1 ();
 FILLCELL_X32 FILLER_278_33 ();
 FILLCELL_X32 FILLER_278_65 ();
 FILLCELL_X32 FILLER_278_97 ();
 FILLCELL_X32 FILLER_278_129 ();
 FILLCELL_X32 FILLER_278_161 ();
 FILLCELL_X32 FILLER_278_193 ();
 FILLCELL_X32 FILLER_278_225 ();
 FILLCELL_X32 FILLER_278_257 ();
 FILLCELL_X32 FILLER_278_289 ();
 FILLCELL_X32 FILLER_278_321 ();
 FILLCELL_X32 FILLER_278_353 ();
 FILLCELL_X32 FILLER_278_385 ();
 FILLCELL_X32 FILLER_278_417 ();
 FILLCELL_X32 FILLER_278_449 ();
 FILLCELL_X32 FILLER_278_481 ();
 FILLCELL_X32 FILLER_278_513 ();
 FILLCELL_X32 FILLER_278_545 ();
 FILLCELL_X32 FILLER_278_577 ();
 FILLCELL_X16 FILLER_278_609 ();
 FILLCELL_X4 FILLER_278_625 ();
 FILLCELL_X2 FILLER_278_629 ();
 FILLCELL_X32 FILLER_278_632 ();
 FILLCELL_X32 FILLER_278_664 ();
 FILLCELL_X32 FILLER_278_696 ();
 FILLCELL_X32 FILLER_278_728 ();
 FILLCELL_X32 FILLER_278_760 ();
 FILLCELL_X32 FILLER_278_792 ();
 FILLCELL_X32 FILLER_278_824 ();
 FILLCELL_X32 FILLER_278_856 ();
 FILLCELL_X32 FILLER_278_888 ();
 FILLCELL_X32 FILLER_278_920 ();
 FILLCELL_X32 FILLER_278_952 ();
 FILLCELL_X32 FILLER_278_984 ();
 FILLCELL_X32 FILLER_278_1016 ();
 FILLCELL_X32 FILLER_278_1048 ();
 FILLCELL_X32 FILLER_278_1080 ();
 FILLCELL_X32 FILLER_278_1112 ();
 FILLCELL_X32 FILLER_278_1144 ();
 FILLCELL_X32 FILLER_278_1176 ();
 FILLCELL_X32 FILLER_278_1208 ();
 FILLCELL_X32 FILLER_278_1240 ();
 FILLCELL_X32 FILLER_278_1272 ();
 FILLCELL_X32 FILLER_278_1304 ();
 FILLCELL_X32 FILLER_278_1336 ();
 FILLCELL_X32 FILLER_278_1368 ();
 FILLCELL_X32 FILLER_278_1400 ();
 FILLCELL_X32 FILLER_278_1432 ();
 FILLCELL_X32 FILLER_278_1464 ();
 FILLCELL_X32 FILLER_278_1496 ();
 FILLCELL_X32 FILLER_278_1528 ();
 FILLCELL_X32 FILLER_278_1560 ();
 FILLCELL_X32 FILLER_278_1592 ();
 FILLCELL_X32 FILLER_278_1624 ();
 FILLCELL_X32 FILLER_278_1656 ();
 FILLCELL_X32 FILLER_278_1688 ();
 FILLCELL_X32 FILLER_278_1720 ();
 FILLCELL_X32 FILLER_278_1752 ();
 FILLCELL_X32 FILLER_278_1784 ();
 FILLCELL_X32 FILLER_278_1816 ();
 FILLCELL_X32 FILLER_278_1848 ();
 FILLCELL_X8 FILLER_278_1880 ();
 FILLCELL_X4 FILLER_278_1888 ();
 FILLCELL_X2 FILLER_278_1892 ();
 FILLCELL_X32 FILLER_278_1895 ();
 FILLCELL_X32 FILLER_278_1927 ();
 FILLCELL_X32 FILLER_278_1959 ();
 FILLCELL_X32 FILLER_278_1991 ();
 FILLCELL_X32 FILLER_278_2023 ();
 FILLCELL_X32 FILLER_278_2055 ();
 FILLCELL_X32 FILLER_278_2087 ();
 FILLCELL_X32 FILLER_278_2119 ();
 FILLCELL_X32 FILLER_278_2151 ();
 FILLCELL_X32 FILLER_278_2183 ();
 FILLCELL_X32 FILLER_278_2215 ();
 FILLCELL_X32 FILLER_278_2247 ();
 FILLCELL_X32 FILLER_278_2279 ();
 FILLCELL_X32 FILLER_278_2311 ();
 FILLCELL_X32 FILLER_278_2343 ();
 FILLCELL_X32 FILLER_278_2375 ();
 FILLCELL_X32 FILLER_278_2407 ();
 FILLCELL_X32 FILLER_278_2439 ();
 FILLCELL_X32 FILLER_278_2471 ();
 FILLCELL_X32 FILLER_278_2503 ();
 FILLCELL_X32 FILLER_278_2535 ();
 FILLCELL_X32 FILLER_278_2567 ();
 FILLCELL_X2 FILLER_278_2599 ();
 FILLCELL_X1 FILLER_278_2601 ();
 FILLCELL_X32 FILLER_279_1 ();
 FILLCELL_X32 FILLER_279_33 ();
 FILLCELL_X32 FILLER_279_65 ();
 FILLCELL_X32 FILLER_279_97 ();
 FILLCELL_X32 FILLER_279_129 ();
 FILLCELL_X32 FILLER_279_161 ();
 FILLCELL_X32 FILLER_279_193 ();
 FILLCELL_X32 FILLER_279_225 ();
 FILLCELL_X32 FILLER_279_257 ();
 FILLCELL_X32 FILLER_279_289 ();
 FILLCELL_X32 FILLER_279_321 ();
 FILLCELL_X32 FILLER_279_353 ();
 FILLCELL_X32 FILLER_279_385 ();
 FILLCELL_X32 FILLER_279_417 ();
 FILLCELL_X32 FILLER_279_449 ();
 FILLCELL_X32 FILLER_279_481 ();
 FILLCELL_X32 FILLER_279_513 ();
 FILLCELL_X32 FILLER_279_545 ();
 FILLCELL_X32 FILLER_279_577 ();
 FILLCELL_X32 FILLER_279_609 ();
 FILLCELL_X32 FILLER_279_641 ();
 FILLCELL_X32 FILLER_279_673 ();
 FILLCELL_X32 FILLER_279_705 ();
 FILLCELL_X32 FILLER_279_737 ();
 FILLCELL_X32 FILLER_279_769 ();
 FILLCELL_X32 FILLER_279_801 ();
 FILLCELL_X32 FILLER_279_833 ();
 FILLCELL_X32 FILLER_279_865 ();
 FILLCELL_X32 FILLER_279_897 ();
 FILLCELL_X32 FILLER_279_929 ();
 FILLCELL_X32 FILLER_279_961 ();
 FILLCELL_X32 FILLER_279_993 ();
 FILLCELL_X32 FILLER_279_1025 ();
 FILLCELL_X32 FILLER_279_1057 ();
 FILLCELL_X32 FILLER_279_1089 ();
 FILLCELL_X32 FILLER_279_1121 ();
 FILLCELL_X32 FILLER_279_1153 ();
 FILLCELL_X32 FILLER_279_1185 ();
 FILLCELL_X32 FILLER_279_1217 ();
 FILLCELL_X8 FILLER_279_1249 ();
 FILLCELL_X4 FILLER_279_1257 ();
 FILLCELL_X2 FILLER_279_1261 ();
 FILLCELL_X32 FILLER_279_1264 ();
 FILLCELL_X32 FILLER_279_1296 ();
 FILLCELL_X32 FILLER_279_1328 ();
 FILLCELL_X32 FILLER_279_1360 ();
 FILLCELL_X32 FILLER_279_1392 ();
 FILLCELL_X32 FILLER_279_1424 ();
 FILLCELL_X32 FILLER_279_1456 ();
 FILLCELL_X32 FILLER_279_1488 ();
 FILLCELL_X32 FILLER_279_1520 ();
 FILLCELL_X32 FILLER_279_1552 ();
 FILLCELL_X32 FILLER_279_1584 ();
 FILLCELL_X32 FILLER_279_1616 ();
 FILLCELL_X32 FILLER_279_1648 ();
 FILLCELL_X32 FILLER_279_1680 ();
 FILLCELL_X32 FILLER_279_1712 ();
 FILLCELL_X32 FILLER_279_1744 ();
 FILLCELL_X32 FILLER_279_1776 ();
 FILLCELL_X32 FILLER_279_1808 ();
 FILLCELL_X32 FILLER_279_1840 ();
 FILLCELL_X32 FILLER_279_1872 ();
 FILLCELL_X32 FILLER_279_1904 ();
 FILLCELL_X32 FILLER_279_1936 ();
 FILLCELL_X32 FILLER_279_1968 ();
 FILLCELL_X32 FILLER_279_2000 ();
 FILLCELL_X32 FILLER_279_2032 ();
 FILLCELL_X32 FILLER_279_2064 ();
 FILLCELL_X32 FILLER_279_2096 ();
 FILLCELL_X32 FILLER_279_2128 ();
 FILLCELL_X32 FILLER_279_2160 ();
 FILLCELL_X32 FILLER_279_2192 ();
 FILLCELL_X32 FILLER_279_2224 ();
 FILLCELL_X32 FILLER_279_2256 ();
 FILLCELL_X32 FILLER_279_2288 ();
 FILLCELL_X32 FILLER_279_2320 ();
 FILLCELL_X32 FILLER_279_2352 ();
 FILLCELL_X32 FILLER_279_2384 ();
 FILLCELL_X32 FILLER_279_2416 ();
 FILLCELL_X32 FILLER_279_2448 ();
 FILLCELL_X32 FILLER_279_2480 ();
 FILLCELL_X8 FILLER_279_2512 ();
 FILLCELL_X4 FILLER_279_2520 ();
 FILLCELL_X2 FILLER_279_2524 ();
 FILLCELL_X32 FILLER_279_2527 ();
 FILLCELL_X32 FILLER_279_2559 ();
 FILLCELL_X8 FILLER_279_2591 ();
 FILLCELL_X2 FILLER_279_2599 ();
 FILLCELL_X1 FILLER_279_2601 ();
 FILLCELL_X32 FILLER_280_1 ();
 FILLCELL_X32 FILLER_280_33 ();
 FILLCELL_X32 FILLER_280_65 ();
 FILLCELL_X32 FILLER_280_97 ();
 FILLCELL_X32 FILLER_280_129 ();
 FILLCELL_X32 FILLER_280_161 ();
 FILLCELL_X32 FILLER_280_193 ();
 FILLCELL_X32 FILLER_280_225 ();
 FILLCELL_X32 FILLER_280_257 ();
 FILLCELL_X32 FILLER_280_289 ();
 FILLCELL_X32 FILLER_280_321 ();
 FILLCELL_X32 FILLER_280_353 ();
 FILLCELL_X32 FILLER_280_385 ();
 FILLCELL_X32 FILLER_280_417 ();
 FILLCELL_X32 FILLER_280_449 ();
 FILLCELL_X32 FILLER_280_481 ();
 FILLCELL_X32 FILLER_280_513 ();
 FILLCELL_X32 FILLER_280_545 ();
 FILLCELL_X32 FILLER_280_577 ();
 FILLCELL_X16 FILLER_280_609 ();
 FILLCELL_X4 FILLER_280_625 ();
 FILLCELL_X2 FILLER_280_629 ();
 FILLCELL_X32 FILLER_280_632 ();
 FILLCELL_X32 FILLER_280_664 ();
 FILLCELL_X32 FILLER_280_696 ();
 FILLCELL_X32 FILLER_280_728 ();
 FILLCELL_X32 FILLER_280_760 ();
 FILLCELL_X32 FILLER_280_792 ();
 FILLCELL_X32 FILLER_280_824 ();
 FILLCELL_X32 FILLER_280_856 ();
 FILLCELL_X32 FILLER_280_888 ();
 FILLCELL_X32 FILLER_280_920 ();
 FILLCELL_X32 FILLER_280_952 ();
 FILLCELL_X32 FILLER_280_984 ();
 FILLCELL_X32 FILLER_280_1016 ();
 FILLCELL_X32 FILLER_280_1048 ();
 FILLCELL_X32 FILLER_280_1080 ();
 FILLCELL_X32 FILLER_280_1112 ();
 FILLCELL_X32 FILLER_280_1144 ();
 FILLCELL_X32 FILLER_280_1176 ();
 FILLCELL_X32 FILLER_280_1208 ();
 FILLCELL_X32 FILLER_280_1240 ();
 FILLCELL_X32 FILLER_280_1272 ();
 FILLCELL_X32 FILLER_280_1304 ();
 FILLCELL_X32 FILLER_280_1336 ();
 FILLCELL_X32 FILLER_280_1368 ();
 FILLCELL_X32 FILLER_280_1400 ();
 FILLCELL_X32 FILLER_280_1432 ();
 FILLCELL_X32 FILLER_280_1464 ();
 FILLCELL_X32 FILLER_280_1496 ();
 FILLCELL_X32 FILLER_280_1528 ();
 FILLCELL_X32 FILLER_280_1560 ();
 FILLCELL_X32 FILLER_280_1592 ();
 FILLCELL_X32 FILLER_280_1624 ();
 FILLCELL_X32 FILLER_280_1656 ();
 FILLCELL_X32 FILLER_280_1688 ();
 FILLCELL_X32 FILLER_280_1720 ();
 FILLCELL_X32 FILLER_280_1752 ();
 FILLCELL_X32 FILLER_280_1784 ();
 FILLCELL_X32 FILLER_280_1816 ();
 FILLCELL_X32 FILLER_280_1848 ();
 FILLCELL_X8 FILLER_280_1880 ();
 FILLCELL_X4 FILLER_280_1888 ();
 FILLCELL_X2 FILLER_280_1892 ();
 FILLCELL_X32 FILLER_280_1895 ();
 FILLCELL_X32 FILLER_280_1927 ();
 FILLCELL_X32 FILLER_280_1959 ();
 FILLCELL_X32 FILLER_280_1991 ();
 FILLCELL_X32 FILLER_280_2023 ();
 FILLCELL_X32 FILLER_280_2055 ();
 FILLCELL_X32 FILLER_280_2087 ();
 FILLCELL_X32 FILLER_280_2119 ();
 FILLCELL_X32 FILLER_280_2151 ();
 FILLCELL_X32 FILLER_280_2183 ();
 FILLCELL_X32 FILLER_280_2215 ();
 FILLCELL_X32 FILLER_280_2247 ();
 FILLCELL_X32 FILLER_280_2279 ();
 FILLCELL_X32 FILLER_280_2311 ();
 FILLCELL_X32 FILLER_280_2343 ();
 FILLCELL_X32 FILLER_280_2375 ();
 FILLCELL_X32 FILLER_280_2407 ();
 FILLCELL_X32 FILLER_280_2439 ();
 FILLCELL_X32 FILLER_280_2471 ();
 FILLCELL_X32 FILLER_280_2503 ();
 FILLCELL_X32 FILLER_280_2535 ();
 FILLCELL_X32 FILLER_280_2567 ();
 FILLCELL_X2 FILLER_280_2599 ();
 FILLCELL_X1 FILLER_280_2601 ();
 FILLCELL_X32 FILLER_281_1 ();
 FILLCELL_X32 FILLER_281_33 ();
 FILLCELL_X32 FILLER_281_65 ();
 FILLCELL_X32 FILLER_281_97 ();
 FILLCELL_X32 FILLER_281_129 ();
 FILLCELL_X32 FILLER_281_161 ();
 FILLCELL_X32 FILLER_281_193 ();
 FILLCELL_X32 FILLER_281_225 ();
 FILLCELL_X32 FILLER_281_257 ();
 FILLCELL_X32 FILLER_281_289 ();
 FILLCELL_X32 FILLER_281_321 ();
 FILLCELL_X32 FILLER_281_353 ();
 FILLCELL_X32 FILLER_281_385 ();
 FILLCELL_X32 FILLER_281_417 ();
 FILLCELL_X32 FILLER_281_449 ();
 FILLCELL_X32 FILLER_281_481 ();
 FILLCELL_X32 FILLER_281_513 ();
 FILLCELL_X32 FILLER_281_545 ();
 FILLCELL_X32 FILLER_281_577 ();
 FILLCELL_X32 FILLER_281_609 ();
 FILLCELL_X32 FILLER_281_641 ();
 FILLCELL_X32 FILLER_281_673 ();
 FILLCELL_X32 FILLER_281_705 ();
 FILLCELL_X32 FILLER_281_737 ();
 FILLCELL_X32 FILLER_281_769 ();
 FILLCELL_X32 FILLER_281_801 ();
 FILLCELL_X32 FILLER_281_833 ();
 FILLCELL_X32 FILLER_281_865 ();
 FILLCELL_X32 FILLER_281_897 ();
 FILLCELL_X32 FILLER_281_929 ();
 FILLCELL_X32 FILLER_281_961 ();
 FILLCELL_X32 FILLER_281_993 ();
 FILLCELL_X32 FILLER_281_1025 ();
 FILLCELL_X32 FILLER_281_1057 ();
 FILLCELL_X32 FILLER_281_1089 ();
 FILLCELL_X32 FILLER_281_1121 ();
 FILLCELL_X32 FILLER_281_1153 ();
 FILLCELL_X32 FILLER_281_1185 ();
 FILLCELL_X32 FILLER_281_1217 ();
 FILLCELL_X8 FILLER_281_1249 ();
 FILLCELL_X4 FILLER_281_1257 ();
 FILLCELL_X2 FILLER_281_1261 ();
 FILLCELL_X32 FILLER_281_1264 ();
 FILLCELL_X32 FILLER_281_1296 ();
 FILLCELL_X32 FILLER_281_1328 ();
 FILLCELL_X32 FILLER_281_1360 ();
 FILLCELL_X32 FILLER_281_1392 ();
 FILLCELL_X32 FILLER_281_1424 ();
 FILLCELL_X32 FILLER_281_1456 ();
 FILLCELL_X32 FILLER_281_1488 ();
 FILLCELL_X32 FILLER_281_1520 ();
 FILLCELL_X32 FILLER_281_1552 ();
 FILLCELL_X32 FILLER_281_1584 ();
 FILLCELL_X32 FILLER_281_1616 ();
 FILLCELL_X32 FILLER_281_1648 ();
 FILLCELL_X32 FILLER_281_1680 ();
 FILLCELL_X32 FILLER_281_1712 ();
 FILLCELL_X32 FILLER_281_1744 ();
 FILLCELL_X32 FILLER_281_1776 ();
 FILLCELL_X32 FILLER_281_1808 ();
 FILLCELL_X32 FILLER_281_1840 ();
 FILLCELL_X32 FILLER_281_1872 ();
 FILLCELL_X32 FILLER_281_1904 ();
 FILLCELL_X32 FILLER_281_1936 ();
 FILLCELL_X32 FILLER_281_1968 ();
 FILLCELL_X32 FILLER_281_2000 ();
 FILLCELL_X32 FILLER_281_2032 ();
 FILLCELL_X32 FILLER_281_2064 ();
 FILLCELL_X32 FILLER_281_2096 ();
 FILLCELL_X32 FILLER_281_2128 ();
 FILLCELL_X32 FILLER_281_2160 ();
 FILLCELL_X32 FILLER_281_2192 ();
 FILLCELL_X32 FILLER_281_2224 ();
 FILLCELL_X32 FILLER_281_2256 ();
 FILLCELL_X32 FILLER_281_2288 ();
 FILLCELL_X32 FILLER_281_2320 ();
 FILLCELL_X32 FILLER_281_2352 ();
 FILLCELL_X32 FILLER_281_2384 ();
 FILLCELL_X32 FILLER_281_2416 ();
 FILLCELL_X32 FILLER_281_2448 ();
 FILLCELL_X32 FILLER_281_2480 ();
 FILLCELL_X8 FILLER_281_2512 ();
 FILLCELL_X4 FILLER_281_2520 ();
 FILLCELL_X2 FILLER_281_2524 ();
 FILLCELL_X32 FILLER_281_2527 ();
 FILLCELL_X32 FILLER_281_2559 ();
 FILLCELL_X8 FILLER_281_2591 ();
 FILLCELL_X2 FILLER_281_2599 ();
 FILLCELL_X1 FILLER_281_2601 ();
 FILLCELL_X32 FILLER_282_1 ();
 FILLCELL_X32 FILLER_282_33 ();
 FILLCELL_X32 FILLER_282_65 ();
 FILLCELL_X32 FILLER_282_97 ();
 FILLCELL_X32 FILLER_282_129 ();
 FILLCELL_X32 FILLER_282_161 ();
 FILLCELL_X32 FILLER_282_193 ();
 FILLCELL_X32 FILLER_282_225 ();
 FILLCELL_X32 FILLER_282_257 ();
 FILLCELL_X32 FILLER_282_289 ();
 FILLCELL_X32 FILLER_282_321 ();
 FILLCELL_X32 FILLER_282_353 ();
 FILLCELL_X32 FILLER_282_385 ();
 FILLCELL_X32 FILLER_282_417 ();
 FILLCELL_X32 FILLER_282_449 ();
 FILLCELL_X32 FILLER_282_481 ();
 FILLCELL_X32 FILLER_282_513 ();
 FILLCELL_X32 FILLER_282_545 ();
 FILLCELL_X32 FILLER_282_577 ();
 FILLCELL_X16 FILLER_282_609 ();
 FILLCELL_X4 FILLER_282_625 ();
 FILLCELL_X2 FILLER_282_629 ();
 FILLCELL_X32 FILLER_282_632 ();
 FILLCELL_X32 FILLER_282_664 ();
 FILLCELL_X32 FILLER_282_696 ();
 FILLCELL_X32 FILLER_282_728 ();
 FILLCELL_X32 FILLER_282_760 ();
 FILLCELL_X32 FILLER_282_792 ();
 FILLCELL_X32 FILLER_282_824 ();
 FILLCELL_X32 FILLER_282_856 ();
 FILLCELL_X32 FILLER_282_888 ();
 FILLCELL_X32 FILLER_282_920 ();
 FILLCELL_X32 FILLER_282_952 ();
 FILLCELL_X32 FILLER_282_984 ();
 FILLCELL_X32 FILLER_282_1016 ();
 FILLCELL_X32 FILLER_282_1048 ();
 FILLCELL_X32 FILLER_282_1080 ();
 FILLCELL_X32 FILLER_282_1112 ();
 FILLCELL_X32 FILLER_282_1144 ();
 FILLCELL_X32 FILLER_282_1176 ();
 FILLCELL_X32 FILLER_282_1208 ();
 FILLCELL_X32 FILLER_282_1240 ();
 FILLCELL_X32 FILLER_282_1272 ();
 FILLCELL_X32 FILLER_282_1304 ();
 FILLCELL_X32 FILLER_282_1336 ();
 FILLCELL_X32 FILLER_282_1368 ();
 FILLCELL_X32 FILLER_282_1400 ();
 FILLCELL_X32 FILLER_282_1432 ();
 FILLCELL_X32 FILLER_282_1464 ();
 FILLCELL_X32 FILLER_282_1496 ();
 FILLCELL_X32 FILLER_282_1528 ();
 FILLCELL_X32 FILLER_282_1560 ();
 FILLCELL_X32 FILLER_282_1592 ();
 FILLCELL_X32 FILLER_282_1624 ();
 FILLCELL_X32 FILLER_282_1656 ();
 FILLCELL_X32 FILLER_282_1688 ();
 FILLCELL_X32 FILLER_282_1720 ();
 FILLCELL_X32 FILLER_282_1752 ();
 FILLCELL_X32 FILLER_282_1784 ();
 FILLCELL_X32 FILLER_282_1816 ();
 FILLCELL_X32 FILLER_282_1848 ();
 FILLCELL_X8 FILLER_282_1880 ();
 FILLCELL_X4 FILLER_282_1888 ();
 FILLCELL_X2 FILLER_282_1892 ();
 FILLCELL_X32 FILLER_282_1895 ();
 FILLCELL_X32 FILLER_282_1927 ();
 FILLCELL_X32 FILLER_282_1959 ();
 FILLCELL_X32 FILLER_282_1991 ();
 FILLCELL_X32 FILLER_282_2023 ();
 FILLCELL_X32 FILLER_282_2055 ();
 FILLCELL_X32 FILLER_282_2087 ();
 FILLCELL_X32 FILLER_282_2119 ();
 FILLCELL_X32 FILLER_282_2151 ();
 FILLCELL_X32 FILLER_282_2183 ();
 FILLCELL_X32 FILLER_282_2215 ();
 FILLCELL_X32 FILLER_282_2247 ();
 FILLCELL_X32 FILLER_282_2279 ();
 FILLCELL_X32 FILLER_282_2311 ();
 FILLCELL_X32 FILLER_282_2343 ();
 FILLCELL_X32 FILLER_282_2375 ();
 FILLCELL_X32 FILLER_282_2407 ();
 FILLCELL_X32 FILLER_282_2439 ();
 FILLCELL_X32 FILLER_282_2471 ();
 FILLCELL_X32 FILLER_282_2503 ();
 FILLCELL_X32 FILLER_282_2535 ();
 FILLCELL_X32 FILLER_282_2567 ();
 FILLCELL_X2 FILLER_282_2599 ();
 FILLCELL_X1 FILLER_282_2601 ();
 FILLCELL_X32 FILLER_283_1 ();
 FILLCELL_X32 FILLER_283_33 ();
 FILLCELL_X32 FILLER_283_65 ();
 FILLCELL_X32 FILLER_283_97 ();
 FILLCELL_X32 FILLER_283_129 ();
 FILLCELL_X32 FILLER_283_161 ();
 FILLCELL_X32 FILLER_283_193 ();
 FILLCELL_X32 FILLER_283_225 ();
 FILLCELL_X32 FILLER_283_257 ();
 FILLCELL_X32 FILLER_283_289 ();
 FILLCELL_X32 FILLER_283_321 ();
 FILLCELL_X32 FILLER_283_353 ();
 FILLCELL_X32 FILLER_283_385 ();
 FILLCELL_X32 FILLER_283_417 ();
 FILLCELL_X32 FILLER_283_449 ();
 FILLCELL_X32 FILLER_283_481 ();
 FILLCELL_X32 FILLER_283_513 ();
 FILLCELL_X32 FILLER_283_545 ();
 FILLCELL_X32 FILLER_283_577 ();
 FILLCELL_X32 FILLER_283_609 ();
 FILLCELL_X32 FILLER_283_641 ();
 FILLCELL_X32 FILLER_283_673 ();
 FILLCELL_X32 FILLER_283_705 ();
 FILLCELL_X32 FILLER_283_737 ();
 FILLCELL_X32 FILLER_283_769 ();
 FILLCELL_X32 FILLER_283_801 ();
 FILLCELL_X32 FILLER_283_833 ();
 FILLCELL_X32 FILLER_283_865 ();
 FILLCELL_X32 FILLER_283_897 ();
 FILLCELL_X32 FILLER_283_929 ();
 FILLCELL_X32 FILLER_283_961 ();
 FILLCELL_X32 FILLER_283_993 ();
 FILLCELL_X32 FILLER_283_1025 ();
 FILLCELL_X32 FILLER_283_1057 ();
 FILLCELL_X32 FILLER_283_1089 ();
 FILLCELL_X32 FILLER_283_1121 ();
 FILLCELL_X32 FILLER_283_1153 ();
 FILLCELL_X32 FILLER_283_1185 ();
 FILLCELL_X32 FILLER_283_1217 ();
 FILLCELL_X8 FILLER_283_1249 ();
 FILLCELL_X4 FILLER_283_1257 ();
 FILLCELL_X2 FILLER_283_1261 ();
 FILLCELL_X32 FILLER_283_1264 ();
 FILLCELL_X32 FILLER_283_1296 ();
 FILLCELL_X32 FILLER_283_1328 ();
 FILLCELL_X32 FILLER_283_1360 ();
 FILLCELL_X32 FILLER_283_1392 ();
 FILLCELL_X32 FILLER_283_1424 ();
 FILLCELL_X32 FILLER_283_1456 ();
 FILLCELL_X32 FILLER_283_1488 ();
 FILLCELL_X32 FILLER_283_1520 ();
 FILLCELL_X32 FILLER_283_1552 ();
 FILLCELL_X32 FILLER_283_1584 ();
 FILLCELL_X32 FILLER_283_1616 ();
 FILLCELL_X32 FILLER_283_1648 ();
 FILLCELL_X32 FILLER_283_1680 ();
 FILLCELL_X32 FILLER_283_1712 ();
 FILLCELL_X32 FILLER_283_1744 ();
 FILLCELL_X32 FILLER_283_1776 ();
 FILLCELL_X32 FILLER_283_1808 ();
 FILLCELL_X32 FILLER_283_1840 ();
 FILLCELL_X32 FILLER_283_1872 ();
 FILLCELL_X32 FILLER_283_1904 ();
 FILLCELL_X32 FILLER_283_1936 ();
 FILLCELL_X32 FILLER_283_1968 ();
 FILLCELL_X32 FILLER_283_2000 ();
 FILLCELL_X32 FILLER_283_2032 ();
 FILLCELL_X32 FILLER_283_2064 ();
 FILLCELL_X32 FILLER_283_2096 ();
 FILLCELL_X32 FILLER_283_2128 ();
 FILLCELL_X32 FILLER_283_2160 ();
 FILLCELL_X32 FILLER_283_2192 ();
 FILLCELL_X32 FILLER_283_2224 ();
 FILLCELL_X32 FILLER_283_2256 ();
 FILLCELL_X32 FILLER_283_2288 ();
 FILLCELL_X32 FILLER_283_2320 ();
 FILLCELL_X32 FILLER_283_2352 ();
 FILLCELL_X32 FILLER_283_2384 ();
 FILLCELL_X32 FILLER_283_2416 ();
 FILLCELL_X32 FILLER_283_2448 ();
 FILLCELL_X32 FILLER_283_2480 ();
 FILLCELL_X8 FILLER_283_2512 ();
 FILLCELL_X4 FILLER_283_2520 ();
 FILLCELL_X2 FILLER_283_2524 ();
 FILLCELL_X32 FILLER_283_2527 ();
 FILLCELL_X32 FILLER_283_2559 ();
 FILLCELL_X8 FILLER_283_2591 ();
 FILLCELL_X2 FILLER_283_2599 ();
 FILLCELL_X1 FILLER_283_2601 ();
 FILLCELL_X32 FILLER_284_1 ();
 FILLCELL_X32 FILLER_284_33 ();
 FILLCELL_X32 FILLER_284_65 ();
 FILLCELL_X32 FILLER_284_97 ();
 FILLCELL_X32 FILLER_284_129 ();
 FILLCELL_X32 FILLER_284_161 ();
 FILLCELL_X32 FILLER_284_193 ();
 FILLCELL_X32 FILLER_284_225 ();
 FILLCELL_X32 FILLER_284_257 ();
 FILLCELL_X32 FILLER_284_289 ();
 FILLCELL_X32 FILLER_284_321 ();
 FILLCELL_X32 FILLER_284_353 ();
 FILLCELL_X32 FILLER_284_385 ();
 FILLCELL_X32 FILLER_284_417 ();
 FILLCELL_X32 FILLER_284_449 ();
 FILLCELL_X32 FILLER_284_481 ();
 FILLCELL_X32 FILLER_284_513 ();
 FILLCELL_X32 FILLER_284_545 ();
 FILLCELL_X32 FILLER_284_577 ();
 FILLCELL_X16 FILLER_284_609 ();
 FILLCELL_X4 FILLER_284_625 ();
 FILLCELL_X2 FILLER_284_629 ();
 FILLCELL_X32 FILLER_284_632 ();
 FILLCELL_X32 FILLER_284_664 ();
 FILLCELL_X32 FILLER_284_696 ();
 FILLCELL_X32 FILLER_284_728 ();
 FILLCELL_X32 FILLER_284_760 ();
 FILLCELL_X32 FILLER_284_792 ();
 FILLCELL_X32 FILLER_284_824 ();
 FILLCELL_X32 FILLER_284_856 ();
 FILLCELL_X32 FILLER_284_888 ();
 FILLCELL_X32 FILLER_284_920 ();
 FILLCELL_X32 FILLER_284_952 ();
 FILLCELL_X32 FILLER_284_984 ();
 FILLCELL_X32 FILLER_284_1016 ();
 FILLCELL_X32 FILLER_284_1048 ();
 FILLCELL_X32 FILLER_284_1080 ();
 FILLCELL_X32 FILLER_284_1112 ();
 FILLCELL_X32 FILLER_284_1144 ();
 FILLCELL_X32 FILLER_284_1176 ();
 FILLCELL_X32 FILLER_284_1208 ();
 FILLCELL_X32 FILLER_284_1240 ();
 FILLCELL_X32 FILLER_284_1272 ();
 FILLCELL_X32 FILLER_284_1304 ();
 FILLCELL_X32 FILLER_284_1336 ();
 FILLCELL_X32 FILLER_284_1368 ();
 FILLCELL_X32 FILLER_284_1400 ();
 FILLCELL_X32 FILLER_284_1432 ();
 FILLCELL_X32 FILLER_284_1464 ();
 FILLCELL_X32 FILLER_284_1496 ();
 FILLCELL_X32 FILLER_284_1528 ();
 FILLCELL_X32 FILLER_284_1560 ();
 FILLCELL_X32 FILLER_284_1592 ();
 FILLCELL_X32 FILLER_284_1624 ();
 FILLCELL_X32 FILLER_284_1656 ();
 FILLCELL_X32 FILLER_284_1688 ();
 FILLCELL_X32 FILLER_284_1720 ();
 FILLCELL_X32 FILLER_284_1752 ();
 FILLCELL_X32 FILLER_284_1784 ();
 FILLCELL_X32 FILLER_284_1816 ();
 FILLCELL_X32 FILLER_284_1848 ();
 FILLCELL_X8 FILLER_284_1880 ();
 FILLCELL_X4 FILLER_284_1888 ();
 FILLCELL_X2 FILLER_284_1892 ();
 FILLCELL_X32 FILLER_284_1895 ();
 FILLCELL_X32 FILLER_284_1927 ();
 FILLCELL_X32 FILLER_284_1959 ();
 FILLCELL_X32 FILLER_284_1991 ();
 FILLCELL_X32 FILLER_284_2023 ();
 FILLCELL_X32 FILLER_284_2055 ();
 FILLCELL_X32 FILLER_284_2087 ();
 FILLCELL_X32 FILLER_284_2119 ();
 FILLCELL_X32 FILLER_284_2151 ();
 FILLCELL_X32 FILLER_284_2183 ();
 FILLCELL_X32 FILLER_284_2215 ();
 FILLCELL_X32 FILLER_284_2247 ();
 FILLCELL_X32 FILLER_284_2279 ();
 FILLCELL_X32 FILLER_284_2311 ();
 FILLCELL_X32 FILLER_284_2343 ();
 FILLCELL_X32 FILLER_284_2375 ();
 FILLCELL_X32 FILLER_284_2407 ();
 FILLCELL_X32 FILLER_284_2439 ();
 FILLCELL_X32 FILLER_284_2471 ();
 FILLCELL_X32 FILLER_284_2503 ();
 FILLCELL_X32 FILLER_284_2535 ();
 FILLCELL_X32 FILLER_284_2567 ();
 FILLCELL_X2 FILLER_284_2599 ();
 FILLCELL_X1 FILLER_284_2601 ();
 FILLCELL_X32 FILLER_285_1 ();
 FILLCELL_X32 FILLER_285_33 ();
 FILLCELL_X32 FILLER_285_65 ();
 FILLCELL_X32 FILLER_285_97 ();
 FILLCELL_X32 FILLER_285_129 ();
 FILLCELL_X32 FILLER_285_161 ();
 FILLCELL_X32 FILLER_285_193 ();
 FILLCELL_X32 FILLER_285_225 ();
 FILLCELL_X32 FILLER_285_257 ();
 FILLCELL_X32 FILLER_285_289 ();
 FILLCELL_X32 FILLER_285_321 ();
 FILLCELL_X32 FILLER_285_353 ();
 FILLCELL_X32 FILLER_285_385 ();
 FILLCELL_X32 FILLER_285_417 ();
 FILLCELL_X32 FILLER_285_449 ();
 FILLCELL_X32 FILLER_285_481 ();
 FILLCELL_X32 FILLER_285_513 ();
 FILLCELL_X32 FILLER_285_545 ();
 FILLCELL_X32 FILLER_285_577 ();
 FILLCELL_X32 FILLER_285_609 ();
 FILLCELL_X32 FILLER_285_641 ();
 FILLCELL_X32 FILLER_285_673 ();
 FILLCELL_X32 FILLER_285_705 ();
 FILLCELL_X32 FILLER_285_737 ();
 FILLCELL_X32 FILLER_285_769 ();
 FILLCELL_X32 FILLER_285_801 ();
 FILLCELL_X32 FILLER_285_833 ();
 FILLCELL_X32 FILLER_285_865 ();
 FILLCELL_X32 FILLER_285_897 ();
 FILLCELL_X32 FILLER_285_929 ();
 FILLCELL_X32 FILLER_285_961 ();
 FILLCELL_X32 FILLER_285_993 ();
 FILLCELL_X32 FILLER_285_1025 ();
 FILLCELL_X32 FILLER_285_1057 ();
 FILLCELL_X32 FILLER_285_1089 ();
 FILLCELL_X32 FILLER_285_1121 ();
 FILLCELL_X32 FILLER_285_1153 ();
 FILLCELL_X32 FILLER_285_1185 ();
 FILLCELL_X32 FILLER_285_1217 ();
 FILLCELL_X8 FILLER_285_1249 ();
 FILLCELL_X4 FILLER_285_1257 ();
 FILLCELL_X2 FILLER_285_1261 ();
 FILLCELL_X32 FILLER_285_1264 ();
 FILLCELL_X32 FILLER_285_1296 ();
 FILLCELL_X32 FILLER_285_1328 ();
 FILLCELL_X32 FILLER_285_1360 ();
 FILLCELL_X32 FILLER_285_1392 ();
 FILLCELL_X32 FILLER_285_1424 ();
 FILLCELL_X32 FILLER_285_1456 ();
 FILLCELL_X32 FILLER_285_1488 ();
 FILLCELL_X32 FILLER_285_1520 ();
 FILLCELL_X32 FILLER_285_1552 ();
 FILLCELL_X32 FILLER_285_1584 ();
 FILLCELL_X32 FILLER_285_1616 ();
 FILLCELL_X32 FILLER_285_1648 ();
 FILLCELL_X32 FILLER_285_1680 ();
 FILLCELL_X32 FILLER_285_1712 ();
 FILLCELL_X32 FILLER_285_1744 ();
 FILLCELL_X32 FILLER_285_1776 ();
 FILLCELL_X32 FILLER_285_1808 ();
 FILLCELL_X32 FILLER_285_1840 ();
 FILLCELL_X32 FILLER_285_1872 ();
 FILLCELL_X32 FILLER_285_1904 ();
 FILLCELL_X32 FILLER_285_1936 ();
 FILLCELL_X32 FILLER_285_1968 ();
 FILLCELL_X32 FILLER_285_2000 ();
 FILLCELL_X32 FILLER_285_2032 ();
 FILLCELL_X32 FILLER_285_2064 ();
 FILLCELL_X32 FILLER_285_2096 ();
 FILLCELL_X32 FILLER_285_2128 ();
 FILLCELL_X32 FILLER_285_2160 ();
 FILLCELL_X32 FILLER_285_2192 ();
 FILLCELL_X32 FILLER_285_2224 ();
 FILLCELL_X32 FILLER_285_2256 ();
 FILLCELL_X32 FILLER_285_2288 ();
 FILLCELL_X32 FILLER_285_2320 ();
 FILLCELL_X32 FILLER_285_2352 ();
 FILLCELL_X32 FILLER_285_2384 ();
 FILLCELL_X32 FILLER_285_2416 ();
 FILLCELL_X32 FILLER_285_2448 ();
 FILLCELL_X32 FILLER_285_2480 ();
 FILLCELL_X8 FILLER_285_2512 ();
 FILLCELL_X4 FILLER_285_2520 ();
 FILLCELL_X2 FILLER_285_2524 ();
 FILLCELL_X32 FILLER_285_2527 ();
 FILLCELL_X32 FILLER_285_2559 ();
 FILLCELL_X8 FILLER_285_2591 ();
 FILLCELL_X2 FILLER_285_2599 ();
 FILLCELL_X1 FILLER_285_2601 ();
 FILLCELL_X32 FILLER_286_1 ();
 FILLCELL_X32 FILLER_286_33 ();
 FILLCELL_X32 FILLER_286_65 ();
 FILLCELL_X32 FILLER_286_97 ();
 FILLCELL_X32 FILLER_286_129 ();
 FILLCELL_X32 FILLER_286_161 ();
 FILLCELL_X32 FILLER_286_193 ();
 FILLCELL_X32 FILLER_286_225 ();
 FILLCELL_X32 FILLER_286_257 ();
 FILLCELL_X32 FILLER_286_289 ();
 FILLCELL_X32 FILLER_286_321 ();
 FILLCELL_X32 FILLER_286_353 ();
 FILLCELL_X32 FILLER_286_385 ();
 FILLCELL_X32 FILLER_286_417 ();
 FILLCELL_X32 FILLER_286_449 ();
 FILLCELL_X32 FILLER_286_481 ();
 FILLCELL_X32 FILLER_286_513 ();
 FILLCELL_X32 FILLER_286_545 ();
 FILLCELL_X32 FILLER_286_577 ();
 FILLCELL_X16 FILLER_286_609 ();
 FILLCELL_X4 FILLER_286_625 ();
 FILLCELL_X2 FILLER_286_629 ();
 FILLCELL_X32 FILLER_286_632 ();
 FILLCELL_X32 FILLER_286_664 ();
 FILLCELL_X32 FILLER_286_696 ();
 FILLCELL_X32 FILLER_286_728 ();
 FILLCELL_X32 FILLER_286_760 ();
 FILLCELL_X32 FILLER_286_792 ();
 FILLCELL_X32 FILLER_286_824 ();
 FILLCELL_X32 FILLER_286_856 ();
 FILLCELL_X32 FILLER_286_888 ();
 FILLCELL_X32 FILLER_286_920 ();
 FILLCELL_X32 FILLER_286_952 ();
 FILLCELL_X32 FILLER_286_984 ();
 FILLCELL_X32 FILLER_286_1016 ();
 FILLCELL_X32 FILLER_286_1048 ();
 FILLCELL_X32 FILLER_286_1080 ();
 FILLCELL_X32 FILLER_286_1112 ();
 FILLCELL_X32 FILLER_286_1144 ();
 FILLCELL_X32 FILLER_286_1176 ();
 FILLCELL_X32 FILLER_286_1208 ();
 FILLCELL_X32 FILLER_286_1240 ();
 FILLCELL_X32 FILLER_286_1272 ();
 FILLCELL_X32 FILLER_286_1304 ();
 FILLCELL_X32 FILLER_286_1336 ();
 FILLCELL_X32 FILLER_286_1368 ();
 FILLCELL_X32 FILLER_286_1400 ();
 FILLCELL_X32 FILLER_286_1432 ();
 FILLCELL_X32 FILLER_286_1464 ();
 FILLCELL_X32 FILLER_286_1496 ();
 FILLCELL_X32 FILLER_286_1528 ();
 FILLCELL_X32 FILLER_286_1560 ();
 FILLCELL_X32 FILLER_286_1592 ();
 FILLCELL_X32 FILLER_286_1624 ();
 FILLCELL_X32 FILLER_286_1656 ();
 FILLCELL_X32 FILLER_286_1688 ();
 FILLCELL_X32 FILLER_286_1720 ();
 FILLCELL_X32 FILLER_286_1752 ();
 FILLCELL_X32 FILLER_286_1784 ();
 FILLCELL_X32 FILLER_286_1816 ();
 FILLCELL_X32 FILLER_286_1848 ();
 FILLCELL_X8 FILLER_286_1880 ();
 FILLCELL_X4 FILLER_286_1888 ();
 FILLCELL_X2 FILLER_286_1892 ();
 FILLCELL_X32 FILLER_286_1895 ();
 FILLCELL_X32 FILLER_286_1927 ();
 FILLCELL_X32 FILLER_286_1959 ();
 FILLCELL_X32 FILLER_286_1991 ();
 FILLCELL_X32 FILLER_286_2023 ();
 FILLCELL_X32 FILLER_286_2055 ();
 FILLCELL_X32 FILLER_286_2087 ();
 FILLCELL_X32 FILLER_286_2119 ();
 FILLCELL_X32 FILLER_286_2151 ();
 FILLCELL_X32 FILLER_286_2183 ();
 FILLCELL_X32 FILLER_286_2215 ();
 FILLCELL_X32 FILLER_286_2247 ();
 FILLCELL_X32 FILLER_286_2279 ();
 FILLCELL_X32 FILLER_286_2311 ();
 FILLCELL_X32 FILLER_286_2343 ();
 FILLCELL_X32 FILLER_286_2375 ();
 FILLCELL_X32 FILLER_286_2407 ();
 FILLCELL_X32 FILLER_286_2439 ();
 FILLCELL_X32 FILLER_286_2471 ();
 FILLCELL_X32 FILLER_286_2503 ();
 FILLCELL_X32 FILLER_286_2535 ();
 FILLCELL_X32 FILLER_286_2567 ();
 FILLCELL_X2 FILLER_286_2599 ();
 FILLCELL_X1 FILLER_286_2601 ();
 FILLCELL_X32 FILLER_287_1 ();
 FILLCELL_X32 FILLER_287_33 ();
 FILLCELL_X32 FILLER_287_65 ();
 FILLCELL_X32 FILLER_287_97 ();
 FILLCELL_X32 FILLER_287_129 ();
 FILLCELL_X32 FILLER_287_161 ();
 FILLCELL_X32 FILLER_287_193 ();
 FILLCELL_X32 FILLER_287_225 ();
 FILLCELL_X32 FILLER_287_257 ();
 FILLCELL_X32 FILLER_287_289 ();
 FILLCELL_X32 FILLER_287_321 ();
 FILLCELL_X32 FILLER_287_353 ();
 FILLCELL_X32 FILLER_287_385 ();
 FILLCELL_X32 FILLER_287_417 ();
 FILLCELL_X32 FILLER_287_449 ();
 FILLCELL_X32 FILLER_287_481 ();
 FILLCELL_X32 FILLER_287_513 ();
 FILLCELL_X32 FILLER_287_545 ();
 FILLCELL_X32 FILLER_287_577 ();
 FILLCELL_X32 FILLER_287_609 ();
 FILLCELL_X32 FILLER_287_641 ();
 FILLCELL_X32 FILLER_287_673 ();
 FILLCELL_X32 FILLER_287_705 ();
 FILLCELL_X32 FILLER_287_737 ();
 FILLCELL_X32 FILLER_287_769 ();
 FILLCELL_X32 FILLER_287_801 ();
 FILLCELL_X32 FILLER_287_833 ();
 FILLCELL_X32 FILLER_287_865 ();
 FILLCELL_X32 FILLER_287_897 ();
 FILLCELL_X32 FILLER_287_929 ();
 FILLCELL_X32 FILLER_287_961 ();
 FILLCELL_X32 FILLER_287_993 ();
 FILLCELL_X32 FILLER_287_1025 ();
 FILLCELL_X32 FILLER_287_1057 ();
 FILLCELL_X32 FILLER_287_1089 ();
 FILLCELL_X32 FILLER_287_1121 ();
 FILLCELL_X32 FILLER_287_1153 ();
 FILLCELL_X32 FILLER_287_1185 ();
 FILLCELL_X32 FILLER_287_1217 ();
 FILLCELL_X8 FILLER_287_1249 ();
 FILLCELL_X4 FILLER_287_1257 ();
 FILLCELL_X2 FILLER_287_1261 ();
 FILLCELL_X32 FILLER_287_1264 ();
 FILLCELL_X32 FILLER_287_1296 ();
 FILLCELL_X32 FILLER_287_1328 ();
 FILLCELL_X32 FILLER_287_1360 ();
 FILLCELL_X32 FILLER_287_1392 ();
 FILLCELL_X32 FILLER_287_1424 ();
 FILLCELL_X32 FILLER_287_1456 ();
 FILLCELL_X32 FILLER_287_1488 ();
 FILLCELL_X32 FILLER_287_1520 ();
 FILLCELL_X32 FILLER_287_1552 ();
 FILLCELL_X32 FILLER_287_1584 ();
 FILLCELL_X32 FILLER_287_1616 ();
 FILLCELL_X32 FILLER_287_1648 ();
 FILLCELL_X32 FILLER_287_1680 ();
 FILLCELL_X32 FILLER_287_1712 ();
 FILLCELL_X32 FILLER_287_1744 ();
 FILLCELL_X32 FILLER_287_1776 ();
 FILLCELL_X32 FILLER_287_1808 ();
 FILLCELL_X32 FILLER_287_1840 ();
 FILLCELL_X32 FILLER_287_1872 ();
 FILLCELL_X32 FILLER_287_1904 ();
 FILLCELL_X32 FILLER_287_1936 ();
 FILLCELL_X32 FILLER_287_1968 ();
 FILLCELL_X32 FILLER_287_2000 ();
 FILLCELL_X32 FILLER_287_2032 ();
 FILLCELL_X32 FILLER_287_2064 ();
 FILLCELL_X32 FILLER_287_2096 ();
 FILLCELL_X32 FILLER_287_2128 ();
 FILLCELL_X32 FILLER_287_2160 ();
 FILLCELL_X32 FILLER_287_2192 ();
 FILLCELL_X32 FILLER_287_2224 ();
 FILLCELL_X32 FILLER_287_2256 ();
 FILLCELL_X32 FILLER_287_2288 ();
 FILLCELL_X32 FILLER_287_2320 ();
 FILLCELL_X32 FILLER_287_2352 ();
 FILLCELL_X32 FILLER_287_2384 ();
 FILLCELL_X32 FILLER_287_2416 ();
 FILLCELL_X32 FILLER_287_2448 ();
 FILLCELL_X32 FILLER_287_2480 ();
 FILLCELL_X8 FILLER_287_2512 ();
 FILLCELL_X4 FILLER_287_2520 ();
 FILLCELL_X2 FILLER_287_2524 ();
 FILLCELL_X32 FILLER_287_2527 ();
 FILLCELL_X32 FILLER_287_2559 ();
 FILLCELL_X8 FILLER_287_2591 ();
 FILLCELL_X2 FILLER_287_2599 ();
 FILLCELL_X1 FILLER_287_2601 ();
 FILLCELL_X32 FILLER_288_1 ();
 FILLCELL_X32 FILLER_288_33 ();
 FILLCELL_X32 FILLER_288_65 ();
 FILLCELL_X32 FILLER_288_97 ();
 FILLCELL_X32 FILLER_288_129 ();
 FILLCELL_X32 FILLER_288_161 ();
 FILLCELL_X32 FILLER_288_193 ();
 FILLCELL_X32 FILLER_288_225 ();
 FILLCELL_X32 FILLER_288_257 ();
 FILLCELL_X32 FILLER_288_289 ();
 FILLCELL_X32 FILLER_288_321 ();
 FILLCELL_X32 FILLER_288_353 ();
 FILLCELL_X32 FILLER_288_385 ();
 FILLCELL_X32 FILLER_288_417 ();
 FILLCELL_X32 FILLER_288_449 ();
 FILLCELL_X32 FILLER_288_481 ();
 FILLCELL_X32 FILLER_288_513 ();
 FILLCELL_X32 FILLER_288_545 ();
 FILLCELL_X32 FILLER_288_577 ();
 FILLCELL_X16 FILLER_288_609 ();
 FILLCELL_X4 FILLER_288_625 ();
 FILLCELL_X2 FILLER_288_629 ();
 FILLCELL_X32 FILLER_288_632 ();
 FILLCELL_X32 FILLER_288_664 ();
 FILLCELL_X32 FILLER_288_696 ();
 FILLCELL_X32 FILLER_288_728 ();
 FILLCELL_X32 FILLER_288_760 ();
 FILLCELL_X32 FILLER_288_792 ();
 FILLCELL_X32 FILLER_288_824 ();
 FILLCELL_X32 FILLER_288_856 ();
 FILLCELL_X32 FILLER_288_888 ();
 FILLCELL_X32 FILLER_288_920 ();
 FILLCELL_X32 FILLER_288_952 ();
 FILLCELL_X32 FILLER_288_984 ();
 FILLCELL_X32 FILLER_288_1016 ();
 FILLCELL_X32 FILLER_288_1048 ();
 FILLCELL_X32 FILLER_288_1080 ();
 FILLCELL_X32 FILLER_288_1112 ();
 FILLCELL_X32 FILLER_288_1144 ();
 FILLCELL_X32 FILLER_288_1176 ();
 FILLCELL_X32 FILLER_288_1208 ();
 FILLCELL_X32 FILLER_288_1240 ();
 FILLCELL_X32 FILLER_288_1272 ();
 FILLCELL_X32 FILLER_288_1304 ();
 FILLCELL_X32 FILLER_288_1336 ();
 FILLCELL_X32 FILLER_288_1368 ();
 FILLCELL_X32 FILLER_288_1400 ();
 FILLCELL_X32 FILLER_288_1432 ();
 FILLCELL_X32 FILLER_288_1464 ();
 FILLCELL_X32 FILLER_288_1496 ();
 FILLCELL_X32 FILLER_288_1528 ();
 FILLCELL_X32 FILLER_288_1560 ();
 FILLCELL_X32 FILLER_288_1592 ();
 FILLCELL_X32 FILLER_288_1624 ();
 FILLCELL_X32 FILLER_288_1656 ();
 FILLCELL_X32 FILLER_288_1688 ();
 FILLCELL_X32 FILLER_288_1720 ();
 FILLCELL_X32 FILLER_288_1752 ();
 FILLCELL_X32 FILLER_288_1784 ();
 FILLCELL_X32 FILLER_288_1816 ();
 FILLCELL_X32 FILLER_288_1848 ();
 FILLCELL_X8 FILLER_288_1880 ();
 FILLCELL_X4 FILLER_288_1888 ();
 FILLCELL_X2 FILLER_288_1892 ();
 FILLCELL_X32 FILLER_288_1895 ();
 FILLCELL_X32 FILLER_288_1927 ();
 FILLCELL_X32 FILLER_288_1959 ();
 FILLCELL_X32 FILLER_288_1991 ();
 FILLCELL_X32 FILLER_288_2023 ();
 FILLCELL_X32 FILLER_288_2055 ();
 FILLCELL_X32 FILLER_288_2087 ();
 FILLCELL_X32 FILLER_288_2119 ();
 FILLCELL_X32 FILLER_288_2151 ();
 FILLCELL_X32 FILLER_288_2183 ();
 FILLCELL_X32 FILLER_288_2215 ();
 FILLCELL_X32 FILLER_288_2247 ();
 FILLCELL_X32 FILLER_288_2279 ();
 FILLCELL_X32 FILLER_288_2311 ();
 FILLCELL_X32 FILLER_288_2343 ();
 FILLCELL_X32 FILLER_288_2375 ();
 FILLCELL_X32 FILLER_288_2407 ();
 FILLCELL_X32 FILLER_288_2439 ();
 FILLCELL_X32 FILLER_288_2471 ();
 FILLCELL_X32 FILLER_288_2503 ();
 FILLCELL_X32 FILLER_288_2535 ();
 FILLCELL_X32 FILLER_288_2567 ();
 FILLCELL_X2 FILLER_288_2599 ();
 FILLCELL_X1 FILLER_288_2601 ();
 FILLCELL_X32 FILLER_289_1 ();
 FILLCELL_X32 FILLER_289_33 ();
 FILLCELL_X32 FILLER_289_65 ();
 FILLCELL_X32 FILLER_289_97 ();
 FILLCELL_X32 FILLER_289_129 ();
 FILLCELL_X32 FILLER_289_161 ();
 FILLCELL_X32 FILLER_289_193 ();
 FILLCELL_X32 FILLER_289_225 ();
 FILLCELL_X32 FILLER_289_257 ();
 FILLCELL_X32 FILLER_289_289 ();
 FILLCELL_X32 FILLER_289_321 ();
 FILLCELL_X32 FILLER_289_353 ();
 FILLCELL_X32 FILLER_289_385 ();
 FILLCELL_X32 FILLER_289_417 ();
 FILLCELL_X32 FILLER_289_449 ();
 FILLCELL_X32 FILLER_289_481 ();
 FILLCELL_X32 FILLER_289_513 ();
 FILLCELL_X32 FILLER_289_545 ();
 FILLCELL_X32 FILLER_289_577 ();
 FILLCELL_X32 FILLER_289_609 ();
 FILLCELL_X32 FILLER_289_641 ();
 FILLCELL_X32 FILLER_289_673 ();
 FILLCELL_X32 FILLER_289_705 ();
 FILLCELL_X32 FILLER_289_737 ();
 FILLCELL_X32 FILLER_289_769 ();
 FILLCELL_X32 FILLER_289_801 ();
 FILLCELL_X32 FILLER_289_833 ();
 FILLCELL_X32 FILLER_289_865 ();
 FILLCELL_X32 FILLER_289_897 ();
 FILLCELL_X32 FILLER_289_929 ();
 FILLCELL_X32 FILLER_289_961 ();
 FILLCELL_X32 FILLER_289_993 ();
 FILLCELL_X32 FILLER_289_1025 ();
 FILLCELL_X32 FILLER_289_1057 ();
 FILLCELL_X32 FILLER_289_1089 ();
 FILLCELL_X32 FILLER_289_1121 ();
 FILLCELL_X32 FILLER_289_1153 ();
 FILLCELL_X32 FILLER_289_1185 ();
 FILLCELL_X32 FILLER_289_1217 ();
 FILLCELL_X8 FILLER_289_1249 ();
 FILLCELL_X4 FILLER_289_1257 ();
 FILLCELL_X2 FILLER_289_1261 ();
 FILLCELL_X32 FILLER_289_1264 ();
 FILLCELL_X32 FILLER_289_1296 ();
 FILLCELL_X32 FILLER_289_1328 ();
 FILLCELL_X32 FILLER_289_1360 ();
 FILLCELL_X32 FILLER_289_1392 ();
 FILLCELL_X32 FILLER_289_1424 ();
 FILLCELL_X32 FILLER_289_1456 ();
 FILLCELL_X32 FILLER_289_1488 ();
 FILLCELL_X32 FILLER_289_1520 ();
 FILLCELL_X32 FILLER_289_1552 ();
 FILLCELL_X32 FILLER_289_1584 ();
 FILLCELL_X32 FILLER_289_1616 ();
 FILLCELL_X32 FILLER_289_1648 ();
 FILLCELL_X32 FILLER_289_1680 ();
 FILLCELL_X32 FILLER_289_1712 ();
 FILLCELL_X32 FILLER_289_1744 ();
 FILLCELL_X32 FILLER_289_1776 ();
 FILLCELL_X32 FILLER_289_1808 ();
 FILLCELL_X32 FILLER_289_1840 ();
 FILLCELL_X32 FILLER_289_1872 ();
 FILLCELL_X32 FILLER_289_1904 ();
 FILLCELL_X32 FILLER_289_1936 ();
 FILLCELL_X32 FILLER_289_1968 ();
 FILLCELL_X32 FILLER_289_2000 ();
 FILLCELL_X32 FILLER_289_2032 ();
 FILLCELL_X32 FILLER_289_2064 ();
 FILLCELL_X32 FILLER_289_2096 ();
 FILLCELL_X32 FILLER_289_2128 ();
 FILLCELL_X32 FILLER_289_2160 ();
 FILLCELL_X32 FILLER_289_2192 ();
 FILLCELL_X32 FILLER_289_2224 ();
 FILLCELL_X32 FILLER_289_2256 ();
 FILLCELL_X32 FILLER_289_2288 ();
 FILLCELL_X32 FILLER_289_2320 ();
 FILLCELL_X32 FILLER_289_2352 ();
 FILLCELL_X32 FILLER_289_2384 ();
 FILLCELL_X32 FILLER_289_2416 ();
 FILLCELL_X32 FILLER_289_2448 ();
 FILLCELL_X32 FILLER_289_2480 ();
 FILLCELL_X8 FILLER_289_2512 ();
 FILLCELL_X4 FILLER_289_2520 ();
 FILLCELL_X2 FILLER_289_2524 ();
 FILLCELL_X32 FILLER_289_2527 ();
 FILLCELL_X32 FILLER_289_2559 ();
 FILLCELL_X8 FILLER_289_2591 ();
 FILLCELL_X2 FILLER_289_2599 ();
 FILLCELL_X1 FILLER_289_2601 ();
 FILLCELL_X32 FILLER_290_1 ();
 FILLCELL_X32 FILLER_290_33 ();
 FILLCELL_X32 FILLER_290_65 ();
 FILLCELL_X32 FILLER_290_97 ();
 FILLCELL_X32 FILLER_290_129 ();
 FILLCELL_X32 FILLER_290_161 ();
 FILLCELL_X32 FILLER_290_193 ();
 FILLCELL_X32 FILLER_290_225 ();
 FILLCELL_X32 FILLER_290_257 ();
 FILLCELL_X32 FILLER_290_289 ();
 FILLCELL_X32 FILLER_290_321 ();
 FILLCELL_X32 FILLER_290_353 ();
 FILLCELL_X32 FILLER_290_385 ();
 FILLCELL_X32 FILLER_290_417 ();
 FILLCELL_X32 FILLER_290_449 ();
 FILLCELL_X32 FILLER_290_481 ();
 FILLCELL_X32 FILLER_290_513 ();
 FILLCELL_X32 FILLER_290_545 ();
 FILLCELL_X32 FILLER_290_577 ();
 FILLCELL_X16 FILLER_290_609 ();
 FILLCELL_X4 FILLER_290_625 ();
 FILLCELL_X2 FILLER_290_629 ();
 FILLCELL_X32 FILLER_290_632 ();
 FILLCELL_X32 FILLER_290_664 ();
 FILLCELL_X32 FILLER_290_696 ();
 FILLCELL_X32 FILLER_290_728 ();
 FILLCELL_X32 FILLER_290_760 ();
 FILLCELL_X32 FILLER_290_792 ();
 FILLCELL_X32 FILLER_290_824 ();
 FILLCELL_X32 FILLER_290_856 ();
 FILLCELL_X32 FILLER_290_888 ();
 FILLCELL_X32 FILLER_290_920 ();
 FILLCELL_X32 FILLER_290_952 ();
 FILLCELL_X32 FILLER_290_984 ();
 FILLCELL_X32 FILLER_290_1016 ();
 FILLCELL_X32 FILLER_290_1048 ();
 FILLCELL_X32 FILLER_290_1080 ();
 FILLCELL_X32 FILLER_290_1112 ();
 FILLCELL_X32 FILLER_290_1144 ();
 FILLCELL_X32 FILLER_290_1176 ();
 FILLCELL_X32 FILLER_290_1208 ();
 FILLCELL_X32 FILLER_290_1240 ();
 FILLCELL_X32 FILLER_290_1272 ();
 FILLCELL_X32 FILLER_290_1304 ();
 FILLCELL_X32 FILLER_290_1336 ();
 FILLCELL_X32 FILLER_290_1368 ();
 FILLCELL_X32 FILLER_290_1400 ();
 FILLCELL_X32 FILLER_290_1432 ();
 FILLCELL_X32 FILLER_290_1464 ();
 FILLCELL_X32 FILLER_290_1496 ();
 FILLCELL_X32 FILLER_290_1528 ();
 FILLCELL_X32 FILLER_290_1560 ();
 FILLCELL_X32 FILLER_290_1592 ();
 FILLCELL_X32 FILLER_290_1624 ();
 FILLCELL_X32 FILLER_290_1656 ();
 FILLCELL_X32 FILLER_290_1688 ();
 FILLCELL_X32 FILLER_290_1720 ();
 FILLCELL_X32 FILLER_290_1752 ();
 FILLCELL_X32 FILLER_290_1784 ();
 FILLCELL_X32 FILLER_290_1816 ();
 FILLCELL_X32 FILLER_290_1848 ();
 FILLCELL_X8 FILLER_290_1880 ();
 FILLCELL_X4 FILLER_290_1888 ();
 FILLCELL_X2 FILLER_290_1892 ();
 FILLCELL_X32 FILLER_290_1895 ();
 FILLCELL_X32 FILLER_290_1927 ();
 FILLCELL_X32 FILLER_290_1959 ();
 FILLCELL_X32 FILLER_290_1991 ();
 FILLCELL_X32 FILLER_290_2023 ();
 FILLCELL_X32 FILLER_290_2055 ();
 FILLCELL_X32 FILLER_290_2087 ();
 FILLCELL_X32 FILLER_290_2119 ();
 FILLCELL_X32 FILLER_290_2151 ();
 FILLCELL_X32 FILLER_290_2183 ();
 FILLCELL_X32 FILLER_290_2215 ();
 FILLCELL_X32 FILLER_290_2247 ();
 FILLCELL_X32 FILLER_290_2279 ();
 FILLCELL_X32 FILLER_290_2311 ();
 FILLCELL_X32 FILLER_290_2343 ();
 FILLCELL_X32 FILLER_290_2375 ();
 FILLCELL_X32 FILLER_290_2407 ();
 FILLCELL_X32 FILLER_290_2439 ();
 FILLCELL_X32 FILLER_290_2471 ();
 FILLCELL_X32 FILLER_290_2503 ();
 FILLCELL_X32 FILLER_290_2535 ();
 FILLCELL_X32 FILLER_290_2567 ();
 FILLCELL_X2 FILLER_290_2599 ();
 FILLCELL_X1 FILLER_290_2601 ();
 FILLCELL_X32 FILLER_291_1 ();
 FILLCELL_X32 FILLER_291_33 ();
 FILLCELL_X32 FILLER_291_65 ();
 FILLCELL_X32 FILLER_291_97 ();
 FILLCELL_X32 FILLER_291_129 ();
 FILLCELL_X32 FILLER_291_161 ();
 FILLCELL_X32 FILLER_291_193 ();
 FILLCELL_X32 FILLER_291_225 ();
 FILLCELL_X32 FILLER_291_257 ();
 FILLCELL_X32 FILLER_291_289 ();
 FILLCELL_X32 FILLER_291_321 ();
 FILLCELL_X32 FILLER_291_353 ();
 FILLCELL_X32 FILLER_291_385 ();
 FILLCELL_X32 FILLER_291_417 ();
 FILLCELL_X32 FILLER_291_449 ();
 FILLCELL_X32 FILLER_291_481 ();
 FILLCELL_X32 FILLER_291_513 ();
 FILLCELL_X32 FILLER_291_545 ();
 FILLCELL_X32 FILLER_291_577 ();
 FILLCELL_X32 FILLER_291_609 ();
 FILLCELL_X32 FILLER_291_641 ();
 FILLCELL_X32 FILLER_291_673 ();
 FILLCELL_X32 FILLER_291_705 ();
 FILLCELL_X32 FILLER_291_737 ();
 FILLCELL_X32 FILLER_291_769 ();
 FILLCELL_X32 FILLER_291_801 ();
 FILLCELL_X32 FILLER_291_833 ();
 FILLCELL_X32 FILLER_291_865 ();
 FILLCELL_X32 FILLER_291_897 ();
 FILLCELL_X32 FILLER_291_929 ();
 FILLCELL_X32 FILLER_291_961 ();
 FILLCELL_X32 FILLER_291_993 ();
 FILLCELL_X32 FILLER_291_1025 ();
 FILLCELL_X32 FILLER_291_1057 ();
 FILLCELL_X32 FILLER_291_1089 ();
 FILLCELL_X32 FILLER_291_1121 ();
 FILLCELL_X32 FILLER_291_1153 ();
 FILLCELL_X32 FILLER_291_1185 ();
 FILLCELL_X32 FILLER_291_1217 ();
 FILLCELL_X8 FILLER_291_1249 ();
 FILLCELL_X4 FILLER_291_1257 ();
 FILLCELL_X2 FILLER_291_1261 ();
 FILLCELL_X32 FILLER_291_1264 ();
 FILLCELL_X32 FILLER_291_1296 ();
 FILLCELL_X32 FILLER_291_1328 ();
 FILLCELL_X32 FILLER_291_1360 ();
 FILLCELL_X32 FILLER_291_1392 ();
 FILLCELL_X32 FILLER_291_1424 ();
 FILLCELL_X32 FILLER_291_1456 ();
 FILLCELL_X32 FILLER_291_1488 ();
 FILLCELL_X32 FILLER_291_1520 ();
 FILLCELL_X32 FILLER_291_1552 ();
 FILLCELL_X32 FILLER_291_1584 ();
 FILLCELL_X32 FILLER_291_1616 ();
 FILLCELL_X32 FILLER_291_1648 ();
 FILLCELL_X32 FILLER_291_1680 ();
 FILLCELL_X32 FILLER_291_1712 ();
 FILLCELL_X32 FILLER_291_1744 ();
 FILLCELL_X32 FILLER_291_1776 ();
 FILLCELL_X32 FILLER_291_1808 ();
 FILLCELL_X32 FILLER_291_1840 ();
 FILLCELL_X32 FILLER_291_1872 ();
 FILLCELL_X32 FILLER_291_1904 ();
 FILLCELL_X32 FILLER_291_1936 ();
 FILLCELL_X32 FILLER_291_1968 ();
 FILLCELL_X32 FILLER_291_2000 ();
 FILLCELL_X32 FILLER_291_2032 ();
 FILLCELL_X32 FILLER_291_2064 ();
 FILLCELL_X32 FILLER_291_2096 ();
 FILLCELL_X32 FILLER_291_2128 ();
 FILLCELL_X32 FILLER_291_2160 ();
 FILLCELL_X32 FILLER_291_2192 ();
 FILLCELL_X32 FILLER_291_2224 ();
 FILLCELL_X32 FILLER_291_2256 ();
 FILLCELL_X32 FILLER_291_2288 ();
 FILLCELL_X32 FILLER_291_2320 ();
 FILLCELL_X32 FILLER_291_2352 ();
 FILLCELL_X32 FILLER_291_2384 ();
 FILLCELL_X32 FILLER_291_2416 ();
 FILLCELL_X32 FILLER_291_2448 ();
 FILLCELL_X32 FILLER_291_2480 ();
 FILLCELL_X8 FILLER_291_2512 ();
 FILLCELL_X4 FILLER_291_2520 ();
 FILLCELL_X2 FILLER_291_2524 ();
 FILLCELL_X32 FILLER_291_2527 ();
 FILLCELL_X32 FILLER_291_2559 ();
 FILLCELL_X8 FILLER_291_2591 ();
 FILLCELL_X2 FILLER_291_2599 ();
 FILLCELL_X1 FILLER_291_2601 ();
 FILLCELL_X32 FILLER_292_1 ();
 FILLCELL_X32 FILLER_292_33 ();
 FILLCELL_X32 FILLER_292_65 ();
 FILLCELL_X32 FILLER_292_97 ();
 FILLCELL_X32 FILLER_292_129 ();
 FILLCELL_X32 FILLER_292_161 ();
 FILLCELL_X32 FILLER_292_193 ();
 FILLCELL_X32 FILLER_292_225 ();
 FILLCELL_X32 FILLER_292_257 ();
 FILLCELL_X32 FILLER_292_289 ();
 FILLCELL_X32 FILLER_292_321 ();
 FILLCELL_X32 FILLER_292_353 ();
 FILLCELL_X32 FILLER_292_385 ();
 FILLCELL_X32 FILLER_292_417 ();
 FILLCELL_X32 FILLER_292_449 ();
 FILLCELL_X32 FILLER_292_481 ();
 FILLCELL_X32 FILLER_292_513 ();
 FILLCELL_X32 FILLER_292_545 ();
 FILLCELL_X32 FILLER_292_577 ();
 FILLCELL_X16 FILLER_292_609 ();
 FILLCELL_X4 FILLER_292_625 ();
 FILLCELL_X2 FILLER_292_629 ();
 FILLCELL_X32 FILLER_292_632 ();
 FILLCELL_X32 FILLER_292_664 ();
 FILLCELL_X32 FILLER_292_696 ();
 FILLCELL_X32 FILLER_292_728 ();
 FILLCELL_X32 FILLER_292_760 ();
 FILLCELL_X32 FILLER_292_792 ();
 FILLCELL_X32 FILLER_292_824 ();
 FILLCELL_X32 FILLER_292_856 ();
 FILLCELL_X32 FILLER_292_888 ();
 FILLCELL_X32 FILLER_292_920 ();
 FILLCELL_X32 FILLER_292_952 ();
 FILLCELL_X32 FILLER_292_984 ();
 FILLCELL_X32 FILLER_292_1016 ();
 FILLCELL_X32 FILLER_292_1048 ();
 FILLCELL_X32 FILLER_292_1080 ();
 FILLCELL_X32 FILLER_292_1112 ();
 FILLCELL_X32 FILLER_292_1144 ();
 FILLCELL_X32 FILLER_292_1176 ();
 FILLCELL_X32 FILLER_292_1208 ();
 FILLCELL_X32 FILLER_292_1240 ();
 FILLCELL_X32 FILLER_292_1272 ();
 FILLCELL_X32 FILLER_292_1304 ();
 FILLCELL_X32 FILLER_292_1336 ();
 FILLCELL_X32 FILLER_292_1368 ();
 FILLCELL_X32 FILLER_292_1400 ();
 FILLCELL_X32 FILLER_292_1432 ();
 FILLCELL_X32 FILLER_292_1464 ();
 FILLCELL_X32 FILLER_292_1496 ();
 FILLCELL_X32 FILLER_292_1528 ();
 FILLCELL_X32 FILLER_292_1560 ();
 FILLCELL_X32 FILLER_292_1592 ();
 FILLCELL_X32 FILLER_292_1624 ();
 FILLCELL_X32 FILLER_292_1656 ();
 FILLCELL_X32 FILLER_292_1688 ();
 FILLCELL_X32 FILLER_292_1720 ();
 FILLCELL_X32 FILLER_292_1752 ();
 FILLCELL_X32 FILLER_292_1784 ();
 FILLCELL_X32 FILLER_292_1816 ();
 FILLCELL_X32 FILLER_292_1848 ();
 FILLCELL_X8 FILLER_292_1880 ();
 FILLCELL_X4 FILLER_292_1888 ();
 FILLCELL_X2 FILLER_292_1892 ();
 FILLCELL_X32 FILLER_292_1895 ();
 FILLCELL_X32 FILLER_292_1927 ();
 FILLCELL_X32 FILLER_292_1959 ();
 FILLCELL_X32 FILLER_292_1991 ();
 FILLCELL_X32 FILLER_292_2023 ();
 FILLCELL_X32 FILLER_292_2055 ();
 FILLCELL_X32 FILLER_292_2087 ();
 FILLCELL_X32 FILLER_292_2119 ();
 FILLCELL_X32 FILLER_292_2151 ();
 FILLCELL_X32 FILLER_292_2183 ();
 FILLCELL_X32 FILLER_292_2215 ();
 FILLCELL_X32 FILLER_292_2247 ();
 FILLCELL_X32 FILLER_292_2279 ();
 FILLCELL_X32 FILLER_292_2311 ();
 FILLCELL_X32 FILLER_292_2343 ();
 FILLCELL_X32 FILLER_292_2375 ();
 FILLCELL_X32 FILLER_292_2407 ();
 FILLCELL_X32 FILLER_292_2439 ();
 FILLCELL_X32 FILLER_292_2471 ();
 FILLCELL_X32 FILLER_292_2503 ();
 FILLCELL_X32 FILLER_292_2535 ();
 FILLCELL_X32 FILLER_292_2567 ();
 FILLCELL_X2 FILLER_292_2599 ();
 FILLCELL_X1 FILLER_292_2601 ();
 FILLCELL_X32 FILLER_293_1 ();
 FILLCELL_X32 FILLER_293_33 ();
 FILLCELL_X32 FILLER_293_65 ();
 FILLCELL_X32 FILLER_293_97 ();
 FILLCELL_X32 FILLER_293_129 ();
 FILLCELL_X32 FILLER_293_161 ();
 FILLCELL_X32 FILLER_293_193 ();
 FILLCELL_X32 FILLER_293_225 ();
 FILLCELL_X32 FILLER_293_257 ();
 FILLCELL_X32 FILLER_293_289 ();
 FILLCELL_X32 FILLER_293_321 ();
 FILLCELL_X32 FILLER_293_353 ();
 FILLCELL_X32 FILLER_293_385 ();
 FILLCELL_X32 FILLER_293_417 ();
 FILLCELL_X32 FILLER_293_449 ();
 FILLCELL_X32 FILLER_293_481 ();
 FILLCELL_X32 FILLER_293_513 ();
 FILLCELL_X32 FILLER_293_545 ();
 FILLCELL_X32 FILLER_293_577 ();
 FILLCELL_X32 FILLER_293_609 ();
 FILLCELL_X32 FILLER_293_641 ();
 FILLCELL_X32 FILLER_293_673 ();
 FILLCELL_X32 FILLER_293_705 ();
 FILLCELL_X32 FILLER_293_737 ();
 FILLCELL_X32 FILLER_293_769 ();
 FILLCELL_X32 FILLER_293_801 ();
 FILLCELL_X32 FILLER_293_833 ();
 FILLCELL_X32 FILLER_293_865 ();
 FILLCELL_X32 FILLER_293_897 ();
 FILLCELL_X32 FILLER_293_929 ();
 FILLCELL_X32 FILLER_293_961 ();
 FILLCELL_X32 FILLER_293_993 ();
 FILLCELL_X32 FILLER_293_1025 ();
 FILLCELL_X32 FILLER_293_1057 ();
 FILLCELL_X32 FILLER_293_1089 ();
 FILLCELL_X32 FILLER_293_1121 ();
 FILLCELL_X32 FILLER_293_1153 ();
 FILLCELL_X32 FILLER_293_1185 ();
 FILLCELL_X32 FILLER_293_1217 ();
 FILLCELL_X8 FILLER_293_1249 ();
 FILLCELL_X4 FILLER_293_1257 ();
 FILLCELL_X2 FILLER_293_1261 ();
 FILLCELL_X32 FILLER_293_1264 ();
 FILLCELL_X32 FILLER_293_1296 ();
 FILLCELL_X32 FILLER_293_1328 ();
 FILLCELL_X32 FILLER_293_1360 ();
 FILLCELL_X32 FILLER_293_1392 ();
 FILLCELL_X32 FILLER_293_1424 ();
 FILLCELL_X32 FILLER_293_1456 ();
 FILLCELL_X32 FILLER_293_1488 ();
 FILLCELL_X32 FILLER_293_1520 ();
 FILLCELL_X32 FILLER_293_1552 ();
 FILLCELL_X32 FILLER_293_1584 ();
 FILLCELL_X32 FILLER_293_1616 ();
 FILLCELL_X32 FILLER_293_1648 ();
 FILLCELL_X32 FILLER_293_1680 ();
 FILLCELL_X32 FILLER_293_1712 ();
 FILLCELL_X32 FILLER_293_1744 ();
 FILLCELL_X32 FILLER_293_1776 ();
 FILLCELL_X32 FILLER_293_1808 ();
 FILLCELL_X32 FILLER_293_1840 ();
 FILLCELL_X32 FILLER_293_1872 ();
 FILLCELL_X32 FILLER_293_1904 ();
 FILLCELL_X32 FILLER_293_1936 ();
 FILLCELL_X32 FILLER_293_1968 ();
 FILLCELL_X32 FILLER_293_2000 ();
 FILLCELL_X32 FILLER_293_2032 ();
 FILLCELL_X32 FILLER_293_2064 ();
 FILLCELL_X32 FILLER_293_2096 ();
 FILLCELL_X32 FILLER_293_2128 ();
 FILLCELL_X32 FILLER_293_2160 ();
 FILLCELL_X32 FILLER_293_2192 ();
 FILLCELL_X32 FILLER_293_2224 ();
 FILLCELL_X32 FILLER_293_2256 ();
 FILLCELL_X32 FILLER_293_2288 ();
 FILLCELL_X32 FILLER_293_2320 ();
 FILLCELL_X32 FILLER_293_2352 ();
 FILLCELL_X32 FILLER_293_2384 ();
 FILLCELL_X32 FILLER_293_2416 ();
 FILLCELL_X32 FILLER_293_2448 ();
 FILLCELL_X32 FILLER_293_2480 ();
 FILLCELL_X8 FILLER_293_2512 ();
 FILLCELL_X4 FILLER_293_2520 ();
 FILLCELL_X2 FILLER_293_2524 ();
 FILLCELL_X32 FILLER_293_2527 ();
 FILLCELL_X32 FILLER_293_2559 ();
 FILLCELL_X8 FILLER_293_2591 ();
 FILLCELL_X2 FILLER_293_2599 ();
 FILLCELL_X1 FILLER_293_2601 ();
 FILLCELL_X32 FILLER_294_1 ();
 FILLCELL_X32 FILLER_294_33 ();
 FILLCELL_X32 FILLER_294_65 ();
 FILLCELL_X32 FILLER_294_97 ();
 FILLCELL_X32 FILLER_294_129 ();
 FILLCELL_X32 FILLER_294_161 ();
 FILLCELL_X32 FILLER_294_193 ();
 FILLCELL_X32 FILLER_294_225 ();
 FILLCELL_X32 FILLER_294_257 ();
 FILLCELL_X32 FILLER_294_289 ();
 FILLCELL_X32 FILLER_294_321 ();
 FILLCELL_X32 FILLER_294_353 ();
 FILLCELL_X32 FILLER_294_385 ();
 FILLCELL_X32 FILLER_294_417 ();
 FILLCELL_X32 FILLER_294_449 ();
 FILLCELL_X32 FILLER_294_481 ();
 FILLCELL_X32 FILLER_294_513 ();
 FILLCELL_X32 FILLER_294_545 ();
 FILLCELL_X32 FILLER_294_577 ();
 FILLCELL_X16 FILLER_294_609 ();
 FILLCELL_X4 FILLER_294_625 ();
 FILLCELL_X2 FILLER_294_629 ();
 FILLCELL_X32 FILLER_294_632 ();
 FILLCELL_X32 FILLER_294_664 ();
 FILLCELL_X32 FILLER_294_696 ();
 FILLCELL_X32 FILLER_294_728 ();
 FILLCELL_X32 FILLER_294_760 ();
 FILLCELL_X32 FILLER_294_792 ();
 FILLCELL_X32 FILLER_294_824 ();
 FILLCELL_X32 FILLER_294_856 ();
 FILLCELL_X32 FILLER_294_888 ();
 FILLCELL_X32 FILLER_294_920 ();
 FILLCELL_X32 FILLER_294_952 ();
 FILLCELL_X32 FILLER_294_984 ();
 FILLCELL_X32 FILLER_294_1016 ();
 FILLCELL_X32 FILLER_294_1048 ();
 FILLCELL_X32 FILLER_294_1080 ();
 FILLCELL_X32 FILLER_294_1112 ();
 FILLCELL_X32 FILLER_294_1144 ();
 FILLCELL_X32 FILLER_294_1176 ();
 FILLCELL_X32 FILLER_294_1208 ();
 FILLCELL_X32 FILLER_294_1240 ();
 FILLCELL_X32 FILLER_294_1272 ();
 FILLCELL_X32 FILLER_294_1304 ();
 FILLCELL_X32 FILLER_294_1336 ();
 FILLCELL_X32 FILLER_294_1368 ();
 FILLCELL_X32 FILLER_294_1400 ();
 FILLCELL_X32 FILLER_294_1432 ();
 FILLCELL_X32 FILLER_294_1464 ();
 FILLCELL_X32 FILLER_294_1496 ();
 FILLCELL_X32 FILLER_294_1528 ();
 FILLCELL_X32 FILLER_294_1560 ();
 FILLCELL_X32 FILLER_294_1592 ();
 FILLCELL_X32 FILLER_294_1624 ();
 FILLCELL_X32 FILLER_294_1656 ();
 FILLCELL_X32 FILLER_294_1688 ();
 FILLCELL_X32 FILLER_294_1720 ();
 FILLCELL_X32 FILLER_294_1752 ();
 FILLCELL_X32 FILLER_294_1784 ();
 FILLCELL_X32 FILLER_294_1816 ();
 FILLCELL_X32 FILLER_294_1848 ();
 FILLCELL_X8 FILLER_294_1880 ();
 FILLCELL_X4 FILLER_294_1888 ();
 FILLCELL_X2 FILLER_294_1892 ();
 FILLCELL_X32 FILLER_294_1895 ();
 FILLCELL_X32 FILLER_294_1927 ();
 FILLCELL_X32 FILLER_294_1959 ();
 FILLCELL_X32 FILLER_294_1991 ();
 FILLCELL_X32 FILLER_294_2023 ();
 FILLCELL_X32 FILLER_294_2055 ();
 FILLCELL_X32 FILLER_294_2087 ();
 FILLCELL_X32 FILLER_294_2119 ();
 FILLCELL_X32 FILLER_294_2151 ();
 FILLCELL_X32 FILLER_294_2183 ();
 FILLCELL_X32 FILLER_294_2215 ();
 FILLCELL_X32 FILLER_294_2247 ();
 FILLCELL_X32 FILLER_294_2279 ();
 FILLCELL_X32 FILLER_294_2311 ();
 FILLCELL_X32 FILLER_294_2343 ();
 FILLCELL_X32 FILLER_294_2375 ();
 FILLCELL_X32 FILLER_294_2407 ();
 FILLCELL_X32 FILLER_294_2439 ();
 FILLCELL_X32 FILLER_294_2471 ();
 FILLCELL_X32 FILLER_294_2503 ();
 FILLCELL_X32 FILLER_294_2535 ();
 FILLCELL_X32 FILLER_294_2567 ();
 FILLCELL_X2 FILLER_294_2599 ();
 FILLCELL_X1 FILLER_294_2601 ();
 FILLCELL_X32 FILLER_295_1 ();
 FILLCELL_X32 FILLER_295_33 ();
 FILLCELL_X32 FILLER_295_65 ();
 FILLCELL_X32 FILLER_295_97 ();
 FILLCELL_X32 FILLER_295_129 ();
 FILLCELL_X32 FILLER_295_161 ();
 FILLCELL_X32 FILLER_295_193 ();
 FILLCELL_X32 FILLER_295_225 ();
 FILLCELL_X32 FILLER_295_257 ();
 FILLCELL_X32 FILLER_295_289 ();
 FILLCELL_X32 FILLER_295_321 ();
 FILLCELL_X32 FILLER_295_353 ();
 FILLCELL_X32 FILLER_295_385 ();
 FILLCELL_X32 FILLER_295_417 ();
 FILLCELL_X32 FILLER_295_449 ();
 FILLCELL_X32 FILLER_295_481 ();
 FILLCELL_X32 FILLER_295_513 ();
 FILLCELL_X32 FILLER_295_545 ();
 FILLCELL_X32 FILLER_295_577 ();
 FILLCELL_X32 FILLER_295_609 ();
 FILLCELL_X32 FILLER_295_641 ();
 FILLCELL_X32 FILLER_295_673 ();
 FILLCELL_X32 FILLER_295_705 ();
 FILLCELL_X32 FILLER_295_737 ();
 FILLCELL_X32 FILLER_295_769 ();
 FILLCELL_X32 FILLER_295_801 ();
 FILLCELL_X32 FILLER_295_833 ();
 FILLCELL_X32 FILLER_295_865 ();
 FILLCELL_X32 FILLER_295_897 ();
 FILLCELL_X32 FILLER_295_929 ();
 FILLCELL_X32 FILLER_295_961 ();
 FILLCELL_X32 FILLER_295_993 ();
 FILLCELL_X32 FILLER_295_1025 ();
 FILLCELL_X32 FILLER_295_1057 ();
 FILLCELL_X32 FILLER_295_1089 ();
 FILLCELL_X32 FILLER_295_1121 ();
 FILLCELL_X32 FILLER_295_1153 ();
 FILLCELL_X32 FILLER_295_1185 ();
 FILLCELL_X32 FILLER_295_1217 ();
 FILLCELL_X8 FILLER_295_1249 ();
 FILLCELL_X4 FILLER_295_1257 ();
 FILLCELL_X2 FILLER_295_1261 ();
 FILLCELL_X32 FILLER_295_1264 ();
 FILLCELL_X32 FILLER_295_1296 ();
 FILLCELL_X32 FILLER_295_1328 ();
 FILLCELL_X32 FILLER_295_1360 ();
 FILLCELL_X32 FILLER_295_1392 ();
 FILLCELL_X32 FILLER_295_1424 ();
 FILLCELL_X32 FILLER_295_1456 ();
 FILLCELL_X32 FILLER_295_1488 ();
 FILLCELL_X32 FILLER_295_1520 ();
 FILLCELL_X32 FILLER_295_1552 ();
 FILLCELL_X32 FILLER_295_1584 ();
 FILLCELL_X32 FILLER_295_1616 ();
 FILLCELL_X32 FILLER_295_1648 ();
 FILLCELL_X32 FILLER_295_1680 ();
 FILLCELL_X32 FILLER_295_1712 ();
 FILLCELL_X32 FILLER_295_1744 ();
 FILLCELL_X32 FILLER_295_1776 ();
 FILLCELL_X32 FILLER_295_1808 ();
 FILLCELL_X32 FILLER_295_1840 ();
 FILLCELL_X32 FILLER_295_1872 ();
 FILLCELL_X32 FILLER_295_1904 ();
 FILLCELL_X32 FILLER_295_1936 ();
 FILLCELL_X32 FILLER_295_1968 ();
 FILLCELL_X32 FILLER_295_2000 ();
 FILLCELL_X32 FILLER_295_2032 ();
 FILLCELL_X32 FILLER_295_2064 ();
 FILLCELL_X32 FILLER_295_2096 ();
 FILLCELL_X32 FILLER_295_2128 ();
 FILLCELL_X32 FILLER_295_2160 ();
 FILLCELL_X32 FILLER_295_2192 ();
 FILLCELL_X32 FILLER_295_2224 ();
 FILLCELL_X32 FILLER_295_2256 ();
 FILLCELL_X32 FILLER_295_2288 ();
 FILLCELL_X32 FILLER_295_2320 ();
 FILLCELL_X32 FILLER_295_2352 ();
 FILLCELL_X32 FILLER_295_2384 ();
 FILLCELL_X32 FILLER_295_2416 ();
 FILLCELL_X32 FILLER_295_2448 ();
 FILLCELL_X32 FILLER_295_2480 ();
 FILLCELL_X8 FILLER_295_2512 ();
 FILLCELL_X4 FILLER_295_2520 ();
 FILLCELL_X2 FILLER_295_2524 ();
 FILLCELL_X32 FILLER_295_2527 ();
 FILLCELL_X32 FILLER_295_2559 ();
 FILLCELL_X8 FILLER_295_2591 ();
 FILLCELL_X2 FILLER_295_2599 ();
 FILLCELL_X1 FILLER_295_2601 ();
 FILLCELL_X32 FILLER_296_1 ();
 FILLCELL_X32 FILLER_296_33 ();
 FILLCELL_X32 FILLER_296_65 ();
 FILLCELL_X32 FILLER_296_97 ();
 FILLCELL_X32 FILLER_296_129 ();
 FILLCELL_X32 FILLER_296_161 ();
 FILLCELL_X32 FILLER_296_193 ();
 FILLCELL_X32 FILLER_296_225 ();
 FILLCELL_X32 FILLER_296_257 ();
 FILLCELL_X32 FILLER_296_289 ();
 FILLCELL_X32 FILLER_296_321 ();
 FILLCELL_X32 FILLER_296_353 ();
 FILLCELL_X32 FILLER_296_385 ();
 FILLCELL_X32 FILLER_296_417 ();
 FILLCELL_X32 FILLER_296_449 ();
 FILLCELL_X32 FILLER_296_481 ();
 FILLCELL_X32 FILLER_296_513 ();
 FILLCELL_X32 FILLER_296_545 ();
 FILLCELL_X32 FILLER_296_577 ();
 FILLCELL_X16 FILLER_296_609 ();
 FILLCELL_X4 FILLER_296_625 ();
 FILLCELL_X2 FILLER_296_629 ();
 FILLCELL_X32 FILLER_296_632 ();
 FILLCELL_X32 FILLER_296_664 ();
 FILLCELL_X32 FILLER_296_696 ();
 FILLCELL_X32 FILLER_296_728 ();
 FILLCELL_X32 FILLER_296_760 ();
 FILLCELL_X32 FILLER_296_792 ();
 FILLCELL_X32 FILLER_296_824 ();
 FILLCELL_X32 FILLER_296_856 ();
 FILLCELL_X32 FILLER_296_888 ();
 FILLCELL_X32 FILLER_296_920 ();
 FILLCELL_X32 FILLER_296_952 ();
 FILLCELL_X32 FILLER_296_984 ();
 FILLCELL_X32 FILLER_296_1016 ();
 FILLCELL_X32 FILLER_296_1048 ();
 FILLCELL_X32 FILLER_296_1080 ();
 FILLCELL_X32 FILLER_296_1112 ();
 FILLCELL_X32 FILLER_296_1144 ();
 FILLCELL_X32 FILLER_296_1176 ();
 FILLCELL_X32 FILLER_296_1208 ();
 FILLCELL_X32 FILLER_296_1240 ();
 FILLCELL_X32 FILLER_296_1272 ();
 FILLCELL_X32 FILLER_296_1304 ();
 FILLCELL_X32 FILLER_296_1336 ();
 FILLCELL_X32 FILLER_296_1368 ();
 FILLCELL_X32 FILLER_296_1400 ();
 FILLCELL_X32 FILLER_296_1432 ();
 FILLCELL_X32 FILLER_296_1464 ();
 FILLCELL_X32 FILLER_296_1496 ();
 FILLCELL_X32 FILLER_296_1528 ();
 FILLCELL_X32 FILLER_296_1560 ();
 FILLCELL_X32 FILLER_296_1592 ();
 FILLCELL_X32 FILLER_296_1624 ();
 FILLCELL_X32 FILLER_296_1656 ();
 FILLCELL_X32 FILLER_296_1688 ();
 FILLCELL_X32 FILLER_296_1720 ();
 FILLCELL_X32 FILLER_296_1752 ();
 FILLCELL_X32 FILLER_296_1784 ();
 FILLCELL_X32 FILLER_296_1816 ();
 FILLCELL_X32 FILLER_296_1848 ();
 FILLCELL_X8 FILLER_296_1880 ();
 FILLCELL_X4 FILLER_296_1888 ();
 FILLCELL_X2 FILLER_296_1892 ();
 FILLCELL_X32 FILLER_296_1895 ();
 FILLCELL_X32 FILLER_296_1927 ();
 FILLCELL_X32 FILLER_296_1959 ();
 FILLCELL_X32 FILLER_296_1991 ();
 FILLCELL_X32 FILLER_296_2023 ();
 FILLCELL_X32 FILLER_296_2055 ();
 FILLCELL_X32 FILLER_296_2087 ();
 FILLCELL_X32 FILLER_296_2119 ();
 FILLCELL_X32 FILLER_296_2151 ();
 FILLCELL_X32 FILLER_296_2183 ();
 FILLCELL_X32 FILLER_296_2215 ();
 FILLCELL_X32 FILLER_296_2247 ();
 FILLCELL_X32 FILLER_296_2279 ();
 FILLCELL_X32 FILLER_296_2311 ();
 FILLCELL_X32 FILLER_296_2343 ();
 FILLCELL_X32 FILLER_296_2375 ();
 FILLCELL_X32 FILLER_296_2407 ();
 FILLCELL_X32 FILLER_296_2439 ();
 FILLCELL_X32 FILLER_296_2471 ();
 FILLCELL_X32 FILLER_296_2503 ();
 FILLCELL_X32 FILLER_296_2535 ();
 FILLCELL_X32 FILLER_296_2567 ();
 FILLCELL_X2 FILLER_296_2599 ();
 FILLCELL_X1 FILLER_296_2601 ();
 FILLCELL_X32 FILLER_297_1 ();
 FILLCELL_X32 FILLER_297_33 ();
 FILLCELL_X32 FILLER_297_65 ();
 FILLCELL_X32 FILLER_297_97 ();
 FILLCELL_X32 FILLER_297_129 ();
 FILLCELL_X32 FILLER_297_161 ();
 FILLCELL_X32 FILLER_297_193 ();
 FILLCELL_X32 FILLER_297_225 ();
 FILLCELL_X32 FILLER_297_257 ();
 FILLCELL_X32 FILLER_297_289 ();
 FILLCELL_X32 FILLER_297_321 ();
 FILLCELL_X32 FILLER_297_353 ();
 FILLCELL_X32 FILLER_297_385 ();
 FILLCELL_X32 FILLER_297_417 ();
 FILLCELL_X32 FILLER_297_449 ();
 FILLCELL_X32 FILLER_297_481 ();
 FILLCELL_X32 FILLER_297_513 ();
 FILLCELL_X32 FILLER_297_545 ();
 FILLCELL_X32 FILLER_297_577 ();
 FILLCELL_X32 FILLER_297_609 ();
 FILLCELL_X32 FILLER_297_641 ();
 FILLCELL_X32 FILLER_297_673 ();
 FILLCELL_X32 FILLER_297_705 ();
 FILLCELL_X32 FILLER_297_737 ();
 FILLCELL_X32 FILLER_297_769 ();
 FILLCELL_X32 FILLER_297_801 ();
 FILLCELL_X32 FILLER_297_833 ();
 FILLCELL_X32 FILLER_297_865 ();
 FILLCELL_X32 FILLER_297_897 ();
 FILLCELL_X32 FILLER_297_929 ();
 FILLCELL_X32 FILLER_297_961 ();
 FILLCELL_X32 FILLER_297_993 ();
 FILLCELL_X32 FILLER_297_1025 ();
 FILLCELL_X32 FILLER_297_1057 ();
 FILLCELL_X32 FILLER_297_1089 ();
 FILLCELL_X32 FILLER_297_1121 ();
 FILLCELL_X32 FILLER_297_1153 ();
 FILLCELL_X32 FILLER_297_1185 ();
 FILLCELL_X32 FILLER_297_1217 ();
 FILLCELL_X8 FILLER_297_1249 ();
 FILLCELL_X4 FILLER_297_1257 ();
 FILLCELL_X2 FILLER_297_1261 ();
 FILLCELL_X32 FILLER_297_1264 ();
 FILLCELL_X32 FILLER_297_1296 ();
 FILLCELL_X32 FILLER_297_1328 ();
 FILLCELL_X32 FILLER_297_1360 ();
 FILLCELL_X32 FILLER_297_1392 ();
 FILLCELL_X32 FILLER_297_1424 ();
 FILLCELL_X32 FILLER_297_1456 ();
 FILLCELL_X32 FILLER_297_1488 ();
 FILLCELL_X32 FILLER_297_1520 ();
 FILLCELL_X32 FILLER_297_1552 ();
 FILLCELL_X32 FILLER_297_1584 ();
 FILLCELL_X32 FILLER_297_1616 ();
 FILLCELL_X32 FILLER_297_1648 ();
 FILLCELL_X32 FILLER_297_1680 ();
 FILLCELL_X32 FILLER_297_1712 ();
 FILLCELL_X32 FILLER_297_1744 ();
 FILLCELL_X32 FILLER_297_1776 ();
 FILLCELL_X32 FILLER_297_1808 ();
 FILLCELL_X32 FILLER_297_1840 ();
 FILLCELL_X32 FILLER_297_1872 ();
 FILLCELL_X32 FILLER_297_1904 ();
 FILLCELL_X32 FILLER_297_1936 ();
 FILLCELL_X32 FILLER_297_1968 ();
 FILLCELL_X32 FILLER_297_2000 ();
 FILLCELL_X32 FILLER_297_2032 ();
 FILLCELL_X32 FILLER_297_2064 ();
 FILLCELL_X32 FILLER_297_2096 ();
 FILLCELL_X32 FILLER_297_2128 ();
 FILLCELL_X32 FILLER_297_2160 ();
 FILLCELL_X32 FILLER_297_2192 ();
 FILLCELL_X32 FILLER_297_2224 ();
 FILLCELL_X32 FILLER_297_2256 ();
 FILLCELL_X32 FILLER_297_2288 ();
 FILLCELL_X32 FILLER_297_2320 ();
 FILLCELL_X32 FILLER_297_2352 ();
 FILLCELL_X32 FILLER_297_2384 ();
 FILLCELL_X32 FILLER_297_2416 ();
 FILLCELL_X32 FILLER_297_2448 ();
 FILLCELL_X32 FILLER_297_2480 ();
 FILLCELL_X8 FILLER_297_2512 ();
 FILLCELL_X4 FILLER_297_2520 ();
 FILLCELL_X2 FILLER_297_2524 ();
 FILLCELL_X32 FILLER_297_2527 ();
 FILLCELL_X32 FILLER_297_2559 ();
 FILLCELL_X8 FILLER_297_2591 ();
 FILLCELL_X2 FILLER_297_2599 ();
 FILLCELL_X1 FILLER_297_2601 ();
 FILLCELL_X32 FILLER_298_1 ();
 FILLCELL_X32 FILLER_298_33 ();
 FILLCELL_X32 FILLER_298_65 ();
 FILLCELL_X32 FILLER_298_97 ();
 FILLCELL_X32 FILLER_298_129 ();
 FILLCELL_X32 FILLER_298_161 ();
 FILLCELL_X32 FILLER_298_193 ();
 FILLCELL_X32 FILLER_298_225 ();
 FILLCELL_X32 FILLER_298_257 ();
 FILLCELL_X32 FILLER_298_289 ();
 FILLCELL_X32 FILLER_298_321 ();
 FILLCELL_X32 FILLER_298_353 ();
 FILLCELL_X32 FILLER_298_385 ();
 FILLCELL_X32 FILLER_298_417 ();
 FILLCELL_X32 FILLER_298_449 ();
 FILLCELL_X32 FILLER_298_481 ();
 FILLCELL_X32 FILLER_298_513 ();
 FILLCELL_X32 FILLER_298_545 ();
 FILLCELL_X32 FILLER_298_577 ();
 FILLCELL_X16 FILLER_298_609 ();
 FILLCELL_X4 FILLER_298_625 ();
 FILLCELL_X2 FILLER_298_629 ();
 FILLCELL_X32 FILLER_298_632 ();
 FILLCELL_X32 FILLER_298_664 ();
 FILLCELL_X32 FILLER_298_696 ();
 FILLCELL_X32 FILLER_298_728 ();
 FILLCELL_X32 FILLER_298_760 ();
 FILLCELL_X32 FILLER_298_792 ();
 FILLCELL_X32 FILLER_298_824 ();
 FILLCELL_X32 FILLER_298_856 ();
 FILLCELL_X32 FILLER_298_888 ();
 FILLCELL_X32 FILLER_298_920 ();
 FILLCELL_X32 FILLER_298_952 ();
 FILLCELL_X32 FILLER_298_984 ();
 FILLCELL_X32 FILLER_298_1016 ();
 FILLCELL_X32 FILLER_298_1048 ();
 FILLCELL_X32 FILLER_298_1080 ();
 FILLCELL_X32 FILLER_298_1112 ();
 FILLCELL_X32 FILLER_298_1144 ();
 FILLCELL_X32 FILLER_298_1176 ();
 FILLCELL_X32 FILLER_298_1208 ();
 FILLCELL_X32 FILLER_298_1240 ();
 FILLCELL_X32 FILLER_298_1272 ();
 FILLCELL_X32 FILLER_298_1304 ();
 FILLCELL_X32 FILLER_298_1336 ();
 FILLCELL_X32 FILLER_298_1368 ();
 FILLCELL_X32 FILLER_298_1400 ();
 FILLCELL_X32 FILLER_298_1432 ();
 FILLCELL_X32 FILLER_298_1464 ();
 FILLCELL_X32 FILLER_298_1496 ();
 FILLCELL_X32 FILLER_298_1528 ();
 FILLCELL_X32 FILLER_298_1560 ();
 FILLCELL_X32 FILLER_298_1592 ();
 FILLCELL_X32 FILLER_298_1624 ();
 FILLCELL_X32 FILLER_298_1656 ();
 FILLCELL_X32 FILLER_298_1688 ();
 FILLCELL_X32 FILLER_298_1720 ();
 FILLCELL_X32 FILLER_298_1752 ();
 FILLCELL_X32 FILLER_298_1784 ();
 FILLCELL_X32 FILLER_298_1816 ();
 FILLCELL_X32 FILLER_298_1848 ();
 FILLCELL_X8 FILLER_298_1880 ();
 FILLCELL_X4 FILLER_298_1888 ();
 FILLCELL_X2 FILLER_298_1892 ();
 FILLCELL_X32 FILLER_298_1895 ();
 FILLCELL_X32 FILLER_298_1927 ();
 FILLCELL_X32 FILLER_298_1959 ();
 FILLCELL_X32 FILLER_298_1991 ();
 FILLCELL_X32 FILLER_298_2023 ();
 FILLCELL_X32 FILLER_298_2055 ();
 FILLCELL_X32 FILLER_298_2087 ();
 FILLCELL_X32 FILLER_298_2119 ();
 FILLCELL_X32 FILLER_298_2151 ();
 FILLCELL_X32 FILLER_298_2183 ();
 FILLCELL_X32 FILLER_298_2215 ();
 FILLCELL_X32 FILLER_298_2247 ();
 FILLCELL_X32 FILLER_298_2279 ();
 FILLCELL_X32 FILLER_298_2311 ();
 FILLCELL_X32 FILLER_298_2343 ();
 FILLCELL_X32 FILLER_298_2375 ();
 FILLCELL_X32 FILLER_298_2407 ();
 FILLCELL_X32 FILLER_298_2439 ();
 FILLCELL_X32 FILLER_298_2471 ();
 FILLCELL_X32 FILLER_298_2503 ();
 FILLCELL_X32 FILLER_298_2535 ();
 FILLCELL_X32 FILLER_298_2567 ();
 FILLCELL_X2 FILLER_298_2599 ();
 FILLCELL_X1 FILLER_298_2601 ();
 FILLCELL_X32 FILLER_299_1 ();
 FILLCELL_X32 FILLER_299_33 ();
 FILLCELL_X32 FILLER_299_65 ();
 FILLCELL_X32 FILLER_299_97 ();
 FILLCELL_X32 FILLER_299_129 ();
 FILLCELL_X32 FILLER_299_161 ();
 FILLCELL_X32 FILLER_299_193 ();
 FILLCELL_X32 FILLER_299_225 ();
 FILLCELL_X32 FILLER_299_257 ();
 FILLCELL_X32 FILLER_299_289 ();
 FILLCELL_X32 FILLER_299_321 ();
 FILLCELL_X32 FILLER_299_353 ();
 FILLCELL_X32 FILLER_299_385 ();
 FILLCELL_X32 FILLER_299_417 ();
 FILLCELL_X32 FILLER_299_449 ();
 FILLCELL_X32 FILLER_299_481 ();
 FILLCELL_X32 FILLER_299_513 ();
 FILLCELL_X32 FILLER_299_545 ();
 FILLCELL_X32 FILLER_299_577 ();
 FILLCELL_X32 FILLER_299_609 ();
 FILLCELL_X32 FILLER_299_641 ();
 FILLCELL_X32 FILLER_299_673 ();
 FILLCELL_X32 FILLER_299_705 ();
 FILLCELL_X32 FILLER_299_737 ();
 FILLCELL_X32 FILLER_299_769 ();
 FILLCELL_X32 FILLER_299_801 ();
 FILLCELL_X32 FILLER_299_833 ();
 FILLCELL_X32 FILLER_299_865 ();
 FILLCELL_X32 FILLER_299_897 ();
 FILLCELL_X32 FILLER_299_929 ();
 FILLCELL_X32 FILLER_299_961 ();
 FILLCELL_X32 FILLER_299_993 ();
 FILLCELL_X32 FILLER_299_1025 ();
 FILLCELL_X32 FILLER_299_1057 ();
 FILLCELL_X32 FILLER_299_1089 ();
 FILLCELL_X32 FILLER_299_1121 ();
 FILLCELL_X32 FILLER_299_1153 ();
 FILLCELL_X32 FILLER_299_1185 ();
 FILLCELL_X32 FILLER_299_1217 ();
 FILLCELL_X8 FILLER_299_1249 ();
 FILLCELL_X4 FILLER_299_1257 ();
 FILLCELL_X2 FILLER_299_1261 ();
 FILLCELL_X32 FILLER_299_1264 ();
 FILLCELL_X32 FILLER_299_1296 ();
 FILLCELL_X32 FILLER_299_1328 ();
 FILLCELL_X32 FILLER_299_1360 ();
 FILLCELL_X32 FILLER_299_1392 ();
 FILLCELL_X32 FILLER_299_1424 ();
 FILLCELL_X32 FILLER_299_1456 ();
 FILLCELL_X32 FILLER_299_1488 ();
 FILLCELL_X32 FILLER_299_1520 ();
 FILLCELL_X32 FILLER_299_1552 ();
 FILLCELL_X32 FILLER_299_1584 ();
 FILLCELL_X32 FILLER_299_1616 ();
 FILLCELL_X32 FILLER_299_1648 ();
 FILLCELL_X32 FILLER_299_1680 ();
 FILLCELL_X32 FILLER_299_1712 ();
 FILLCELL_X32 FILLER_299_1744 ();
 FILLCELL_X32 FILLER_299_1776 ();
 FILLCELL_X32 FILLER_299_1808 ();
 FILLCELL_X32 FILLER_299_1840 ();
 FILLCELL_X32 FILLER_299_1872 ();
 FILLCELL_X32 FILLER_299_1904 ();
 FILLCELL_X32 FILLER_299_1936 ();
 FILLCELL_X32 FILLER_299_1968 ();
 FILLCELL_X32 FILLER_299_2000 ();
 FILLCELL_X32 FILLER_299_2032 ();
 FILLCELL_X32 FILLER_299_2064 ();
 FILLCELL_X32 FILLER_299_2096 ();
 FILLCELL_X32 FILLER_299_2128 ();
 FILLCELL_X32 FILLER_299_2160 ();
 FILLCELL_X32 FILLER_299_2192 ();
 FILLCELL_X32 FILLER_299_2224 ();
 FILLCELL_X32 FILLER_299_2256 ();
 FILLCELL_X32 FILLER_299_2288 ();
 FILLCELL_X32 FILLER_299_2320 ();
 FILLCELL_X32 FILLER_299_2352 ();
 FILLCELL_X32 FILLER_299_2384 ();
 FILLCELL_X32 FILLER_299_2416 ();
 FILLCELL_X32 FILLER_299_2448 ();
 FILLCELL_X32 FILLER_299_2480 ();
 FILLCELL_X8 FILLER_299_2512 ();
 FILLCELL_X4 FILLER_299_2520 ();
 FILLCELL_X2 FILLER_299_2524 ();
 FILLCELL_X32 FILLER_299_2527 ();
 FILLCELL_X32 FILLER_299_2559 ();
 FILLCELL_X8 FILLER_299_2591 ();
 FILLCELL_X2 FILLER_299_2599 ();
 FILLCELL_X1 FILLER_299_2601 ();
 FILLCELL_X32 FILLER_300_1 ();
 FILLCELL_X32 FILLER_300_33 ();
 FILLCELL_X32 FILLER_300_65 ();
 FILLCELL_X32 FILLER_300_97 ();
 FILLCELL_X32 FILLER_300_129 ();
 FILLCELL_X32 FILLER_300_161 ();
 FILLCELL_X32 FILLER_300_193 ();
 FILLCELL_X32 FILLER_300_225 ();
 FILLCELL_X32 FILLER_300_257 ();
 FILLCELL_X32 FILLER_300_289 ();
 FILLCELL_X32 FILLER_300_321 ();
 FILLCELL_X32 FILLER_300_353 ();
 FILLCELL_X32 FILLER_300_385 ();
 FILLCELL_X32 FILLER_300_417 ();
 FILLCELL_X32 FILLER_300_449 ();
 FILLCELL_X32 FILLER_300_481 ();
 FILLCELL_X32 FILLER_300_513 ();
 FILLCELL_X32 FILLER_300_545 ();
 FILLCELL_X32 FILLER_300_577 ();
 FILLCELL_X16 FILLER_300_609 ();
 FILLCELL_X4 FILLER_300_625 ();
 FILLCELL_X2 FILLER_300_629 ();
 FILLCELL_X32 FILLER_300_632 ();
 FILLCELL_X32 FILLER_300_664 ();
 FILLCELL_X32 FILLER_300_696 ();
 FILLCELL_X32 FILLER_300_728 ();
 FILLCELL_X32 FILLER_300_760 ();
 FILLCELL_X32 FILLER_300_792 ();
 FILLCELL_X32 FILLER_300_824 ();
 FILLCELL_X32 FILLER_300_856 ();
 FILLCELL_X32 FILLER_300_888 ();
 FILLCELL_X32 FILLER_300_920 ();
 FILLCELL_X32 FILLER_300_952 ();
 FILLCELL_X32 FILLER_300_984 ();
 FILLCELL_X32 FILLER_300_1016 ();
 FILLCELL_X32 FILLER_300_1048 ();
 FILLCELL_X32 FILLER_300_1080 ();
 FILLCELL_X32 FILLER_300_1112 ();
 FILLCELL_X32 FILLER_300_1144 ();
 FILLCELL_X32 FILLER_300_1176 ();
 FILLCELL_X32 FILLER_300_1208 ();
 FILLCELL_X32 FILLER_300_1240 ();
 FILLCELL_X32 FILLER_300_1272 ();
 FILLCELL_X32 FILLER_300_1304 ();
 FILLCELL_X32 FILLER_300_1336 ();
 FILLCELL_X32 FILLER_300_1368 ();
 FILLCELL_X32 FILLER_300_1400 ();
 FILLCELL_X32 FILLER_300_1432 ();
 FILLCELL_X32 FILLER_300_1464 ();
 FILLCELL_X32 FILLER_300_1496 ();
 FILLCELL_X32 FILLER_300_1528 ();
 FILLCELL_X32 FILLER_300_1560 ();
 FILLCELL_X32 FILLER_300_1592 ();
 FILLCELL_X32 FILLER_300_1624 ();
 FILLCELL_X32 FILLER_300_1656 ();
 FILLCELL_X32 FILLER_300_1688 ();
 FILLCELL_X32 FILLER_300_1720 ();
 FILLCELL_X32 FILLER_300_1752 ();
 FILLCELL_X32 FILLER_300_1784 ();
 FILLCELL_X32 FILLER_300_1816 ();
 FILLCELL_X32 FILLER_300_1848 ();
 FILLCELL_X8 FILLER_300_1880 ();
 FILLCELL_X4 FILLER_300_1888 ();
 FILLCELL_X2 FILLER_300_1892 ();
 FILLCELL_X32 FILLER_300_1895 ();
 FILLCELL_X32 FILLER_300_1927 ();
 FILLCELL_X32 FILLER_300_1959 ();
 FILLCELL_X32 FILLER_300_1991 ();
 FILLCELL_X32 FILLER_300_2023 ();
 FILLCELL_X32 FILLER_300_2055 ();
 FILLCELL_X32 FILLER_300_2087 ();
 FILLCELL_X32 FILLER_300_2119 ();
 FILLCELL_X32 FILLER_300_2151 ();
 FILLCELL_X32 FILLER_300_2183 ();
 FILLCELL_X32 FILLER_300_2215 ();
 FILLCELL_X32 FILLER_300_2247 ();
 FILLCELL_X32 FILLER_300_2279 ();
 FILLCELL_X32 FILLER_300_2311 ();
 FILLCELL_X32 FILLER_300_2343 ();
 FILLCELL_X32 FILLER_300_2375 ();
 FILLCELL_X32 FILLER_300_2407 ();
 FILLCELL_X32 FILLER_300_2439 ();
 FILLCELL_X32 FILLER_300_2471 ();
 FILLCELL_X32 FILLER_300_2503 ();
 FILLCELL_X32 FILLER_300_2535 ();
 FILLCELL_X32 FILLER_300_2567 ();
 FILLCELL_X2 FILLER_300_2599 ();
 FILLCELL_X1 FILLER_300_2601 ();
 FILLCELL_X32 FILLER_301_1 ();
 FILLCELL_X32 FILLER_301_33 ();
 FILLCELL_X32 FILLER_301_65 ();
 FILLCELL_X32 FILLER_301_97 ();
 FILLCELL_X32 FILLER_301_129 ();
 FILLCELL_X32 FILLER_301_161 ();
 FILLCELL_X32 FILLER_301_193 ();
 FILLCELL_X32 FILLER_301_225 ();
 FILLCELL_X32 FILLER_301_257 ();
 FILLCELL_X32 FILLER_301_289 ();
 FILLCELL_X32 FILLER_301_321 ();
 FILLCELL_X32 FILLER_301_353 ();
 FILLCELL_X32 FILLER_301_385 ();
 FILLCELL_X32 FILLER_301_417 ();
 FILLCELL_X32 FILLER_301_449 ();
 FILLCELL_X32 FILLER_301_481 ();
 FILLCELL_X32 FILLER_301_513 ();
 FILLCELL_X32 FILLER_301_545 ();
 FILLCELL_X32 FILLER_301_577 ();
 FILLCELL_X32 FILLER_301_609 ();
 FILLCELL_X32 FILLER_301_641 ();
 FILLCELL_X32 FILLER_301_673 ();
 FILLCELL_X32 FILLER_301_705 ();
 FILLCELL_X32 FILLER_301_737 ();
 FILLCELL_X32 FILLER_301_769 ();
 FILLCELL_X32 FILLER_301_801 ();
 FILLCELL_X32 FILLER_301_833 ();
 FILLCELL_X32 FILLER_301_865 ();
 FILLCELL_X32 FILLER_301_897 ();
 FILLCELL_X32 FILLER_301_929 ();
 FILLCELL_X32 FILLER_301_961 ();
 FILLCELL_X32 FILLER_301_993 ();
 FILLCELL_X32 FILLER_301_1025 ();
 FILLCELL_X32 FILLER_301_1057 ();
 FILLCELL_X32 FILLER_301_1089 ();
 FILLCELL_X32 FILLER_301_1121 ();
 FILLCELL_X32 FILLER_301_1153 ();
 FILLCELL_X32 FILLER_301_1185 ();
 FILLCELL_X32 FILLER_301_1217 ();
 FILLCELL_X8 FILLER_301_1249 ();
 FILLCELL_X4 FILLER_301_1257 ();
 FILLCELL_X2 FILLER_301_1261 ();
 FILLCELL_X32 FILLER_301_1264 ();
 FILLCELL_X32 FILLER_301_1296 ();
 FILLCELL_X32 FILLER_301_1328 ();
 FILLCELL_X32 FILLER_301_1360 ();
 FILLCELL_X32 FILLER_301_1392 ();
 FILLCELL_X32 FILLER_301_1424 ();
 FILLCELL_X32 FILLER_301_1456 ();
 FILLCELL_X32 FILLER_301_1488 ();
 FILLCELL_X32 FILLER_301_1520 ();
 FILLCELL_X32 FILLER_301_1552 ();
 FILLCELL_X32 FILLER_301_1584 ();
 FILLCELL_X32 FILLER_301_1616 ();
 FILLCELL_X32 FILLER_301_1648 ();
 FILLCELL_X32 FILLER_301_1680 ();
 FILLCELL_X32 FILLER_301_1712 ();
 FILLCELL_X32 FILLER_301_1744 ();
 FILLCELL_X32 FILLER_301_1776 ();
 FILLCELL_X32 FILLER_301_1808 ();
 FILLCELL_X32 FILLER_301_1840 ();
 FILLCELL_X32 FILLER_301_1872 ();
 FILLCELL_X32 FILLER_301_1904 ();
 FILLCELL_X32 FILLER_301_1936 ();
 FILLCELL_X32 FILLER_301_1968 ();
 FILLCELL_X32 FILLER_301_2000 ();
 FILLCELL_X32 FILLER_301_2032 ();
 FILLCELL_X32 FILLER_301_2064 ();
 FILLCELL_X32 FILLER_301_2096 ();
 FILLCELL_X32 FILLER_301_2128 ();
 FILLCELL_X32 FILLER_301_2160 ();
 FILLCELL_X32 FILLER_301_2192 ();
 FILLCELL_X32 FILLER_301_2224 ();
 FILLCELL_X32 FILLER_301_2256 ();
 FILLCELL_X32 FILLER_301_2288 ();
 FILLCELL_X32 FILLER_301_2320 ();
 FILLCELL_X32 FILLER_301_2352 ();
 FILLCELL_X32 FILLER_301_2384 ();
 FILLCELL_X32 FILLER_301_2416 ();
 FILLCELL_X32 FILLER_301_2448 ();
 FILLCELL_X32 FILLER_301_2480 ();
 FILLCELL_X8 FILLER_301_2512 ();
 FILLCELL_X4 FILLER_301_2520 ();
 FILLCELL_X2 FILLER_301_2524 ();
 FILLCELL_X32 FILLER_301_2527 ();
 FILLCELL_X32 FILLER_301_2559 ();
 FILLCELL_X8 FILLER_301_2591 ();
 FILLCELL_X2 FILLER_301_2599 ();
 FILLCELL_X1 FILLER_301_2601 ();
 FILLCELL_X32 FILLER_302_1 ();
 FILLCELL_X32 FILLER_302_33 ();
 FILLCELL_X32 FILLER_302_65 ();
 FILLCELL_X32 FILLER_302_97 ();
 FILLCELL_X32 FILLER_302_129 ();
 FILLCELL_X32 FILLER_302_161 ();
 FILLCELL_X32 FILLER_302_193 ();
 FILLCELL_X32 FILLER_302_225 ();
 FILLCELL_X32 FILLER_302_257 ();
 FILLCELL_X32 FILLER_302_289 ();
 FILLCELL_X32 FILLER_302_321 ();
 FILLCELL_X32 FILLER_302_353 ();
 FILLCELL_X32 FILLER_302_385 ();
 FILLCELL_X32 FILLER_302_417 ();
 FILLCELL_X32 FILLER_302_449 ();
 FILLCELL_X32 FILLER_302_481 ();
 FILLCELL_X32 FILLER_302_513 ();
 FILLCELL_X32 FILLER_302_545 ();
 FILLCELL_X32 FILLER_302_577 ();
 FILLCELL_X16 FILLER_302_609 ();
 FILLCELL_X4 FILLER_302_625 ();
 FILLCELL_X2 FILLER_302_629 ();
 FILLCELL_X32 FILLER_302_632 ();
 FILLCELL_X32 FILLER_302_664 ();
 FILLCELL_X32 FILLER_302_696 ();
 FILLCELL_X32 FILLER_302_728 ();
 FILLCELL_X32 FILLER_302_760 ();
 FILLCELL_X32 FILLER_302_792 ();
 FILLCELL_X32 FILLER_302_824 ();
 FILLCELL_X32 FILLER_302_856 ();
 FILLCELL_X32 FILLER_302_888 ();
 FILLCELL_X32 FILLER_302_920 ();
 FILLCELL_X32 FILLER_302_952 ();
 FILLCELL_X32 FILLER_302_984 ();
 FILLCELL_X32 FILLER_302_1016 ();
 FILLCELL_X32 FILLER_302_1048 ();
 FILLCELL_X32 FILLER_302_1080 ();
 FILLCELL_X32 FILLER_302_1112 ();
 FILLCELL_X32 FILLER_302_1144 ();
 FILLCELL_X32 FILLER_302_1176 ();
 FILLCELL_X32 FILLER_302_1208 ();
 FILLCELL_X32 FILLER_302_1240 ();
 FILLCELL_X32 FILLER_302_1272 ();
 FILLCELL_X32 FILLER_302_1304 ();
 FILLCELL_X32 FILLER_302_1336 ();
 FILLCELL_X32 FILLER_302_1368 ();
 FILLCELL_X32 FILLER_302_1400 ();
 FILLCELL_X32 FILLER_302_1432 ();
 FILLCELL_X32 FILLER_302_1464 ();
 FILLCELL_X32 FILLER_302_1496 ();
 FILLCELL_X32 FILLER_302_1528 ();
 FILLCELL_X32 FILLER_302_1560 ();
 FILLCELL_X32 FILLER_302_1592 ();
 FILLCELL_X32 FILLER_302_1624 ();
 FILLCELL_X32 FILLER_302_1656 ();
 FILLCELL_X32 FILLER_302_1688 ();
 FILLCELL_X32 FILLER_302_1720 ();
 FILLCELL_X32 FILLER_302_1752 ();
 FILLCELL_X32 FILLER_302_1784 ();
 FILLCELL_X32 FILLER_302_1816 ();
 FILLCELL_X32 FILLER_302_1848 ();
 FILLCELL_X8 FILLER_302_1880 ();
 FILLCELL_X4 FILLER_302_1888 ();
 FILLCELL_X2 FILLER_302_1892 ();
 FILLCELL_X32 FILLER_302_1895 ();
 FILLCELL_X32 FILLER_302_1927 ();
 FILLCELL_X32 FILLER_302_1959 ();
 FILLCELL_X32 FILLER_302_1991 ();
 FILLCELL_X32 FILLER_302_2023 ();
 FILLCELL_X32 FILLER_302_2055 ();
 FILLCELL_X32 FILLER_302_2087 ();
 FILLCELL_X32 FILLER_302_2119 ();
 FILLCELL_X32 FILLER_302_2151 ();
 FILLCELL_X32 FILLER_302_2183 ();
 FILLCELL_X32 FILLER_302_2215 ();
 FILLCELL_X32 FILLER_302_2247 ();
 FILLCELL_X32 FILLER_302_2279 ();
 FILLCELL_X32 FILLER_302_2311 ();
 FILLCELL_X32 FILLER_302_2343 ();
 FILLCELL_X32 FILLER_302_2375 ();
 FILLCELL_X32 FILLER_302_2407 ();
 FILLCELL_X32 FILLER_302_2439 ();
 FILLCELL_X32 FILLER_302_2471 ();
 FILLCELL_X32 FILLER_302_2503 ();
 FILLCELL_X32 FILLER_302_2535 ();
 FILLCELL_X32 FILLER_302_2567 ();
 FILLCELL_X2 FILLER_302_2599 ();
 FILLCELL_X1 FILLER_302_2601 ();
 FILLCELL_X32 FILLER_303_1 ();
 FILLCELL_X32 FILLER_303_33 ();
 FILLCELL_X32 FILLER_303_65 ();
 FILLCELL_X32 FILLER_303_97 ();
 FILLCELL_X32 FILLER_303_129 ();
 FILLCELL_X32 FILLER_303_161 ();
 FILLCELL_X32 FILLER_303_193 ();
 FILLCELL_X32 FILLER_303_225 ();
 FILLCELL_X32 FILLER_303_257 ();
 FILLCELL_X32 FILLER_303_289 ();
 FILLCELL_X32 FILLER_303_321 ();
 FILLCELL_X32 FILLER_303_353 ();
 FILLCELL_X32 FILLER_303_385 ();
 FILLCELL_X32 FILLER_303_417 ();
 FILLCELL_X32 FILLER_303_449 ();
 FILLCELL_X32 FILLER_303_481 ();
 FILLCELL_X32 FILLER_303_513 ();
 FILLCELL_X32 FILLER_303_545 ();
 FILLCELL_X32 FILLER_303_577 ();
 FILLCELL_X32 FILLER_303_609 ();
 FILLCELL_X32 FILLER_303_641 ();
 FILLCELL_X32 FILLER_303_673 ();
 FILLCELL_X32 FILLER_303_705 ();
 FILLCELL_X32 FILLER_303_737 ();
 FILLCELL_X32 FILLER_303_769 ();
 FILLCELL_X32 FILLER_303_801 ();
 FILLCELL_X32 FILLER_303_833 ();
 FILLCELL_X32 FILLER_303_865 ();
 FILLCELL_X32 FILLER_303_897 ();
 FILLCELL_X32 FILLER_303_929 ();
 FILLCELL_X32 FILLER_303_961 ();
 FILLCELL_X32 FILLER_303_993 ();
 FILLCELL_X32 FILLER_303_1025 ();
 FILLCELL_X32 FILLER_303_1057 ();
 FILLCELL_X32 FILLER_303_1089 ();
 FILLCELL_X32 FILLER_303_1121 ();
 FILLCELL_X32 FILLER_303_1153 ();
 FILLCELL_X32 FILLER_303_1185 ();
 FILLCELL_X32 FILLER_303_1217 ();
 FILLCELL_X8 FILLER_303_1249 ();
 FILLCELL_X4 FILLER_303_1257 ();
 FILLCELL_X2 FILLER_303_1261 ();
 FILLCELL_X32 FILLER_303_1264 ();
 FILLCELL_X32 FILLER_303_1296 ();
 FILLCELL_X32 FILLER_303_1328 ();
 FILLCELL_X32 FILLER_303_1360 ();
 FILLCELL_X32 FILLER_303_1392 ();
 FILLCELL_X32 FILLER_303_1424 ();
 FILLCELL_X32 FILLER_303_1456 ();
 FILLCELL_X32 FILLER_303_1488 ();
 FILLCELL_X32 FILLER_303_1520 ();
 FILLCELL_X32 FILLER_303_1552 ();
 FILLCELL_X32 FILLER_303_1584 ();
 FILLCELL_X32 FILLER_303_1616 ();
 FILLCELL_X32 FILLER_303_1648 ();
 FILLCELL_X32 FILLER_303_1680 ();
 FILLCELL_X32 FILLER_303_1712 ();
 FILLCELL_X32 FILLER_303_1744 ();
 FILLCELL_X32 FILLER_303_1776 ();
 FILLCELL_X32 FILLER_303_1808 ();
 FILLCELL_X32 FILLER_303_1840 ();
 FILLCELL_X32 FILLER_303_1872 ();
 FILLCELL_X32 FILLER_303_1904 ();
 FILLCELL_X32 FILLER_303_1936 ();
 FILLCELL_X32 FILLER_303_1968 ();
 FILLCELL_X32 FILLER_303_2000 ();
 FILLCELL_X32 FILLER_303_2032 ();
 FILLCELL_X32 FILLER_303_2064 ();
 FILLCELL_X32 FILLER_303_2096 ();
 FILLCELL_X32 FILLER_303_2128 ();
 FILLCELL_X32 FILLER_303_2160 ();
 FILLCELL_X32 FILLER_303_2192 ();
 FILLCELL_X32 FILLER_303_2224 ();
 FILLCELL_X32 FILLER_303_2256 ();
 FILLCELL_X32 FILLER_303_2288 ();
 FILLCELL_X32 FILLER_303_2320 ();
 FILLCELL_X32 FILLER_303_2352 ();
 FILLCELL_X32 FILLER_303_2384 ();
 FILLCELL_X32 FILLER_303_2416 ();
 FILLCELL_X32 FILLER_303_2448 ();
 FILLCELL_X32 FILLER_303_2480 ();
 FILLCELL_X8 FILLER_303_2512 ();
 FILLCELL_X4 FILLER_303_2520 ();
 FILLCELL_X2 FILLER_303_2524 ();
 FILLCELL_X32 FILLER_303_2527 ();
 FILLCELL_X32 FILLER_303_2559 ();
 FILLCELL_X8 FILLER_303_2591 ();
 FILLCELL_X2 FILLER_303_2599 ();
 FILLCELL_X1 FILLER_303_2601 ();
 FILLCELL_X32 FILLER_304_1 ();
 FILLCELL_X32 FILLER_304_33 ();
 FILLCELL_X32 FILLER_304_65 ();
 FILLCELL_X32 FILLER_304_97 ();
 FILLCELL_X32 FILLER_304_129 ();
 FILLCELL_X32 FILLER_304_161 ();
 FILLCELL_X32 FILLER_304_193 ();
 FILLCELL_X32 FILLER_304_225 ();
 FILLCELL_X32 FILLER_304_257 ();
 FILLCELL_X32 FILLER_304_289 ();
 FILLCELL_X32 FILLER_304_321 ();
 FILLCELL_X32 FILLER_304_353 ();
 FILLCELL_X32 FILLER_304_385 ();
 FILLCELL_X32 FILLER_304_417 ();
 FILLCELL_X32 FILLER_304_449 ();
 FILLCELL_X32 FILLER_304_481 ();
 FILLCELL_X32 FILLER_304_513 ();
 FILLCELL_X32 FILLER_304_545 ();
 FILLCELL_X32 FILLER_304_577 ();
 FILLCELL_X16 FILLER_304_609 ();
 FILLCELL_X4 FILLER_304_625 ();
 FILLCELL_X2 FILLER_304_629 ();
 FILLCELL_X32 FILLER_304_632 ();
 FILLCELL_X32 FILLER_304_664 ();
 FILLCELL_X32 FILLER_304_696 ();
 FILLCELL_X32 FILLER_304_728 ();
 FILLCELL_X32 FILLER_304_760 ();
 FILLCELL_X32 FILLER_304_792 ();
 FILLCELL_X32 FILLER_304_824 ();
 FILLCELL_X32 FILLER_304_856 ();
 FILLCELL_X32 FILLER_304_888 ();
 FILLCELL_X32 FILLER_304_920 ();
 FILLCELL_X32 FILLER_304_952 ();
 FILLCELL_X32 FILLER_304_984 ();
 FILLCELL_X32 FILLER_304_1016 ();
 FILLCELL_X32 FILLER_304_1048 ();
 FILLCELL_X32 FILLER_304_1080 ();
 FILLCELL_X32 FILLER_304_1112 ();
 FILLCELL_X32 FILLER_304_1144 ();
 FILLCELL_X32 FILLER_304_1176 ();
 FILLCELL_X32 FILLER_304_1208 ();
 FILLCELL_X32 FILLER_304_1240 ();
 FILLCELL_X32 FILLER_304_1272 ();
 FILLCELL_X32 FILLER_304_1304 ();
 FILLCELL_X32 FILLER_304_1336 ();
 FILLCELL_X32 FILLER_304_1368 ();
 FILLCELL_X32 FILLER_304_1400 ();
 FILLCELL_X32 FILLER_304_1432 ();
 FILLCELL_X32 FILLER_304_1464 ();
 FILLCELL_X32 FILLER_304_1496 ();
 FILLCELL_X32 FILLER_304_1528 ();
 FILLCELL_X32 FILLER_304_1560 ();
 FILLCELL_X32 FILLER_304_1592 ();
 FILLCELL_X32 FILLER_304_1624 ();
 FILLCELL_X32 FILLER_304_1656 ();
 FILLCELL_X32 FILLER_304_1688 ();
 FILLCELL_X32 FILLER_304_1720 ();
 FILLCELL_X32 FILLER_304_1752 ();
 FILLCELL_X32 FILLER_304_1784 ();
 FILLCELL_X32 FILLER_304_1816 ();
 FILLCELL_X32 FILLER_304_1848 ();
 FILLCELL_X8 FILLER_304_1880 ();
 FILLCELL_X4 FILLER_304_1888 ();
 FILLCELL_X2 FILLER_304_1892 ();
 FILLCELL_X32 FILLER_304_1895 ();
 FILLCELL_X32 FILLER_304_1927 ();
 FILLCELL_X32 FILLER_304_1959 ();
 FILLCELL_X32 FILLER_304_1991 ();
 FILLCELL_X32 FILLER_304_2023 ();
 FILLCELL_X32 FILLER_304_2055 ();
 FILLCELL_X32 FILLER_304_2087 ();
 FILLCELL_X32 FILLER_304_2119 ();
 FILLCELL_X32 FILLER_304_2151 ();
 FILLCELL_X32 FILLER_304_2183 ();
 FILLCELL_X32 FILLER_304_2215 ();
 FILLCELL_X32 FILLER_304_2247 ();
 FILLCELL_X32 FILLER_304_2279 ();
 FILLCELL_X32 FILLER_304_2311 ();
 FILLCELL_X32 FILLER_304_2343 ();
 FILLCELL_X32 FILLER_304_2375 ();
 FILLCELL_X32 FILLER_304_2407 ();
 FILLCELL_X32 FILLER_304_2439 ();
 FILLCELL_X32 FILLER_304_2471 ();
 FILLCELL_X32 FILLER_304_2503 ();
 FILLCELL_X32 FILLER_304_2535 ();
 FILLCELL_X32 FILLER_304_2567 ();
 FILLCELL_X2 FILLER_304_2599 ();
 FILLCELL_X1 FILLER_304_2601 ();
 FILLCELL_X32 FILLER_305_1 ();
 FILLCELL_X32 FILLER_305_33 ();
 FILLCELL_X32 FILLER_305_65 ();
 FILLCELL_X32 FILLER_305_97 ();
 FILLCELL_X32 FILLER_305_129 ();
 FILLCELL_X32 FILLER_305_161 ();
 FILLCELL_X32 FILLER_305_193 ();
 FILLCELL_X32 FILLER_305_225 ();
 FILLCELL_X32 FILLER_305_257 ();
 FILLCELL_X32 FILLER_305_289 ();
 FILLCELL_X32 FILLER_305_321 ();
 FILLCELL_X32 FILLER_305_353 ();
 FILLCELL_X32 FILLER_305_385 ();
 FILLCELL_X32 FILLER_305_417 ();
 FILLCELL_X32 FILLER_305_449 ();
 FILLCELL_X32 FILLER_305_481 ();
 FILLCELL_X32 FILLER_305_513 ();
 FILLCELL_X32 FILLER_305_545 ();
 FILLCELL_X32 FILLER_305_577 ();
 FILLCELL_X32 FILLER_305_609 ();
 FILLCELL_X32 FILLER_305_641 ();
 FILLCELL_X32 FILLER_305_673 ();
 FILLCELL_X32 FILLER_305_705 ();
 FILLCELL_X32 FILLER_305_737 ();
 FILLCELL_X32 FILLER_305_769 ();
 FILLCELL_X32 FILLER_305_801 ();
 FILLCELL_X32 FILLER_305_833 ();
 FILLCELL_X32 FILLER_305_865 ();
 FILLCELL_X32 FILLER_305_897 ();
 FILLCELL_X32 FILLER_305_929 ();
 FILLCELL_X32 FILLER_305_961 ();
 FILLCELL_X32 FILLER_305_993 ();
 FILLCELL_X32 FILLER_305_1025 ();
 FILLCELL_X32 FILLER_305_1057 ();
 FILLCELL_X32 FILLER_305_1089 ();
 FILLCELL_X32 FILLER_305_1121 ();
 FILLCELL_X32 FILLER_305_1153 ();
 FILLCELL_X32 FILLER_305_1185 ();
 FILLCELL_X32 FILLER_305_1217 ();
 FILLCELL_X8 FILLER_305_1249 ();
 FILLCELL_X4 FILLER_305_1257 ();
 FILLCELL_X2 FILLER_305_1261 ();
 FILLCELL_X32 FILLER_305_1264 ();
 FILLCELL_X32 FILLER_305_1296 ();
 FILLCELL_X32 FILLER_305_1328 ();
 FILLCELL_X32 FILLER_305_1360 ();
 FILLCELL_X32 FILLER_305_1392 ();
 FILLCELL_X32 FILLER_305_1424 ();
 FILLCELL_X32 FILLER_305_1456 ();
 FILLCELL_X32 FILLER_305_1488 ();
 FILLCELL_X32 FILLER_305_1520 ();
 FILLCELL_X32 FILLER_305_1552 ();
 FILLCELL_X32 FILLER_305_1584 ();
 FILLCELL_X32 FILLER_305_1616 ();
 FILLCELL_X32 FILLER_305_1648 ();
 FILLCELL_X32 FILLER_305_1680 ();
 FILLCELL_X32 FILLER_305_1712 ();
 FILLCELL_X32 FILLER_305_1744 ();
 FILLCELL_X32 FILLER_305_1776 ();
 FILLCELL_X32 FILLER_305_1808 ();
 FILLCELL_X32 FILLER_305_1840 ();
 FILLCELL_X32 FILLER_305_1872 ();
 FILLCELL_X32 FILLER_305_1904 ();
 FILLCELL_X32 FILLER_305_1936 ();
 FILLCELL_X32 FILLER_305_1968 ();
 FILLCELL_X32 FILLER_305_2000 ();
 FILLCELL_X32 FILLER_305_2032 ();
 FILLCELL_X32 FILLER_305_2064 ();
 FILLCELL_X32 FILLER_305_2096 ();
 FILLCELL_X32 FILLER_305_2128 ();
 FILLCELL_X32 FILLER_305_2160 ();
 FILLCELL_X32 FILLER_305_2192 ();
 FILLCELL_X32 FILLER_305_2224 ();
 FILLCELL_X32 FILLER_305_2256 ();
 FILLCELL_X32 FILLER_305_2288 ();
 FILLCELL_X32 FILLER_305_2320 ();
 FILLCELL_X32 FILLER_305_2352 ();
 FILLCELL_X32 FILLER_305_2384 ();
 FILLCELL_X32 FILLER_305_2416 ();
 FILLCELL_X32 FILLER_305_2448 ();
 FILLCELL_X32 FILLER_305_2480 ();
 FILLCELL_X8 FILLER_305_2512 ();
 FILLCELL_X4 FILLER_305_2520 ();
 FILLCELL_X2 FILLER_305_2524 ();
 FILLCELL_X32 FILLER_305_2527 ();
 FILLCELL_X32 FILLER_305_2559 ();
 FILLCELL_X8 FILLER_305_2591 ();
 FILLCELL_X2 FILLER_305_2599 ();
 FILLCELL_X1 FILLER_305_2601 ();
 FILLCELL_X32 FILLER_306_1 ();
 FILLCELL_X32 FILLER_306_33 ();
 FILLCELL_X32 FILLER_306_65 ();
 FILLCELL_X32 FILLER_306_97 ();
 FILLCELL_X32 FILLER_306_129 ();
 FILLCELL_X32 FILLER_306_161 ();
 FILLCELL_X32 FILLER_306_193 ();
 FILLCELL_X32 FILLER_306_225 ();
 FILLCELL_X32 FILLER_306_257 ();
 FILLCELL_X32 FILLER_306_289 ();
 FILLCELL_X32 FILLER_306_321 ();
 FILLCELL_X32 FILLER_306_353 ();
 FILLCELL_X32 FILLER_306_385 ();
 FILLCELL_X32 FILLER_306_417 ();
 FILLCELL_X32 FILLER_306_449 ();
 FILLCELL_X32 FILLER_306_481 ();
 FILLCELL_X32 FILLER_306_513 ();
 FILLCELL_X32 FILLER_306_545 ();
 FILLCELL_X32 FILLER_306_577 ();
 FILLCELL_X16 FILLER_306_609 ();
 FILLCELL_X4 FILLER_306_625 ();
 FILLCELL_X2 FILLER_306_629 ();
 FILLCELL_X32 FILLER_306_632 ();
 FILLCELL_X32 FILLER_306_664 ();
 FILLCELL_X32 FILLER_306_696 ();
 FILLCELL_X32 FILLER_306_728 ();
 FILLCELL_X32 FILLER_306_760 ();
 FILLCELL_X32 FILLER_306_792 ();
 FILLCELL_X32 FILLER_306_824 ();
 FILLCELL_X32 FILLER_306_856 ();
 FILLCELL_X32 FILLER_306_888 ();
 FILLCELL_X32 FILLER_306_920 ();
 FILLCELL_X32 FILLER_306_952 ();
 FILLCELL_X32 FILLER_306_984 ();
 FILLCELL_X32 FILLER_306_1016 ();
 FILLCELL_X32 FILLER_306_1048 ();
 FILLCELL_X32 FILLER_306_1080 ();
 FILLCELL_X32 FILLER_306_1112 ();
 FILLCELL_X32 FILLER_306_1144 ();
 FILLCELL_X32 FILLER_306_1176 ();
 FILLCELL_X32 FILLER_306_1208 ();
 FILLCELL_X32 FILLER_306_1240 ();
 FILLCELL_X32 FILLER_306_1272 ();
 FILLCELL_X32 FILLER_306_1304 ();
 FILLCELL_X32 FILLER_306_1336 ();
 FILLCELL_X32 FILLER_306_1368 ();
 FILLCELL_X32 FILLER_306_1400 ();
 FILLCELL_X32 FILLER_306_1432 ();
 FILLCELL_X32 FILLER_306_1464 ();
 FILLCELL_X32 FILLER_306_1496 ();
 FILLCELL_X32 FILLER_306_1528 ();
 FILLCELL_X32 FILLER_306_1560 ();
 FILLCELL_X32 FILLER_306_1592 ();
 FILLCELL_X32 FILLER_306_1624 ();
 FILLCELL_X32 FILLER_306_1656 ();
 FILLCELL_X32 FILLER_306_1688 ();
 FILLCELL_X32 FILLER_306_1720 ();
 FILLCELL_X32 FILLER_306_1752 ();
 FILLCELL_X32 FILLER_306_1784 ();
 FILLCELL_X32 FILLER_306_1816 ();
 FILLCELL_X32 FILLER_306_1848 ();
 FILLCELL_X8 FILLER_306_1880 ();
 FILLCELL_X4 FILLER_306_1888 ();
 FILLCELL_X2 FILLER_306_1892 ();
 FILLCELL_X32 FILLER_306_1895 ();
 FILLCELL_X32 FILLER_306_1927 ();
 FILLCELL_X32 FILLER_306_1959 ();
 FILLCELL_X32 FILLER_306_1991 ();
 FILLCELL_X32 FILLER_306_2023 ();
 FILLCELL_X32 FILLER_306_2055 ();
 FILLCELL_X32 FILLER_306_2087 ();
 FILLCELL_X32 FILLER_306_2119 ();
 FILLCELL_X32 FILLER_306_2151 ();
 FILLCELL_X32 FILLER_306_2183 ();
 FILLCELL_X32 FILLER_306_2215 ();
 FILLCELL_X32 FILLER_306_2247 ();
 FILLCELL_X32 FILLER_306_2279 ();
 FILLCELL_X32 FILLER_306_2311 ();
 FILLCELL_X32 FILLER_306_2343 ();
 FILLCELL_X32 FILLER_306_2375 ();
 FILLCELL_X32 FILLER_306_2407 ();
 FILLCELL_X32 FILLER_306_2439 ();
 FILLCELL_X32 FILLER_306_2471 ();
 FILLCELL_X32 FILLER_306_2503 ();
 FILLCELL_X32 FILLER_306_2535 ();
 FILLCELL_X32 FILLER_306_2567 ();
 FILLCELL_X2 FILLER_306_2599 ();
 FILLCELL_X1 FILLER_306_2601 ();
 FILLCELL_X32 FILLER_307_1 ();
 FILLCELL_X32 FILLER_307_33 ();
 FILLCELL_X32 FILLER_307_65 ();
 FILLCELL_X32 FILLER_307_97 ();
 FILLCELL_X32 FILLER_307_129 ();
 FILLCELL_X32 FILLER_307_161 ();
 FILLCELL_X32 FILLER_307_193 ();
 FILLCELL_X32 FILLER_307_225 ();
 FILLCELL_X32 FILLER_307_257 ();
 FILLCELL_X32 FILLER_307_289 ();
 FILLCELL_X32 FILLER_307_321 ();
 FILLCELL_X32 FILLER_307_353 ();
 FILLCELL_X32 FILLER_307_385 ();
 FILLCELL_X32 FILLER_307_417 ();
 FILLCELL_X32 FILLER_307_449 ();
 FILLCELL_X32 FILLER_307_481 ();
 FILLCELL_X32 FILLER_307_513 ();
 FILLCELL_X32 FILLER_307_545 ();
 FILLCELL_X32 FILLER_307_577 ();
 FILLCELL_X32 FILLER_307_609 ();
 FILLCELL_X32 FILLER_307_641 ();
 FILLCELL_X32 FILLER_307_673 ();
 FILLCELL_X32 FILLER_307_705 ();
 FILLCELL_X32 FILLER_307_737 ();
 FILLCELL_X32 FILLER_307_769 ();
 FILLCELL_X32 FILLER_307_801 ();
 FILLCELL_X32 FILLER_307_833 ();
 FILLCELL_X32 FILLER_307_865 ();
 FILLCELL_X32 FILLER_307_897 ();
 FILLCELL_X32 FILLER_307_929 ();
 FILLCELL_X32 FILLER_307_961 ();
 FILLCELL_X32 FILLER_307_993 ();
 FILLCELL_X32 FILLER_307_1025 ();
 FILLCELL_X32 FILLER_307_1057 ();
 FILLCELL_X32 FILLER_307_1089 ();
 FILLCELL_X32 FILLER_307_1121 ();
 FILLCELL_X32 FILLER_307_1153 ();
 FILLCELL_X32 FILLER_307_1185 ();
 FILLCELL_X32 FILLER_307_1217 ();
 FILLCELL_X8 FILLER_307_1249 ();
 FILLCELL_X4 FILLER_307_1257 ();
 FILLCELL_X2 FILLER_307_1261 ();
 FILLCELL_X32 FILLER_307_1264 ();
 FILLCELL_X32 FILLER_307_1296 ();
 FILLCELL_X32 FILLER_307_1328 ();
 FILLCELL_X32 FILLER_307_1360 ();
 FILLCELL_X32 FILLER_307_1392 ();
 FILLCELL_X32 FILLER_307_1424 ();
 FILLCELL_X32 FILLER_307_1456 ();
 FILLCELL_X32 FILLER_307_1488 ();
 FILLCELL_X32 FILLER_307_1520 ();
 FILLCELL_X32 FILLER_307_1552 ();
 FILLCELL_X32 FILLER_307_1584 ();
 FILLCELL_X32 FILLER_307_1616 ();
 FILLCELL_X32 FILLER_307_1648 ();
 FILLCELL_X32 FILLER_307_1680 ();
 FILLCELL_X32 FILLER_307_1712 ();
 FILLCELL_X32 FILLER_307_1744 ();
 FILLCELL_X32 FILLER_307_1776 ();
 FILLCELL_X32 FILLER_307_1808 ();
 FILLCELL_X32 FILLER_307_1840 ();
 FILLCELL_X32 FILLER_307_1872 ();
 FILLCELL_X32 FILLER_307_1904 ();
 FILLCELL_X32 FILLER_307_1936 ();
 FILLCELL_X32 FILLER_307_1968 ();
 FILLCELL_X32 FILLER_307_2000 ();
 FILLCELL_X32 FILLER_307_2032 ();
 FILLCELL_X32 FILLER_307_2064 ();
 FILLCELL_X32 FILLER_307_2096 ();
 FILLCELL_X32 FILLER_307_2128 ();
 FILLCELL_X32 FILLER_307_2160 ();
 FILLCELL_X32 FILLER_307_2192 ();
 FILLCELL_X32 FILLER_307_2224 ();
 FILLCELL_X32 FILLER_307_2256 ();
 FILLCELL_X32 FILLER_307_2288 ();
 FILLCELL_X32 FILLER_307_2320 ();
 FILLCELL_X32 FILLER_307_2352 ();
 FILLCELL_X32 FILLER_307_2384 ();
 FILLCELL_X32 FILLER_307_2416 ();
 FILLCELL_X32 FILLER_307_2448 ();
 FILLCELL_X32 FILLER_307_2480 ();
 FILLCELL_X8 FILLER_307_2512 ();
 FILLCELL_X4 FILLER_307_2520 ();
 FILLCELL_X2 FILLER_307_2524 ();
 FILLCELL_X32 FILLER_307_2527 ();
 FILLCELL_X32 FILLER_307_2559 ();
 FILLCELL_X8 FILLER_307_2591 ();
 FILLCELL_X2 FILLER_307_2599 ();
 FILLCELL_X1 FILLER_307_2601 ();
 FILLCELL_X32 FILLER_308_1 ();
 FILLCELL_X32 FILLER_308_33 ();
 FILLCELL_X32 FILLER_308_65 ();
 FILLCELL_X32 FILLER_308_97 ();
 FILLCELL_X32 FILLER_308_129 ();
 FILLCELL_X32 FILLER_308_161 ();
 FILLCELL_X32 FILLER_308_193 ();
 FILLCELL_X32 FILLER_308_225 ();
 FILLCELL_X32 FILLER_308_257 ();
 FILLCELL_X32 FILLER_308_289 ();
 FILLCELL_X32 FILLER_308_321 ();
 FILLCELL_X32 FILLER_308_353 ();
 FILLCELL_X32 FILLER_308_385 ();
 FILLCELL_X32 FILLER_308_417 ();
 FILLCELL_X32 FILLER_308_449 ();
 FILLCELL_X32 FILLER_308_481 ();
 FILLCELL_X32 FILLER_308_513 ();
 FILLCELL_X32 FILLER_308_545 ();
 FILLCELL_X32 FILLER_308_577 ();
 FILLCELL_X16 FILLER_308_609 ();
 FILLCELL_X4 FILLER_308_625 ();
 FILLCELL_X2 FILLER_308_629 ();
 FILLCELL_X32 FILLER_308_632 ();
 FILLCELL_X32 FILLER_308_664 ();
 FILLCELL_X32 FILLER_308_696 ();
 FILLCELL_X32 FILLER_308_728 ();
 FILLCELL_X32 FILLER_308_760 ();
 FILLCELL_X32 FILLER_308_792 ();
 FILLCELL_X32 FILLER_308_824 ();
 FILLCELL_X32 FILLER_308_856 ();
 FILLCELL_X32 FILLER_308_888 ();
 FILLCELL_X32 FILLER_308_920 ();
 FILLCELL_X32 FILLER_308_952 ();
 FILLCELL_X32 FILLER_308_984 ();
 FILLCELL_X32 FILLER_308_1016 ();
 FILLCELL_X32 FILLER_308_1048 ();
 FILLCELL_X32 FILLER_308_1080 ();
 FILLCELL_X32 FILLER_308_1112 ();
 FILLCELL_X32 FILLER_308_1144 ();
 FILLCELL_X32 FILLER_308_1176 ();
 FILLCELL_X32 FILLER_308_1208 ();
 FILLCELL_X32 FILLER_308_1240 ();
 FILLCELL_X32 FILLER_308_1272 ();
 FILLCELL_X32 FILLER_308_1304 ();
 FILLCELL_X32 FILLER_308_1336 ();
 FILLCELL_X32 FILLER_308_1368 ();
 FILLCELL_X32 FILLER_308_1400 ();
 FILLCELL_X32 FILLER_308_1432 ();
 FILLCELL_X32 FILLER_308_1464 ();
 FILLCELL_X32 FILLER_308_1496 ();
 FILLCELL_X32 FILLER_308_1528 ();
 FILLCELL_X32 FILLER_308_1560 ();
 FILLCELL_X32 FILLER_308_1592 ();
 FILLCELL_X32 FILLER_308_1624 ();
 FILLCELL_X32 FILLER_308_1656 ();
 FILLCELL_X32 FILLER_308_1688 ();
 FILLCELL_X32 FILLER_308_1720 ();
 FILLCELL_X32 FILLER_308_1752 ();
 FILLCELL_X32 FILLER_308_1784 ();
 FILLCELL_X32 FILLER_308_1816 ();
 FILLCELL_X32 FILLER_308_1848 ();
 FILLCELL_X8 FILLER_308_1880 ();
 FILLCELL_X4 FILLER_308_1888 ();
 FILLCELL_X2 FILLER_308_1892 ();
 FILLCELL_X32 FILLER_308_1895 ();
 FILLCELL_X32 FILLER_308_1927 ();
 FILLCELL_X32 FILLER_308_1959 ();
 FILLCELL_X32 FILLER_308_1991 ();
 FILLCELL_X32 FILLER_308_2023 ();
 FILLCELL_X32 FILLER_308_2055 ();
 FILLCELL_X32 FILLER_308_2087 ();
 FILLCELL_X32 FILLER_308_2119 ();
 FILLCELL_X32 FILLER_308_2151 ();
 FILLCELL_X32 FILLER_308_2183 ();
 FILLCELL_X32 FILLER_308_2215 ();
 FILLCELL_X32 FILLER_308_2247 ();
 FILLCELL_X32 FILLER_308_2279 ();
 FILLCELL_X32 FILLER_308_2311 ();
 FILLCELL_X32 FILLER_308_2343 ();
 FILLCELL_X32 FILLER_308_2375 ();
 FILLCELL_X32 FILLER_308_2407 ();
 FILLCELL_X32 FILLER_308_2439 ();
 FILLCELL_X32 FILLER_308_2471 ();
 FILLCELL_X32 FILLER_308_2503 ();
 FILLCELL_X32 FILLER_308_2535 ();
 FILLCELL_X32 FILLER_308_2567 ();
 FILLCELL_X2 FILLER_308_2599 ();
 FILLCELL_X1 FILLER_308_2601 ();
 FILLCELL_X32 FILLER_309_1 ();
 FILLCELL_X32 FILLER_309_33 ();
 FILLCELL_X32 FILLER_309_65 ();
 FILLCELL_X32 FILLER_309_97 ();
 FILLCELL_X32 FILLER_309_129 ();
 FILLCELL_X32 FILLER_309_161 ();
 FILLCELL_X32 FILLER_309_193 ();
 FILLCELL_X32 FILLER_309_225 ();
 FILLCELL_X32 FILLER_309_257 ();
 FILLCELL_X32 FILLER_309_289 ();
 FILLCELL_X32 FILLER_309_321 ();
 FILLCELL_X32 FILLER_309_353 ();
 FILLCELL_X32 FILLER_309_385 ();
 FILLCELL_X32 FILLER_309_417 ();
 FILLCELL_X32 FILLER_309_449 ();
 FILLCELL_X32 FILLER_309_481 ();
 FILLCELL_X32 FILLER_309_513 ();
 FILLCELL_X32 FILLER_309_545 ();
 FILLCELL_X32 FILLER_309_577 ();
 FILLCELL_X32 FILLER_309_609 ();
 FILLCELL_X32 FILLER_309_641 ();
 FILLCELL_X32 FILLER_309_673 ();
 FILLCELL_X32 FILLER_309_705 ();
 FILLCELL_X32 FILLER_309_737 ();
 FILLCELL_X32 FILLER_309_769 ();
 FILLCELL_X32 FILLER_309_801 ();
 FILLCELL_X32 FILLER_309_833 ();
 FILLCELL_X32 FILLER_309_865 ();
 FILLCELL_X32 FILLER_309_897 ();
 FILLCELL_X32 FILLER_309_929 ();
 FILLCELL_X32 FILLER_309_961 ();
 FILLCELL_X32 FILLER_309_993 ();
 FILLCELL_X32 FILLER_309_1025 ();
 FILLCELL_X32 FILLER_309_1057 ();
 FILLCELL_X32 FILLER_309_1089 ();
 FILLCELL_X32 FILLER_309_1121 ();
 FILLCELL_X32 FILLER_309_1153 ();
 FILLCELL_X32 FILLER_309_1185 ();
 FILLCELL_X32 FILLER_309_1217 ();
 FILLCELL_X8 FILLER_309_1249 ();
 FILLCELL_X4 FILLER_309_1257 ();
 FILLCELL_X2 FILLER_309_1261 ();
 FILLCELL_X32 FILLER_309_1264 ();
 FILLCELL_X32 FILLER_309_1296 ();
 FILLCELL_X32 FILLER_309_1328 ();
 FILLCELL_X32 FILLER_309_1360 ();
 FILLCELL_X32 FILLER_309_1392 ();
 FILLCELL_X32 FILLER_309_1424 ();
 FILLCELL_X32 FILLER_309_1456 ();
 FILLCELL_X32 FILLER_309_1488 ();
 FILLCELL_X32 FILLER_309_1520 ();
 FILLCELL_X32 FILLER_309_1552 ();
 FILLCELL_X32 FILLER_309_1584 ();
 FILLCELL_X32 FILLER_309_1616 ();
 FILLCELL_X32 FILLER_309_1648 ();
 FILLCELL_X32 FILLER_309_1680 ();
 FILLCELL_X32 FILLER_309_1712 ();
 FILLCELL_X32 FILLER_309_1744 ();
 FILLCELL_X32 FILLER_309_1776 ();
 FILLCELL_X32 FILLER_309_1808 ();
 FILLCELL_X32 FILLER_309_1840 ();
 FILLCELL_X32 FILLER_309_1872 ();
 FILLCELL_X32 FILLER_309_1904 ();
 FILLCELL_X32 FILLER_309_1936 ();
 FILLCELL_X32 FILLER_309_1968 ();
 FILLCELL_X32 FILLER_309_2000 ();
 FILLCELL_X32 FILLER_309_2032 ();
 FILLCELL_X32 FILLER_309_2064 ();
 FILLCELL_X32 FILLER_309_2096 ();
 FILLCELL_X32 FILLER_309_2128 ();
 FILLCELL_X32 FILLER_309_2160 ();
 FILLCELL_X32 FILLER_309_2192 ();
 FILLCELL_X32 FILLER_309_2224 ();
 FILLCELL_X32 FILLER_309_2256 ();
 FILLCELL_X32 FILLER_309_2288 ();
 FILLCELL_X32 FILLER_309_2320 ();
 FILLCELL_X32 FILLER_309_2352 ();
 FILLCELL_X32 FILLER_309_2384 ();
 FILLCELL_X32 FILLER_309_2416 ();
 FILLCELL_X32 FILLER_309_2448 ();
 FILLCELL_X32 FILLER_309_2480 ();
 FILLCELL_X8 FILLER_309_2512 ();
 FILLCELL_X4 FILLER_309_2520 ();
 FILLCELL_X2 FILLER_309_2524 ();
 FILLCELL_X32 FILLER_309_2527 ();
 FILLCELL_X32 FILLER_309_2559 ();
 FILLCELL_X8 FILLER_309_2591 ();
 FILLCELL_X2 FILLER_309_2599 ();
 FILLCELL_X1 FILLER_309_2601 ();
 FILLCELL_X32 FILLER_310_1 ();
 FILLCELL_X32 FILLER_310_33 ();
 FILLCELL_X32 FILLER_310_65 ();
 FILLCELL_X32 FILLER_310_97 ();
 FILLCELL_X32 FILLER_310_129 ();
 FILLCELL_X32 FILLER_310_161 ();
 FILLCELL_X32 FILLER_310_193 ();
 FILLCELL_X32 FILLER_310_225 ();
 FILLCELL_X32 FILLER_310_257 ();
 FILLCELL_X32 FILLER_310_289 ();
 FILLCELL_X32 FILLER_310_321 ();
 FILLCELL_X32 FILLER_310_353 ();
 FILLCELL_X32 FILLER_310_385 ();
 FILLCELL_X32 FILLER_310_417 ();
 FILLCELL_X32 FILLER_310_449 ();
 FILLCELL_X32 FILLER_310_481 ();
 FILLCELL_X32 FILLER_310_513 ();
 FILLCELL_X32 FILLER_310_545 ();
 FILLCELL_X32 FILLER_310_577 ();
 FILLCELL_X16 FILLER_310_609 ();
 FILLCELL_X4 FILLER_310_625 ();
 FILLCELL_X2 FILLER_310_629 ();
 FILLCELL_X32 FILLER_310_632 ();
 FILLCELL_X32 FILLER_310_664 ();
 FILLCELL_X32 FILLER_310_696 ();
 FILLCELL_X32 FILLER_310_728 ();
 FILLCELL_X32 FILLER_310_760 ();
 FILLCELL_X32 FILLER_310_792 ();
 FILLCELL_X32 FILLER_310_824 ();
 FILLCELL_X32 FILLER_310_856 ();
 FILLCELL_X32 FILLER_310_888 ();
 FILLCELL_X32 FILLER_310_920 ();
 FILLCELL_X32 FILLER_310_952 ();
 FILLCELL_X32 FILLER_310_984 ();
 FILLCELL_X32 FILLER_310_1016 ();
 FILLCELL_X32 FILLER_310_1048 ();
 FILLCELL_X32 FILLER_310_1080 ();
 FILLCELL_X32 FILLER_310_1112 ();
 FILLCELL_X32 FILLER_310_1144 ();
 FILLCELL_X32 FILLER_310_1176 ();
 FILLCELL_X32 FILLER_310_1208 ();
 FILLCELL_X32 FILLER_310_1240 ();
 FILLCELL_X32 FILLER_310_1272 ();
 FILLCELL_X32 FILLER_310_1304 ();
 FILLCELL_X32 FILLER_310_1336 ();
 FILLCELL_X32 FILLER_310_1368 ();
 FILLCELL_X32 FILLER_310_1400 ();
 FILLCELL_X32 FILLER_310_1432 ();
 FILLCELL_X32 FILLER_310_1464 ();
 FILLCELL_X32 FILLER_310_1496 ();
 FILLCELL_X32 FILLER_310_1528 ();
 FILLCELL_X32 FILLER_310_1560 ();
 FILLCELL_X32 FILLER_310_1592 ();
 FILLCELL_X32 FILLER_310_1624 ();
 FILLCELL_X32 FILLER_310_1656 ();
 FILLCELL_X32 FILLER_310_1688 ();
 FILLCELL_X32 FILLER_310_1720 ();
 FILLCELL_X32 FILLER_310_1752 ();
 FILLCELL_X32 FILLER_310_1784 ();
 FILLCELL_X32 FILLER_310_1816 ();
 FILLCELL_X32 FILLER_310_1848 ();
 FILLCELL_X8 FILLER_310_1880 ();
 FILLCELL_X4 FILLER_310_1888 ();
 FILLCELL_X2 FILLER_310_1892 ();
 FILLCELL_X32 FILLER_310_1895 ();
 FILLCELL_X32 FILLER_310_1927 ();
 FILLCELL_X32 FILLER_310_1959 ();
 FILLCELL_X32 FILLER_310_1991 ();
 FILLCELL_X32 FILLER_310_2023 ();
 FILLCELL_X32 FILLER_310_2055 ();
 FILLCELL_X32 FILLER_310_2087 ();
 FILLCELL_X32 FILLER_310_2119 ();
 FILLCELL_X32 FILLER_310_2151 ();
 FILLCELL_X32 FILLER_310_2183 ();
 FILLCELL_X32 FILLER_310_2215 ();
 FILLCELL_X32 FILLER_310_2247 ();
 FILLCELL_X32 FILLER_310_2279 ();
 FILLCELL_X32 FILLER_310_2311 ();
 FILLCELL_X32 FILLER_310_2343 ();
 FILLCELL_X32 FILLER_310_2375 ();
 FILLCELL_X32 FILLER_310_2407 ();
 FILLCELL_X32 FILLER_310_2439 ();
 FILLCELL_X32 FILLER_310_2471 ();
 FILLCELL_X32 FILLER_310_2503 ();
 FILLCELL_X32 FILLER_310_2535 ();
 FILLCELL_X32 FILLER_310_2567 ();
 FILLCELL_X2 FILLER_310_2599 ();
 FILLCELL_X1 FILLER_310_2601 ();
 FILLCELL_X32 FILLER_311_1 ();
 FILLCELL_X32 FILLER_311_33 ();
 FILLCELL_X32 FILLER_311_65 ();
 FILLCELL_X32 FILLER_311_97 ();
 FILLCELL_X32 FILLER_311_129 ();
 FILLCELL_X32 FILLER_311_161 ();
 FILLCELL_X32 FILLER_311_193 ();
 FILLCELL_X32 FILLER_311_225 ();
 FILLCELL_X32 FILLER_311_257 ();
 FILLCELL_X32 FILLER_311_289 ();
 FILLCELL_X32 FILLER_311_321 ();
 FILLCELL_X32 FILLER_311_353 ();
 FILLCELL_X32 FILLER_311_385 ();
 FILLCELL_X32 FILLER_311_417 ();
 FILLCELL_X32 FILLER_311_449 ();
 FILLCELL_X32 FILLER_311_481 ();
 FILLCELL_X32 FILLER_311_513 ();
 FILLCELL_X32 FILLER_311_545 ();
 FILLCELL_X32 FILLER_311_577 ();
 FILLCELL_X32 FILLER_311_609 ();
 FILLCELL_X32 FILLER_311_641 ();
 FILLCELL_X32 FILLER_311_673 ();
 FILLCELL_X32 FILLER_311_705 ();
 FILLCELL_X32 FILLER_311_737 ();
 FILLCELL_X32 FILLER_311_769 ();
 FILLCELL_X32 FILLER_311_801 ();
 FILLCELL_X32 FILLER_311_833 ();
 FILLCELL_X32 FILLER_311_865 ();
 FILLCELL_X32 FILLER_311_897 ();
 FILLCELL_X32 FILLER_311_929 ();
 FILLCELL_X32 FILLER_311_961 ();
 FILLCELL_X32 FILLER_311_993 ();
 FILLCELL_X32 FILLER_311_1025 ();
 FILLCELL_X32 FILLER_311_1057 ();
 FILLCELL_X32 FILLER_311_1089 ();
 FILLCELL_X32 FILLER_311_1121 ();
 FILLCELL_X32 FILLER_311_1153 ();
 FILLCELL_X32 FILLER_311_1185 ();
 FILLCELL_X32 FILLER_311_1217 ();
 FILLCELL_X8 FILLER_311_1249 ();
 FILLCELL_X4 FILLER_311_1257 ();
 FILLCELL_X2 FILLER_311_1261 ();
 FILLCELL_X32 FILLER_311_1264 ();
 FILLCELL_X32 FILLER_311_1296 ();
 FILLCELL_X32 FILLER_311_1328 ();
 FILLCELL_X32 FILLER_311_1360 ();
 FILLCELL_X32 FILLER_311_1392 ();
 FILLCELL_X32 FILLER_311_1424 ();
 FILLCELL_X32 FILLER_311_1456 ();
 FILLCELL_X32 FILLER_311_1488 ();
 FILLCELL_X32 FILLER_311_1520 ();
 FILLCELL_X32 FILLER_311_1552 ();
 FILLCELL_X32 FILLER_311_1584 ();
 FILLCELL_X32 FILLER_311_1616 ();
 FILLCELL_X32 FILLER_311_1648 ();
 FILLCELL_X32 FILLER_311_1680 ();
 FILLCELL_X32 FILLER_311_1712 ();
 FILLCELL_X32 FILLER_311_1744 ();
 FILLCELL_X32 FILLER_311_1776 ();
 FILLCELL_X32 FILLER_311_1808 ();
 FILLCELL_X32 FILLER_311_1840 ();
 FILLCELL_X32 FILLER_311_1872 ();
 FILLCELL_X32 FILLER_311_1904 ();
 FILLCELL_X32 FILLER_311_1936 ();
 FILLCELL_X32 FILLER_311_1968 ();
 FILLCELL_X32 FILLER_311_2000 ();
 FILLCELL_X32 FILLER_311_2032 ();
 FILLCELL_X32 FILLER_311_2064 ();
 FILLCELL_X32 FILLER_311_2096 ();
 FILLCELL_X32 FILLER_311_2128 ();
 FILLCELL_X32 FILLER_311_2160 ();
 FILLCELL_X32 FILLER_311_2192 ();
 FILLCELL_X32 FILLER_311_2224 ();
 FILLCELL_X32 FILLER_311_2256 ();
 FILLCELL_X32 FILLER_311_2288 ();
 FILLCELL_X32 FILLER_311_2320 ();
 FILLCELL_X32 FILLER_311_2352 ();
 FILLCELL_X32 FILLER_311_2384 ();
 FILLCELL_X32 FILLER_311_2416 ();
 FILLCELL_X32 FILLER_311_2448 ();
 FILLCELL_X32 FILLER_311_2480 ();
 FILLCELL_X8 FILLER_311_2512 ();
 FILLCELL_X4 FILLER_311_2520 ();
 FILLCELL_X2 FILLER_311_2524 ();
 FILLCELL_X32 FILLER_311_2527 ();
 FILLCELL_X32 FILLER_311_2559 ();
 FILLCELL_X8 FILLER_311_2591 ();
 FILLCELL_X2 FILLER_311_2599 ();
 FILLCELL_X1 FILLER_311_2601 ();
 FILLCELL_X32 FILLER_312_1 ();
 FILLCELL_X32 FILLER_312_33 ();
 FILLCELL_X32 FILLER_312_65 ();
 FILLCELL_X32 FILLER_312_97 ();
 FILLCELL_X32 FILLER_312_129 ();
 FILLCELL_X32 FILLER_312_161 ();
 FILLCELL_X32 FILLER_312_193 ();
 FILLCELL_X32 FILLER_312_225 ();
 FILLCELL_X32 FILLER_312_257 ();
 FILLCELL_X32 FILLER_312_289 ();
 FILLCELL_X32 FILLER_312_321 ();
 FILLCELL_X32 FILLER_312_353 ();
 FILLCELL_X32 FILLER_312_385 ();
 FILLCELL_X32 FILLER_312_417 ();
 FILLCELL_X32 FILLER_312_449 ();
 FILLCELL_X32 FILLER_312_481 ();
 FILLCELL_X32 FILLER_312_513 ();
 FILLCELL_X32 FILLER_312_545 ();
 FILLCELL_X32 FILLER_312_577 ();
 FILLCELL_X16 FILLER_312_609 ();
 FILLCELL_X4 FILLER_312_625 ();
 FILLCELL_X2 FILLER_312_629 ();
 FILLCELL_X32 FILLER_312_632 ();
 FILLCELL_X32 FILLER_312_664 ();
 FILLCELL_X32 FILLER_312_696 ();
 FILLCELL_X32 FILLER_312_728 ();
 FILLCELL_X32 FILLER_312_760 ();
 FILLCELL_X32 FILLER_312_792 ();
 FILLCELL_X32 FILLER_312_824 ();
 FILLCELL_X32 FILLER_312_856 ();
 FILLCELL_X32 FILLER_312_888 ();
 FILLCELL_X32 FILLER_312_920 ();
 FILLCELL_X32 FILLER_312_952 ();
 FILLCELL_X32 FILLER_312_984 ();
 FILLCELL_X32 FILLER_312_1016 ();
 FILLCELL_X32 FILLER_312_1048 ();
 FILLCELL_X32 FILLER_312_1080 ();
 FILLCELL_X32 FILLER_312_1112 ();
 FILLCELL_X32 FILLER_312_1144 ();
 FILLCELL_X32 FILLER_312_1176 ();
 FILLCELL_X32 FILLER_312_1208 ();
 FILLCELL_X32 FILLER_312_1240 ();
 FILLCELL_X32 FILLER_312_1272 ();
 FILLCELL_X32 FILLER_312_1304 ();
 FILLCELL_X32 FILLER_312_1336 ();
 FILLCELL_X32 FILLER_312_1368 ();
 FILLCELL_X32 FILLER_312_1400 ();
 FILLCELL_X32 FILLER_312_1432 ();
 FILLCELL_X32 FILLER_312_1464 ();
 FILLCELL_X32 FILLER_312_1496 ();
 FILLCELL_X32 FILLER_312_1528 ();
 FILLCELL_X32 FILLER_312_1560 ();
 FILLCELL_X32 FILLER_312_1592 ();
 FILLCELL_X32 FILLER_312_1624 ();
 FILLCELL_X32 FILLER_312_1656 ();
 FILLCELL_X32 FILLER_312_1688 ();
 FILLCELL_X32 FILLER_312_1720 ();
 FILLCELL_X32 FILLER_312_1752 ();
 FILLCELL_X32 FILLER_312_1784 ();
 FILLCELL_X32 FILLER_312_1816 ();
 FILLCELL_X32 FILLER_312_1848 ();
 FILLCELL_X8 FILLER_312_1880 ();
 FILLCELL_X4 FILLER_312_1888 ();
 FILLCELL_X2 FILLER_312_1892 ();
 FILLCELL_X32 FILLER_312_1895 ();
 FILLCELL_X32 FILLER_312_1927 ();
 FILLCELL_X32 FILLER_312_1959 ();
 FILLCELL_X32 FILLER_312_1991 ();
 FILLCELL_X32 FILLER_312_2023 ();
 FILLCELL_X32 FILLER_312_2055 ();
 FILLCELL_X32 FILLER_312_2087 ();
 FILLCELL_X32 FILLER_312_2119 ();
 FILLCELL_X32 FILLER_312_2151 ();
 FILLCELL_X32 FILLER_312_2183 ();
 FILLCELL_X32 FILLER_312_2215 ();
 FILLCELL_X32 FILLER_312_2247 ();
 FILLCELL_X32 FILLER_312_2279 ();
 FILLCELL_X32 FILLER_312_2311 ();
 FILLCELL_X32 FILLER_312_2343 ();
 FILLCELL_X32 FILLER_312_2375 ();
 FILLCELL_X32 FILLER_312_2407 ();
 FILLCELL_X32 FILLER_312_2439 ();
 FILLCELL_X32 FILLER_312_2471 ();
 FILLCELL_X32 FILLER_312_2503 ();
 FILLCELL_X32 FILLER_312_2535 ();
 FILLCELL_X32 FILLER_312_2567 ();
 FILLCELL_X2 FILLER_312_2599 ();
 FILLCELL_X1 FILLER_312_2601 ();
 FILLCELL_X32 FILLER_313_1 ();
 FILLCELL_X32 FILLER_313_33 ();
 FILLCELL_X32 FILLER_313_65 ();
 FILLCELL_X32 FILLER_313_97 ();
 FILLCELL_X32 FILLER_313_129 ();
 FILLCELL_X32 FILLER_313_161 ();
 FILLCELL_X32 FILLER_313_193 ();
 FILLCELL_X32 FILLER_313_225 ();
 FILLCELL_X32 FILLER_313_257 ();
 FILLCELL_X32 FILLER_313_289 ();
 FILLCELL_X32 FILLER_313_321 ();
 FILLCELL_X32 FILLER_313_353 ();
 FILLCELL_X32 FILLER_313_385 ();
 FILLCELL_X32 FILLER_313_417 ();
 FILLCELL_X32 FILLER_313_449 ();
 FILLCELL_X32 FILLER_313_481 ();
 FILLCELL_X32 FILLER_313_513 ();
 FILLCELL_X32 FILLER_313_545 ();
 FILLCELL_X32 FILLER_313_577 ();
 FILLCELL_X32 FILLER_313_609 ();
 FILLCELL_X32 FILLER_313_641 ();
 FILLCELL_X32 FILLER_313_673 ();
 FILLCELL_X32 FILLER_313_705 ();
 FILLCELL_X32 FILLER_313_737 ();
 FILLCELL_X32 FILLER_313_769 ();
 FILLCELL_X32 FILLER_313_801 ();
 FILLCELL_X32 FILLER_313_833 ();
 FILLCELL_X32 FILLER_313_865 ();
 FILLCELL_X32 FILLER_313_897 ();
 FILLCELL_X32 FILLER_313_929 ();
 FILLCELL_X32 FILLER_313_961 ();
 FILLCELL_X32 FILLER_313_993 ();
 FILLCELL_X32 FILLER_313_1025 ();
 FILLCELL_X32 FILLER_313_1057 ();
 FILLCELL_X32 FILLER_313_1089 ();
 FILLCELL_X32 FILLER_313_1121 ();
 FILLCELL_X32 FILLER_313_1153 ();
 FILLCELL_X32 FILLER_313_1185 ();
 FILLCELL_X32 FILLER_313_1217 ();
 FILLCELL_X8 FILLER_313_1249 ();
 FILLCELL_X4 FILLER_313_1257 ();
 FILLCELL_X2 FILLER_313_1261 ();
 FILLCELL_X32 FILLER_313_1264 ();
 FILLCELL_X32 FILLER_313_1296 ();
 FILLCELL_X32 FILLER_313_1328 ();
 FILLCELL_X32 FILLER_313_1360 ();
 FILLCELL_X32 FILLER_313_1392 ();
 FILLCELL_X32 FILLER_313_1424 ();
 FILLCELL_X32 FILLER_313_1456 ();
 FILLCELL_X32 FILLER_313_1488 ();
 FILLCELL_X32 FILLER_313_1520 ();
 FILLCELL_X32 FILLER_313_1552 ();
 FILLCELL_X32 FILLER_313_1584 ();
 FILLCELL_X32 FILLER_313_1616 ();
 FILLCELL_X32 FILLER_313_1648 ();
 FILLCELL_X32 FILLER_313_1680 ();
 FILLCELL_X32 FILLER_313_1712 ();
 FILLCELL_X32 FILLER_313_1744 ();
 FILLCELL_X32 FILLER_313_1776 ();
 FILLCELL_X32 FILLER_313_1808 ();
 FILLCELL_X32 FILLER_313_1840 ();
 FILLCELL_X32 FILLER_313_1872 ();
 FILLCELL_X32 FILLER_313_1904 ();
 FILLCELL_X32 FILLER_313_1936 ();
 FILLCELL_X32 FILLER_313_1968 ();
 FILLCELL_X32 FILLER_313_2000 ();
 FILLCELL_X32 FILLER_313_2032 ();
 FILLCELL_X32 FILLER_313_2064 ();
 FILLCELL_X32 FILLER_313_2096 ();
 FILLCELL_X32 FILLER_313_2128 ();
 FILLCELL_X32 FILLER_313_2160 ();
 FILLCELL_X32 FILLER_313_2192 ();
 FILLCELL_X32 FILLER_313_2224 ();
 FILLCELL_X32 FILLER_313_2256 ();
 FILLCELL_X32 FILLER_313_2288 ();
 FILLCELL_X32 FILLER_313_2320 ();
 FILLCELL_X32 FILLER_313_2352 ();
 FILLCELL_X32 FILLER_313_2384 ();
 FILLCELL_X32 FILLER_313_2416 ();
 FILLCELL_X32 FILLER_313_2448 ();
 FILLCELL_X32 FILLER_313_2480 ();
 FILLCELL_X8 FILLER_313_2512 ();
 FILLCELL_X4 FILLER_313_2520 ();
 FILLCELL_X2 FILLER_313_2524 ();
 FILLCELL_X32 FILLER_313_2527 ();
 FILLCELL_X32 FILLER_313_2559 ();
 FILLCELL_X8 FILLER_313_2591 ();
 FILLCELL_X2 FILLER_313_2599 ();
 FILLCELL_X1 FILLER_313_2601 ();
 FILLCELL_X32 FILLER_314_1 ();
 FILLCELL_X32 FILLER_314_33 ();
 FILLCELL_X32 FILLER_314_65 ();
 FILLCELL_X32 FILLER_314_97 ();
 FILLCELL_X32 FILLER_314_129 ();
 FILLCELL_X32 FILLER_314_161 ();
 FILLCELL_X32 FILLER_314_193 ();
 FILLCELL_X32 FILLER_314_225 ();
 FILLCELL_X32 FILLER_314_257 ();
 FILLCELL_X32 FILLER_314_289 ();
 FILLCELL_X32 FILLER_314_321 ();
 FILLCELL_X32 FILLER_314_353 ();
 FILLCELL_X32 FILLER_314_385 ();
 FILLCELL_X32 FILLER_314_417 ();
 FILLCELL_X32 FILLER_314_449 ();
 FILLCELL_X32 FILLER_314_481 ();
 FILLCELL_X32 FILLER_314_513 ();
 FILLCELL_X32 FILLER_314_545 ();
 FILLCELL_X32 FILLER_314_577 ();
 FILLCELL_X16 FILLER_314_609 ();
 FILLCELL_X4 FILLER_314_625 ();
 FILLCELL_X2 FILLER_314_629 ();
 FILLCELL_X32 FILLER_314_632 ();
 FILLCELL_X32 FILLER_314_664 ();
 FILLCELL_X32 FILLER_314_696 ();
 FILLCELL_X32 FILLER_314_728 ();
 FILLCELL_X32 FILLER_314_760 ();
 FILLCELL_X32 FILLER_314_792 ();
 FILLCELL_X32 FILLER_314_824 ();
 FILLCELL_X32 FILLER_314_856 ();
 FILLCELL_X32 FILLER_314_888 ();
 FILLCELL_X32 FILLER_314_920 ();
 FILLCELL_X32 FILLER_314_952 ();
 FILLCELL_X32 FILLER_314_984 ();
 FILLCELL_X32 FILLER_314_1016 ();
 FILLCELL_X32 FILLER_314_1048 ();
 FILLCELL_X32 FILLER_314_1080 ();
 FILLCELL_X32 FILLER_314_1112 ();
 FILLCELL_X32 FILLER_314_1144 ();
 FILLCELL_X32 FILLER_314_1176 ();
 FILLCELL_X32 FILLER_314_1208 ();
 FILLCELL_X32 FILLER_314_1240 ();
 FILLCELL_X32 FILLER_314_1272 ();
 FILLCELL_X32 FILLER_314_1304 ();
 FILLCELL_X32 FILLER_314_1336 ();
 FILLCELL_X32 FILLER_314_1368 ();
 FILLCELL_X32 FILLER_314_1400 ();
 FILLCELL_X32 FILLER_314_1432 ();
 FILLCELL_X32 FILLER_314_1464 ();
 FILLCELL_X32 FILLER_314_1496 ();
 FILLCELL_X32 FILLER_314_1528 ();
 FILLCELL_X32 FILLER_314_1560 ();
 FILLCELL_X32 FILLER_314_1592 ();
 FILLCELL_X32 FILLER_314_1624 ();
 FILLCELL_X32 FILLER_314_1656 ();
 FILLCELL_X32 FILLER_314_1688 ();
 FILLCELL_X32 FILLER_314_1720 ();
 FILLCELL_X32 FILLER_314_1752 ();
 FILLCELL_X32 FILLER_314_1784 ();
 FILLCELL_X32 FILLER_314_1816 ();
 FILLCELL_X32 FILLER_314_1848 ();
 FILLCELL_X8 FILLER_314_1880 ();
 FILLCELL_X4 FILLER_314_1888 ();
 FILLCELL_X2 FILLER_314_1892 ();
 FILLCELL_X32 FILLER_314_1895 ();
 FILLCELL_X32 FILLER_314_1927 ();
 FILLCELL_X32 FILLER_314_1959 ();
 FILLCELL_X32 FILLER_314_1991 ();
 FILLCELL_X32 FILLER_314_2023 ();
 FILLCELL_X32 FILLER_314_2055 ();
 FILLCELL_X32 FILLER_314_2087 ();
 FILLCELL_X32 FILLER_314_2119 ();
 FILLCELL_X32 FILLER_314_2151 ();
 FILLCELL_X32 FILLER_314_2183 ();
 FILLCELL_X32 FILLER_314_2215 ();
 FILLCELL_X32 FILLER_314_2247 ();
 FILLCELL_X32 FILLER_314_2279 ();
 FILLCELL_X32 FILLER_314_2311 ();
 FILLCELL_X32 FILLER_314_2343 ();
 FILLCELL_X32 FILLER_314_2375 ();
 FILLCELL_X32 FILLER_314_2407 ();
 FILLCELL_X32 FILLER_314_2439 ();
 FILLCELL_X32 FILLER_314_2471 ();
 FILLCELL_X32 FILLER_314_2503 ();
 FILLCELL_X32 FILLER_314_2535 ();
 FILLCELL_X32 FILLER_314_2567 ();
 FILLCELL_X2 FILLER_314_2599 ();
 FILLCELL_X1 FILLER_314_2601 ();
 FILLCELL_X32 FILLER_315_1 ();
 FILLCELL_X32 FILLER_315_33 ();
 FILLCELL_X32 FILLER_315_65 ();
 FILLCELL_X32 FILLER_315_97 ();
 FILLCELL_X32 FILLER_315_129 ();
 FILLCELL_X32 FILLER_315_161 ();
 FILLCELL_X32 FILLER_315_193 ();
 FILLCELL_X32 FILLER_315_225 ();
 FILLCELL_X32 FILLER_315_257 ();
 FILLCELL_X32 FILLER_315_289 ();
 FILLCELL_X32 FILLER_315_321 ();
 FILLCELL_X32 FILLER_315_353 ();
 FILLCELL_X32 FILLER_315_385 ();
 FILLCELL_X32 FILLER_315_417 ();
 FILLCELL_X32 FILLER_315_449 ();
 FILLCELL_X32 FILLER_315_481 ();
 FILLCELL_X32 FILLER_315_513 ();
 FILLCELL_X32 FILLER_315_545 ();
 FILLCELL_X32 FILLER_315_577 ();
 FILLCELL_X32 FILLER_315_609 ();
 FILLCELL_X32 FILLER_315_641 ();
 FILLCELL_X32 FILLER_315_673 ();
 FILLCELL_X32 FILLER_315_705 ();
 FILLCELL_X32 FILLER_315_737 ();
 FILLCELL_X32 FILLER_315_769 ();
 FILLCELL_X32 FILLER_315_801 ();
 FILLCELL_X32 FILLER_315_833 ();
 FILLCELL_X32 FILLER_315_865 ();
 FILLCELL_X32 FILLER_315_897 ();
 FILLCELL_X32 FILLER_315_929 ();
 FILLCELL_X32 FILLER_315_961 ();
 FILLCELL_X32 FILLER_315_993 ();
 FILLCELL_X32 FILLER_315_1025 ();
 FILLCELL_X32 FILLER_315_1057 ();
 FILLCELL_X32 FILLER_315_1089 ();
 FILLCELL_X32 FILLER_315_1121 ();
 FILLCELL_X32 FILLER_315_1153 ();
 FILLCELL_X32 FILLER_315_1185 ();
 FILLCELL_X32 FILLER_315_1217 ();
 FILLCELL_X8 FILLER_315_1249 ();
 FILLCELL_X4 FILLER_315_1257 ();
 FILLCELL_X2 FILLER_315_1261 ();
 FILLCELL_X32 FILLER_315_1264 ();
 FILLCELL_X32 FILLER_315_1296 ();
 FILLCELL_X32 FILLER_315_1328 ();
 FILLCELL_X32 FILLER_315_1360 ();
 FILLCELL_X32 FILLER_315_1392 ();
 FILLCELL_X32 FILLER_315_1424 ();
 FILLCELL_X32 FILLER_315_1456 ();
 FILLCELL_X32 FILLER_315_1488 ();
 FILLCELL_X32 FILLER_315_1520 ();
 FILLCELL_X32 FILLER_315_1552 ();
 FILLCELL_X32 FILLER_315_1584 ();
 FILLCELL_X32 FILLER_315_1616 ();
 FILLCELL_X32 FILLER_315_1648 ();
 FILLCELL_X32 FILLER_315_1680 ();
 FILLCELL_X32 FILLER_315_1712 ();
 FILLCELL_X32 FILLER_315_1744 ();
 FILLCELL_X32 FILLER_315_1776 ();
 FILLCELL_X32 FILLER_315_1808 ();
 FILLCELL_X32 FILLER_315_1840 ();
 FILLCELL_X32 FILLER_315_1872 ();
 FILLCELL_X32 FILLER_315_1904 ();
 FILLCELL_X32 FILLER_315_1936 ();
 FILLCELL_X32 FILLER_315_1968 ();
 FILLCELL_X32 FILLER_315_2000 ();
 FILLCELL_X32 FILLER_315_2032 ();
 FILLCELL_X32 FILLER_315_2064 ();
 FILLCELL_X32 FILLER_315_2096 ();
 FILLCELL_X32 FILLER_315_2128 ();
 FILLCELL_X32 FILLER_315_2160 ();
 FILLCELL_X32 FILLER_315_2192 ();
 FILLCELL_X32 FILLER_315_2224 ();
 FILLCELL_X32 FILLER_315_2256 ();
 FILLCELL_X32 FILLER_315_2288 ();
 FILLCELL_X32 FILLER_315_2320 ();
 FILLCELL_X32 FILLER_315_2352 ();
 FILLCELL_X32 FILLER_315_2384 ();
 FILLCELL_X32 FILLER_315_2416 ();
 FILLCELL_X32 FILLER_315_2448 ();
 FILLCELL_X32 FILLER_315_2480 ();
 FILLCELL_X8 FILLER_315_2512 ();
 FILLCELL_X4 FILLER_315_2520 ();
 FILLCELL_X2 FILLER_315_2524 ();
 FILLCELL_X32 FILLER_315_2527 ();
 FILLCELL_X32 FILLER_315_2559 ();
 FILLCELL_X8 FILLER_315_2591 ();
 FILLCELL_X2 FILLER_315_2599 ();
 FILLCELL_X1 FILLER_315_2601 ();
 FILLCELL_X32 FILLER_316_1 ();
 FILLCELL_X32 FILLER_316_33 ();
 FILLCELL_X32 FILLER_316_65 ();
 FILLCELL_X32 FILLER_316_97 ();
 FILLCELL_X32 FILLER_316_129 ();
 FILLCELL_X32 FILLER_316_161 ();
 FILLCELL_X32 FILLER_316_193 ();
 FILLCELL_X32 FILLER_316_225 ();
 FILLCELL_X32 FILLER_316_257 ();
 FILLCELL_X32 FILLER_316_289 ();
 FILLCELL_X32 FILLER_316_321 ();
 FILLCELL_X32 FILLER_316_353 ();
 FILLCELL_X32 FILLER_316_385 ();
 FILLCELL_X32 FILLER_316_417 ();
 FILLCELL_X32 FILLER_316_449 ();
 FILLCELL_X32 FILLER_316_481 ();
 FILLCELL_X32 FILLER_316_513 ();
 FILLCELL_X32 FILLER_316_545 ();
 FILLCELL_X32 FILLER_316_577 ();
 FILLCELL_X16 FILLER_316_609 ();
 FILLCELL_X4 FILLER_316_625 ();
 FILLCELL_X2 FILLER_316_629 ();
 FILLCELL_X32 FILLER_316_632 ();
 FILLCELL_X32 FILLER_316_664 ();
 FILLCELL_X32 FILLER_316_696 ();
 FILLCELL_X32 FILLER_316_728 ();
 FILLCELL_X32 FILLER_316_760 ();
 FILLCELL_X32 FILLER_316_792 ();
 FILLCELL_X32 FILLER_316_824 ();
 FILLCELL_X32 FILLER_316_856 ();
 FILLCELL_X32 FILLER_316_888 ();
 FILLCELL_X32 FILLER_316_920 ();
 FILLCELL_X32 FILLER_316_952 ();
 FILLCELL_X32 FILLER_316_984 ();
 FILLCELL_X32 FILLER_316_1016 ();
 FILLCELL_X32 FILLER_316_1048 ();
 FILLCELL_X32 FILLER_316_1080 ();
 FILLCELL_X32 FILLER_316_1112 ();
 FILLCELL_X32 FILLER_316_1144 ();
 FILLCELL_X32 FILLER_316_1176 ();
 FILLCELL_X32 FILLER_316_1208 ();
 FILLCELL_X32 FILLER_316_1240 ();
 FILLCELL_X32 FILLER_316_1272 ();
 FILLCELL_X32 FILLER_316_1304 ();
 FILLCELL_X32 FILLER_316_1336 ();
 FILLCELL_X32 FILLER_316_1368 ();
 FILLCELL_X32 FILLER_316_1400 ();
 FILLCELL_X32 FILLER_316_1432 ();
 FILLCELL_X32 FILLER_316_1464 ();
 FILLCELL_X32 FILLER_316_1496 ();
 FILLCELL_X32 FILLER_316_1528 ();
 FILLCELL_X32 FILLER_316_1560 ();
 FILLCELL_X32 FILLER_316_1592 ();
 FILLCELL_X32 FILLER_316_1624 ();
 FILLCELL_X32 FILLER_316_1656 ();
 FILLCELL_X32 FILLER_316_1688 ();
 FILLCELL_X32 FILLER_316_1720 ();
 FILLCELL_X32 FILLER_316_1752 ();
 FILLCELL_X32 FILLER_316_1784 ();
 FILLCELL_X32 FILLER_316_1816 ();
 FILLCELL_X32 FILLER_316_1848 ();
 FILLCELL_X8 FILLER_316_1880 ();
 FILLCELL_X4 FILLER_316_1888 ();
 FILLCELL_X2 FILLER_316_1892 ();
 FILLCELL_X32 FILLER_316_1895 ();
 FILLCELL_X32 FILLER_316_1927 ();
 FILLCELL_X32 FILLER_316_1959 ();
 FILLCELL_X32 FILLER_316_1991 ();
 FILLCELL_X32 FILLER_316_2023 ();
 FILLCELL_X32 FILLER_316_2055 ();
 FILLCELL_X32 FILLER_316_2087 ();
 FILLCELL_X32 FILLER_316_2119 ();
 FILLCELL_X32 FILLER_316_2151 ();
 FILLCELL_X32 FILLER_316_2183 ();
 FILLCELL_X32 FILLER_316_2215 ();
 FILLCELL_X32 FILLER_316_2247 ();
 FILLCELL_X32 FILLER_316_2279 ();
 FILLCELL_X32 FILLER_316_2311 ();
 FILLCELL_X32 FILLER_316_2343 ();
 FILLCELL_X32 FILLER_316_2375 ();
 FILLCELL_X32 FILLER_316_2407 ();
 FILLCELL_X32 FILLER_316_2439 ();
 FILLCELL_X32 FILLER_316_2471 ();
 FILLCELL_X32 FILLER_316_2503 ();
 FILLCELL_X32 FILLER_316_2535 ();
 FILLCELL_X32 FILLER_316_2567 ();
 FILLCELL_X2 FILLER_316_2599 ();
 FILLCELL_X1 FILLER_316_2601 ();
 FILLCELL_X32 FILLER_317_1 ();
 FILLCELL_X32 FILLER_317_33 ();
 FILLCELL_X32 FILLER_317_65 ();
 FILLCELL_X32 FILLER_317_97 ();
 FILLCELL_X32 FILLER_317_129 ();
 FILLCELL_X32 FILLER_317_161 ();
 FILLCELL_X32 FILLER_317_193 ();
 FILLCELL_X32 FILLER_317_225 ();
 FILLCELL_X32 FILLER_317_257 ();
 FILLCELL_X32 FILLER_317_289 ();
 FILLCELL_X32 FILLER_317_321 ();
 FILLCELL_X32 FILLER_317_353 ();
 FILLCELL_X32 FILLER_317_385 ();
 FILLCELL_X32 FILLER_317_417 ();
 FILLCELL_X32 FILLER_317_449 ();
 FILLCELL_X32 FILLER_317_481 ();
 FILLCELL_X32 FILLER_317_513 ();
 FILLCELL_X32 FILLER_317_545 ();
 FILLCELL_X32 FILLER_317_577 ();
 FILLCELL_X32 FILLER_317_609 ();
 FILLCELL_X32 FILLER_317_641 ();
 FILLCELL_X32 FILLER_317_673 ();
 FILLCELL_X32 FILLER_317_705 ();
 FILLCELL_X32 FILLER_317_737 ();
 FILLCELL_X32 FILLER_317_769 ();
 FILLCELL_X32 FILLER_317_801 ();
 FILLCELL_X32 FILLER_317_833 ();
 FILLCELL_X32 FILLER_317_865 ();
 FILLCELL_X32 FILLER_317_897 ();
 FILLCELL_X32 FILLER_317_929 ();
 FILLCELL_X32 FILLER_317_961 ();
 FILLCELL_X32 FILLER_317_993 ();
 FILLCELL_X32 FILLER_317_1025 ();
 FILLCELL_X32 FILLER_317_1057 ();
 FILLCELL_X32 FILLER_317_1089 ();
 FILLCELL_X32 FILLER_317_1121 ();
 FILLCELL_X32 FILLER_317_1153 ();
 FILLCELL_X32 FILLER_317_1185 ();
 FILLCELL_X32 FILLER_317_1217 ();
 FILLCELL_X8 FILLER_317_1249 ();
 FILLCELL_X4 FILLER_317_1257 ();
 FILLCELL_X2 FILLER_317_1261 ();
 FILLCELL_X32 FILLER_317_1264 ();
 FILLCELL_X32 FILLER_317_1296 ();
 FILLCELL_X32 FILLER_317_1328 ();
 FILLCELL_X32 FILLER_317_1360 ();
 FILLCELL_X32 FILLER_317_1392 ();
 FILLCELL_X32 FILLER_317_1424 ();
 FILLCELL_X32 FILLER_317_1456 ();
 FILLCELL_X32 FILLER_317_1488 ();
 FILLCELL_X32 FILLER_317_1520 ();
 FILLCELL_X32 FILLER_317_1552 ();
 FILLCELL_X32 FILLER_317_1584 ();
 FILLCELL_X32 FILLER_317_1616 ();
 FILLCELL_X32 FILLER_317_1648 ();
 FILLCELL_X32 FILLER_317_1680 ();
 FILLCELL_X32 FILLER_317_1712 ();
 FILLCELL_X32 FILLER_317_1744 ();
 FILLCELL_X32 FILLER_317_1776 ();
 FILLCELL_X32 FILLER_317_1808 ();
 FILLCELL_X32 FILLER_317_1840 ();
 FILLCELL_X32 FILLER_317_1872 ();
 FILLCELL_X32 FILLER_317_1904 ();
 FILLCELL_X32 FILLER_317_1936 ();
 FILLCELL_X32 FILLER_317_1968 ();
 FILLCELL_X32 FILLER_317_2000 ();
 FILLCELL_X32 FILLER_317_2032 ();
 FILLCELL_X32 FILLER_317_2064 ();
 FILLCELL_X32 FILLER_317_2096 ();
 FILLCELL_X32 FILLER_317_2128 ();
 FILLCELL_X32 FILLER_317_2160 ();
 FILLCELL_X32 FILLER_317_2192 ();
 FILLCELL_X32 FILLER_317_2224 ();
 FILLCELL_X32 FILLER_317_2256 ();
 FILLCELL_X32 FILLER_317_2288 ();
 FILLCELL_X32 FILLER_317_2320 ();
 FILLCELL_X32 FILLER_317_2352 ();
 FILLCELL_X32 FILLER_317_2384 ();
 FILLCELL_X32 FILLER_317_2416 ();
 FILLCELL_X32 FILLER_317_2448 ();
 FILLCELL_X32 FILLER_317_2480 ();
 FILLCELL_X8 FILLER_317_2512 ();
 FILLCELL_X4 FILLER_317_2520 ();
 FILLCELL_X2 FILLER_317_2524 ();
 FILLCELL_X32 FILLER_317_2527 ();
 FILLCELL_X32 FILLER_317_2559 ();
 FILLCELL_X8 FILLER_317_2591 ();
 FILLCELL_X2 FILLER_317_2599 ();
 FILLCELL_X1 FILLER_317_2601 ();
 FILLCELL_X32 FILLER_318_1 ();
 FILLCELL_X32 FILLER_318_33 ();
 FILLCELL_X32 FILLER_318_65 ();
 FILLCELL_X32 FILLER_318_97 ();
 FILLCELL_X32 FILLER_318_129 ();
 FILLCELL_X32 FILLER_318_161 ();
 FILLCELL_X32 FILLER_318_193 ();
 FILLCELL_X32 FILLER_318_225 ();
 FILLCELL_X32 FILLER_318_257 ();
 FILLCELL_X32 FILLER_318_289 ();
 FILLCELL_X32 FILLER_318_321 ();
 FILLCELL_X32 FILLER_318_353 ();
 FILLCELL_X32 FILLER_318_385 ();
 FILLCELL_X32 FILLER_318_417 ();
 FILLCELL_X32 FILLER_318_449 ();
 FILLCELL_X32 FILLER_318_481 ();
 FILLCELL_X32 FILLER_318_513 ();
 FILLCELL_X32 FILLER_318_545 ();
 FILLCELL_X32 FILLER_318_577 ();
 FILLCELL_X16 FILLER_318_609 ();
 FILLCELL_X4 FILLER_318_625 ();
 FILLCELL_X2 FILLER_318_629 ();
 FILLCELL_X32 FILLER_318_632 ();
 FILLCELL_X32 FILLER_318_664 ();
 FILLCELL_X32 FILLER_318_696 ();
 FILLCELL_X32 FILLER_318_728 ();
 FILLCELL_X32 FILLER_318_760 ();
 FILLCELL_X32 FILLER_318_792 ();
 FILLCELL_X32 FILLER_318_824 ();
 FILLCELL_X32 FILLER_318_856 ();
 FILLCELL_X32 FILLER_318_888 ();
 FILLCELL_X32 FILLER_318_920 ();
 FILLCELL_X32 FILLER_318_952 ();
 FILLCELL_X32 FILLER_318_984 ();
 FILLCELL_X32 FILLER_318_1016 ();
 FILLCELL_X32 FILLER_318_1048 ();
 FILLCELL_X32 FILLER_318_1080 ();
 FILLCELL_X32 FILLER_318_1112 ();
 FILLCELL_X32 FILLER_318_1144 ();
 FILLCELL_X32 FILLER_318_1176 ();
 FILLCELL_X32 FILLER_318_1208 ();
 FILLCELL_X32 FILLER_318_1240 ();
 FILLCELL_X32 FILLER_318_1272 ();
 FILLCELL_X32 FILLER_318_1304 ();
 FILLCELL_X32 FILLER_318_1336 ();
 FILLCELL_X32 FILLER_318_1368 ();
 FILLCELL_X32 FILLER_318_1400 ();
 FILLCELL_X32 FILLER_318_1432 ();
 FILLCELL_X32 FILLER_318_1464 ();
 FILLCELL_X32 FILLER_318_1496 ();
 FILLCELL_X32 FILLER_318_1528 ();
 FILLCELL_X32 FILLER_318_1560 ();
 FILLCELL_X32 FILLER_318_1592 ();
 FILLCELL_X32 FILLER_318_1624 ();
 FILLCELL_X32 FILLER_318_1656 ();
 FILLCELL_X32 FILLER_318_1688 ();
 FILLCELL_X32 FILLER_318_1720 ();
 FILLCELL_X32 FILLER_318_1752 ();
 FILLCELL_X32 FILLER_318_1784 ();
 FILLCELL_X32 FILLER_318_1816 ();
 FILLCELL_X32 FILLER_318_1848 ();
 FILLCELL_X8 FILLER_318_1880 ();
 FILLCELL_X4 FILLER_318_1888 ();
 FILLCELL_X2 FILLER_318_1892 ();
 FILLCELL_X32 FILLER_318_1895 ();
 FILLCELL_X32 FILLER_318_1927 ();
 FILLCELL_X32 FILLER_318_1959 ();
 FILLCELL_X32 FILLER_318_1991 ();
 FILLCELL_X32 FILLER_318_2023 ();
 FILLCELL_X32 FILLER_318_2055 ();
 FILLCELL_X32 FILLER_318_2087 ();
 FILLCELL_X32 FILLER_318_2119 ();
 FILLCELL_X32 FILLER_318_2151 ();
 FILLCELL_X32 FILLER_318_2183 ();
 FILLCELL_X32 FILLER_318_2215 ();
 FILLCELL_X32 FILLER_318_2247 ();
 FILLCELL_X32 FILLER_318_2279 ();
 FILLCELL_X32 FILLER_318_2311 ();
 FILLCELL_X32 FILLER_318_2343 ();
 FILLCELL_X32 FILLER_318_2375 ();
 FILLCELL_X32 FILLER_318_2407 ();
 FILLCELL_X32 FILLER_318_2439 ();
 FILLCELL_X32 FILLER_318_2471 ();
 FILLCELL_X32 FILLER_318_2503 ();
 FILLCELL_X32 FILLER_318_2535 ();
 FILLCELL_X32 FILLER_318_2567 ();
 FILLCELL_X2 FILLER_318_2599 ();
 FILLCELL_X1 FILLER_318_2601 ();
 FILLCELL_X32 FILLER_319_1 ();
 FILLCELL_X32 FILLER_319_33 ();
 FILLCELL_X32 FILLER_319_65 ();
 FILLCELL_X32 FILLER_319_97 ();
 FILLCELL_X32 FILLER_319_129 ();
 FILLCELL_X32 FILLER_319_161 ();
 FILLCELL_X32 FILLER_319_193 ();
 FILLCELL_X32 FILLER_319_225 ();
 FILLCELL_X32 FILLER_319_257 ();
 FILLCELL_X32 FILLER_319_289 ();
 FILLCELL_X32 FILLER_319_321 ();
 FILLCELL_X32 FILLER_319_353 ();
 FILLCELL_X32 FILLER_319_385 ();
 FILLCELL_X32 FILLER_319_417 ();
 FILLCELL_X32 FILLER_319_449 ();
 FILLCELL_X32 FILLER_319_481 ();
 FILLCELL_X32 FILLER_319_513 ();
 FILLCELL_X32 FILLER_319_545 ();
 FILLCELL_X32 FILLER_319_577 ();
 FILLCELL_X32 FILLER_319_609 ();
 FILLCELL_X32 FILLER_319_641 ();
 FILLCELL_X32 FILLER_319_673 ();
 FILLCELL_X32 FILLER_319_705 ();
 FILLCELL_X32 FILLER_319_737 ();
 FILLCELL_X32 FILLER_319_769 ();
 FILLCELL_X32 FILLER_319_801 ();
 FILLCELL_X32 FILLER_319_833 ();
 FILLCELL_X32 FILLER_319_865 ();
 FILLCELL_X32 FILLER_319_897 ();
 FILLCELL_X32 FILLER_319_929 ();
 FILLCELL_X32 FILLER_319_961 ();
 FILLCELL_X32 FILLER_319_993 ();
 FILLCELL_X32 FILLER_319_1025 ();
 FILLCELL_X32 FILLER_319_1057 ();
 FILLCELL_X32 FILLER_319_1089 ();
 FILLCELL_X32 FILLER_319_1121 ();
 FILLCELL_X32 FILLER_319_1153 ();
 FILLCELL_X32 FILLER_319_1185 ();
 FILLCELL_X32 FILLER_319_1217 ();
 FILLCELL_X8 FILLER_319_1249 ();
 FILLCELL_X4 FILLER_319_1257 ();
 FILLCELL_X2 FILLER_319_1261 ();
 FILLCELL_X32 FILLER_319_1264 ();
 FILLCELL_X32 FILLER_319_1296 ();
 FILLCELL_X32 FILLER_319_1328 ();
 FILLCELL_X32 FILLER_319_1360 ();
 FILLCELL_X32 FILLER_319_1392 ();
 FILLCELL_X32 FILLER_319_1424 ();
 FILLCELL_X32 FILLER_319_1456 ();
 FILLCELL_X32 FILLER_319_1488 ();
 FILLCELL_X32 FILLER_319_1520 ();
 FILLCELL_X32 FILLER_319_1552 ();
 FILLCELL_X32 FILLER_319_1584 ();
 FILLCELL_X32 FILLER_319_1616 ();
 FILLCELL_X32 FILLER_319_1648 ();
 FILLCELL_X32 FILLER_319_1680 ();
 FILLCELL_X32 FILLER_319_1712 ();
 FILLCELL_X32 FILLER_319_1744 ();
 FILLCELL_X32 FILLER_319_1776 ();
 FILLCELL_X32 FILLER_319_1808 ();
 FILLCELL_X32 FILLER_319_1840 ();
 FILLCELL_X32 FILLER_319_1872 ();
 FILLCELL_X32 FILLER_319_1904 ();
 FILLCELL_X32 FILLER_319_1936 ();
 FILLCELL_X32 FILLER_319_1968 ();
 FILLCELL_X32 FILLER_319_2000 ();
 FILLCELL_X32 FILLER_319_2032 ();
 FILLCELL_X32 FILLER_319_2064 ();
 FILLCELL_X32 FILLER_319_2096 ();
 FILLCELL_X32 FILLER_319_2128 ();
 FILLCELL_X32 FILLER_319_2160 ();
 FILLCELL_X32 FILLER_319_2192 ();
 FILLCELL_X32 FILLER_319_2224 ();
 FILLCELL_X32 FILLER_319_2256 ();
 FILLCELL_X32 FILLER_319_2288 ();
 FILLCELL_X32 FILLER_319_2320 ();
 FILLCELL_X32 FILLER_319_2352 ();
 FILLCELL_X32 FILLER_319_2384 ();
 FILLCELL_X32 FILLER_319_2416 ();
 FILLCELL_X32 FILLER_319_2448 ();
 FILLCELL_X32 FILLER_319_2480 ();
 FILLCELL_X8 FILLER_319_2512 ();
 FILLCELL_X4 FILLER_319_2520 ();
 FILLCELL_X2 FILLER_319_2524 ();
 FILLCELL_X32 FILLER_319_2527 ();
 FILLCELL_X32 FILLER_319_2559 ();
 FILLCELL_X8 FILLER_319_2591 ();
 FILLCELL_X2 FILLER_319_2599 ();
 FILLCELL_X1 FILLER_319_2601 ();
 FILLCELL_X32 FILLER_320_1 ();
 FILLCELL_X32 FILLER_320_33 ();
 FILLCELL_X32 FILLER_320_65 ();
 FILLCELL_X32 FILLER_320_97 ();
 FILLCELL_X32 FILLER_320_129 ();
 FILLCELL_X32 FILLER_320_161 ();
 FILLCELL_X32 FILLER_320_193 ();
 FILLCELL_X32 FILLER_320_225 ();
 FILLCELL_X32 FILLER_320_257 ();
 FILLCELL_X32 FILLER_320_289 ();
 FILLCELL_X32 FILLER_320_321 ();
 FILLCELL_X32 FILLER_320_353 ();
 FILLCELL_X32 FILLER_320_385 ();
 FILLCELL_X32 FILLER_320_417 ();
 FILLCELL_X32 FILLER_320_449 ();
 FILLCELL_X32 FILLER_320_481 ();
 FILLCELL_X32 FILLER_320_513 ();
 FILLCELL_X32 FILLER_320_545 ();
 FILLCELL_X32 FILLER_320_577 ();
 FILLCELL_X16 FILLER_320_609 ();
 FILLCELL_X4 FILLER_320_625 ();
 FILLCELL_X2 FILLER_320_629 ();
 FILLCELL_X32 FILLER_320_632 ();
 FILLCELL_X32 FILLER_320_664 ();
 FILLCELL_X32 FILLER_320_696 ();
 FILLCELL_X32 FILLER_320_728 ();
 FILLCELL_X32 FILLER_320_760 ();
 FILLCELL_X32 FILLER_320_792 ();
 FILLCELL_X32 FILLER_320_824 ();
 FILLCELL_X32 FILLER_320_856 ();
 FILLCELL_X32 FILLER_320_888 ();
 FILLCELL_X32 FILLER_320_920 ();
 FILLCELL_X32 FILLER_320_952 ();
 FILLCELL_X32 FILLER_320_984 ();
 FILLCELL_X32 FILLER_320_1016 ();
 FILLCELL_X32 FILLER_320_1048 ();
 FILLCELL_X32 FILLER_320_1080 ();
 FILLCELL_X32 FILLER_320_1112 ();
 FILLCELL_X32 FILLER_320_1144 ();
 FILLCELL_X32 FILLER_320_1176 ();
 FILLCELL_X32 FILLER_320_1208 ();
 FILLCELL_X32 FILLER_320_1240 ();
 FILLCELL_X32 FILLER_320_1272 ();
 FILLCELL_X32 FILLER_320_1304 ();
 FILLCELL_X32 FILLER_320_1336 ();
 FILLCELL_X32 FILLER_320_1368 ();
 FILLCELL_X32 FILLER_320_1400 ();
 FILLCELL_X32 FILLER_320_1432 ();
 FILLCELL_X32 FILLER_320_1464 ();
 FILLCELL_X32 FILLER_320_1496 ();
 FILLCELL_X32 FILLER_320_1528 ();
 FILLCELL_X32 FILLER_320_1560 ();
 FILLCELL_X32 FILLER_320_1592 ();
 FILLCELL_X32 FILLER_320_1624 ();
 FILLCELL_X32 FILLER_320_1656 ();
 FILLCELL_X32 FILLER_320_1688 ();
 FILLCELL_X32 FILLER_320_1720 ();
 FILLCELL_X32 FILLER_320_1752 ();
 FILLCELL_X32 FILLER_320_1784 ();
 FILLCELL_X32 FILLER_320_1816 ();
 FILLCELL_X32 FILLER_320_1848 ();
 FILLCELL_X8 FILLER_320_1880 ();
 FILLCELL_X4 FILLER_320_1888 ();
 FILLCELL_X2 FILLER_320_1892 ();
 FILLCELL_X32 FILLER_320_1895 ();
 FILLCELL_X32 FILLER_320_1927 ();
 FILLCELL_X32 FILLER_320_1959 ();
 FILLCELL_X32 FILLER_320_1991 ();
 FILLCELL_X32 FILLER_320_2023 ();
 FILLCELL_X32 FILLER_320_2055 ();
 FILLCELL_X32 FILLER_320_2087 ();
 FILLCELL_X32 FILLER_320_2119 ();
 FILLCELL_X32 FILLER_320_2151 ();
 FILLCELL_X32 FILLER_320_2183 ();
 FILLCELL_X32 FILLER_320_2215 ();
 FILLCELL_X32 FILLER_320_2247 ();
 FILLCELL_X32 FILLER_320_2279 ();
 FILLCELL_X32 FILLER_320_2311 ();
 FILLCELL_X32 FILLER_320_2343 ();
 FILLCELL_X32 FILLER_320_2375 ();
 FILLCELL_X32 FILLER_320_2407 ();
 FILLCELL_X32 FILLER_320_2439 ();
 FILLCELL_X32 FILLER_320_2471 ();
 FILLCELL_X32 FILLER_320_2503 ();
 FILLCELL_X32 FILLER_320_2535 ();
 FILLCELL_X32 FILLER_320_2567 ();
 FILLCELL_X2 FILLER_320_2599 ();
 FILLCELL_X1 FILLER_320_2601 ();
 FILLCELL_X32 FILLER_321_1 ();
 FILLCELL_X32 FILLER_321_33 ();
 FILLCELL_X32 FILLER_321_65 ();
 FILLCELL_X32 FILLER_321_97 ();
 FILLCELL_X32 FILLER_321_129 ();
 FILLCELL_X32 FILLER_321_161 ();
 FILLCELL_X32 FILLER_321_193 ();
 FILLCELL_X32 FILLER_321_225 ();
 FILLCELL_X32 FILLER_321_257 ();
 FILLCELL_X32 FILLER_321_289 ();
 FILLCELL_X32 FILLER_321_321 ();
 FILLCELL_X32 FILLER_321_353 ();
 FILLCELL_X32 FILLER_321_385 ();
 FILLCELL_X32 FILLER_321_417 ();
 FILLCELL_X32 FILLER_321_449 ();
 FILLCELL_X32 FILLER_321_481 ();
 FILLCELL_X32 FILLER_321_513 ();
 FILLCELL_X32 FILLER_321_545 ();
 FILLCELL_X32 FILLER_321_577 ();
 FILLCELL_X32 FILLER_321_609 ();
 FILLCELL_X32 FILLER_321_641 ();
 FILLCELL_X32 FILLER_321_673 ();
 FILLCELL_X32 FILLER_321_705 ();
 FILLCELL_X32 FILLER_321_737 ();
 FILLCELL_X32 FILLER_321_769 ();
 FILLCELL_X32 FILLER_321_801 ();
 FILLCELL_X32 FILLER_321_833 ();
 FILLCELL_X32 FILLER_321_865 ();
 FILLCELL_X32 FILLER_321_897 ();
 FILLCELL_X32 FILLER_321_929 ();
 FILLCELL_X32 FILLER_321_961 ();
 FILLCELL_X32 FILLER_321_993 ();
 FILLCELL_X32 FILLER_321_1025 ();
 FILLCELL_X32 FILLER_321_1057 ();
 FILLCELL_X32 FILLER_321_1089 ();
 FILLCELL_X32 FILLER_321_1121 ();
 FILLCELL_X32 FILLER_321_1153 ();
 FILLCELL_X32 FILLER_321_1185 ();
 FILLCELL_X32 FILLER_321_1217 ();
 FILLCELL_X8 FILLER_321_1249 ();
 FILLCELL_X4 FILLER_321_1257 ();
 FILLCELL_X2 FILLER_321_1261 ();
 FILLCELL_X32 FILLER_321_1264 ();
 FILLCELL_X32 FILLER_321_1296 ();
 FILLCELL_X32 FILLER_321_1328 ();
 FILLCELL_X32 FILLER_321_1360 ();
 FILLCELL_X32 FILLER_321_1392 ();
 FILLCELL_X32 FILLER_321_1424 ();
 FILLCELL_X32 FILLER_321_1456 ();
 FILLCELL_X32 FILLER_321_1488 ();
 FILLCELL_X32 FILLER_321_1520 ();
 FILLCELL_X32 FILLER_321_1552 ();
 FILLCELL_X32 FILLER_321_1584 ();
 FILLCELL_X32 FILLER_321_1616 ();
 FILLCELL_X32 FILLER_321_1648 ();
 FILLCELL_X32 FILLER_321_1680 ();
 FILLCELL_X32 FILLER_321_1712 ();
 FILLCELL_X32 FILLER_321_1744 ();
 FILLCELL_X32 FILLER_321_1776 ();
 FILLCELL_X32 FILLER_321_1808 ();
 FILLCELL_X32 FILLER_321_1840 ();
 FILLCELL_X32 FILLER_321_1872 ();
 FILLCELL_X32 FILLER_321_1904 ();
 FILLCELL_X32 FILLER_321_1936 ();
 FILLCELL_X32 FILLER_321_1968 ();
 FILLCELL_X32 FILLER_321_2000 ();
 FILLCELL_X32 FILLER_321_2032 ();
 FILLCELL_X32 FILLER_321_2064 ();
 FILLCELL_X32 FILLER_321_2096 ();
 FILLCELL_X32 FILLER_321_2128 ();
 FILLCELL_X32 FILLER_321_2160 ();
 FILLCELL_X32 FILLER_321_2192 ();
 FILLCELL_X32 FILLER_321_2224 ();
 FILLCELL_X32 FILLER_321_2256 ();
 FILLCELL_X32 FILLER_321_2288 ();
 FILLCELL_X32 FILLER_321_2320 ();
 FILLCELL_X32 FILLER_321_2352 ();
 FILLCELL_X32 FILLER_321_2384 ();
 FILLCELL_X32 FILLER_321_2416 ();
 FILLCELL_X32 FILLER_321_2448 ();
 FILLCELL_X32 FILLER_321_2480 ();
 FILLCELL_X8 FILLER_321_2512 ();
 FILLCELL_X4 FILLER_321_2520 ();
 FILLCELL_X2 FILLER_321_2524 ();
 FILLCELL_X32 FILLER_321_2527 ();
 FILLCELL_X32 FILLER_321_2559 ();
 FILLCELL_X8 FILLER_321_2591 ();
 FILLCELL_X2 FILLER_321_2599 ();
 FILLCELL_X1 FILLER_321_2601 ();
 FILLCELL_X32 FILLER_322_1 ();
 FILLCELL_X32 FILLER_322_33 ();
 FILLCELL_X32 FILLER_322_65 ();
 FILLCELL_X32 FILLER_322_97 ();
 FILLCELL_X32 FILLER_322_129 ();
 FILLCELL_X32 FILLER_322_161 ();
 FILLCELL_X32 FILLER_322_193 ();
 FILLCELL_X32 FILLER_322_225 ();
 FILLCELL_X32 FILLER_322_257 ();
 FILLCELL_X32 FILLER_322_289 ();
 FILLCELL_X32 FILLER_322_321 ();
 FILLCELL_X32 FILLER_322_353 ();
 FILLCELL_X32 FILLER_322_385 ();
 FILLCELL_X32 FILLER_322_417 ();
 FILLCELL_X32 FILLER_322_449 ();
 FILLCELL_X32 FILLER_322_481 ();
 FILLCELL_X32 FILLER_322_513 ();
 FILLCELL_X32 FILLER_322_545 ();
 FILLCELL_X32 FILLER_322_577 ();
 FILLCELL_X16 FILLER_322_609 ();
 FILLCELL_X4 FILLER_322_625 ();
 FILLCELL_X2 FILLER_322_629 ();
 FILLCELL_X32 FILLER_322_632 ();
 FILLCELL_X32 FILLER_322_664 ();
 FILLCELL_X32 FILLER_322_696 ();
 FILLCELL_X32 FILLER_322_728 ();
 FILLCELL_X32 FILLER_322_760 ();
 FILLCELL_X32 FILLER_322_792 ();
 FILLCELL_X32 FILLER_322_824 ();
 FILLCELL_X32 FILLER_322_856 ();
 FILLCELL_X32 FILLER_322_888 ();
 FILLCELL_X32 FILLER_322_920 ();
 FILLCELL_X32 FILLER_322_952 ();
 FILLCELL_X32 FILLER_322_984 ();
 FILLCELL_X32 FILLER_322_1016 ();
 FILLCELL_X32 FILLER_322_1048 ();
 FILLCELL_X32 FILLER_322_1080 ();
 FILLCELL_X32 FILLER_322_1112 ();
 FILLCELL_X32 FILLER_322_1144 ();
 FILLCELL_X32 FILLER_322_1176 ();
 FILLCELL_X32 FILLER_322_1208 ();
 FILLCELL_X32 FILLER_322_1240 ();
 FILLCELL_X32 FILLER_322_1272 ();
 FILLCELL_X32 FILLER_322_1304 ();
 FILLCELL_X32 FILLER_322_1336 ();
 FILLCELL_X32 FILLER_322_1368 ();
 FILLCELL_X32 FILLER_322_1400 ();
 FILLCELL_X32 FILLER_322_1432 ();
 FILLCELL_X32 FILLER_322_1464 ();
 FILLCELL_X32 FILLER_322_1496 ();
 FILLCELL_X32 FILLER_322_1528 ();
 FILLCELL_X32 FILLER_322_1560 ();
 FILLCELL_X32 FILLER_322_1592 ();
 FILLCELL_X32 FILLER_322_1624 ();
 FILLCELL_X32 FILLER_322_1656 ();
 FILLCELL_X32 FILLER_322_1688 ();
 FILLCELL_X32 FILLER_322_1720 ();
 FILLCELL_X32 FILLER_322_1752 ();
 FILLCELL_X32 FILLER_322_1784 ();
 FILLCELL_X32 FILLER_322_1816 ();
 FILLCELL_X32 FILLER_322_1848 ();
 FILLCELL_X8 FILLER_322_1880 ();
 FILLCELL_X4 FILLER_322_1888 ();
 FILLCELL_X2 FILLER_322_1892 ();
 FILLCELL_X32 FILLER_322_1895 ();
 FILLCELL_X32 FILLER_322_1927 ();
 FILLCELL_X32 FILLER_322_1959 ();
 FILLCELL_X32 FILLER_322_1991 ();
 FILLCELL_X32 FILLER_322_2023 ();
 FILLCELL_X32 FILLER_322_2055 ();
 FILLCELL_X32 FILLER_322_2087 ();
 FILLCELL_X32 FILLER_322_2119 ();
 FILLCELL_X32 FILLER_322_2151 ();
 FILLCELL_X32 FILLER_322_2183 ();
 FILLCELL_X32 FILLER_322_2215 ();
 FILLCELL_X32 FILLER_322_2247 ();
 FILLCELL_X32 FILLER_322_2279 ();
 FILLCELL_X32 FILLER_322_2311 ();
 FILLCELL_X32 FILLER_322_2343 ();
 FILLCELL_X32 FILLER_322_2375 ();
 FILLCELL_X32 FILLER_322_2407 ();
 FILLCELL_X32 FILLER_322_2439 ();
 FILLCELL_X32 FILLER_322_2471 ();
 FILLCELL_X32 FILLER_322_2503 ();
 FILLCELL_X32 FILLER_322_2535 ();
 FILLCELL_X32 FILLER_322_2567 ();
 FILLCELL_X2 FILLER_322_2599 ();
 FILLCELL_X1 FILLER_322_2601 ();
 FILLCELL_X32 FILLER_323_1 ();
 FILLCELL_X32 FILLER_323_33 ();
 FILLCELL_X32 FILLER_323_65 ();
 FILLCELL_X32 FILLER_323_97 ();
 FILLCELL_X32 FILLER_323_129 ();
 FILLCELL_X32 FILLER_323_161 ();
 FILLCELL_X32 FILLER_323_193 ();
 FILLCELL_X32 FILLER_323_225 ();
 FILLCELL_X32 FILLER_323_257 ();
 FILLCELL_X32 FILLER_323_289 ();
 FILLCELL_X32 FILLER_323_321 ();
 FILLCELL_X32 FILLER_323_353 ();
 FILLCELL_X32 FILLER_323_385 ();
 FILLCELL_X32 FILLER_323_417 ();
 FILLCELL_X32 FILLER_323_449 ();
 FILLCELL_X32 FILLER_323_481 ();
 FILLCELL_X32 FILLER_323_513 ();
 FILLCELL_X32 FILLER_323_545 ();
 FILLCELL_X32 FILLER_323_577 ();
 FILLCELL_X32 FILLER_323_609 ();
 FILLCELL_X32 FILLER_323_641 ();
 FILLCELL_X32 FILLER_323_673 ();
 FILLCELL_X32 FILLER_323_705 ();
 FILLCELL_X32 FILLER_323_737 ();
 FILLCELL_X32 FILLER_323_769 ();
 FILLCELL_X32 FILLER_323_801 ();
 FILLCELL_X32 FILLER_323_833 ();
 FILLCELL_X32 FILLER_323_865 ();
 FILLCELL_X32 FILLER_323_897 ();
 FILLCELL_X32 FILLER_323_929 ();
 FILLCELL_X32 FILLER_323_961 ();
 FILLCELL_X32 FILLER_323_993 ();
 FILLCELL_X32 FILLER_323_1025 ();
 FILLCELL_X32 FILLER_323_1057 ();
 FILLCELL_X32 FILLER_323_1089 ();
 FILLCELL_X32 FILLER_323_1121 ();
 FILLCELL_X32 FILLER_323_1153 ();
 FILLCELL_X32 FILLER_323_1185 ();
 FILLCELL_X32 FILLER_323_1217 ();
 FILLCELL_X8 FILLER_323_1249 ();
 FILLCELL_X4 FILLER_323_1257 ();
 FILLCELL_X2 FILLER_323_1261 ();
 FILLCELL_X32 FILLER_323_1264 ();
 FILLCELL_X32 FILLER_323_1296 ();
 FILLCELL_X32 FILLER_323_1328 ();
 FILLCELL_X32 FILLER_323_1360 ();
 FILLCELL_X32 FILLER_323_1392 ();
 FILLCELL_X32 FILLER_323_1424 ();
 FILLCELL_X32 FILLER_323_1456 ();
 FILLCELL_X32 FILLER_323_1488 ();
 FILLCELL_X32 FILLER_323_1520 ();
 FILLCELL_X32 FILLER_323_1552 ();
 FILLCELL_X32 FILLER_323_1584 ();
 FILLCELL_X32 FILLER_323_1616 ();
 FILLCELL_X32 FILLER_323_1648 ();
 FILLCELL_X32 FILLER_323_1680 ();
 FILLCELL_X32 FILLER_323_1712 ();
 FILLCELL_X32 FILLER_323_1744 ();
 FILLCELL_X32 FILLER_323_1776 ();
 FILLCELL_X32 FILLER_323_1808 ();
 FILLCELL_X32 FILLER_323_1840 ();
 FILLCELL_X32 FILLER_323_1872 ();
 FILLCELL_X32 FILLER_323_1904 ();
 FILLCELL_X32 FILLER_323_1936 ();
 FILLCELL_X32 FILLER_323_1968 ();
 FILLCELL_X32 FILLER_323_2000 ();
 FILLCELL_X32 FILLER_323_2032 ();
 FILLCELL_X32 FILLER_323_2064 ();
 FILLCELL_X32 FILLER_323_2096 ();
 FILLCELL_X32 FILLER_323_2128 ();
 FILLCELL_X32 FILLER_323_2160 ();
 FILLCELL_X32 FILLER_323_2192 ();
 FILLCELL_X32 FILLER_323_2224 ();
 FILLCELL_X32 FILLER_323_2256 ();
 FILLCELL_X32 FILLER_323_2288 ();
 FILLCELL_X32 FILLER_323_2320 ();
 FILLCELL_X32 FILLER_323_2352 ();
 FILLCELL_X32 FILLER_323_2384 ();
 FILLCELL_X32 FILLER_323_2416 ();
 FILLCELL_X32 FILLER_323_2448 ();
 FILLCELL_X32 FILLER_323_2480 ();
 FILLCELL_X8 FILLER_323_2512 ();
 FILLCELL_X4 FILLER_323_2520 ();
 FILLCELL_X2 FILLER_323_2524 ();
 FILLCELL_X32 FILLER_323_2527 ();
 FILLCELL_X32 FILLER_323_2559 ();
 FILLCELL_X8 FILLER_323_2591 ();
 FILLCELL_X2 FILLER_323_2599 ();
 FILLCELL_X1 FILLER_323_2601 ();
 FILLCELL_X32 FILLER_324_1 ();
 FILLCELL_X32 FILLER_324_33 ();
 FILLCELL_X32 FILLER_324_65 ();
 FILLCELL_X32 FILLER_324_97 ();
 FILLCELL_X32 FILLER_324_129 ();
 FILLCELL_X32 FILLER_324_161 ();
 FILLCELL_X32 FILLER_324_193 ();
 FILLCELL_X32 FILLER_324_225 ();
 FILLCELL_X32 FILLER_324_257 ();
 FILLCELL_X32 FILLER_324_289 ();
 FILLCELL_X32 FILLER_324_321 ();
 FILLCELL_X32 FILLER_324_353 ();
 FILLCELL_X32 FILLER_324_385 ();
 FILLCELL_X32 FILLER_324_417 ();
 FILLCELL_X32 FILLER_324_449 ();
 FILLCELL_X32 FILLER_324_481 ();
 FILLCELL_X32 FILLER_324_513 ();
 FILLCELL_X32 FILLER_324_545 ();
 FILLCELL_X32 FILLER_324_577 ();
 FILLCELL_X16 FILLER_324_609 ();
 FILLCELL_X4 FILLER_324_625 ();
 FILLCELL_X2 FILLER_324_629 ();
 FILLCELL_X32 FILLER_324_632 ();
 FILLCELL_X32 FILLER_324_664 ();
 FILLCELL_X32 FILLER_324_696 ();
 FILLCELL_X32 FILLER_324_728 ();
 FILLCELL_X32 FILLER_324_760 ();
 FILLCELL_X32 FILLER_324_792 ();
 FILLCELL_X32 FILLER_324_824 ();
 FILLCELL_X32 FILLER_324_856 ();
 FILLCELL_X32 FILLER_324_888 ();
 FILLCELL_X32 FILLER_324_920 ();
 FILLCELL_X32 FILLER_324_952 ();
 FILLCELL_X32 FILLER_324_984 ();
 FILLCELL_X32 FILLER_324_1016 ();
 FILLCELL_X32 FILLER_324_1048 ();
 FILLCELL_X32 FILLER_324_1080 ();
 FILLCELL_X32 FILLER_324_1112 ();
 FILLCELL_X32 FILLER_324_1144 ();
 FILLCELL_X32 FILLER_324_1176 ();
 FILLCELL_X32 FILLER_324_1208 ();
 FILLCELL_X32 FILLER_324_1240 ();
 FILLCELL_X32 FILLER_324_1272 ();
 FILLCELL_X32 FILLER_324_1304 ();
 FILLCELL_X32 FILLER_324_1336 ();
 FILLCELL_X32 FILLER_324_1368 ();
 FILLCELL_X32 FILLER_324_1400 ();
 FILLCELL_X32 FILLER_324_1432 ();
 FILLCELL_X32 FILLER_324_1464 ();
 FILLCELL_X32 FILLER_324_1496 ();
 FILLCELL_X32 FILLER_324_1528 ();
 FILLCELL_X32 FILLER_324_1560 ();
 FILLCELL_X32 FILLER_324_1592 ();
 FILLCELL_X32 FILLER_324_1624 ();
 FILLCELL_X32 FILLER_324_1656 ();
 FILLCELL_X32 FILLER_324_1688 ();
 FILLCELL_X32 FILLER_324_1720 ();
 FILLCELL_X32 FILLER_324_1752 ();
 FILLCELL_X32 FILLER_324_1784 ();
 FILLCELL_X32 FILLER_324_1816 ();
 FILLCELL_X32 FILLER_324_1848 ();
 FILLCELL_X8 FILLER_324_1880 ();
 FILLCELL_X4 FILLER_324_1888 ();
 FILLCELL_X2 FILLER_324_1892 ();
 FILLCELL_X32 FILLER_324_1895 ();
 FILLCELL_X32 FILLER_324_1927 ();
 FILLCELL_X32 FILLER_324_1959 ();
 FILLCELL_X32 FILLER_324_1991 ();
 FILLCELL_X32 FILLER_324_2023 ();
 FILLCELL_X32 FILLER_324_2055 ();
 FILLCELL_X32 FILLER_324_2087 ();
 FILLCELL_X32 FILLER_324_2119 ();
 FILLCELL_X32 FILLER_324_2151 ();
 FILLCELL_X32 FILLER_324_2183 ();
 FILLCELL_X32 FILLER_324_2215 ();
 FILLCELL_X32 FILLER_324_2247 ();
 FILLCELL_X32 FILLER_324_2279 ();
 FILLCELL_X32 FILLER_324_2311 ();
 FILLCELL_X32 FILLER_324_2343 ();
 FILLCELL_X32 FILLER_324_2375 ();
 FILLCELL_X32 FILLER_324_2407 ();
 FILLCELL_X32 FILLER_324_2439 ();
 FILLCELL_X32 FILLER_324_2471 ();
 FILLCELL_X32 FILLER_324_2503 ();
 FILLCELL_X32 FILLER_324_2535 ();
 FILLCELL_X32 FILLER_324_2567 ();
 FILLCELL_X2 FILLER_324_2599 ();
 FILLCELL_X1 FILLER_324_2601 ();
 FILLCELL_X32 FILLER_325_1 ();
 FILLCELL_X32 FILLER_325_33 ();
 FILLCELL_X32 FILLER_325_65 ();
 FILLCELL_X32 FILLER_325_97 ();
 FILLCELL_X32 FILLER_325_129 ();
 FILLCELL_X32 FILLER_325_161 ();
 FILLCELL_X32 FILLER_325_193 ();
 FILLCELL_X32 FILLER_325_225 ();
 FILLCELL_X32 FILLER_325_257 ();
 FILLCELL_X32 FILLER_325_289 ();
 FILLCELL_X32 FILLER_325_321 ();
 FILLCELL_X32 FILLER_325_353 ();
 FILLCELL_X32 FILLER_325_385 ();
 FILLCELL_X32 FILLER_325_417 ();
 FILLCELL_X32 FILLER_325_449 ();
 FILLCELL_X32 FILLER_325_481 ();
 FILLCELL_X32 FILLER_325_513 ();
 FILLCELL_X32 FILLER_325_545 ();
 FILLCELL_X32 FILLER_325_577 ();
 FILLCELL_X32 FILLER_325_609 ();
 FILLCELL_X32 FILLER_325_641 ();
 FILLCELL_X32 FILLER_325_673 ();
 FILLCELL_X32 FILLER_325_705 ();
 FILLCELL_X32 FILLER_325_737 ();
 FILLCELL_X32 FILLER_325_769 ();
 FILLCELL_X32 FILLER_325_801 ();
 FILLCELL_X32 FILLER_325_833 ();
 FILLCELL_X32 FILLER_325_865 ();
 FILLCELL_X32 FILLER_325_897 ();
 FILLCELL_X32 FILLER_325_929 ();
 FILLCELL_X32 FILLER_325_961 ();
 FILLCELL_X32 FILLER_325_993 ();
 FILLCELL_X32 FILLER_325_1025 ();
 FILLCELL_X32 FILLER_325_1057 ();
 FILLCELL_X32 FILLER_325_1089 ();
 FILLCELL_X32 FILLER_325_1121 ();
 FILLCELL_X32 FILLER_325_1153 ();
 FILLCELL_X32 FILLER_325_1185 ();
 FILLCELL_X32 FILLER_325_1217 ();
 FILLCELL_X8 FILLER_325_1249 ();
 FILLCELL_X4 FILLER_325_1257 ();
 FILLCELL_X2 FILLER_325_1261 ();
 FILLCELL_X32 FILLER_325_1264 ();
 FILLCELL_X32 FILLER_325_1296 ();
 FILLCELL_X32 FILLER_325_1328 ();
 FILLCELL_X32 FILLER_325_1360 ();
 FILLCELL_X32 FILLER_325_1392 ();
 FILLCELL_X32 FILLER_325_1424 ();
 FILLCELL_X32 FILLER_325_1456 ();
 FILLCELL_X32 FILLER_325_1488 ();
 FILLCELL_X32 FILLER_325_1520 ();
 FILLCELL_X32 FILLER_325_1552 ();
 FILLCELL_X32 FILLER_325_1584 ();
 FILLCELL_X32 FILLER_325_1616 ();
 FILLCELL_X32 FILLER_325_1648 ();
 FILLCELL_X32 FILLER_325_1680 ();
 FILLCELL_X32 FILLER_325_1712 ();
 FILLCELL_X32 FILLER_325_1744 ();
 FILLCELL_X32 FILLER_325_1776 ();
 FILLCELL_X32 FILLER_325_1808 ();
 FILLCELL_X32 FILLER_325_1840 ();
 FILLCELL_X32 FILLER_325_1872 ();
 FILLCELL_X32 FILLER_325_1904 ();
 FILLCELL_X32 FILLER_325_1936 ();
 FILLCELL_X32 FILLER_325_1968 ();
 FILLCELL_X32 FILLER_325_2000 ();
 FILLCELL_X32 FILLER_325_2032 ();
 FILLCELL_X32 FILLER_325_2064 ();
 FILLCELL_X32 FILLER_325_2096 ();
 FILLCELL_X32 FILLER_325_2128 ();
 FILLCELL_X32 FILLER_325_2160 ();
 FILLCELL_X32 FILLER_325_2192 ();
 FILLCELL_X32 FILLER_325_2224 ();
 FILLCELL_X32 FILLER_325_2256 ();
 FILLCELL_X32 FILLER_325_2288 ();
 FILLCELL_X32 FILLER_325_2320 ();
 FILLCELL_X32 FILLER_325_2352 ();
 FILLCELL_X32 FILLER_325_2384 ();
 FILLCELL_X32 FILLER_325_2416 ();
 FILLCELL_X32 FILLER_325_2448 ();
 FILLCELL_X32 FILLER_325_2480 ();
 FILLCELL_X8 FILLER_325_2512 ();
 FILLCELL_X4 FILLER_325_2520 ();
 FILLCELL_X2 FILLER_325_2524 ();
 FILLCELL_X32 FILLER_325_2527 ();
 FILLCELL_X32 FILLER_325_2559 ();
 FILLCELL_X8 FILLER_325_2591 ();
 FILLCELL_X2 FILLER_325_2599 ();
 FILLCELL_X1 FILLER_325_2601 ();
 FILLCELL_X32 FILLER_326_1 ();
 FILLCELL_X32 FILLER_326_33 ();
 FILLCELL_X32 FILLER_326_65 ();
 FILLCELL_X32 FILLER_326_97 ();
 FILLCELL_X32 FILLER_326_129 ();
 FILLCELL_X32 FILLER_326_161 ();
 FILLCELL_X32 FILLER_326_193 ();
 FILLCELL_X32 FILLER_326_225 ();
 FILLCELL_X32 FILLER_326_257 ();
 FILLCELL_X32 FILLER_326_289 ();
 FILLCELL_X32 FILLER_326_321 ();
 FILLCELL_X32 FILLER_326_353 ();
 FILLCELL_X32 FILLER_326_385 ();
 FILLCELL_X32 FILLER_326_417 ();
 FILLCELL_X32 FILLER_326_449 ();
 FILLCELL_X32 FILLER_326_481 ();
 FILLCELL_X32 FILLER_326_513 ();
 FILLCELL_X32 FILLER_326_545 ();
 FILLCELL_X32 FILLER_326_577 ();
 FILLCELL_X16 FILLER_326_609 ();
 FILLCELL_X4 FILLER_326_625 ();
 FILLCELL_X2 FILLER_326_629 ();
 FILLCELL_X32 FILLER_326_632 ();
 FILLCELL_X32 FILLER_326_664 ();
 FILLCELL_X32 FILLER_326_696 ();
 FILLCELL_X32 FILLER_326_728 ();
 FILLCELL_X32 FILLER_326_760 ();
 FILLCELL_X32 FILLER_326_792 ();
 FILLCELL_X32 FILLER_326_824 ();
 FILLCELL_X32 FILLER_326_856 ();
 FILLCELL_X32 FILLER_326_888 ();
 FILLCELL_X32 FILLER_326_920 ();
 FILLCELL_X32 FILLER_326_952 ();
 FILLCELL_X32 FILLER_326_984 ();
 FILLCELL_X32 FILLER_326_1016 ();
 FILLCELL_X32 FILLER_326_1048 ();
 FILLCELL_X32 FILLER_326_1080 ();
 FILLCELL_X32 FILLER_326_1112 ();
 FILLCELL_X32 FILLER_326_1144 ();
 FILLCELL_X32 FILLER_326_1176 ();
 FILLCELL_X32 FILLER_326_1208 ();
 FILLCELL_X32 FILLER_326_1240 ();
 FILLCELL_X32 FILLER_326_1272 ();
 FILLCELL_X32 FILLER_326_1304 ();
 FILLCELL_X32 FILLER_326_1336 ();
 FILLCELL_X32 FILLER_326_1368 ();
 FILLCELL_X32 FILLER_326_1400 ();
 FILLCELL_X32 FILLER_326_1432 ();
 FILLCELL_X32 FILLER_326_1464 ();
 FILLCELL_X32 FILLER_326_1496 ();
 FILLCELL_X32 FILLER_326_1528 ();
 FILLCELL_X32 FILLER_326_1560 ();
 FILLCELL_X32 FILLER_326_1592 ();
 FILLCELL_X32 FILLER_326_1624 ();
 FILLCELL_X32 FILLER_326_1656 ();
 FILLCELL_X32 FILLER_326_1688 ();
 FILLCELL_X32 FILLER_326_1720 ();
 FILLCELL_X32 FILLER_326_1752 ();
 FILLCELL_X32 FILLER_326_1784 ();
 FILLCELL_X32 FILLER_326_1816 ();
 FILLCELL_X32 FILLER_326_1848 ();
 FILLCELL_X8 FILLER_326_1880 ();
 FILLCELL_X4 FILLER_326_1888 ();
 FILLCELL_X2 FILLER_326_1892 ();
 FILLCELL_X32 FILLER_326_1895 ();
 FILLCELL_X32 FILLER_326_1927 ();
 FILLCELL_X32 FILLER_326_1959 ();
 FILLCELL_X32 FILLER_326_1991 ();
 FILLCELL_X32 FILLER_326_2023 ();
 FILLCELL_X32 FILLER_326_2055 ();
 FILLCELL_X32 FILLER_326_2087 ();
 FILLCELL_X32 FILLER_326_2119 ();
 FILLCELL_X32 FILLER_326_2151 ();
 FILLCELL_X32 FILLER_326_2183 ();
 FILLCELL_X32 FILLER_326_2215 ();
 FILLCELL_X32 FILLER_326_2247 ();
 FILLCELL_X32 FILLER_326_2279 ();
 FILLCELL_X32 FILLER_326_2311 ();
 FILLCELL_X32 FILLER_326_2343 ();
 FILLCELL_X32 FILLER_326_2375 ();
 FILLCELL_X32 FILLER_326_2407 ();
 FILLCELL_X32 FILLER_326_2439 ();
 FILLCELL_X32 FILLER_326_2471 ();
 FILLCELL_X32 FILLER_326_2503 ();
 FILLCELL_X32 FILLER_326_2535 ();
 FILLCELL_X32 FILLER_326_2567 ();
 FILLCELL_X2 FILLER_326_2599 ();
 FILLCELL_X1 FILLER_326_2601 ();
 FILLCELL_X32 FILLER_327_1 ();
 FILLCELL_X32 FILLER_327_33 ();
 FILLCELL_X32 FILLER_327_65 ();
 FILLCELL_X32 FILLER_327_97 ();
 FILLCELL_X32 FILLER_327_129 ();
 FILLCELL_X32 FILLER_327_161 ();
 FILLCELL_X32 FILLER_327_193 ();
 FILLCELL_X32 FILLER_327_225 ();
 FILLCELL_X32 FILLER_327_257 ();
 FILLCELL_X32 FILLER_327_289 ();
 FILLCELL_X32 FILLER_327_321 ();
 FILLCELL_X32 FILLER_327_353 ();
 FILLCELL_X32 FILLER_327_385 ();
 FILLCELL_X32 FILLER_327_417 ();
 FILLCELL_X32 FILLER_327_449 ();
 FILLCELL_X32 FILLER_327_481 ();
 FILLCELL_X32 FILLER_327_513 ();
 FILLCELL_X32 FILLER_327_545 ();
 FILLCELL_X32 FILLER_327_577 ();
 FILLCELL_X32 FILLER_327_609 ();
 FILLCELL_X32 FILLER_327_641 ();
 FILLCELL_X32 FILLER_327_673 ();
 FILLCELL_X32 FILLER_327_705 ();
 FILLCELL_X32 FILLER_327_737 ();
 FILLCELL_X32 FILLER_327_769 ();
 FILLCELL_X32 FILLER_327_801 ();
 FILLCELL_X32 FILLER_327_833 ();
 FILLCELL_X32 FILLER_327_865 ();
 FILLCELL_X32 FILLER_327_897 ();
 FILLCELL_X32 FILLER_327_929 ();
 FILLCELL_X32 FILLER_327_961 ();
 FILLCELL_X32 FILLER_327_993 ();
 FILLCELL_X32 FILLER_327_1025 ();
 FILLCELL_X32 FILLER_327_1057 ();
 FILLCELL_X32 FILLER_327_1089 ();
 FILLCELL_X32 FILLER_327_1121 ();
 FILLCELL_X32 FILLER_327_1153 ();
 FILLCELL_X32 FILLER_327_1185 ();
 FILLCELL_X32 FILLER_327_1217 ();
 FILLCELL_X8 FILLER_327_1249 ();
 FILLCELL_X4 FILLER_327_1257 ();
 FILLCELL_X2 FILLER_327_1261 ();
 FILLCELL_X32 FILLER_327_1264 ();
 FILLCELL_X32 FILLER_327_1296 ();
 FILLCELL_X32 FILLER_327_1328 ();
 FILLCELL_X32 FILLER_327_1360 ();
 FILLCELL_X32 FILLER_327_1392 ();
 FILLCELL_X32 FILLER_327_1424 ();
 FILLCELL_X32 FILLER_327_1456 ();
 FILLCELL_X32 FILLER_327_1488 ();
 FILLCELL_X32 FILLER_327_1520 ();
 FILLCELL_X32 FILLER_327_1552 ();
 FILLCELL_X32 FILLER_327_1584 ();
 FILLCELL_X32 FILLER_327_1616 ();
 FILLCELL_X32 FILLER_327_1648 ();
 FILLCELL_X32 FILLER_327_1680 ();
 FILLCELL_X32 FILLER_327_1712 ();
 FILLCELL_X32 FILLER_327_1744 ();
 FILLCELL_X32 FILLER_327_1776 ();
 FILLCELL_X32 FILLER_327_1808 ();
 FILLCELL_X32 FILLER_327_1840 ();
 FILLCELL_X32 FILLER_327_1872 ();
 FILLCELL_X32 FILLER_327_1904 ();
 FILLCELL_X32 FILLER_327_1936 ();
 FILLCELL_X32 FILLER_327_1968 ();
 FILLCELL_X32 FILLER_327_2000 ();
 FILLCELL_X32 FILLER_327_2032 ();
 FILLCELL_X32 FILLER_327_2064 ();
 FILLCELL_X32 FILLER_327_2096 ();
 FILLCELL_X32 FILLER_327_2128 ();
 FILLCELL_X32 FILLER_327_2160 ();
 FILLCELL_X32 FILLER_327_2192 ();
 FILLCELL_X32 FILLER_327_2224 ();
 FILLCELL_X32 FILLER_327_2256 ();
 FILLCELL_X32 FILLER_327_2288 ();
 FILLCELL_X32 FILLER_327_2320 ();
 FILLCELL_X32 FILLER_327_2352 ();
 FILLCELL_X32 FILLER_327_2384 ();
 FILLCELL_X32 FILLER_327_2416 ();
 FILLCELL_X32 FILLER_327_2448 ();
 FILLCELL_X32 FILLER_327_2480 ();
 FILLCELL_X8 FILLER_327_2512 ();
 FILLCELL_X4 FILLER_327_2520 ();
 FILLCELL_X2 FILLER_327_2524 ();
 FILLCELL_X32 FILLER_327_2527 ();
 FILLCELL_X32 FILLER_327_2559 ();
 FILLCELL_X8 FILLER_327_2591 ();
 FILLCELL_X2 FILLER_327_2599 ();
 FILLCELL_X1 FILLER_327_2601 ();
 FILLCELL_X32 FILLER_328_1 ();
 FILLCELL_X32 FILLER_328_33 ();
 FILLCELL_X32 FILLER_328_65 ();
 FILLCELL_X32 FILLER_328_97 ();
 FILLCELL_X32 FILLER_328_129 ();
 FILLCELL_X32 FILLER_328_161 ();
 FILLCELL_X32 FILLER_328_193 ();
 FILLCELL_X32 FILLER_328_225 ();
 FILLCELL_X32 FILLER_328_257 ();
 FILLCELL_X32 FILLER_328_289 ();
 FILLCELL_X32 FILLER_328_321 ();
 FILLCELL_X32 FILLER_328_353 ();
 FILLCELL_X32 FILLER_328_385 ();
 FILLCELL_X32 FILLER_328_417 ();
 FILLCELL_X32 FILLER_328_449 ();
 FILLCELL_X32 FILLER_328_481 ();
 FILLCELL_X32 FILLER_328_513 ();
 FILLCELL_X32 FILLER_328_545 ();
 FILLCELL_X32 FILLER_328_577 ();
 FILLCELL_X16 FILLER_328_609 ();
 FILLCELL_X4 FILLER_328_625 ();
 FILLCELL_X2 FILLER_328_629 ();
 FILLCELL_X32 FILLER_328_632 ();
 FILLCELL_X32 FILLER_328_664 ();
 FILLCELL_X32 FILLER_328_696 ();
 FILLCELL_X32 FILLER_328_728 ();
 FILLCELL_X32 FILLER_328_760 ();
 FILLCELL_X32 FILLER_328_792 ();
 FILLCELL_X32 FILLER_328_824 ();
 FILLCELL_X32 FILLER_328_856 ();
 FILLCELL_X32 FILLER_328_888 ();
 FILLCELL_X32 FILLER_328_920 ();
 FILLCELL_X32 FILLER_328_952 ();
 FILLCELL_X32 FILLER_328_984 ();
 FILLCELL_X32 FILLER_328_1016 ();
 FILLCELL_X32 FILLER_328_1048 ();
 FILLCELL_X32 FILLER_328_1080 ();
 FILLCELL_X32 FILLER_328_1112 ();
 FILLCELL_X32 FILLER_328_1144 ();
 FILLCELL_X32 FILLER_328_1176 ();
 FILLCELL_X32 FILLER_328_1208 ();
 FILLCELL_X32 FILLER_328_1240 ();
 FILLCELL_X32 FILLER_328_1272 ();
 FILLCELL_X32 FILLER_328_1304 ();
 FILLCELL_X32 FILLER_328_1336 ();
 FILLCELL_X32 FILLER_328_1368 ();
 FILLCELL_X32 FILLER_328_1400 ();
 FILLCELL_X32 FILLER_328_1432 ();
 FILLCELL_X32 FILLER_328_1464 ();
 FILLCELL_X32 FILLER_328_1496 ();
 FILLCELL_X32 FILLER_328_1528 ();
 FILLCELL_X32 FILLER_328_1560 ();
 FILLCELL_X32 FILLER_328_1592 ();
 FILLCELL_X32 FILLER_328_1624 ();
 FILLCELL_X32 FILLER_328_1656 ();
 FILLCELL_X32 FILLER_328_1688 ();
 FILLCELL_X32 FILLER_328_1720 ();
 FILLCELL_X32 FILLER_328_1752 ();
 FILLCELL_X32 FILLER_328_1784 ();
 FILLCELL_X32 FILLER_328_1816 ();
 FILLCELL_X32 FILLER_328_1848 ();
 FILLCELL_X8 FILLER_328_1880 ();
 FILLCELL_X4 FILLER_328_1888 ();
 FILLCELL_X2 FILLER_328_1892 ();
 FILLCELL_X32 FILLER_328_1895 ();
 FILLCELL_X32 FILLER_328_1927 ();
 FILLCELL_X32 FILLER_328_1959 ();
 FILLCELL_X32 FILLER_328_1991 ();
 FILLCELL_X32 FILLER_328_2023 ();
 FILLCELL_X32 FILLER_328_2055 ();
 FILLCELL_X32 FILLER_328_2087 ();
 FILLCELL_X32 FILLER_328_2119 ();
 FILLCELL_X32 FILLER_328_2151 ();
 FILLCELL_X32 FILLER_328_2183 ();
 FILLCELL_X32 FILLER_328_2215 ();
 FILLCELL_X32 FILLER_328_2247 ();
 FILLCELL_X32 FILLER_328_2279 ();
 FILLCELL_X32 FILLER_328_2311 ();
 FILLCELL_X32 FILLER_328_2343 ();
 FILLCELL_X32 FILLER_328_2375 ();
 FILLCELL_X32 FILLER_328_2407 ();
 FILLCELL_X32 FILLER_328_2439 ();
 FILLCELL_X32 FILLER_328_2471 ();
 FILLCELL_X32 FILLER_328_2503 ();
 FILLCELL_X32 FILLER_328_2535 ();
 FILLCELL_X32 FILLER_328_2567 ();
 FILLCELL_X2 FILLER_328_2599 ();
 FILLCELL_X1 FILLER_328_2601 ();
 FILLCELL_X32 FILLER_329_1 ();
 FILLCELL_X32 FILLER_329_33 ();
 FILLCELL_X32 FILLER_329_65 ();
 FILLCELL_X32 FILLER_329_97 ();
 FILLCELL_X32 FILLER_329_129 ();
 FILLCELL_X32 FILLER_329_161 ();
 FILLCELL_X32 FILLER_329_193 ();
 FILLCELL_X32 FILLER_329_225 ();
 FILLCELL_X32 FILLER_329_257 ();
 FILLCELL_X32 FILLER_329_289 ();
 FILLCELL_X32 FILLER_329_321 ();
 FILLCELL_X32 FILLER_329_353 ();
 FILLCELL_X32 FILLER_329_385 ();
 FILLCELL_X32 FILLER_329_417 ();
 FILLCELL_X32 FILLER_329_449 ();
 FILLCELL_X32 FILLER_329_481 ();
 FILLCELL_X32 FILLER_329_513 ();
 FILLCELL_X32 FILLER_329_545 ();
 FILLCELL_X32 FILLER_329_577 ();
 FILLCELL_X32 FILLER_329_609 ();
 FILLCELL_X32 FILLER_329_641 ();
 FILLCELL_X32 FILLER_329_673 ();
 FILLCELL_X32 FILLER_329_705 ();
 FILLCELL_X32 FILLER_329_737 ();
 FILLCELL_X32 FILLER_329_769 ();
 FILLCELL_X32 FILLER_329_801 ();
 FILLCELL_X32 FILLER_329_833 ();
 FILLCELL_X32 FILLER_329_865 ();
 FILLCELL_X32 FILLER_329_897 ();
 FILLCELL_X32 FILLER_329_929 ();
 FILLCELL_X32 FILLER_329_961 ();
 FILLCELL_X32 FILLER_329_993 ();
 FILLCELL_X32 FILLER_329_1025 ();
 FILLCELL_X32 FILLER_329_1057 ();
 FILLCELL_X32 FILLER_329_1089 ();
 FILLCELL_X32 FILLER_329_1121 ();
 FILLCELL_X32 FILLER_329_1153 ();
 FILLCELL_X32 FILLER_329_1185 ();
 FILLCELL_X32 FILLER_329_1217 ();
 FILLCELL_X8 FILLER_329_1249 ();
 FILLCELL_X4 FILLER_329_1257 ();
 FILLCELL_X2 FILLER_329_1261 ();
 FILLCELL_X32 FILLER_329_1264 ();
 FILLCELL_X32 FILLER_329_1296 ();
 FILLCELL_X32 FILLER_329_1328 ();
 FILLCELL_X32 FILLER_329_1360 ();
 FILLCELL_X32 FILLER_329_1392 ();
 FILLCELL_X32 FILLER_329_1424 ();
 FILLCELL_X32 FILLER_329_1456 ();
 FILLCELL_X32 FILLER_329_1488 ();
 FILLCELL_X32 FILLER_329_1520 ();
 FILLCELL_X32 FILLER_329_1552 ();
 FILLCELL_X32 FILLER_329_1584 ();
 FILLCELL_X32 FILLER_329_1616 ();
 FILLCELL_X32 FILLER_329_1648 ();
 FILLCELL_X32 FILLER_329_1680 ();
 FILLCELL_X32 FILLER_329_1712 ();
 FILLCELL_X32 FILLER_329_1744 ();
 FILLCELL_X32 FILLER_329_1776 ();
 FILLCELL_X32 FILLER_329_1808 ();
 FILLCELL_X32 FILLER_329_1840 ();
 FILLCELL_X32 FILLER_329_1872 ();
 FILLCELL_X32 FILLER_329_1904 ();
 FILLCELL_X32 FILLER_329_1936 ();
 FILLCELL_X32 FILLER_329_1968 ();
 FILLCELL_X32 FILLER_329_2000 ();
 FILLCELL_X32 FILLER_329_2032 ();
 FILLCELL_X32 FILLER_329_2064 ();
 FILLCELL_X32 FILLER_329_2096 ();
 FILLCELL_X32 FILLER_329_2128 ();
 FILLCELL_X32 FILLER_329_2160 ();
 FILLCELL_X32 FILLER_329_2192 ();
 FILLCELL_X32 FILLER_329_2224 ();
 FILLCELL_X32 FILLER_329_2256 ();
 FILLCELL_X32 FILLER_329_2288 ();
 FILLCELL_X32 FILLER_329_2320 ();
 FILLCELL_X32 FILLER_329_2352 ();
 FILLCELL_X32 FILLER_329_2384 ();
 FILLCELL_X32 FILLER_329_2416 ();
 FILLCELL_X32 FILLER_329_2448 ();
 FILLCELL_X32 FILLER_329_2480 ();
 FILLCELL_X8 FILLER_329_2512 ();
 FILLCELL_X4 FILLER_329_2520 ();
 FILLCELL_X2 FILLER_329_2524 ();
 FILLCELL_X32 FILLER_329_2527 ();
 FILLCELL_X32 FILLER_329_2559 ();
 FILLCELL_X8 FILLER_329_2591 ();
 FILLCELL_X2 FILLER_329_2599 ();
 FILLCELL_X1 FILLER_329_2601 ();
 FILLCELL_X32 FILLER_330_1 ();
 FILLCELL_X32 FILLER_330_33 ();
 FILLCELL_X32 FILLER_330_65 ();
 FILLCELL_X32 FILLER_330_97 ();
 FILLCELL_X32 FILLER_330_129 ();
 FILLCELL_X32 FILLER_330_161 ();
 FILLCELL_X32 FILLER_330_193 ();
 FILLCELL_X32 FILLER_330_225 ();
 FILLCELL_X32 FILLER_330_257 ();
 FILLCELL_X32 FILLER_330_289 ();
 FILLCELL_X32 FILLER_330_321 ();
 FILLCELL_X32 FILLER_330_353 ();
 FILLCELL_X32 FILLER_330_385 ();
 FILLCELL_X32 FILLER_330_417 ();
 FILLCELL_X32 FILLER_330_449 ();
 FILLCELL_X32 FILLER_330_481 ();
 FILLCELL_X32 FILLER_330_513 ();
 FILLCELL_X32 FILLER_330_545 ();
 FILLCELL_X32 FILLER_330_577 ();
 FILLCELL_X16 FILLER_330_609 ();
 FILLCELL_X4 FILLER_330_625 ();
 FILLCELL_X2 FILLER_330_629 ();
 FILLCELL_X32 FILLER_330_632 ();
 FILLCELL_X32 FILLER_330_664 ();
 FILLCELL_X32 FILLER_330_696 ();
 FILLCELL_X32 FILLER_330_728 ();
 FILLCELL_X32 FILLER_330_760 ();
 FILLCELL_X32 FILLER_330_792 ();
 FILLCELL_X32 FILLER_330_824 ();
 FILLCELL_X32 FILLER_330_856 ();
 FILLCELL_X32 FILLER_330_888 ();
 FILLCELL_X32 FILLER_330_920 ();
 FILLCELL_X32 FILLER_330_952 ();
 FILLCELL_X32 FILLER_330_984 ();
 FILLCELL_X32 FILLER_330_1016 ();
 FILLCELL_X32 FILLER_330_1048 ();
 FILLCELL_X32 FILLER_330_1080 ();
 FILLCELL_X32 FILLER_330_1112 ();
 FILLCELL_X32 FILLER_330_1144 ();
 FILLCELL_X32 FILLER_330_1176 ();
 FILLCELL_X32 FILLER_330_1208 ();
 FILLCELL_X32 FILLER_330_1240 ();
 FILLCELL_X32 FILLER_330_1272 ();
 FILLCELL_X32 FILLER_330_1304 ();
 FILLCELL_X32 FILLER_330_1336 ();
 FILLCELL_X32 FILLER_330_1368 ();
 FILLCELL_X32 FILLER_330_1400 ();
 FILLCELL_X32 FILLER_330_1432 ();
 FILLCELL_X32 FILLER_330_1464 ();
 FILLCELL_X32 FILLER_330_1496 ();
 FILLCELL_X32 FILLER_330_1528 ();
 FILLCELL_X32 FILLER_330_1560 ();
 FILLCELL_X32 FILLER_330_1592 ();
 FILLCELL_X32 FILLER_330_1624 ();
 FILLCELL_X32 FILLER_330_1656 ();
 FILLCELL_X32 FILLER_330_1688 ();
 FILLCELL_X32 FILLER_330_1720 ();
 FILLCELL_X32 FILLER_330_1752 ();
 FILLCELL_X32 FILLER_330_1784 ();
 FILLCELL_X32 FILLER_330_1816 ();
 FILLCELL_X32 FILLER_330_1848 ();
 FILLCELL_X8 FILLER_330_1880 ();
 FILLCELL_X4 FILLER_330_1888 ();
 FILLCELL_X2 FILLER_330_1892 ();
 FILLCELL_X32 FILLER_330_1895 ();
 FILLCELL_X32 FILLER_330_1927 ();
 FILLCELL_X32 FILLER_330_1959 ();
 FILLCELL_X32 FILLER_330_1991 ();
 FILLCELL_X32 FILLER_330_2023 ();
 FILLCELL_X32 FILLER_330_2055 ();
 FILLCELL_X32 FILLER_330_2087 ();
 FILLCELL_X32 FILLER_330_2119 ();
 FILLCELL_X32 FILLER_330_2151 ();
 FILLCELL_X32 FILLER_330_2183 ();
 FILLCELL_X32 FILLER_330_2215 ();
 FILLCELL_X32 FILLER_330_2247 ();
 FILLCELL_X32 FILLER_330_2279 ();
 FILLCELL_X32 FILLER_330_2311 ();
 FILLCELL_X32 FILLER_330_2343 ();
 FILLCELL_X32 FILLER_330_2375 ();
 FILLCELL_X32 FILLER_330_2407 ();
 FILLCELL_X32 FILLER_330_2439 ();
 FILLCELL_X32 FILLER_330_2471 ();
 FILLCELL_X32 FILLER_330_2503 ();
 FILLCELL_X32 FILLER_330_2535 ();
 FILLCELL_X32 FILLER_330_2567 ();
 FILLCELL_X2 FILLER_330_2599 ();
 FILLCELL_X1 FILLER_330_2601 ();
 FILLCELL_X32 FILLER_331_1 ();
 FILLCELL_X32 FILLER_331_33 ();
 FILLCELL_X32 FILLER_331_65 ();
 FILLCELL_X32 FILLER_331_97 ();
 FILLCELL_X32 FILLER_331_129 ();
 FILLCELL_X32 FILLER_331_161 ();
 FILLCELL_X32 FILLER_331_193 ();
 FILLCELL_X32 FILLER_331_225 ();
 FILLCELL_X32 FILLER_331_257 ();
 FILLCELL_X32 FILLER_331_289 ();
 FILLCELL_X32 FILLER_331_321 ();
 FILLCELL_X32 FILLER_331_353 ();
 FILLCELL_X32 FILLER_331_385 ();
 FILLCELL_X32 FILLER_331_417 ();
 FILLCELL_X32 FILLER_331_449 ();
 FILLCELL_X32 FILLER_331_481 ();
 FILLCELL_X32 FILLER_331_513 ();
 FILLCELL_X32 FILLER_331_545 ();
 FILLCELL_X32 FILLER_331_577 ();
 FILLCELL_X32 FILLER_331_609 ();
 FILLCELL_X32 FILLER_331_641 ();
 FILLCELL_X32 FILLER_331_673 ();
 FILLCELL_X32 FILLER_331_705 ();
 FILLCELL_X32 FILLER_331_737 ();
 FILLCELL_X32 FILLER_331_769 ();
 FILLCELL_X32 FILLER_331_801 ();
 FILLCELL_X32 FILLER_331_833 ();
 FILLCELL_X32 FILLER_331_865 ();
 FILLCELL_X32 FILLER_331_897 ();
 FILLCELL_X32 FILLER_331_929 ();
 FILLCELL_X32 FILLER_331_961 ();
 FILLCELL_X32 FILLER_331_993 ();
 FILLCELL_X32 FILLER_331_1025 ();
 FILLCELL_X32 FILLER_331_1057 ();
 FILLCELL_X32 FILLER_331_1089 ();
 FILLCELL_X32 FILLER_331_1121 ();
 FILLCELL_X32 FILLER_331_1153 ();
 FILLCELL_X32 FILLER_331_1185 ();
 FILLCELL_X32 FILLER_331_1217 ();
 FILLCELL_X8 FILLER_331_1249 ();
 FILLCELL_X4 FILLER_331_1257 ();
 FILLCELL_X2 FILLER_331_1261 ();
 FILLCELL_X32 FILLER_331_1264 ();
 FILLCELL_X32 FILLER_331_1296 ();
 FILLCELL_X32 FILLER_331_1328 ();
 FILLCELL_X32 FILLER_331_1360 ();
 FILLCELL_X32 FILLER_331_1392 ();
 FILLCELL_X32 FILLER_331_1424 ();
 FILLCELL_X32 FILLER_331_1456 ();
 FILLCELL_X32 FILLER_331_1488 ();
 FILLCELL_X32 FILLER_331_1520 ();
 FILLCELL_X32 FILLER_331_1552 ();
 FILLCELL_X32 FILLER_331_1584 ();
 FILLCELL_X32 FILLER_331_1616 ();
 FILLCELL_X32 FILLER_331_1648 ();
 FILLCELL_X32 FILLER_331_1680 ();
 FILLCELL_X32 FILLER_331_1712 ();
 FILLCELL_X32 FILLER_331_1744 ();
 FILLCELL_X32 FILLER_331_1776 ();
 FILLCELL_X32 FILLER_331_1808 ();
 FILLCELL_X32 FILLER_331_1840 ();
 FILLCELL_X32 FILLER_331_1872 ();
 FILLCELL_X32 FILLER_331_1904 ();
 FILLCELL_X32 FILLER_331_1936 ();
 FILLCELL_X32 FILLER_331_1968 ();
 FILLCELL_X32 FILLER_331_2000 ();
 FILLCELL_X32 FILLER_331_2032 ();
 FILLCELL_X32 FILLER_331_2064 ();
 FILLCELL_X32 FILLER_331_2096 ();
 FILLCELL_X32 FILLER_331_2128 ();
 FILLCELL_X32 FILLER_331_2160 ();
 FILLCELL_X32 FILLER_331_2192 ();
 FILLCELL_X32 FILLER_331_2224 ();
 FILLCELL_X32 FILLER_331_2256 ();
 FILLCELL_X32 FILLER_331_2288 ();
 FILLCELL_X32 FILLER_331_2320 ();
 FILLCELL_X32 FILLER_331_2352 ();
 FILLCELL_X32 FILLER_331_2384 ();
 FILLCELL_X32 FILLER_331_2416 ();
 FILLCELL_X32 FILLER_331_2448 ();
 FILLCELL_X32 FILLER_331_2480 ();
 FILLCELL_X8 FILLER_331_2512 ();
 FILLCELL_X4 FILLER_331_2520 ();
 FILLCELL_X2 FILLER_331_2524 ();
 FILLCELL_X32 FILLER_331_2527 ();
 FILLCELL_X32 FILLER_331_2559 ();
 FILLCELL_X8 FILLER_331_2591 ();
 FILLCELL_X2 FILLER_331_2599 ();
 FILLCELL_X1 FILLER_331_2601 ();
 FILLCELL_X32 FILLER_332_1 ();
 FILLCELL_X32 FILLER_332_33 ();
 FILLCELL_X32 FILLER_332_65 ();
 FILLCELL_X32 FILLER_332_97 ();
 FILLCELL_X32 FILLER_332_129 ();
 FILLCELL_X32 FILLER_332_161 ();
 FILLCELL_X32 FILLER_332_193 ();
 FILLCELL_X32 FILLER_332_225 ();
 FILLCELL_X32 FILLER_332_257 ();
 FILLCELL_X32 FILLER_332_289 ();
 FILLCELL_X32 FILLER_332_321 ();
 FILLCELL_X32 FILLER_332_353 ();
 FILLCELL_X32 FILLER_332_385 ();
 FILLCELL_X32 FILLER_332_417 ();
 FILLCELL_X32 FILLER_332_449 ();
 FILLCELL_X32 FILLER_332_481 ();
 FILLCELL_X32 FILLER_332_513 ();
 FILLCELL_X32 FILLER_332_545 ();
 FILLCELL_X32 FILLER_332_577 ();
 FILLCELL_X16 FILLER_332_609 ();
 FILLCELL_X4 FILLER_332_625 ();
 FILLCELL_X2 FILLER_332_629 ();
 FILLCELL_X32 FILLER_332_632 ();
 FILLCELL_X32 FILLER_332_664 ();
 FILLCELL_X32 FILLER_332_696 ();
 FILLCELL_X32 FILLER_332_728 ();
 FILLCELL_X32 FILLER_332_760 ();
 FILLCELL_X32 FILLER_332_792 ();
 FILLCELL_X32 FILLER_332_824 ();
 FILLCELL_X32 FILLER_332_856 ();
 FILLCELL_X32 FILLER_332_888 ();
 FILLCELL_X32 FILLER_332_920 ();
 FILLCELL_X32 FILLER_332_952 ();
 FILLCELL_X32 FILLER_332_984 ();
 FILLCELL_X32 FILLER_332_1016 ();
 FILLCELL_X32 FILLER_332_1048 ();
 FILLCELL_X32 FILLER_332_1080 ();
 FILLCELL_X32 FILLER_332_1112 ();
 FILLCELL_X32 FILLER_332_1144 ();
 FILLCELL_X32 FILLER_332_1176 ();
 FILLCELL_X32 FILLER_332_1208 ();
 FILLCELL_X32 FILLER_332_1240 ();
 FILLCELL_X32 FILLER_332_1272 ();
 FILLCELL_X32 FILLER_332_1304 ();
 FILLCELL_X32 FILLER_332_1336 ();
 FILLCELL_X32 FILLER_332_1368 ();
 FILLCELL_X32 FILLER_332_1400 ();
 FILLCELL_X32 FILLER_332_1432 ();
 FILLCELL_X32 FILLER_332_1464 ();
 FILLCELL_X32 FILLER_332_1496 ();
 FILLCELL_X32 FILLER_332_1528 ();
 FILLCELL_X32 FILLER_332_1560 ();
 FILLCELL_X32 FILLER_332_1592 ();
 FILLCELL_X32 FILLER_332_1624 ();
 FILLCELL_X32 FILLER_332_1656 ();
 FILLCELL_X32 FILLER_332_1688 ();
 FILLCELL_X32 FILLER_332_1720 ();
 FILLCELL_X32 FILLER_332_1752 ();
 FILLCELL_X32 FILLER_332_1784 ();
 FILLCELL_X32 FILLER_332_1816 ();
 FILLCELL_X32 FILLER_332_1848 ();
 FILLCELL_X8 FILLER_332_1880 ();
 FILLCELL_X4 FILLER_332_1888 ();
 FILLCELL_X2 FILLER_332_1892 ();
 FILLCELL_X32 FILLER_332_1895 ();
 FILLCELL_X32 FILLER_332_1927 ();
 FILLCELL_X32 FILLER_332_1959 ();
 FILLCELL_X32 FILLER_332_1991 ();
 FILLCELL_X32 FILLER_332_2023 ();
 FILLCELL_X32 FILLER_332_2055 ();
 FILLCELL_X32 FILLER_332_2087 ();
 FILLCELL_X32 FILLER_332_2119 ();
 FILLCELL_X32 FILLER_332_2151 ();
 FILLCELL_X32 FILLER_332_2183 ();
 FILLCELL_X32 FILLER_332_2215 ();
 FILLCELL_X32 FILLER_332_2247 ();
 FILLCELL_X32 FILLER_332_2279 ();
 FILLCELL_X32 FILLER_332_2311 ();
 FILLCELL_X32 FILLER_332_2343 ();
 FILLCELL_X32 FILLER_332_2375 ();
 FILLCELL_X32 FILLER_332_2407 ();
 FILLCELL_X32 FILLER_332_2439 ();
 FILLCELL_X32 FILLER_332_2471 ();
 FILLCELL_X32 FILLER_332_2503 ();
 FILLCELL_X32 FILLER_332_2535 ();
 FILLCELL_X32 FILLER_332_2567 ();
 FILLCELL_X2 FILLER_332_2599 ();
 FILLCELL_X1 FILLER_332_2601 ();
 FILLCELL_X32 FILLER_333_1 ();
 FILLCELL_X32 FILLER_333_33 ();
 FILLCELL_X32 FILLER_333_65 ();
 FILLCELL_X32 FILLER_333_97 ();
 FILLCELL_X32 FILLER_333_129 ();
 FILLCELL_X32 FILLER_333_161 ();
 FILLCELL_X32 FILLER_333_193 ();
 FILLCELL_X32 FILLER_333_225 ();
 FILLCELL_X32 FILLER_333_257 ();
 FILLCELL_X32 FILLER_333_289 ();
 FILLCELL_X32 FILLER_333_321 ();
 FILLCELL_X32 FILLER_333_353 ();
 FILLCELL_X32 FILLER_333_385 ();
 FILLCELL_X32 FILLER_333_417 ();
 FILLCELL_X32 FILLER_333_449 ();
 FILLCELL_X32 FILLER_333_481 ();
 FILLCELL_X32 FILLER_333_513 ();
 FILLCELL_X32 FILLER_333_545 ();
 FILLCELL_X32 FILLER_333_577 ();
 FILLCELL_X32 FILLER_333_609 ();
 FILLCELL_X32 FILLER_333_641 ();
 FILLCELL_X32 FILLER_333_673 ();
 FILLCELL_X32 FILLER_333_705 ();
 FILLCELL_X32 FILLER_333_737 ();
 FILLCELL_X32 FILLER_333_769 ();
 FILLCELL_X32 FILLER_333_801 ();
 FILLCELL_X32 FILLER_333_833 ();
 FILLCELL_X32 FILLER_333_865 ();
 FILLCELL_X32 FILLER_333_897 ();
 FILLCELL_X32 FILLER_333_929 ();
 FILLCELL_X32 FILLER_333_961 ();
 FILLCELL_X32 FILLER_333_993 ();
 FILLCELL_X32 FILLER_333_1025 ();
 FILLCELL_X32 FILLER_333_1057 ();
 FILLCELL_X32 FILLER_333_1089 ();
 FILLCELL_X32 FILLER_333_1121 ();
 FILLCELL_X32 FILLER_333_1153 ();
 FILLCELL_X32 FILLER_333_1185 ();
 FILLCELL_X32 FILLER_333_1217 ();
 FILLCELL_X8 FILLER_333_1249 ();
 FILLCELL_X4 FILLER_333_1257 ();
 FILLCELL_X2 FILLER_333_1261 ();
 FILLCELL_X32 FILLER_333_1264 ();
 FILLCELL_X32 FILLER_333_1296 ();
 FILLCELL_X32 FILLER_333_1328 ();
 FILLCELL_X32 FILLER_333_1360 ();
 FILLCELL_X32 FILLER_333_1392 ();
 FILLCELL_X32 FILLER_333_1424 ();
 FILLCELL_X32 FILLER_333_1456 ();
 FILLCELL_X32 FILLER_333_1488 ();
 FILLCELL_X32 FILLER_333_1520 ();
 FILLCELL_X32 FILLER_333_1552 ();
 FILLCELL_X32 FILLER_333_1584 ();
 FILLCELL_X32 FILLER_333_1616 ();
 FILLCELL_X32 FILLER_333_1648 ();
 FILLCELL_X32 FILLER_333_1680 ();
 FILLCELL_X32 FILLER_333_1712 ();
 FILLCELL_X32 FILLER_333_1744 ();
 FILLCELL_X32 FILLER_333_1776 ();
 FILLCELL_X32 FILLER_333_1808 ();
 FILLCELL_X32 FILLER_333_1840 ();
 FILLCELL_X32 FILLER_333_1872 ();
 FILLCELL_X32 FILLER_333_1904 ();
 FILLCELL_X32 FILLER_333_1936 ();
 FILLCELL_X32 FILLER_333_1968 ();
 FILLCELL_X32 FILLER_333_2000 ();
 FILLCELL_X32 FILLER_333_2032 ();
 FILLCELL_X32 FILLER_333_2064 ();
 FILLCELL_X32 FILLER_333_2096 ();
 FILLCELL_X32 FILLER_333_2128 ();
 FILLCELL_X32 FILLER_333_2160 ();
 FILLCELL_X32 FILLER_333_2192 ();
 FILLCELL_X32 FILLER_333_2224 ();
 FILLCELL_X32 FILLER_333_2256 ();
 FILLCELL_X32 FILLER_333_2288 ();
 FILLCELL_X32 FILLER_333_2320 ();
 FILLCELL_X32 FILLER_333_2352 ();
 FILLCELL_X32 FILLER_333_2384 ();
 FILLCELL_X32 FILLER_333_2416 ();
 FILLCELL_X32 FILLER_333_2448 ();
 FILLCELL_X32 FILLER_333_2480 ();
 FILLCELL_X8 FILLER_333_2512 ();
 FILLCELL_X4 FILLER_333_2520 ();
 FILLCELL_X2 FILLER_333_2524 ();
 FILLCELL_X32 FILLER_333_2527 ();
 FILLCELL_X32 FILLER_333_2559 ();
 FILLCELL_X8 FILLER_333_2591 ();
 FILLCELL_X2 FILLER_333_2599 ();
 FILLCELL_X1 FILLER_333_2601 ();
 FILLCELL_X32 FILLER_334_1 ();
 FILLCELL_X32 FILLER_334_33 ();
 FILLCELL_X32 FILLER_334_65 ();
 FILLCELL_X32 FILLER_334_97 ();
 FILLCELL_X32 FILLER_334_129 ();
 FILLCELL_X32 FILLER_334_161 ();
 FILLCELL_X32 FILLER_334_193 ();
 FILLCELL_X32 FILLER_334_225 ();
 FILLCELL_X32 FILLER_334_257 ();
 FILLCELL_X32 FILLER_334_289 ();
 FILLCELL_X32 FILLER_334_321 ();
 FILLCELL_X32 FILLER_334_353 ();
 FILLCELL_X32 FILLER_334_385 ();
 FILLCELL_X32 FILLER_334_417 ();
 FILLCELL_X32 FILLER_334_449 ();
 FILLCELL_X32 FILLER_334_481 ();
 FILLCELL_X32 FILLER_334_513 ();
 FILLCELL_X32 FILLER_334_545 ();
 FILLCELL_X32 FILLER_334_577 ();
 FILLCELL_X16 FILLER_334_609 ();
 FILLCELL_X4 FILLER_334_625 ();
 FILLCELL_X2 FILLER_334_629 ();
 FILLCELL_X32 FILLER_334_632 ();
 FILLCELL_X32 FILLER_334_664 ();
 FILLCELL_X32 FILLER_334_696 ();
 FILLCELL_X32 FILLER_334_728 ();
 FILLCELL_X32 FILLER_334_760 ();
 FILLCELL_X32 FILLER_334_792 ();
 FILLCELL_X32 FILLER_334_824 ();
 FILLCELL_X32 FILLER_334_856 ();
 FILLCELL_X32 FILLER_334_888 ();
 FILLCELL_X32 FILLER_334_920 ();
 FILLCELL_X32 FILLER_334_952 ();
 FILLCELL_X32 FILLER_334_984 ();
 FILLCELL_X32 FILLER_334_1016 ();
 FILLCELL_X32 FILLER_334_1048 ();
 FILLCELL_X32 FILLER_334_1080 ();
 FILLCELL_X32 FILLER_334_1112 ();
 FILLCELL_X32 FILLER_334_1144 ();
 FILLCELL_X32 FILLER_334_1176 ();
 FILLCELL_X32 FILLER_334_1208 ();
 FILLCELL_X32 FILLER_334_1240 ();
 FILLCELL_X32 FILLER_334_1272 ();
 FILLCELL_X32 FILLER_334_1304 ();
 FILLCELL_X32 FILLER_334_1336 ();
 FILLCELL_X32 FILLER_334_1368 ();
 FILLCELL_X32 FILLER_334_1400 ();
 FILLCELL_X32 FILLER_334_1432 ();
 FILLCELL_X32 FILLER_334_1464 ();
 FILLCELL_X32 FILLER_334_1496 ();
 FILLCELL_X32 FILLER_334_1528 ();
 FILLCELL_X32 FILLER_334_1560 ();
 FILLCELL_X32 FILLER_334_1592 ();
 FILLCELL_X32 FILLER_334_1624 ();
 FILLCELL_X32 FILLER_334_1656 ();
 FILLCELL_X32 FILLER_334_1688 ();
 FILLCELL_X32 FILLER_334_1720 ();
 FILLCELL_X32 FILLER_334_1752 ();
 FILLCELL_X32 FILLER_334_1784 ();
 FILLCELL_X32 FILLER_334_1816 ();
 FILLCELL_X32 FILLER_334_1848 ();
 FILLCELL_X8 FILLER_334_1880 ();
 FILLCELL_X4 FILLER_334_1888 ();
 FILLCELL_X2 FILLER_334_1892 ();
 FILLCELL_X32 FILLER_334_1895 ();
 FILLCELL_X32 FILLER_334_1927 ();
 FILLCELL_X32 FILLER_334_1959 ();
 FILLCELL_X32 FILLER_334_1991 ();
 FILLCELL_X32 FILLER_334_2023 ();
 FILLCELL_X32 FILLER_334_2055 ();
 FILLCELL_X32 FILLER_334_2087 ();
 FILLCELL_X32 FILLER_334_2119 ();
 FILLCELL_X32 FILLER_334_2151 ();
 FILLCELL_X32 FILLER_334_2183 ();
 FILLCELL_X32 FILLER_334_2215 ();
 FILLCELL_X32 FILLER_334_2247 ();
 FILLCELL_X32 FILLER_334_2279 ();
 FILLCELL_X32 FILLER_334_2311 ();
 FILLCELL_X32 FILLER_334_2343 ();
 FILLCELL_X32 FILLER_334_2375 ();
 FILLCELL_X32 FILLER_334_2407 ();
 FILLCELL_X32 FILLER_334_2439 ();
 FILLCELL_X32 FILLER_334_2471 ();
 FILLCELL_X32 FILLER_334_2503 ();
 FILLCELL_X32 FILLER_334_2535 ();
 FILLCELL_X32 FILLER_334_2567 ();
 FILLCELL_X2 FILLER_334_2599 ();
 FILLCELL_X1 FILLER_334_2601 ();
 FILLCELL_X32 FILLER_335_1 ();
 FILLCELL_X32 FILLER_335_33 ();
 FILLCELL_X32 FILLER_335_65 ();
 FILLCELL_X32 FILLER_335_97 ();
 FILLCELL_X32 FILLER_335_129 ();
 FILLCELL_X32 FILLER_335_161 ();
 FILLCELL_X32 FILLER_335_193 ();
 FILLCELL_X32 FILLER_335_225 ();
 FILLCELL_X32 FILLER_335_257 ();
 FILLCELL_X32 FILLER_335_289 ();
 FILLCELL_X32 FILLER_335_321 ();
 FILLCELL_X32 FILLER_335_353 ();
 FILLCELL_X32 FILLER_335_385 ();
 FILLCELL_X32 FILLER_335_417 ();
 FILLCELL_X32 FILLER_335_449 ();
 FILLCELL_X32 FILLER_335_481 ();
 FILLCELL_X32 FILLER_335_513 ();
 FILLCELL_X32 FILLER_335_545 ();
 FILLCELL_X32 FILLER_335_577 ();
 FILLCELL_X32 FILLER_335_609 ();
 FILLCELL_X32 FILLER_335_641 ();
 FILLCELL_X32 FILLER_335_673 ();
 FILLCELL_X32 FILLER_335_705 ();
 FILLCELL_X32 FILLER_335_737 ();
 FILLCELL_X32 FILLER_335_769 ();
 FILLCELL_X32 FILLER_335_801 ();
 FILLCELL_X32 FILLER_335_833 ();
 FILLCELL_X32 FILLER_335_865 ();
 FILLCELL_X32 FILLER_335_897 ();
 FILLCELL_X32 FILLER_335_929 ();
 FILLCELL_X32 FILLER_335_961 ();
 FILLCELL_X32 FILLER_335_993 ();
 FILLCELL_X32 FILLER_335_1025 ();
 FILLCELL_X32 FILLER_335_1057 ();
 FILLCELL_X32 FILLER_335_1089 ();
 FILLCELL_X32 FILLER_335_1121 ();
 FILLCELL_X32 FILLER_335_1153 ();
 FILLCELL_X32 FILLER_335_1185 ();
 FILLCELL_X32 FILLER_335_1217 ();
 FILLCELL_X8 FILLER_335_1249 ();
 FILLCELL_X4 FILLER_335_1257 ();
 FILLCELL_X2 FILLER_335_1261 ();
 FILLCELL_X32 FILLER_335_1264 ();
 FILLCELL_X32 FILLER_335_1296 ();
 FILLCELL_X32 FILLER_335_1328 ();
 FILLCELL_X32 FILLER_335_1360 ();
 FILLCELL_X32 FILLER_335_1392 ();
 FILLCELL_X32 FILLER_335_1424 ();
 FILLCELL_X32 FILLER_335_1456 ();
 FILLCELL_X32 FILLER_335_1488 ();
 FILLCELL_X32 FILLER_335_1520 ();
 FILLCELL_X32 FILLER_335_1552 ();
 FILLCELL_X32 FILLER_335_1584 ();
 FILLCELL_X32 FILLER_335_1616 ();
 FILLCELL_X32 FILLER_335_1648 ();
 FILLCELL_X32 FILLER_335_1680 ();
 FILLCELL_X32 FILLER_335_1712 ();
 FILLCELL_X32 FILLER_335_1744 ();
 FILLCELL_X32 FILLER_335_1776 ();
 FILLCELL_X32 FILLER_335_1808 ();
 FILLCELL_X32 FILLER_335_1840 ();
 FILLCELL_X32 FILLER_335_1872 ();
 FILLCELL_X32 FILLER_335_1904 ();
 FILLCELL_X32 FILLER_335_1936 ();
 FILLCELL_X32 FILLER_335_1968 ();
 FILLCELL_X32 FILLER_335_2000 ();
 FILLCELL_X32 FILLER_335_2032 ();
 FILLCELL_X32 FILLER_335_2064 ();
 FILLCELL_X32 FILLER_335_2096 ();
 FILLCELL_X32 FILLER_335_2128 ();
 FILLCELL_X32 FILLER_335_2160 ();
 FILLCELL_X32 FILLER_335_2192 ();
 FILLCELL_X32 FILLER_335_2224 ();
 FILLCELL_X32 FILLER_335_2256 ();
 FILLCELL_X32 FILLER_335_2288 ();
 FILLCELL_X32 FILLER_335_2320 ();
 FILLCELL_X32 FILLER_335_2352 ();
 FILLCELL_X32 FILLER_335_2384 ();
 FILLCELL_X32 FILLER_335_2416 ();
 FILLCELL_X32 FILLER_335_2448 ();
 FILLCELL_X32 FILLER_335_2480 ();
 FILLCELL_X8 FILLER_335_2512 ();
 FILLCELL_X4 FILLER_335_2520 ();
 FILLCELL_X2 FILLER_335_2524 ();
 FILLCELL_X32 FILLER_335_2527 ();
 FILLCELL_X32 FILLER_335_2559 ();
 FILLCELL_X8 FILLER_335_2591 ();
 FILLCELL_X2 FILLER_335_2599 ();
 FILLCELL_X1 FILLER_335_2601 ();
 FILLCELL_X32 FILLER_336_1 ();
 FILLCELL_X32 FILLER_336_33 ();
 FILLCELL_X32 FILLER_336_65 ();
 FILLCELL_X32 FILLER_336_97 ();
 FILLCELL_X32 FILLER_336_129 ();
 FILLCELL_X32 FILLER_336_161 ();
 FILLCELL_X32 FILLER_336_193 ();
 FILLCELL_X32 FILLER_336_225 ();
 FILLCELL_X32 FILLER_336_257 ();
 FILLCELL_X32 FILLER_336_289 ();
 FILLCELL_X32 FILLER_336_321 ();
 FILLCELL_X32 FILLER_336_353 ();
 FILLCELL_X32 FILLER_336_385 ();
 FILLCELL_X32 FILLER_336_417 ();
 FILLCELL_X32 FILLER_336_449 ();
 FILLCELL_X32 FILLER_336_481 ();
 FILLCELL_X32 FILLER_336_513 ();
 FILLCELL_X32 FILLER_336_545 ();
 FILLCELL_X32 FILLER_336_577 ();
 FILLCELL_X16 FILLER_336_609 ();
 FILLCELL_X4 FILLER_336_625 ();
 FILLCELL_X2 FILLER_336_629 ();
 FILLCELL_X32 FILLER_336_632 ();
 FILLCELL_X32 FILLER_336_664 ();
 FILLCELL_X32 FILLER_336_696 ();
 FILLCELL_X32 FILLER_336_728 ();
 FILLCELL_X32 FILLER_336_760 ();
 FILLCELL_X32 FILLER_336_792 ();
 FILLCELL_X32 FILLER_336_824 ();
 FILLCELL_X32 FILLER_336_856 ();
 FILLCELL_X32 FILLER_336_888 ();
 FILLCELL_X32 FILLER_336_920 ();
 FILLCELL_X32 FILLER_336_952 ();
 FILLCELL_X32 FILLER_336_984 ();
 FILLCELL_X32 FILLER_336_1016 ();
 FILLCELL_X32 FILLER_336_1048 ();
 FILLCELL_X32 FILLER_336_1080 ();
 FILLCELL_X32 FILLER_336_1112 ();
 FILLCELL_X32 FILLER_336_1144 ();
 FILLCELL_X32 FILLER_336_1176 ();
 FILLCELL_X32 FILLER_336_1208 ();
 FILLCELL_X32 FILLER_336_1240 ();
 FILLCELL_X32 FILLER_336_1272 ();
 FILLCELL_X32 FILLER_336_1304 ();
 FILLCELL_X32 FILLER_336_1336 ();
 FILLCELL_X32 FILLER_336_1368 ();
 FILLCELL_X32 FILLER_336_1400 ();
 FILLCELL_X32 FILLER_336_1432 ();
 FILLCELL_X32 FILLER_336_1464 ();
 FILLCELL_X32 FILLER_336_1496 ();
 FILLCELL_X32 FILLER_336_1528 ();
 FILLCELL_X32 FILLER_336_1560 ();
 FILLCELL_X32 FILLER_336_1592 ();
 FILLCELL_X32 FILLER_336_1624 ();
 FILLCELL_X32 FILLER_336_1656 ();
 FILLCELL_X32 FILLER_336_1688 ();
 FILLCELL_X32 FILLER_336_1720 ();
 FILLCELL_X32 FILLER_336_1752 ();
 FILLCELL_X32 FILLER_336_1784 ();
 FILLCELL_X32 FILLER_336_1816 ();
 FILLCELL_X32 FILLER_336_1848 ();
 FILLCELL_X8 FILLER_336_1880 ();
 FILLCELL_X4 FILLER_336_1888 ();
 FILLCELL_X2 FILLER_336_1892 ();
 FILLCELL_X32 FILLER_336_1895 ();
 FILLCELL_X32 FILLER_336_1927 ();
 FILLCELL_X32 FILLER_336_1959 ();
 FILLCELL_X32 FILLER_336_1991 ();
 FILLCELL_X32 FILLER_336_2023 ();
 FILLCELL_X32 FILLER_336_2055 ();
 FILLCELL_X32 FILLER_336_2087 ();
 FILLCELL_X32 FILLER_336_2119 ();
 FILLCELL_X32 FILLER_336_2151 ();
 FILLCELL_X32 FILLER_336_2183 ();
 FILLCELL_X32 FILLER_336_2215 ();
 FILLCELL_X32 FILLER_336_2247 ();
 FILLCELL_X32 FILLER_336_2279 ();
 FILLCELL_X32 FILLER_336_2311 ();
 FILLCELL_X32 FILLER_336_2343 ();
 FILLCELL_X32 FILLER_336_2375 ();
 FILLCELL_X32 FILLER_336_2407 ();
 FILLCELL_X32 FILLER_336_2439 ();
 FILLCELL_X32 FILLER_336_2471 ();
 FILLCELL_X32 FILLER_336_2503 ();
 FILLCELL_X32 FILLER_336_2535 ();
 FILLCELL_X32 FILLER_336_2567 ();
 FILLCELL_X2 FILLER_336_2599 ();
 FILLCELL_X1 FILLER_336_2601 ();
 FILLCELL_X32 FILLER_337_1 ();
 FILLCELL_X32 FILLER_337_33 ();
 FILLCELL_X32 FILLER_337_65 ();
 FILLCELL_X32 FILLER_337_97 ();
 FILLCELL_X32 FILLER_337_129 ();
 FILLCELL_X32 FILLER_337_161 ();
 FILLCELL_X32 FILLER_337_193 ();
 FILLCELL_X32 FILLER_337_225 ();
 FILLCELL_X32 FILLER_337_257 ();
 FILLCELL_X32 FILLER_337_289 ();
 FILLCELL_X32 FILLER_337_321 ();
 FILLCELL_X32 FILLER_337_353 ();
 FILLCELL_X32 FILLER_337_385 ();
 FILLCELL_X32 FILLER_337_417 ();
 FILLCELL_X32 FILLER_337_449 ();
 FILLCELL_X32 FILLER_337_481 ();
 FILLCELL_X32 FILLER_337_513 ();
 FILLCELL_X32 FILLER_337_545 ();
 FILLCELL_X32 FILLER_337_577 ();
 FILLCELL_X32 FILLER_337_609 ();
 FILLCELL_X32 FILLER_337_641 ();
 FILLCELL_X32 FILLER_337_673 ();
 FILLCELL_X32 FILLER_337_705 ();
 FILLCELL_X32 FILLER_337_737 ();
 FILLCELL_X32 FILLER_337_769 ();
 FILLCELL_X32 FILLER_337_801 ();
 FILLCELL_X32 FILLER_337_833 ();
 FILLCELL_X32 FILLER_337_865 ();
 FILLCELL_X32 FILLER_337_897 ();
 FILLCELL_X32 FILLER_337_929 ();
 FILLCELL_X32 FILLER_337_961 ();
 FILLCELL_X32 FILLER_337_993 ();
 FILLCELL_X32 FILLER_337_1025 ();
 FILLCELL_X32 FILLER_337_1057 ();
 FILLCELL_X32 FILLER_337_1089 ();
 FILLCELL_X32 FILLER_337_1121 ();
 FILLCELL_X32 FILLER_337_1153 ();
 FILLCELL_X32 FILLER_337_1185 ();
 FILLCELL_X32 FILLER_337_1217 ();
 FILLCELL_X8 FILLER_337_1249 ();
 FILLCELL_X4 FILLER_337_1257 ();
 FILLCELL_X2 FILLER_337_1261 ();
 FILLCELL_X32 FILLER_337_1264 ();
 FILLCELL_X32 FILLER_337_1296 ();
 FILLCELL_X32 FILLER_337_1328 ();
 FILLCELL_X32 FILLER_337_1360 ();
 FILLCELL_X32 FILLER_337_1392 ();
 FILLCELL_X32 FILLER_337_1424 ();
 FILLCELL_X32 FILLER_337_1456 ();
 FILLCELL_X32 FILLER_337_1488 ();
 FILLCELL_X32 FILLER_337_1520 ();
 FILLCELL_X32 FILLER_337_1552 ();
 FILLCELL_X32 FILLER_337_1584 ();
 FILLCELL_X32 FILLER_337_1616 ();
 FILLCELL_X32 FILLER_337_1648 ();
 FILLCELL_X32 FILLER_337_1680 ();
 FILLCELL_X32 FILLER_337_1712 ();
 FILLCELL_X32 FILLER_337_1744 ();
 FILLCELL_X32 FILLER_337_1776 ();
 FILLCELL_X32 FILLER_337_1808 ();
 FILLCELL_X32 FILLER_337_1840 ();
 FILLCELL_X32 FILLER_337_1872 ();
 FILLCELL_X32 FILLER_337_1904 ();
 FILLCELL_X32 FILLER_337_1936 ();
 FILLCELL_X32 FILLER_337_1968 ();
 FILLCELL_X32 FILLER_337_2000 ();
 FILLCELL_X32 FILLER_337_2032 ();
 FILLCELL_X32 FILLER_337_2064 ();
 FILLCELL_X32 FILLER_337_2096 ();
 FILLCELL_X32 FILLER_337_2128 ();
 FILLCELL_X32 FILLER_337_2160 ();
 FILLCELL_X32 FILLER_337_2192 ();
 FILLCELL_X32 FILLER_337_2224 ();
 FILLCELL_X32 FILLER_337_2256 ();
 FILLCELL_X32 FILLER_337_2288 ();
 FILLCELL_X32 FILLER_337_2320 ();
 FILLCELL_X32 FILLER_337_2352 ();
 FILLCELL_X32 FILLER_337_2384 ();
 FILLCELL_X32 FILLER_337_2416 ();
 FILLCELL_X32 FILLER_337_2448 ();
 FILLCELL_X32 FILLER_337_2480 ();
 FILLCELL_X8 FILLER_337_2512 ();
 FILLCELL_X4 FILLER_337_2520 ();
 FILLCELL_X2 FILLER_337_2524 ();
 FILLCELL_X32 FILLER_337_2527 ();
 FILLCELL_X32 FILLER_337_2559 ();
 FILLCELL_X8 FILLER_337_2591 ();
 FILLCELL_X2 FILLER_337_2599 ();
 FILLCELL_X1 FILLER_337_2601 ();
 FILLCELL_X32 FILLER_338_1 ();
 FILLCELL_X32 FILLER_338_33 ();
 FILLCELL_X32 FILLER_338_65 ();
 FILLCELL_X32 FILLER_338_97 ();
 FILLCELL_X32 FILLER_338_129 ();
 FILLCELL_X32 FILLER_338_161 ();
 FILLCELL_X32 FILLER_338_193 ();
 FILLCELL_X32 FILLER_338_225 ();
 FILLCELL_X32 FILLER_338_257 ();
 FILLCELL_X32 FILLER_338_289 ();
 FILLCELL_X32 FILLER_338_321 ();
 FILLCELL_X32 FILLER_338_353 ();
 FILLCELL_X32 FILLER_338_385 ();
 FILLCELL_X32 FILLER_338_417 ();
 FILLCELL_X32 FILLER_338_449 ();
 FILLCELL_X32 FILLER_338_481 ();
 FILLCELL_X32 FILLER_338_513 ();
 FILLCELL_X32 FILLER_338_545 ();
 FILLCELL_X32 FILLER_338_577 ();
 FILLCELL_X16 FILLER_338_609 ();
 FILLCELL_X4 FILLER_338_625 ();
 FILLCELL_X2 FILLER_338_629 ();
 FILLCELL_X32 FILLER_338_632 ();
 FILLCELL_X32 FILLER_338_664 ();
 FILLCELL_X32 FILLER_338_696 ();
 FILLCELL_X32 FILLER_338_728 ();
 FILLCELL_X32 FILLER_338_760 ();
 FILLCELL_X32 FILLER_338_792 ();
 FILLCELL_X32 FILLER_338_824 ();
 FILLCELL_X32 FILLER_338_856 ();
 FILLCELL_X32 FILLER_338_888 ();
 FILLCELL_X32 FILLER_338_920 ();
 FILLCELL_X32 FILLER_338_952 ();
 FILLCELL_X32 FILLER_338_984 ();
 FILLCELL_X32 FILLER_338_1016 ();
 FILLCELL_X32 FILLER_338_1048 ();
 FILLCELL_X32 FILLER_338_1080 ();
 FILLCELL_X32 FILLER_338_1112 ();
 FILLCELL_X32 FILLER_338_1144 ();
 FILLCELL_X32 FILLER_338_1176 ();
 FILLCELL_X32 FILLER_338_1208 ();
 FILLCELL_X32 FILLER_338_1240 ();
 FILLCELL_X32 FILLER_338_1272 ();
 FILLCELL_X32 FILLER_338_1304 ();
 FILLCELL_X32 FILLER_338_1336 ();
 FILLCELL_X32 FILLER_338_1368 ();
 FILLCELL_X32 FILLER_338_1400 ();
 FILLCELL_X32 FILLER_338_1432 ();
 FILLCELL_X32 FILLER_338_1464 ();
 FILLCELL_X32 FILLER_338_1496 ();
 FILLCELL_X32 FILLER_338_1528 ();
 FILLCELL_X32 FILLER_338_1560 ();
 FILLCELL_X32 FILLER_338_1592 ();
 FILLCELL_X32 FILLER_338_1624 ();
 FILLCELL_X32 FILLER_338_1656 ();
 FILLCELL_X32 FILLER_338_1688 ();
 FILLCELL_X32 FILLER_338_1720 ();
 FILLCELL_X32 FILLER_338_1752 ();
 FILLCELL_X32 FILLER_338_1784 ();
 FILLCELL_X32 FILLER_338_1816 ();
 FILLCELL_X32 FILLER_338_1848 ();
 FILLCELL_X8 FILLER_338_1880 ();
 FILLCELL_X4 FILLER_338_1888 ();
 FILLCELL_X2 FILLER_338_1892 ();
 FILLCELL_X32 FILLER_338_1895 ();
 FILLCELL_X32 FILLER_338_1927 ();
 FILLCELL_X32 FILLER_338_1959 ();
 FILLCELL_X32 FILLER_338_1991 ();
 FILLCELL_X32 FILLER_338_2023 ();
 FILLCELL_X32 FILLER_338_2055 ();
 FILLCELL_X32 FILLER_338_2087 ();
 FILLCELL_X32 FILLER_338_2119 ();
 FILLCELL_X32 FILLER_338_2151 ();
 FILLCELL_X32 FILLER_338_2183 ();
 FILLCELL_X32 FILLER_338_2215 ();
 FILLCELL_X32 FILLER_338_2247 ();
 FILLCELL_X32 FILLER_338_2279 ();
 FILLCELL_X32 FILLER_338_2311 ();
 FILLCELL_X32 FILLER_338_2343 ();
 FILLCELL_X32 FILLER_338_2375 ();
 FILLCELL_X32 FILLER_338_2407 ();
 FILLCELL_X32 FILLER_338_2439 ();
 FILLCELL_X32 FILLER_338_2471 ();
 FILLCELL_X32 FILLER_338_2503 ();
 FILLCELL_X32 FILLER_338_2535 ();
 FILLCELL_X32 FILLER_338_2567 ();
 FILLCELL_X2 FILLER_338_2599 ();
 FILLCELL_X1 FILLER_338_2601 ();
 FILLCELL_X32 FILLER_339_1 ();
 FILLCELL_X32 FILLER_339_33 ();
 FILLCELL_X32 FILLER_339_65 ();
 FILLCELL_X32 FILLER_339_97 ();
 FILLCELL_X32 FILLER_339_129 ();
 FILLCELL_X32 FILLER_339_161 ();
 FILLCELL_X32 FILLER_339_193 ();
 FILLCELL_X32 FILLER_339_225 ();
 FILLCELL_X32 FILLER_339_257 ();
 FILLCELL_X32 FILLER_339_289 ();
 FILLCELL_X32 FILLER_339_321 ();
 FILLCELL_X32 FILLER_339_353 ();
 FILLCELL_X32 FILLER_339_385 ();
 FILLCELL_X32 FILLER_339_417 ();
 FILLCELL_X32 FILLER_339_449 ();
 FILLCELL_X32 FILLER_339_481 ();
 FILLCELL_X32 FILLER_339_513 ();
 FILLCELL_X32 FILLER_339_545 ();
 FILLCELL_X32 FILLER_339_577 ();
 FILLCELL_X32 FILLER_339_609 ();
 FILLCELL_X32 FILLER_339_641 ();
 FILLCELL_X32 FILLER_339_673 ();
 FILLCELL_X32 FILLER_339_705 ();
 FILLCELL_X32 FILLER_339_737 ();
 FILLCELL_X32 FILLER_339_769 ();
 FILLCELL_X32 FILLER_339_801 ();
 FILLCELL_X32 FILLER_339_833 ();
 FILLCELL_X32 FILLER_339_865 ();
 FILLCELL_X32 FILLER_339_897 ();
 FILLCELL_X32 FILLER_339_929 ();
 FILLCELL_X32 FILLER_339_961 ();
 FILLCELL_X32 FILLER_339_993 ();
 FILLCELL_X32 FILLER_339_1025 ();
 FILLCELL_X32 FILLER_339_1057 ();
 FILLCELL_X32 FILLER_339_1089 ();
 FILLCELL_X32 FILLER_339_1121 ();
 FILLCELL_X32 FILLER_339_1153 ();
 FILLCELL_X32 FILLER_339_1185 ();
 FILLCELL_X32 FILLER_339_1217 ();
 FILLCELL_X8 FILLER_339_1249 ();
 FILLCELL_X4 FILLER_339_1257 ();
 FILLCELL_X2 FILLER_339_1261 ();
 FILLCELL_X32 FILLER_339_1264 ();
 FILLCELL_X32 FILLER_339_1296 ();
 FILLCELL_X32 FILLER_339_1328 ();
 FILLCELL_X32 FILLER_339_1360 ();
 FILLCELL_X32 FILLER_339_1392 ();
 FILLCELL_X32 FILLER_339_1424 ();
 FILLCELL_X32 FILLER_339_1456 ();
 FILLCELL_X32 FILLER_339_1488 ();
 FILLCELL_X32 FILLER_339_1520 ();
 FILLCELL_X32 FILLER_339_1552 ();
 FILLCELL_X32 FILLER_339_1584 ();
 FILLCELL_X32 FILLER_339_1616 ();
 FILLCELL_X32 FILLER_339_1648 ();
 FILLCELL_X32 FILLER_339_1680 ();
 FILLCELL_X32 FILLER_339_1712 ();
 FILLCELL_X32 FILLER_339_1744 ();
 FILLCELL_X32 FILLER_339_1776 ();
 FILLCELL_X32 FILLER_339_1808 ();
 FILLCELL_X32 FILLER_339_1840 ();
 FILLCELL_X32 FILLER_339_1872 ();
 FILLCELL_X32 FILLER_339_1904 ();
 FILLCELL_X32 FILLER_339_1936 ();
 FILLCELL_X32 FILLER_339_1968 ();
 FILLCELL_X32 FILLER_339_2000 ();
 FILLCELL_X32 FILLER_339_2032 ();
 FILLCELL_X32 FILLER_339_2064 ();
 FILLCELL_X32 FILLER_339_2096 ();
 FILLCELL_X32 FILLER_339_2128 ();
 FILLCELL_X32 FILLER_339_2160 ();
 FILLCELL_X32 FILLER_339_2192 ();
 FILLCELL_X32 FILLER_339_2224 ();
 FILLCELL_X32 FILLER_339_2256 ();
 FILLCELL_X32 FILLER_339_2288 ();
 FILLCELL_X32 FILLER_339_2320 ();
 FILLCELL_X32 FILLER_339_2352 ();
 FILLCELL_X32 FILLER_339_2384 ();
 FILLCELL_X32 FILLER_339_2416 ();
 FILLCELL_X32 FILLER_339_2448 ();
 FILLCELL_X32 FILLER_339_2480 ();
 FILLCELL_X8 FILLER_339_2512 ();
 FILLCELL_X4 FILLER_339_2520 ();
 FILLCELL_X2 FILLER_339_2524 ();
 FILLCELL_X32 FILLER_339_2527 ();
 FILLCELL_X32 FILLER_339_2559 ();
 FILLCELL_X8 FILLER_339_2591 ();
 FILLCELL_X2 FILLER_339_2599 ();
 FILLCELL_X1 FILLER_339_2601 ();
 FILLCELL_X32 FILLER_340_1 ();
 FILLCELL_X32 FILLER_340_33 ();
 FILLCELL_X32 FILLER_340_65 ();
 FILLCELL_X32 FILLER_340_97 ();
 FILLCELL_X32 FILLER_340_129 ();
 FILLCELL_X32 FILLER_340_161 ();
 FILLCELL_X32 FILLER_340_193 ();
 FILLCELL_X32 FILLER_340_225 ();
 FILLCELL_X32 FILLER_340_257 ();
 FILLCELL_X32 FILLER_340_289 ();
 FILLCELL_X32 FILLER_340_321 ();
 FILLCELL_X32 FILLER_340_353 ();
 FILLCELL_X32 FILLER_340_385 ();
 FILLCELL_X32 FILLER_340_417 ();
 FILLCELL_X32 FILLER_340_449 ();
 FILLCELL_X32 FILLER_340_481 ();
 FILLCELL_X32 FILLER_340_513 ();
 FILLCELL_X32 FILLER_340_545 ();
 FILLCELL_X32 FILLER_340_577 ();
 FILLCELL_X16 FILLER_340_609 ();
 FILLCELL_X4 FILLER_340_625 ();
 FILLCELL_X2 FILLER_340_629 ();
 FILLCELL_X32 FILLER_340_632 ();
 FILLCELL_X32 FILLER_340_664 ();
 FILLCELL_X32 FILLER_340_696 ();
 FILLCELL_X32 FILLER_340_728 ();
 FILLCELL_X32 FILLER_340_760 ();
 FILLCELL_X32 FILLER_340_792 ();
 FILLCELL_X32 FILLER_340_824 ();
 FILLCELL_X32 FILLER_340_856 ();
 FILLCELL_X32 FILLER_340_888 ();
 FILLCELL_X32 FILLER_340_920 ();
 FILLCELL_X32 FILLER_340_952 ();
 FILLCELL_X32 FILLER_340_984 ();
 FILLCELL_X32 FILLER_340_1016 ();
 FILLCELL_X32 FILLER_340_1048 ();
 FILLCELL_X32 FILLER_340_1080 ();
 FILLCELL_X32 FILLER_340_1112 ();
 FILLCELL_X32 FILLER_340_1144 ();
 FILLCELL_X32 FILLER_340_1176 ();
 FILLCELL_X32 FILLER_340_1208 ();
 FILLCELL_X32 FILLER_340_1240 ();
 FILLCELL_X32 FILLER_340_1272 ();
 FILLCELL_X32 FILLER_340_1304 ();
 FILLCELL_X32 FILLER_340_1336 ();
 FILLCELL_X32 FILLER_340_1368 ();
 FILLCELL_X32 FILLER_340_1400 ();
 FILLCELL_X32 FILLER_340_1432 ();
 FILLCELL_X32 FILLER_340_1464 ();
 FILLCELL_X32 FILLER_340_1496 ();
 FILLCELL_X32 FILLER_340_1528 ();
 FILLCELL_X32 FILLER_340_1560 ();
 FILLCELL_X32 FILLER_340_1592 ();
 FILLCELL_X32 FILLER_340_1624 ();
 FILLCELL_X32 FILLER_340_1656 ();
 FILLCELL_X32 FILLER_340_1688 ();
 FILLCELL_X32 FILLER_340_1720 ();
 FILLCELL_X32 FILLER_340_1752 ();
 FILLCELL_X32 FILLER_340_1784 ();
 FILLCELL_X32 FILLER_340_1816 ();
 FILLCELL_X32 FILLER_340_1848 ();
 FILLCELL_X8 FILLER_340_1880 ();
 FILLCELL_X4 FILLER_340_1888 ();
 FILLCELL_X2 FILLER_340_1892 ();
 FILLCELL_X32 FILLER_340_1895 ();
 FILLCELL_X32 FILLER_340_1927 ();
 FILLCELL_X32 FILLER_340_1959 ();
 FILLCELL_X32 FILLER_340_1991 ();
 FILLCELL_X32 FILLER_340_2023 ();
 FILLCELL_X32 FILLER_340_2055 ();
 FILLCELL_X32 FILLER_340_2087 ();
 FILLCELL_X32 FILLER_340_2119 ();
 FILLCELL_X32 FILLER_340_2151 ();
 FILLCELL_X32 FILLER_340_2183 ();
 FILLCELL_X32 FILLER_340_2215 ();
 FILLCELL_X32 FILLER_340_2247 ();
 FILLCELL_X32 FILLER_340_2279 ();
 FILLCELL_X32 FILLER_340_2311 ();
 FILLCELL_X32 FILLER_340_2343 ();
 FILLCELL_X32 FILLER_340_2375 ();
 FILLCELL_X32 FILLER_340_2407 ();
 FILLCELL_X32 FILLER_340_2439 ();
 FILLCELL_X32 FILLER_340_2471 ();
 FILLCELL_X32 FILLER_340_2503 ();
 FILLCELL_X32 FILLER_340_2535 ();
 FILLCELL_X32 FILLER_340_2567 ();
 FILLCELL_X2 FILLER_340_2599 ();
 FILLCELL_X1 FILLER_340_2601 ();
 FILLCELL_X32 FILLER_341_1 ();
 FILLCELL_X32 FILLER_341_33 ();
 FILLCELL_X32 FILLER_341_65 ();
 FILLCELL_X32 FILLER_341_97 ();
 FILLCELL_X32 FILLER_341_129 ();
 FILLCELL_X32 FILLER_341_161 ();
 FILLCELL_X32 FILLER_341_193 ();
 FILLCELL_X32 FILLER_341_225 ();
 FILLCELL_X32 FILLER_341_257 ();
 FILLCELL_X32 FILLER_341_289 ();
 FILLCELL_X32 FILLER_341_321 ();
 FILLCELL_X32 FILLER_341_353 ();
 FILLCELL_X32 FILLER_341_385 ();
 FILLCELL_X32 FILLER_341_417 ();
 FILLCELL_X32 FILLER_341_449 ();
 FILLCELL_X32 FILLER_341_481 ();
 FILLCELL_X32 FILLER_341_513 ();
 FILLCELL_X32 FILLER_341_545 ();
 FILLCELL_X32 FILLER_341_577 ();
 FILLCELL_X32 FILLER_341_609 ();
 FILLCELL_X32 FILLER_341_641 ();
 FILLCELL_X32 FILLER_341_673 ();
 FILLCELL_X32 FILLER_341_705 ();
 FILLCELL_X32 FILLER_341_737 ();
 FILLCELL_X32 FILLER_341_769 ();
 FILLCELL_X32 FILLER_341_801 ();
 FILLCELL_X32 FILLER_341_833 ();
 FILLCELL_X32 FILLER_341_865 ();
 FILLCELL_X32 FILLER_341_897 ();
 FILLCELL_X32 FILLER_341_929 ();
 FILLCELL_X32 FILLER_341_961 ();
 FILLCELL_X32 FILLER_341_993 ();
 FILLCELL_X32 FILLER_341_1025 ();
 FILLCELL_X32 FILLER_341_1057 ();
 FILLCELL_X32 FILLER_341_1089 ();
 FILLCELL_X32 FILLER_341_1121 ();
 FILLCELL_X32 FILLER_341_1153 ();
 FILLCELL_X32 FILLER_341_1185 ();
 FILLCELL_X32 FILLER_341_1217 ();
 FILLCELL_X8 FILLER_341_1249 ();
 FILLCELL_X4 FILLER_341_1257 ();
 FILLCELL_X2 FILLER_341_1261 ();
 FILLCELL_X32 FILLER_341_1264 ();
 FILLCELL_X32 FILLER_341_1296 ();
 FILLCELL_X32 FILLER_341_1328 ();
 FILLCELL_X32 FILLER_341_1360 ();
 FILLCELL_X32 FILLER_341_1392 ();
 FILLCELL_X32 FILLER_341_1424 ();
 FILLCELL_X32 FILLER_341_1456 ();
 FILLCELL_X32 FILLER_341_1488 ();
 FILLCELL_X32 FILLER_341_1520 ();
 FILLCELL_X32 FILLER_341_1552 ();
 FILLCELL_X32 FILLER_341_1584 ();
 FILLCELL_X32 FILLER_341_1616 ();
 FILLCELL_X32 FILLER_341_1648 ();
 FILLCELL_X32 FILLER_341_1680 ();
 FILLCELL_X32 FILLER_341_1712 ();
 FILLCELL_X32 FILLER_341_1744 ();
 FILLCELL_X32 FILLER_341_1776 ();
 FILLCELL_X32 FILLER_341_1808 ();
 FILLCELL_X32 FILLER_341_1840 ();
 FILLCELL_X32 FILLER_341_1872 ();
 FILLCELL_X32 FILLER_341_1904 ();
 FILLCELL_X32 FILLER_341_1936 ();
 FILLCELL_X32 FILLER_341_1968 ();
 FILLCELL_X32 FILLER_341_2000 ();
 FILLCELL_X32 FILLER_341_2032 ();
 FILLCELL_X32 FILLER_341_2064 ();
 FILLCELL_X32 FILLER_341_2096 ();
 FILLCELL_X32 FILLER_341_2128 ();
 FILLCELL_X32 FILLER_341_2160 ();
 FILLCELL_X32 FILLER_341_2192 ();
 FILLCELL_X32 FILLER_341_2224 ();
 FILLCELL_X32 FILLER_341_2256 ();
 FILLCELL_X32 FILLER_341_2288 ();
 FILLCELL_X32 FILLER_341_2320 ();
 FILLCELL_X32 FILLER_341_2352 ();
 FILLCELL_X32 FILLER_341_2384 ();
 FILLCELL_X32 FILLER_341_2416 ();
 FILLCELL_X32 FILLER_341_2448 ();
 FILLCELL_X32 FILLER_341_2480 ();
 FILLCELL_X8 FILLER_341_2512 ();
 FILLCELL_X4 FILLER_341_2520 ();
 FILLCELL_X2 FILLER_341_2524 ();
 FILLCELL_X32 FILLER_341_2527 ();
 FILLCELL_X32 FILLER_341_2559 ();
 FILLCELL_X8 FILLER_341_2591 ();
 FILLCELL_X2 FILLER_341_2599 ();
 FILLCELL_X1 FILLER_341_2601 ();
 FILLCELL_X32 FILLER_342_1 ();
 FILLCELL_X32 FILLER_342_33 ();
 FILLCELL_X32 FILLER_342_65 ();
 FILLCELL_X32 FILLER_342_97 ();
 FILLCELL_X32 FILLER_342_129 ();
 FILLCELL_X32 FILLER_342_161 ();
 FILLCELL_X32 FILLER_342_193 ();
 FILLCELL_X32 FILLER_342_225 ();
 FILLCELL_X32 FILLER_342_257 ();
 FILLCELL_X32 FILLER_342_289 ();
 FILLCELL_X32 FILLER_342_321 ();
 FILLCELL_X32 FILLER_342_353 ();
 FILLCELL_X32 FILLER_342_385 ();
 FILLCELL_X32 FILLER_342_417 ();
 FILLCELL_X32 FILLER_342_449 ();
 FILLCELL_X32 FILLER_342_481 ();
 FILLCELL_X32 FILLER_342_513 ();
 FILLCELL_X32 FILLER_342_545 ();
 FILLCELL_X32 FILLER_342_577 ();
 FILLCELL_X16 FILLER_342_609 ();
 FILLCELL_X4 FILLER_342_625 ();
 FILLCELL_X2 FILLER_342_629 ();
 FILLCELL_X32 FILLER_342_632 ();
 FILLCELL_X32 FILLER_342_664 ();
 FILLCELL_X32 FILLER_342_696 ();
 FILLCELL_X32 FILLER_342_728 ();
 FILLCELL_X32 FILLER_342_760 ();
 FILLCELL_X32 FILLER_342_792 ();
 FILLCELL_X32 FILLER_342_824 ();
 FILLCELL_X32 FILLER_342_856 ();
 FILLCELL_X32 FILLER_342_888 ();
 FILLCELL_X32 FILLER_342_920 ();
 FILLCELL_X32 FILLER_342_952 ();
 FILLCELL_X32 FILLER_342_984 ();
 FILLCELL_X32 FILLER_342_1016 ();
 FILLCELL_X32 FILLER_342_1048 ();
 FILLCELL_X32 FILLER_342_1080 ();
 FILLCELL_X32 FILLER_342_1112 ();
 FILLCELL_X32 FILLER_342_1144 ();
 FILLCELL_X32 FILLER_342_1176 ();
 FILLCELL_X32 FILLER_342_1208 ();
 FILLCELL_X32 FILLER_342_1240 ();
 FILLCELL_X32 FILLER_342_1272 ();
 FILLCELL_X32 FILLER_342_1304 ();
 FILLCELL_X32 FILLER_342_1336 ();
 FILLCELL_X32 FILLER_342_1368 ();
 FILLCELL_X32 FILLER_342_1400 ();
 FILLCELL_X32 FILLER_342_1432 ();
 FILLCELL_X32 FILLER_342_1464 ();
 FILLCELL_X32 FILLER_342_1496 ();
 FILLCELL_X32 FILLER_342_1528 ();
 FILLCELL_X32 FILLER_342_1560 ();
 FILLCELL_X32 FILLER_342_1592 ();
 FILLCELL_X32 FILLER_342_1624 ();
 FILLCELL_X32 FILLER_342_1656 ();
 FILLCELL_X32 FILLER_342_1688 ();
 FILLCELL_X32 FILLER_342_1720 ();
 FILLCELL_X32 FILLER_342_1752 ();
 FILLCELL_X32 FILLER_342_1784 ();
 FILLCELL_X32 FILLER_342_1816 ();
 FILLCELL_X32 FILLER_342_1848 ();
 FILLCELL_X8 FILLER_342_1880 ();
 FILLCELL_X4 FILLER_342_1888 ();
 FILLCELL_X2 FILLER_342_1892 ();
 FILLCELL_X32 FILLER_342_1895 ();
 FILLCELL_X32 FILLER_342_1927 ();
 FILLCELL_X32 FILLER_342_1959 ();
 FILLCELL_X32 FILLER_342_1991 ();
 FILLCELL_X32 FILLER_342_2023 ();
 FILLCELL_X32 FILLER_342_2055 ();
 FILLCELL_X32 FILLER_342_2087 ();
 FILLCELL_X32 FILLER_342_2119 ();
 FILLCELL_X32 FILLER_342_2151 ();
 FILLCELL_X32 FILLER_342_2183 ();
 FILLCELL_X32 FILLER_342_2215 ();
 FILLCELL_X32 FILLER_342_2247 ();
 FILLCELL_X32 FILLER_342_2279 ();
 FILLCELL_X32 FILLER_342_2311 ();
 FILLCELL_X32 FILLER_342_2343 ();
 FILLCELL_X32 FILLER_342_2375 ();
 FILLCELL_X32 FILLER_342_2407 ();
 FILLCELL_X32 FILLER_342_2439 ();
 FILLCELL_X32 FILLER_342_2471 ();
 FILLCELL_X32 FILLER_342_2503 ();
 FILLCELL_X32 FILLER_342_2535 ();
 FILLCELL_X32 FILLER_342_2567 ();
 FILLCELL_X2 FILLER_342_2599 ();
 FILLCELL_X1 FILLER_342_2601 ();
 FILLCELL_X32 FILLER_343_1 ();
 FILLCELL_X32 FILLER_343_33 ();
 FILLCELL_X32 FILLER_343_65 ();
 FILLCELL_X32 FILLER_343_97 ();
 FILLCELL_X32 FILLER_343_129 ();
 FILLCELL_X32 FILLER_343_161 ();
 FILLCELL_X32 FILLER_343_193 ();
 FILLCELL_X32 FILLER_343_225 ();
 FILLCELL_X32 FILLER_343_257 ();
 FILLCELL_X32 FILLER_343_289 ();
 FILLCELL_X32 FILLER_343_321 ();
 FILLCELL_X32 FILLER_343_353 ();
 FILLCELL_X32 FILLER_343_385 ();
 FILLCELL_X32 FILLER_343_417 ();
 FILLCELL_X32 FILLER_343_449 ();
 FILLCELL_X32 FILLER_343_481 ();
 FILLCELL_X32 FILLER_343_513 ();
 FILLCELL_X32 FILLER_343_545 ();
 FILLCELL_X32 FILLER_343_577 ();
 FILLCELL_X32 FILLER_343_609 ();
 FILLCELL_X32 FILLER_343_641 ();
 FILLCELL_X32 FILLER_343_673 ();
 FILLCELL_X32 FILLER_343_705 ();
 FILLCELL_X32 FILLER_343_737 ();
 FILLCELL_X32 FILLER_343_769 ();
 FILLCELL_X32 FILLER_343_801 ();
 FILLCELL_X32 FILLER_343_833 ();
 FILLCELL_X32 FILLER_343_865 ();
 FILLCELL_X32 FILLER_343_897 ();
 FILLCELL_X32 FILLER_343_929 ();
 FILLCELL_X32 FILLER_343_961 ();
 FILLCELL_X32 FILLER_343_993 ();
 FILLCELL_X32 FILLER_343_1025 ();
 FILLCELL_X32 FILLER_343_1057 ();
 FILLCELL_X32 FILLER_343_1089 ();
 FILLCELL_X32 FILLER_343_1121 ();
 FILLCELL_X32 FILLER_343_1153 ();
 FILLCELL_X32 FILLER_343_1185 ();
 FILLCELL_X32 FILLER_343_1217 ();
 FILLCELL_X8 FILLER_343_1249 ();
 FILLCELL_X4 FILLER_343_1257 ();
 FILLCELL_X2 FILLER_343_1261 ();
 FILLCELL_X32 FILLER_343_1264 ();
 FILLCELL_X32 FILLER_343_1296 ();
 FILLCELL_X32 FILLER_343_1328 ();
 FILLCELL_X32 FILLER_343_1360 ();
 FILLCELL_X32 FILLER_343_1392 ();
 FILLCELL_X32 FILLER_343_1424 ();
 FILLCELL_X32 FILLER_343_1456 ();
 FILLCELL_X32 FILLER_343_1488 ();
 FILLCELL_X32 FILLER_343_1520 ();
 FILLCELL_X32 FILLER_343_1552 ();
 FILLCELL_X32 FILLER_343_1584 ();
 FILLCELL_X32 FILLER_343_1616 ();
 FILLCELL_X32 FILLER_343_1648 ();
 FILLCELL_X32 FILLER_343_1680 ();
 FILLCELL_X32 FILLER_343_1712 ();
 FILLCELL_X32 FILLER_343_1744 ();
 FILLCELL_X32 FILLER_343_1776 ();
 FILLCELL_X32 FILLER_343_1808 ();
 FILLCELL_X32 FILLER_343_1840 ();
 FILLCELL_X32 FILLER_343_1872 ();
 FILLCELL_X32 FILLER_343_1904 ();
 FILLCELL_X32 FILLER_343_1936 ();
 FILLCELL_X32 FILLER_343_1968 ();
 FILLCELL_X32 FILLER_343_2000 ();
 FILLCELL_X32 FILLER_343_2032 ();
 FILLCELL_X32 FILLER_343_2064 ();
 FILLCELL_X32 FILLER_343_2096 ();
 FILLCELL_X32 FILLER_343_2128 ();
 FILLCELL_X32 FILLER_343_2160 ();
 FILLCELL_X32 FILLER_343_2192 ();
 FILLCELL_X32 FILLER_343_2224 ();
 FILLCELL_X32 FILLER_343_2256 ();
 FILLCELL_X32 FILLER_343_2288 ();
 FILLCELL_X32 FILLER_343_2320 ();
 FILLCELL_X32 FILLER_343_2352 ();
 FILLCELL_X32 FILLER_343_2384 ();
 FILLCELL_X32 FILLER_343_2416 ();
 FILLCELL_X32 FILLER_343_2448 ();
 FILLCELL_X32 FILLER_343_2480 ();
 FILLCELL_X8 FILLER_343_2512 ();
 FILLCELL_X4 FILLER_343_2520 ();
 FILLCELL_X2 FILLER_343_2524 ();
 FILLCELL_X32 FILLER_343_2527 ();
 FILLCELL_X32 FILLER_343_2559 ();
 FILLCELL_X8 FILLER_343_2591 ();
 FILLCELL_X2 FILLER_343_2599 ();
 FILLCELL_X1 FILLER_343_2601 ();
 FILLCELL_X32 FILLER_344_1 ();
 FILLCELL_X32 FILLER_344_33 ();
 FILLCELL_X32 FILLER_344_65 ();
 FILLCELL_X32 FILLER_344_97 ();
 FILLCELL_X32 FILLER_344_129 ();
 FILLCELL_X32 FILLER_344_161 ();
 FILLCELL_X32 FILLER_344_193 ();
 FILLCELL_X32 FILLER_344_225 ();
 FILLCELL_X32 FILLER_344_257 ();
 FILLCELL_X32 FILLER_344_289 ();
 FILLCELL_X32 FILLER_344_321 ();
 FILLCELL_X32 FILLER_344_353 ();
 FILLCELL_X32 FILLER_344_385 ();
 FILLCELL_X32 FILLER_344_417 ();
 FILLCELL_X32 FILLER_344_449 ();
 FILLCELL_X32 FILLER_344_481 ();
 FILLCELL_X32 FILLER_344_513 ();
 FILLCELL_X32 FILLER_344_545 ();
 FILLCELL_X32 FILLER_344_577 ();
 FILLCELL_X16 FILLER_344_609 ();
 FILLCELL_X4 FILLER_344_625 ();
 FILLCELL_X2 FILLER_344_629 ();
 FILLCELL_X32 FILLER_344_632 ();
 FILLCELL_X32 FILLER_344_664 ();
 FILLCELL_X32 FILLER_344_696 ();
 FILLCELL_X32 FILLER_344_728 ();
 FILLCELL_X32 FILLER_344_760 ();
 FILLCELL_X32 FILLER_344_792 ();
 FILLCELL_X32 FILLER_344_824 ();
 FILLCELL_X32 FILLER_344_856 ();
 FILLCELL_X32 FILLER_344_888 ();
 FILLCELL_X32 FILLER_344_920 ();
 FILLCELL_X32 FILLER_344_952 ();
 FILLCELL_X32 FILLER_344_984 ();
 FILLCELL_X32 FILLER_344_1016 ();
 FILLCELL_X32 FILLER_344_1048 ();
 FILLCELL_X32 FILLER_344_1080 ();
 FILLCELL_X32 FILLER_344_1112 ();
 FILLCELL_X32 FILLER_344_1144 ();
 FILLCELL_X32 FILLER_344_1176 ();
 FILLCELL_X32 FILLER_344_1208 ();
 FILLCELL_X32 FILLER_344_1240 ();
 FILLCELL_X32 FILLER_344_1272 ();
 FILLCELL_X32 FILLER_344_1304 ();
 FILLCELL_X32 FILLER_344_1336 ();
 FILLCELL_X32 FILLER_344_1368 ();
 FILLCELL_X32 FILLER_344_1400 ();
 FILLCELL_X32 FILLER_344_1432 ();
 FILLCELL_X32 FILLER_344_1464 ();
 FILLCELL_X32 FILLER_344_1496 ();
 FILLCELL_X32 FILLER_344_1528 ();
 FILLCELL_X32 FILLER_344_1560 ();
 FILLCELL_X32 FILLER_344_1592 ();
 FILLCELL_X32 FILLER_344_1624 ();
 FILLCELL_X32 FILLER_344_1656 ();
 FILLCELL_X32 FILLER_344_1688 ();
 FILLCELL_X32 FILLER_344_1720 ();
 FILLCELL_X32 FILLER_344_1752 ();
 FILLCELL_X32 FILLER_344_1784 ();
 FILLCELL_X32 FILLER_344_1816 ();
 FILLCELL_X32 FILLER_344_1848 ();
 FILLCELL_X8 FILLER_344_1880 ();
 FILLCELL_X4 FILLER_344_1888 ();
 FILLCELL_X2 FILLER_344_1892 ();
 FILLCELL_X32 FILLER_344_1895 ();
 FILLCELL_X32 FILLER_344_1927 ();
 FILLCELL_X32 FILLER_344_1959 ();
 FILLCELL_X32 FILLER_344_1991 ();
 FILLCELL_X32 FILLER_344_2023 ();
 FILLCELL_X32 FILLER_344_2055 ();
 FILLCELL_X32 FILLER_344_2087 ();
 FILLCELL_X32 FILLER_344_2119 ();
 FILLCELL_X32 FILLER_344_2151 ();
 FILLCELL_X32 FILLER_344_2183 ();
 FILLCELL_X32 FILLER_344_2215 ();
 FILLCELL_X32 FILLER_344_2247 ();
 FILLCELL_X32 FILLER_344_2279 ();
 FILLCELL_X32 FILLER_344_2311 ();
 FILLCELL_X32 FILLER_344_2343 ();
 FILLCELL_X32 FILLER_344_2375 ();
 FILLCELL_X32 FILLER_344_2407 ();
 FILLCELL_X32 FILLER_344_2439 ();
 FILLCELL_X32 FILLER_344_2471 ();
 FILLCELL_X32 FILLER_344_2503 ();
 FILLCELL_X32 FILLER_344_2535 ();
 FILLCELL_X32 FILLER_344_2567 ();
 FILLCELL_X2 FILLER_344_2599 ();
 FILLCELL_X1 FILLER_344_2601 ();
 FILLCELL_X32 FILLER_345_1 ();
 FILLCELL_X32 FILLER_345_33 ();
 FILLCELL_X32 FILLER_345_65 ();
 FILLCELL_X32 FILLER_345_97 ();
 FILLCELL_X32 FILLER_345_129 ();
 FILLCELL_X32 FILLER_345_161 ();
 FILLCELL_X32 FILLER_345_193 ();
 FILLCELL_X32 FILLER_345_225 ();
 FILLCELL_X32 FILLER_345_257 ();
 FILLCELL_X32 FILLER_345_289 ();
 FILLCELL_X32 FILLER_345_321 ();
 FILLCELL_X32 FILLER_345_353 ();
 FILLCELL_X32 FILLER_345_385 ();
 FILLCELL_X32 FILLER_345_417 ();
 FILLCELL_X32 FILLER_345_449 ();
 FILLCELL_X32 FILLER_345_481 ();
 FILLCELL_X32 FILLER_345_513 ();
 FILLCELL_X32 FILLER_345_545 ();
 FILLCELL_X32 FILLER_345_577 ();
 FILLCELL_X32 FILLER_345_609 ();
 FILLCELL_X32 FILLER_345_641 ();
 FILLCELL_X32 FILLER_345_673 ();
 FILLCELL_X32 FILLER_345_705 ();
 FILLCELL_X32 FILLER_345_737 ();
 FILLCELL_X32 FILLER_345_769 ();
 FILLCELL_X32 FILLER_345_801 ();
 FILLCELL_X32 FILLER_345_833 ();
 FILLCELL_X32 FILLER_345_865 ();
 FILLCELL_X32 FILLER_345_897 ();
 FILLCELL_X32 FILLER_345_929 ();
 FILLCELL_X32 FILLER_345_961 ();
 FILLCELL_X32 FILLER_345_993 ();
 FILLCELL_X32 FILLER_345_1025 ();
 FILLCELL_X32 FILLER_345_1057 ();
 FILLCELL_X32 FILLER_345_1089 ();
 FILLCELL_X32 FILLER_345_1121 ();
 FILLCELL_X32 FILLER_345_1153 ();
 FILLCELL_X32 FILLER_345_1185 ();
 FILLCELL_X32 FILLER_345_1217 ();
 FILLCELL_X8 FILLER_345_1249 ();
 FILLCELL_X4 FILLER_345_1257 ();
 FILLCELL_X2 FILLER_345_1261 ();
 FILLCELL_X32 FILLER_345_1264 ();
 FILLCELL_X32 FILLER_345_1296 ();
 FILLCELL_X32 FILLER_345_1328 ();
 FILLCELL_X32 FILLER_345_1360 ();
 FILLCELL_X32 FILLER_345_1392 ();
 FILLCELL_X32 FILLER_345_1424 ();
 FILLCELL_X32 FILLER_345_1456 ();
 FILLCELL_X32 FILLER_345_1488 ();
 FILLCELL_X32 FILLER_345_1520 ();
 FILLCELL_X32 FILLER_345_1552 ();
 FILLCELL_X32 FILLER_345_1584 ();
 FILLCELL_X32 FILLER_345_1616 ();
 FILLCELL_X32 FILLER_345_1648 ();
 FILLCELL_X32 FILLER_345_1680 ();
 FILLCELL_X32 FILLER_345_1712 ();
 FILLCELL_X32 FILLER_345_1744 ();
 FILLCELL_X32 FILLER_345_1776 ();
 FILLCELL_X32 FILLER_345_1808 ();
 FILLCELL_X32 FILLER_345_1840 ();
 FILLCELL_X32 FILLER_345_1872 ();
 FILLCELL_X32 FILLER_345_1904 ();
 FILLCELL_X32 FILLER_345_1936 ();
 FILLCELL_X32 FILLER_345_1968 ();
 FILLCELL_X32 FILLER_345_2000 ();
 FILLCELL_X32 FILLER_345_2032 ();
 FILLCELL_X32 FILLER_345_2064 ();
 FILLCELL_X32 FILLER_345_2096 ();
 FILLCELL_X32 FILLER_345_2128 ();
 FILLCELL_X32 FILLER_345_2160 ();
 FILLCELL_X32 FILLER_345_2192 ();
 FILLCELL_X32 FILLER_345_2224 ();
 FILLCELL_X32 FILLER_345_2256 ();
 FILLCELL_X32 FILLER_345_2288 ();
 FILLCELL_X32 FILLER_345_2320 ();
 FILLCELL_X32 FILLER_345_2352 ();
 FILLCELL_X32 FILLER_345_2384 ();
 FILLCELL_X32 FILLER_345_2416 ();
 FILLCELL_X32 FILLER_345_2448 ();
 FILLCELL_X32 FILLER_345_2480 ();
 FILLCELL_X8 FILLER_345_2512 ();
 FILLCELL_X4 FILLER_345_2520 ();
 FILLCELL_X2 FILLER_345_2524 ();
 FILLCELL_X32 FILLER_345_2527 ();
 FILLCELL_X32 FILLER_345_2559 ();
 FILLCELL_X8 FILLER_345_2591 ();
 FILLCELL_X2 FILLER_345_2599 ();
 FILLCELL_X1 FILLER_345_2601 ();
 FILLCELL_X32 FILLER_346_1 ();
 FILLCELL_X32 FILLER_346_33 ();
 FILLCELL_X32 FILLER_346_65 ();
 FILLCELL_X32 FILLER_346_97 ();
 FILLCELL_X32 FILLER_346_129 ();
 FILLCELL_X32 FILLER_346_161 ();
 FILLCELL_X32 FILLER_346_193 ();
 FILLCELL_X32 FILLER_346_225 ();
 FILLCELL_X32 FILLER_346_257 ();
 FILLCELL_X32 FILLER_346_289 ();
 FILLCELL_X32 FILLER_346_321 ();
 FILLCELL_X32 FILLER_346_353 ();
 FILLCELL_X32 FILLER_346_385 ();
 FILLCELL_X32 FILLER_346_417 ();
 FILLCELL_X32 FILLER_346_449 ();
 FILLCELL_X32 FILLER_346_481 ();
 FILLCELL_X32 FILLER_346_513 ();
 FILLCELL_X32 FILLER_346_545 ();
 FILLCELL_X32 FILLER_346_577 ();
 FILLCELL_X16 FILLER_346_609 ();
 FILLCELL_X4 FILLER_346_625 ();
 FILLCELL_X2 FILLER_346_629 ();
 FILLCELL_X32 FILLER_346_632 ();
 FILLCELL_X32 FILLER_346_664 ();
 FILLCELL_X32 FILLER_346_696 ();
 FILLCELL_X32 FILLER_346_728 ();
 FILLCELL_X32 FILLER_346_760 ();
 FILLCELL_X32 FILLER_346_792 ();
 FILLCELL_X32 FILLER_346_824 ();
 FILLCELL_X32 FILLER_346_856 ();
 FILLCELL_X32 FILLER_346_888 ();
 FILLCELL_X32 FILLER_346_920 ();
 FILLCELL_X32 FILLER_346_952 ();
 FILLCELL_X32 FILLER_346_984 ();
 FILLCELL_X32 FILLER_346_1016 ();
 FILLCELL_X32 FILLER_346_1048 ();
 FILLCELL_X32 FILLER_346_1080 ();
 FILLCELL_X32 FILLER_346_1112 ();
 FILLCELL_X32 FILLER_346_1144 ();
 FILLCELL_X32 FILLER_346_1176 ();
 FILLCELL_X32 FILLER_346_1208 ();
 FILLCELL_X32 FILLER_346_1240 ();
 FILLCELL_X32 FILLER_346_1272 ();
 FILLCELL_X32 FILLER_346_1304 ();
 FILLCELL_X32 FILLER_346_1336 ();
 FILLCELL_X32 FILLER_346_1368 ();
 FILLCELL_X32 FILLER_346_1400 ();
 FILLCELL_X32 FILLER_346_1432 ();
 FILLCELL_X32 FILLER_346_1464 ();
 FILLCELL_X32 FILLER_346_1496 ();
 FILLCELL_X32 FILLER_346_1528 ();
 FILLCELL_X32 FILLER_346_1560 ();
 FILLCELL_X32 FILLER_346_1592 ();
 FILLCELL_X32 FILLER_346_1624 ();
 FILLCELL_X32 FILLER_346_1656 ();
 FILLCELL_X32 FILLER_346_1688 ();
 FILLCELL_X32 FILLER_346_1720 ();
 FILLCELL_X32 FILLER_346_1752 ();
 FILLCELL_X32 FILLER_346_1784 ();
 FILLCELL_X32 FILLER_346_1816 ();
 FILLCELL_X32 FILLER_346_1848 ();
 FILLCELL_X8 FILLER_346_1880 ();
 FILLCELL_X4 FILLER_346_1888 ();
 FILLCELL_X2 FILLER_346_1892 ();
 FILLCELL_X32 FILLER_346_1895 ();
 FILLCELL_X32 FILLER_346_1927 ();
 FILLCELL_X32 FILLER_346_1959 ();
 FILLCELL_X32 FILLER_346_1991 ();
 FILLCELL_X32 FILLER_346_2023 ();
 FILLCELL_X32 FILLER_346_2055 ();
 FILLCELL_X32 FILLER_346_2087 ();
 FILLCELL_X32 FILLER_346_2119 ();
 FILLCELL_X32 FILLER_346_2151 ();
 FILLCELL_X32 FILLER_346_2183 ();
 FILLCELL_X32 FILLER_346_2215 ();
 FILLCELL_X32 FILLER_346_2247 ();
 FILLCELL_X32 FILLER_346_2279 ();
 FILLCELL_X32 FILLER_346_2311 ();
 FILLCELL_X32 FILLER_346_2343 ();
 FILLCELL_X32 FILLER_346_2375 ();
 FILLCELL_X32 FILLER_346_2407 ();
 FILLCELL_X32 FILLER_346_2439 ();
 FILLCELL_X32 FILLER_346_2471 ();
 FILLCELL_X32 FILLER_346_2503 ();
 FILLCELL_X32 FILLER_346_2535 ();
 FILLCELL_X32 FILLER_346_2567 ();
 FILLCELL_X2 FILLER_346_2599 ();
 FILLCELL_X1 FILLER_346_2601 ();
 FILLCELL_X32 FILLER_347_1 ();
 FILLCELL_X32 FILLER_347_33 ();
 FILLCELL_X32 FILLER_347_65 ();
 FILLCELL_X32 FILLER_347_97 ();
 FILLCELL_X32 FILLER_347_129 ();
 FILLCELL_X32 FILLER_347_161 ();
 FILLCELL_X32 FILLER_347_193 ();
 FILLCELL_X32 FILLER_347_225 ();
 FILLCELL_X32 FILLER_347_257 ();
 FILLCELL_X32 FILLER_347_289 ();
 FILLCELL_X32 FILLER_347_321 ();
 FILLCELL_X32 FILLER_347_353 ();
 FILLCELL_X32 FILLER_347_385 ();
 FILLCELL_X32 FILLER_347_417 ();
 FILLCELL_X32 FILLER_347_449 ();
 FILLCELL_X32 FILLER_347_481 ();
 FILLCELL_X32 FILLER_347_513 ();
 FILLCELL_X32 FILLER_347_545 ();
 FILLCELL_X32 FILLER_347_577 ();
 FILLCELL_X32 FILLER_347_609 ();
 FILLCELL_X32 FILLER_347_641 ();
 FILLCELL_X32 FILLER_347_673 ();
 FILLCELL_X32 FILLER_347_705 ();
 FILLCELL_X32 FILLER_347_737 ();
 FILLCELL_X32 FILLER_347_769 ();
 FILLCELL_X32 FILLER_347_801 ();
 FILLCELL_X32 FILLER_347_833 ();
 FILLCELL_X32 FILLER_347_865 ();
 FILLCELL_X32 FILLER_347_897 ();
 FILLCELL_X32 FILLER_347_929 ();
 FILLCELL_X32 FILLER_347_961 ();
 FILLCELL_X32 FILLER_347_993 ();
 FILLCELL_X32 FILLER_347_1025 ();
 FILLCELL_X32 FILLER_347_1057 ();
 FILLCELL_X32 FILLER_347_1089 ();
 FILLCELL_X32 FILLER_347_1121 ();
 FILLCELL_X32 FILLER_347_1153 ();
 FILLCELL_X32 FILLER_347_1185 ();
 FILLCELL_X32 FILLER_347_1217 ();
 FILLCELL_X8 FILLER_347_1249 ();
 FILLCELL_X4 FILLER_347_1257 ();
 FILLCELL_X2 FILLER_347_1261 ();
 FILLCELL_X32 FILLER_347_1264 ();
 FILLCELL_X32 FILLER_347_1296 ();
 FILLCELL_X32 FILLER_347_1328 ();
 FILLCELL_X32 FILLER_347_1360 ();
 FILLCELL_X32 FILLER_347_1392 ();
 FILLCELL_X32 FILLER_347_1424 ();
 FILLCELL_X32 FILLER_347_1456 ();
 FILLCELL_X32 FILLER_347_1488 ();
 FILLCELL_X32 FILLER_347_1520 ();
 FILLCELL_X32 FILLER_347_1552 ();
 FILLCELL_X32 FILLER_347_1584 ();
 FILLCELL_X32 FILLER_347_1616 ();
 FILLCELL_X32 FILLER_347_1648 ();
 FILLCELL_X32 FILLER_347_1680 ();
 FILLCELL_X32 FILLER_347_1712 ();
 FILLCELL_X32 FILLER_347_1744 ();
 FILLCELL_X32 FILLER_347_1776 ();
 FILLCELL_X32 FILLER_347_1808 ();
 FILLCELL_X32 FILLER_347_1840 ();
 FILLCELL_X32 FILLER_347_1872 ();
 FILLCELL_X32 FILLER_347_1904 ();
 FILLCELL_X32 FILLER_347_1936 ();
 FILLCELL_X32 FILLER_347_1968 ();
 FILLCELL_X32 FILLER_347_2000 ();
 FILLCELL_X32 FILLER_347_2032 ();
 FILLCELL_X32 FILLER_347_2064 ();
 FILLCELL_X32 FILLER_347_2096 ();
 FILLCELL_X32 FILLER_347_2128 ();
 FILLCELL_X32 FILLER_347_2160 ();
 FILLCELL_X32 FILLER_347_2192 ();
 FILLCELL_X32 FILLER_347_2224 ();
 FILLCELL_X32 FILLER_347_2256 ();
 FILLCELL_X32 FILLER_347_2288 ();
 FILLCELL_X32 FILLER_347_2320 ();
 FILLCELL_X32 FILLER_347_2352 ();
 FILLCELL_X32 FILLER_347_2384 ();
 FILLCELL_X32 FILLER_347_2416 ();
 FILLCELL_X32 FILLER_347_2448 ();
 FILLCELL_X32 FILLER_347_2480 ();
 FILLCELL_X8 FILLER_347_2512 ();
 FILLCELL_X4 FILLER_347_2520 ();
 FILLCELL_X2 FILLER_347_2524 ();
 FILLCELL_X32 FILLER_347_2527 ();
 FILLCELL_X32 FILLER_347_2559 ();
 FILLCELL_X8 FILLER_347_2591 ();
 FILLCELL_X2 FILLER_347_2599 ();
 FILLCELL_X1 FILLER_347_2601 ();
 FILLCELL_X32 FILLER_348_1 ();
 FILLCELL_X32 FILLER_348_33 ();
 FILLCELL_X32 FILLER_348_65 ();
 FILLCELL_X32 FILLER_348_97 ();
 FILLCELL_X32 FILLER_348_129 ();
 FILLCELL_X32 FILLER_348_161 ();
 FILLCELL_X32 FILLER_348_193 ();
 FILLCELL_X32 FILLER_348_225 ();
 FILLCELL_X32 FILLER_348_257 ();
 FILLCELL_X32 FILLER_348_289 ();
 FILLCELL_X32 FILLER_348_321 ();
 FILLCELL_X32 FILLER_348_353 ();
 FILLCELL_X32 FILLER_348_385 ();
 FILLCELL_X32 FILLER_348_417 ();
 FILLCELL_X32 FILLER_348_449 ();
 FILLCELL_X32 FILLER_348_481 ();
 FILLCELL_X32 FILLER_348_513 ();
 FILLCELL_X32 FILLER_348_545 ();
 FILLCELL_X32 FILLER_348_577 ();
 FILLCELL_X16 FILLER_348_609 ();
 FILLCELL_X4 FILLER_348_625 ();
 FILLCELL_X2 FILLER_348_629 ();
 FILLCELL_X32 FILLER_348_632 ();
 FILLCELL_X32 FILLER_348_664 ();
 FILLCELL_X32 FILLER_348_696 ();
 FILLCELL_X32 FILLER_348_728 ();
 FILLCELL_X32 FILLER_348_760 ();
 FILLCELL_X32 FILLER_348_792 ();
 FILLCELL_X32 FILLER_348_824 ();
 FILLCELL_X32 FILLER_348_856 ();
 FILLCELL_X32 FILLER_348_888 ();
 FILLCELL_X32 FILLER_348_920 ();
 FILLCELL_X32 FILLER_348_952 ();
 FILLCELL_X32 FILLER_348_984 ();
 FILLCELL_X32 FILLER_348_1016 ();
 FILLCELL_X32 FILLER_348_1048 ();
 FILLCELL_X32 FILLER_348_1080 ();
 FILLCELL_X32 FILLER_348_1112 ();
 FILLCELL_X32 FILLER_348_1144 ();
 FILLCELL_X32 FILLER_348_1176 ();
 FILLCELL_X32 FILLER_348_1208 ();
 FILLCELL_X32 FILLER_348_1240 ();
 FILLCELL_X32 FILLER_348_1272 ();
 FILLCELL_X32 FILLER_348_1304 ();
 FILLCELL_X32 FILLER_348_1336 ();
 FILLCELL_X32 FILLER_348_1368 ();
 FILLCELL_X32 FILLER_348_1400 ();
 FILLCELL_X32 FILLER_348_1432 ();
 FILLCELL_X32 FILLER_348_1464 ();
 FILLCELL_X32 FILLER_348_1496 ();
 FILLCELL_X32 FILLER_348_1528 ();
 FILLCELL_X32 FILLER_348_1560 ();
 FILLCELL_X32 FILLER_348_1592 ();
 FILLCELL_X32 FILLER_348_1624 ();
 FILLCELL_X32 FILLER_348_1656 ();
 FILLCELL_X32 FILLER_348_1688 ();
 FILLCELL_X32 FILLER_348_1720 ();
 FILLCELL_X32 FILLER_348_1752 ();
 FILLCELL_X32 FILLER_348_1784 ();
 FILLCELL_X32 FILLER_348_1816 ();
 FILLCELL_X32 FILLER_348_1848 ();
 FILLCELL_X8 FILLER_348_1880 ();
 FILLCELL_X4 FILLER_348_1888 ();
 FILLCELL_X2 FILLER_348_1892 ();
 FILLCELL_X32 FILLER_348_1895 ();
 FILLCELL_X32 FILLER_348_1927 ();
 FILLCELL_X32 FILLER_348_1959 ();
 FILLCELL_X32 FILLER_348_1991 ();
 FILLCELL_X32 FILLER_348_2023 ();
 FILLCELL_X32 FILLER_348_2055 ();
 FILLCELL_X32 FILLER_348_2087 ();
 FILLCELL_X32 FILLER_348_2119 ();
 FILLCELL_X32 FILLER_348_2151 ();
 FILLCELL_X32 FILLER_348_2183 ();
 FILLCELL_X32 FILLER_348_2215 ();
 FILLCELL_X32 FILLER_348_2247 ();
 FILLCELL_X32 FILLER_348_2279 ();
 FILLCELL_X32 FILLER_348_2311 ();
 FILLCELL_X32 FILLER_348_2343 ();
 FILLCELL_X32 FILLER_348_2375 ();
 FILLCELL_X32 FILLER_348_2407 ();
 FILLCELL_X32 FILLER_348_2439 ();
 FILLCELL_X32 FILLER_348_2471 ();
 FILLCELL_X32 FILLER_348_2503 ();
 FILLCELL_X32 FILLER_348_2535 ();
 FILLCELL_X32 FILLER_348_2567 ();
 FILLCELL_X2 FILLER_348_2599 ();
 FILLCELL_X1 FILLER_348_2601 ();
 FILLCELL_X32 FILLER_349_1 ();
 FILLCELL_X32 FILLER_349_33 ();
 FILLCELL_X32 FILLER_349_65 ();
 FILLCELL_X32 FILLER_349_97 ();
 FILLCELL_X32 FILLER_349_129 ();
 FILLCELL_X32 FILLER_349_161 ();
 FILLCELL_X32 FILLER_349_193 ();
 FILLCELL_X32 FILLER_349_225 ();
 FILLCELL_X32 FILLER_349_257 ();
 FILLCELL_X32 FILLER_349_289 ();
 FILLCELL_X32 FILLER_349_321 ();
 FILLCELL_X32 FILLER_349_353 ();
 FILLCELL_X32 FILLER_349_385 ();
 FILLCELL_X32 FILLER_349_417 ();
 FILLCELL_X32 FILLER_349_449 ();
 FILLCELL_X32 FILLER_349_481 ();
 FILLCELL_X32 FILLER_349_513 ();
 FILLCELL_X32 FILLER_349_545 ();
 FILLCELL_X32 FILLER_349_577 ();
 FILLCELL_X32 FILLER_349_609 ();
 FILLCELL_X32 FILLER_349_641 ();
 FILLCELL_X32 FILLER_349_673 ();
 FILLCELL_X32 FILLER_349_705 ();
 FILLCELL_X32 FILLER_349_737 ();
 FILLCELL_X32 FILLER_349_769 ();
 FILLCELL_X32 FILLER_349_801 ();
 FILLCELL_X32 FILLER_349_833 ();
 FILLCELL_X32 FILLER_349_865 ();
 FILLCELL_X32 FILLER_349_897 ();
 FILLCELL_X32 FILLER_349_929 ();
 FILLCELL_X32 FILLER_349_961 ();
 FILLCELL_X32 FILLER_349_993 ();
 FILLCELL_X32 FILLER_349_1025 ();
 FILLCELL_X32 FILLER_349_1057 ();
 FILLCELL_X32 FILLER_349_1089 ();
 FILLCELL_X32 FILLER_349_1121 ();
 FILLCELL_X32 FILLER_349_1153 ();
 FILLCELL_X32 FILLER_349_1185 ();
 FILLCELL_X32 FILLER_349_1217 ();
 FILLCELL_X8 FILLER_349_1249 ();
 FILLCELL_X4 FILLER_349_1257 ();
 FILLCELL_X2 FILLER_349_1261 ();
 FILLCELL_X32 FILLER_349_1264 ();
 FILLCELL_X32 FILLER_349_1296 ();
 FILLCELL_X32 FILLER_349_1328 ();
 FILLCELL_X32 FILLER_349_1360 ();
 FILLCELL_X32 FILLER_349_1392 ();
 FILLCELL_X32 FILLER_349_1424 ();
 FILLCELL_X32 FILLER_349_1456 ();
 FILLCELL_X32 FILLER_349_1488 ();
 FILLCELL_X32 FILLER_349_1520 ();
 FILLCELL_X32 FILLER_349_1552 ();
 FILLCELL_X32 FILLER_349_1584 ();
 FILLCELL_X32 FILLER_349_1616 ();
 FILLCELL_X32 FILLER_349_1648 ();
 FILLCELL_X32 FILLER_349_1680 ();
 FILLCELL_X32 FILLER_349_1712 ();
 FILLCELL_X32 FILLER_349_1744 ();
 FILLCELL_X32 FILLER_349_1776 ();
 FILLCELL_X32 FILLER_349_1808 ();
 FILLCELL_X32 FILLER_349_1840 ();
 FILLCELL_X32 FILLER_349_1872 ();
 FILLCELL_X32 FILLER_349_1904 ();
 FILLCELL_X32 FILLER_349_1936 ();
 FILLCELL_X32 FILLER_349_1968 ();
 FILLCELL_X32 FILLER_349_2000 ();
 FILLCELL_X32 FILLER_349_2032 ();
 FILLCELL_X32 FILLER_349_2064 ();
 FILLCELL_X32 FILLER_349_2096 ();
 FILLCELL_X32 FILLER_349_2128 ();
 FILLCELL_X32 FILLER_349_2160 ();
 FILLCELL_X32 FILLER_349_2192 ();
 FILLCELL_X32 FILLER_349_2224 ();
 FILLCELL_X32 FILLER_349_2256 ();
 FILLCELL_X32 FILLER_349_2288 ();
 FILLCELL_X32 FILLER_349_2320 ();
 FILLCELL_X32 FILLER_349_2352 ();
 FILLCELL_X32 FILLER_349_2384 ();
 FILLCELL_X32 FILLER_349_2416 ();
 FILLCELL_X32 FILLER_349_2448 ();
 FILLCELL_X32 FILLER_349_2480 ();
 FILLCELL_X8 FILLER_349_2512 ();
 FILLCELL_X4 FILLER_349_2520 ();
 FILLCELL_X2 FILLER_349_2524 ();
 FILLCELL_X32 FILLER_349_2527 ();
 FILLCELL_X32 FILLER_349_2559 ();
 FILLCELL_X8 FILLER_349_2591 ();
 FILLCELL_X2 FILLER_349_2599 ();
 FILLCELL_X1 FILLER_349_2601 ();
 FILLCELL_X32 FILLER_350_1 ();
 FILLCELL_X32 FILLER_350_33 ();
 FILLCELL_X32 FILLER_350_65 ();
 FILLCELL_X32 FILLER_350_97 ();
 FILLCELL_X32 FILLER_350_129 ();
 FILLCELL_X32 FILLER_350_161 ();
 FILLCELL_X32 FILLER_350_193 ();
 FILLCELL_X32 FILLER_350_225 ();
 FILLCELL_X32 FILLER_350_257 ();
 FILLCELL_X32 FILLER_350_289 ();
 FILLCELL_X32 FILLER_350_321 ();
 FILLCELL_X32 FILLER_350_353 ();
 FILLCELL_X32 FILLER_350_385 ();
 FILLCELL_X32 FILLER_350_417 ();
 FILLCELL_X32 FILLER_350_449 ();
 FILLCELL_X32 FILLER_350_481 ();
 FILLCELL_X32 FILLER_350_513 ();
 FILLCELL_X32 FILLER_350_545 ();
 FILLCELL_X32 FILLER_350_577 ();
 FILLCELL_X16 FILLER_350_609 ();
 FILLCELL_X4 FILLER_350_625 ();
 FILLCELL_X2 FILLER_350_629 ();
 FILLCELL_X32 FILLER_350_632 ();
 FILLCELL_X32 FILLER_350_664 ();
 FILLCELL_X32 FILLER_350_696 ();
 FILLCELL_X32 FILLER_350_728 ();
 FILLCELL_X32 FILLER_350_760 ();
 FILLCELL_X32 FILLER_350_792 ();
 FILLCELL_X32 FILLER_350_824 ();
 FILLCELL_X32 FILLER_350_856 ();
 FILLCELL_X32 FILLER_350_888 ();
 FILLCELL_X32 FILLER_350_920 ();
 FILLCELL_X32 FILLER_350_952 ();
 FILLCELL_X32 FILLER_350_984 ();
 FILLCELL_X32 FILLER_350_1016 ();
 FILLCELL_X32 FILLER_350_1048 ();
 FILLCELL_X32 FILLER_350_1080 ();
 FILLCELL_X32 FILLER_350_1112 ();
 FILLCELL_X32 FILLER_350_1144 ();
 FILLCELL_X32 FILLER_350_1176 ();
 FILLCELL_X32 FILLER_350_1208 ();
 FILLCELL_X32 FILLER_350_1240 ();
 FILLCELL_X16 FILLER_350_1272 ();
 FILLCELL_X1 FILLER_350_1288 ();
 FILLCELL_X32 FILLER_350_1292 ();
 FILLCELL_X32 FILLER_350_1324 ();
 FILLCELL_X32 FILLER_350_1356 ();
 FILLCELL_X32 FILLER_350_1388 ();
 FILLCELL_X32 FILLER_350_1420 ();
 FILLCELL_X32 FILLER_350_1452 ();
 FILLCELL_X32 FILLER_350_1484 ();
 FILLCELL_X32 FILLER_350_1516 ();
 FILLCELL_X32 FILLER_350_1548 ();
 FILLCELL_X32 FILLER_350_1580 ();
 FILLCELL_X32 FILLER_350_1612 ();
 FILLCELL_X32 FILLER_350_1644 ();
 FILLCELL_X32 FILLER_350_1676 ();
 FILLCELL_X32 FILLER_350_1708 ();
 FILLCELL_X32 FILLER_350_1740 ();
 FILLCELL_X32 FILLER_350_1772 ();
 FILLCELL_X32 FILLER_350_1804 ();
 FILLCELL_X32 FILLER_350_1836 ();
 FILLCELL_X16 FILLER_350_1868 ();
 FILLCELL_X8 FILLER_350_1884 ();
 FILLCELL_X2 FILLER_350_1892 ();
 FILLCELL_X32 FILLER_350_1895 ();
 FILLCELL_X32 FILLER_350_1927 ();
 FILLCELL_X32 FILLER_350_1959 ();
 FILLCELL_X32 FILLER_350_1991 ();
 FILLCELL_X32 FILLER_350_2023 ();
 FILLCELL_X32 FILLER_350_2055 ();
 FILLCELL_X32 FILLER_350_2087 ();
 FILLCELL_X32 FILLER_350_2119 ();
 FILLCELL_X32 FILLER_350_2151 ();
 FILLCELL_X32 FILLER_350_2183 ();
 FILLCELL_X32 FILLER_350_2215 ();
 FILLCELL_X32 FILLER_350_2247 ();
 FILLCELL_X32 FILLER_350_2279 ();
 FILLCELL_X32 FILLER_350_2311 ();
 FILLCELL_X32 FILLER_350_2343 ();
 FILLCELL_X32 FILLER_350_2375 ();
 FILLCELL_X32 FILLER_350_2407 ();
 FILLCELL_X32 FILLER_350_2439 ();
 FILLCELL_X32 FILLER_350_2471 ();
 FILLCELL_X32 FILLER_350_2503 ();
 FILLCELL_X32 FILLER_350_2535 ();
 FILLCELL_X32 FILLER_350_2567 ();
 FILLCELL_X2 FILLER_350_2599 ();
 FILLCELL_X1 FILLER_350_2601 ();
 FILLCELL_X32 FILLER_351_1 ();
 FILLCELL_X32 FILLER_351_33 ();
 FILLCELL_X32 FILLER_351_65 ();
 FILLCELL_X32 FILLER_351_97 ();
 FILLCELL_X32 FILLER_351_129 ();
 FILLCELL_X32 FILLER_351_161 ();
 FILLCELL_X32 FILLER_351_193 ();
 FILLCELL_X32 FILLER_351_225 ();
 FILLCELL_X32 FILLER_351_257 ();
 FILLCELL_X32 FILLER_351_289 ();
 FILLCELL_X32 FILLER_351_321 ();
 FILLCELL_X32 FILLER_351_353 ();
 FILLCELL_X32 FILLER_351_385 ();
 FILLCELL_X32 FILLER_351_417 ();
 FILLCELL_X32 FILLER_351_449 ();
 FILLCELL_X32 FILLER_351_481 ();
 FILLCELL_X32 FILLER_351_513 ();
 FILLCELL_X32 FILLER_351_545 ();
 FILLCELL_X32 FILLER_351_577 ();
 FILLCELL_X32 FILLER_351_609 ();
 FILLCELL_X32 FILLER_351_641 ();
 FILLCELL_X32 FILLER_351_673 ();
 FILLCELL_X32 FILLER_351_705 ();
 FILLCELL_X32 FILLER_351_737 ();
 FILLCELL_X32 FILLER_351_769 ();
 FILLCELL_X32 FILLER_351_801 ();
 FILLCELL_X32 FILLER_351_833 ();
 FILLCELL_X32 FILLER_351_865 ();
 FILLCELL_X32 FILLER_351_897 ();
 FILLCELL_X32 FILLER_351_929 ();
 FILLCELL_X32 FILLER_351_961 ();
 FILLCELL_X32 FILLER_351_993 ();
 FILLCELL_X32 FILLER_351_1025 ();
 FILLCELL_X32 FILLER_351_1057 ();
 FILLCELL_X32 FILLER_351_1089 ();
 FILLCELL_X32 FILLER_351_1121 ();
 FILLCELL_X32 FILLER_351_1153 ();
 FILLCELL_X32 FILLER_351_1185 ();
 FILLCELL_X16 FILLER_351_1217 ();
 FILLCELL_X2 FILLER_351_1233 ();
 FILLCELL_X8 FILLER_351_1237 ();
 FILLCELL_X4 FILLER_351_1245 ();
 FILLCELL_X1 FILLER_351_1249 ();
 FILLCELL_X8 FILLER_351_1253 ();
 FILLCELL_X2 FILLER_351_1261 ();
 FILLCELL_X16 FILLER_351_1264 ();
 FILLCELL_X4 FILLER_351_1280 ();
 FILLCELL_X2 FILLER_351_1284 ();
 FILLCELL_X32 FILLER_351_1289 ();
 FILLCELL_X32 FILLER_351_1321 ();
 FILLCELL_X32 FILLER_351_1353 ();
 FILLCELL_X32 FILLER_351_1385 ();
 FILLCELL_X32 FILLER_351_1417 ();
 FILLCELL_X32 FILLER_351_1449 ();
 FILLCELL_X32 FILLER_351_1481 ();
 FILLCELL_X32 FILLER_351_1513 ();
 FILLCELL_X32 FILLER_351_1545 ();
 FILLCELL_X32 FILLER_351_1577 ();
 FILLCELL_X32 FILLER_351_1609 ();
 FILLCELL_X32 FILLER_351_1641 ();
 FILLCELL_X32 FILLER_351_1673 ();
 FILLCELL_X32 FILLER_351_1705 ();
 FILLCELL_X32 FILLER_351_1737 ();
 FILLCELL_X32 FILLER_351_1769 ();
 FILLCELL_X32 FILLER_351_1801 ();
 FILLCELL_X32 FILLER_351_1833 ();
 FILLCELL_X32 FILLER_351_1865 ();
 FILLCELL_X32 FILLER_351_1897 ();
 FILLCELL_X32 FILLER_351_1929 ();
 FILLCELL_X32 FILLER_351_1961 ();
 FILLCELL_X32 FILLER_351_1993 ();
 FILLCELL_X32 FILLER_351_2025 ();
 FILLCELL_X32 FILLER_351_2057 ();
 FILLCELL_X32 FILLER_351_2089 ();
 FILLCELL_X32 FILLER_351_2121 ();
 FILLCELL_X32 FILLER_351_2153 ();
 FILLCELL_X32 FILLER_351_2185 ();
 FILLCELL_X32 FILLER_351_2217 ();
 FILLCELL_X32 FILLER_351_2249 ();
 FILLCELL_X32 FILLER_351_2281 ();
 FILLCELL_X32 FILLER_351_2313 ();
 FILLCELL_X32 FILLER_351_2345 ();
 FILLCELL_X32 FILLER_351_2377 ();
 FILLCELL_X32 FILLER_351_2409 ();
 FILLCELL_X32 FILLER_351_2441 ();
 FILLCELL_X32 FILLER_351_2473 ();
 FILLCELL_X16 FILLER_351_2505 ();
 FILLCELL_X4 FILLER_351_2521 ();
 FILLCELL_X1 FILLER_351_2525 ();
 FILLCELL_X32 FILLER_351_2527 ();
 FILLCELL_X32 FILLER_351_2559 ();
 FILLCELL_X8 FILLER_351_2591 ();
 FILLCELL_X2 FILLER_351_2599 ();
 FILLCELL_X1 FILLER_351_2601 ();
 FILLCELL_X32 FILLER_352_1 ();
 FILLCELL_X32 FILLER_352_33 ();
 FILLCELL_X32 FILLER_352_65 ();
 FILLCELL_X32 FILLER_352_97 ();
 FILLCELL_X32 FILLER_352_129 ();
 FILLCELL_X32 FILLER_352_161 ();
 FILLCELL_X32 FILLER_352_193 ();
 FILLCELL_X32 FILLER_352_225 ();
 FILLCELL_X32 FILLER_352_257 ();
 FILLCELL_X32 FILLER_352_289 ();
 FILLCELL_X32 FILLER_352_321 ();
 FILLCELL_X32 FILLER_352_353 ();
 FILLCELL_X32 FILLER_352_385 ();
 FILLCELL_X32 FILLER_352_417 ();
 FILLCELL_X32 FILLER_352_449 ();
 FILLCELL_X32 FILLER_352_481 ();
 FILLCELL_X32 FILLER_352_513 ();
 FILLCELL_X32 FILLER_352_545 ();
 FILLCELL_X32 FILLER_352_577 ();
 FILLCELL_X16 FILLER_352_609 ();
 FILLCELL_X4 FILLER_352_625 ();
 FILLCELL_X2 FILLER_352_629 ();
 FILLCELL_X32 FILLER_352_632 ();
 FILLCELL_X32 FILLER_352_664 ();
 FILLCELL_X32 FILLER_352_696 ();
 FILLCELL_X32 FILLER_352_728 ();
 FILLCELL_X32 FILLER_352_760 ();
 FILLCELL_X32 FILLER_352_792 ();
 FILLCELL_X32 FILLER_352_824 ();
 FILLCELL_X32 FILLER_352_856 ();
 FILLCELL_X32 FILLER_352_888 ();
 FILLCELL_X32 FILLER_352_920 ();
 FILLCELL_X32 FILLER_352_952 ();
 FILLCELL_X32 FILLER_352_984 ();
 FILLCELL_X32 FILLER_352_1016 ();
 FILLCELL_X32 FILLER_352_1048 ();
 FILLCELL_X32 FILLER_352_1080 ();
 FILLCELL_X32 FILLER_352_1112 ();
 FILLCELL_X32 FILLER_352_1144 ();
 FILLCELL_X32 FILLER_352_1176 ();
 FILLCELL_X16 FILLER_352_1208 ();
 FILLCELL_X4 FILLER_352_1224 ();
 FILLCELL_X1 FILLER_352_1228 ();
 FILLCELL_X16 FILLER_352_1232 ();
 FILLCELL_X2 FILLER_352_1248 ();
 FILLCELL_X8 FILLER_352_1253 ();
 FILLCELL_X1 FILLER_352_1261 ();
 FILLCELL_X32 FILLER_352_1263 ();
 FILLCELL_X32 FILLER_352_1295 ();
 FILLCELL_X32 FILLER_352_1327 ();
 FILLCELL_X32 FILLER_352_1359 ();
 FILLCELL_X32 FILLER_352_1391 ();
 FILLCELL_X32 FILLER_352_1423 ();
 FILLCELL_X32 FILLER_352_1455 ();
 FILLCELL_X32 FILLER_352_1487 ();
 FILLCELL_X32 FILLER_352_1519 ();
 FILLCELL_X32 FILLER_352_1551 ();
 FILLCELL_X32 FILLER_352_1583 ();
 FILLCELL_X32 FILLER_352_1615 ();
 FILLCELL_X32 FILLER_352_1647 ();
 FILLCELL_X32 FILLER_352_1679 ();
 FILLCELL_X32 FILLER_352_1711 ();
 FILLCELL_X32 FILLER_352_1743 ();
 FILLCELL_X32 FILLER_352_1775 ();
 FILLCELL_X32 FILLER_352_1807 ();
 FILLCELL_X32 FILLER_352_1839 ();
 FILLCELL_X16 FILLER_352_1871 ();
 FILLCELL_X4 FILLER_352_1887 ();
 FILLCELL_X2 FILLER_352_1891 ();
 FILLCELL_X32 FILLER_352_1894 ();
 FILLCELL_X32 FILLER_352_1926 ();
 FILLCELL_X32 FILLER_352_1958 ();
 FILLCELL_X32 FILLER_352_1990 ();
 FILLCELL_X32 FILLER_352_2022 ();
 FILLCELL_X32 FILLER_352_2054 ();
 FILLCELL_X32 FILLER_352_2086 ();
 FILLCELL_X32 FILLER_352_2118 ();
 FILLCELL_X32 FILLER_352_2150 ();
 FILLCELL_X32 FILLER_352_2182 ();
 FILLCELL_X32 FILLER_352_2214 ();
 FILLCELL_X32 FILLER_352_2246 ();
 FILLCELL_X32 FILLER_352_2278 ();
 FILLCELL_X32 FILLER_352_2310 ();
 FILLCELL_X32 FILLER_352_2342 ();
 FILLCELL_X32 FILLER_352_2374 ();
 FILLCELL_X32 FILLER_352_2406 ();
 FILLCELL_X32 FILLER_352_2438 ();
 FILLCELL_X32 FILLER_352_2470 ();
 FILLCELL_X16 FILLER_352_2502 ();
 FILLCELL_X4 FILLER_352_2518 ();
 FILLCELL_X2 FILLER_352_2522 ();
 FILLCELL_X32 FILLER_352_2525 ();
 FILLCELL_X32 FILLER_352_2557 ();
 FILLCELL_X8 FILLER_352_2589 ();
 FILLCELL_X4 FILLER_352_2597 ();
 FILLCELL_X1 FILLER_352_2601 ();
endmodule
