module shadow_register (clk,
    main_load_en,
    rst_n,
    shadow_capture_en,
    shadow_load_en,
    use_shadow_out,
    main_data_in,
    main_data_out,
    shadow_data_in,
    shadow_data_out);
 input clk;
 input main_load_en;
 input rst_n;
 input shadow_capture_en;
 input shadow_load_en;
 input use_shadow_out;
 input [31:0] main_data_in;
 output [31:0] main_data_out;
 input [31:0] shadow_data_in;
 output [31:0] shadow_data_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire \main_reg[0] ;
 wire \main_reg[10] ;
 wire \main_reg[11] ;
 wire \main_reg[12] ;
 wire \main_reg[13] ;
 wire \main_reg[14] ;
 wire \main_reg[15] ;
 wire \main_reg[16] ;
 wire \main_reg[17] ;
 wire \main_reg[18] ;
 wire \main_reg[19] ;
 wire \main_reg[1] ;
 wire \main_reg[20] ;
 wire \main_reg[21] ;
 wire \main_reg[22] ;
 wire \main_reg[23] ;
 wire \main_reg[24] ;
 wire \main_reg[25] ;
 wire \main_reg[26] ;
 wire \main_reg[27] ;
 wire \main_reg[28] ;
 wire \main_reg[29] ;
 wire \main_reg[2] ;
 wire \main_reg[30] ;
 wire \main_reg[31] ;
 wire \main_reg[3] ;
 wire \main_reg[4] ;
 wire \main_reg[5] ;
 wire \main_reg[6] ;
 wire \main_reg[7] ;
 wire \main_reg[8] ;
 wire \main_reg[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net130;

 sky130_fd_sc_hd__buf_6 _147_ (.A(main_load_en),
    .X(_064_));
 sky130_fd_sc_hd__buf_8 _148_ (.A(_064_),
    .X(_065_));
 sky130_fd_sc_hd__mux2_1 _149_ (.A0(\main_reg[0] ),
    .A1(net2),
    .S(_065_),
    .X(_000_));
 sky130_fd_sc_hd__mux2_1 _150_ (.A0(\main_reg[10] ),
    .A1(net3),
    .S(_065_),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _151_ (.A0(\main_reg[11] ),
    .A1(net4),
    .S(_065_),
    .X(_002_));
 sky130_fd_sc_hd__mux2_1 _152_ (.A0(\main_reg[12] ),
    .A1(net5),
    .S(_065_),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _153_ (.A0(\main_reg[13] ),
    .A1(net6),
    .S(_065_),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _154_ (.A0(\main_reg[14] ),
    .A1(net7),
    .S(_065_),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _155_ (.A0(\main_reg[15] ),
    .A1(net8),
    .S(_065_),
    .X(_006_));
 sky130_fd_sc_hd__mux2_1 _156_ (.A0(\main_reg[16] ),
    .A1(net9),
    .S(_065_),
    .X(_007_));
 sky130_fd_sc_hd__mux2_1 _157_ (.A0(\main_reg[17] ),
    .A1(net10),
    .S(_065_),
    .X(_008_));
 sky130_fd_sc_hd__mux2_1 _158_ (.A0(\main_reg[18] ),
    .A1(net11),
    .S(_065_),
    .X(_009_));
 sky130_fd_sc_hd__buf_8 _159_ (.A(_064_),
    .X(_066_));
 sky130_fd_sc_hd__mux2_1 _160_ (.A0(\main_reg[19] ),
    .A1(net12),
    .S(_066_),
    .X(_010_));
 sky130_fd_sc_hd__mux2_1 _161_ (.A0(\main_reg[1] ),
    .A1(net13),
    .S(_066_),
    .X(_011_));
 sky130_fd_sc_hd__mux2_1 _162_ (.A0(\main_reg[20] ),
    .A1(net14),
    .S(_066_),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _163_ (.A0(\main_reg[21] ),
    .A1(net15),
    .S(_066_),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _164_ (.A0(\main_reg[22] ),
    .A1(net16),
    .S(_066_),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _165_ (.A0(\main_reg[23] ),
    .A1(net17),
    .S(_066_),
    .X(_015_));
 sky130_fd_sc_hd__mux2_1 _166_ (.A0(\main_reg[24] ),
    .A1(net18),
    .S(_066_),
    .X(_016_));
 sky130_fd_sc_hd__mux2_1 _167_ (.A0(\main_reg[25] ),
    .A1(net19),
    .S(_066_),
    .X(_017_));
 sky130_fd_sc_hd__mux2_1 _168_ (.A0(\main_reg[26] ),
    .A1(net20),
    .S(_066_),
    .X(_018_));
 sky130_fd_sc_hd__mux2_1 _169_ (.A0(\main_reg[27] ),
    .A1(net21),
    .S(_066_),
    .X(_019_));
 sky130_fd_sc_hd__buf_8 _170_ (.A(_064_),
    .X(_067_));
 sky130_fd_sc_hd__mux2_1 _171_ (.A0(\main_reg[28] ),
    .A1(net22),
    .S(_067_),
    .X(_020_));
 sky130_fd_sc_hd__mux2_1 _172_ (.A0(\main_reg[29] ),
    .A1(net23),
    .S(_067_),
    .X(_021_));
 sky130_fd_sc_hd__mux2_1 _173_ (.A0(\main_reg[2] ),
    .A1(net24),
    .S(_067_),
    .X(_022_));
 sky130_fd_sc_hd__mux2_1 _174_ (.A0(\main_reg[30] ),
    .A1(net25),
    .S(_067_),
    .X(_023_));
 sky130_fd_sc_hd__mux2_1 _175_ (.A0(\main_reg[31] ),
    .A1(net26),
    .S(_067_),
    .X(_024_));
 sky130_fd_sc_hd__mux2_1 _176_ (.A0(\main_reg[3] ),
    .A1(net27),
    .S(_067_),
    .X(_025_));
 sky130_fd_sc_hd__mux2_1 _177_ (.A0(\main_reg[4] ),
    .A1(net28),
    .S(_067_),
    .X(_026_));
 sky130_fd_sc_hd__mux2_1 _178_ (.A0(\main_reg[5] ),
    .A1(net29),
    .S(_067_),
    .X(_027_));
 sky130_fd_sc_hd__mux2_1 _179_ (.A0(\main_reg[6] ),
    .A1(net30),
    .S(_067_),
    .X(_028_));
 sky130_fd_sc_hd__mux2_1 _180_ (.A0(\main_reg[7] ),
    .A1(net31),
    .S(_067_),
    .X(_029_));
 sky130_fd_sc_hd__mux2_1 _181_ (.A0(\main_reg[8] ),
    .A1(net32),
    .S(_064_),
    .X(_030_));
 sky130_fd_sc_hd__mux2_1 _182_ (.A0(\main_reg[9] ),
    .A1(net33),
    .S(_064_),
    .X(_031_));
 sky130_fd_sc_hd__buf_2 _183_ (.A(shadow_capture_en),
    .X(_068_));
 sky130_fd_sc_hd__buf_2 _184_ (.A(_068_),
    .X(_069_));
 sky130_fd_sc_hd__buf_6 _185_ (.A(shadow_load_en),
    .X(_070_));
 sky130_fd_sc_hd__buf_8 _186_ (.A(_070_),
    .X(_071_));
 sky130_fd_sc_hd__mux2i_1 _187_ (.A0(net98),
    .A1(net34),
    .S(_071_),
    .Y(_072_));
 sky130_fd_sc_hd__buf_2 _188_ (.A(_068_),
    .X(_073_));
 sky130_fd_sc_hd__nand2_1 _189_ (.A(_073_),
    .B(\main_reg[0] ),
    .Y(_074_));
 sky130_fd_sc_hd__o21ai_0 _190_ (.A1(_069_),
    .A2(_072_),
    .B1(_074_),
    .Y(_032_));
 sky130_fd_sc_hd__mux2i_1 _191_ (.A0(net99),
    .A1(net35),
    .S(_071_),
    .Y(_075_));
 sky130_fd_sc_hd__nand2_1 _192_ (.A(_073_),
    .B(\main_reg[10] ),
    .Y(_076_));
 sky130_fd_sc_hd__o21ai_0 _193_ (.A1(_069_),
    .A2(_075_),
    .B1(_076_),
    .Y(_033_));
 sky130_fd_sc_hd__mux2i_1 _194_ (.A0(net100),
    .A1(net36),
    .S(_071_),
    .Y(_077_));
 sky130_fd_sc_hd__nand2_1 _195_ (.A(_073_),
    .B(\main_reg[11] ),
    .Y(_078_));
 sky130_fd_sc_hd__o21ai_0 _196_ (.A1(_069_),
    .A2(_077_),
    .B1(_078_),
    .Y(_034_));
 sky130_fd_sc_hd__mux2i_1 _197_ (.A0(net101),
    .A1(net37),
    .S(_071_),
    .Y(_079_));
 sky130_fd_sc_hd__nand2_1 _198_ (.A(_073_),
    .B(\main_reg[12] ),
    .Y(_080_));
 sky130_fd_sc_hd__o21ai_0 _199_ (.A1(_069_),
    .A2(_079_),
    .B1(_080_),
    .Y(_035_));
 sky130_fd_sc_hd__mux2i_1 _200_ (.A0(net102),
    .A1(net38),
    .S(_071_),
    .Y(_081_));
 sky130_fd_sc_hd__nand2_1 _201_ (.A(_073_),
    .B(\main_reg[13] ),
    .Y(_082_));
 sky130_fd_sc_hd__o21ai_0 _202_ (.A1(_069_),
    .A2(_081_),
    .B1(_082_),
    .Y(_036_));
 sky130_fd_sc_hd__mux2i_1 _203_ (.A0(net103),
    .A1(net39),
    .S(_071_),
    .Y(_083_));
 sky130_fd_sc_hd__nand2_1 _204_ (.A(_073_),
    .B(\main_reg[14] ),
    .Y(_084_));
 sky130_fd_sc_hd__o21ai_0 _205_ (.A1(_069_),
    .A2(_083_),
    .B1(_084_),
    .Y(_037_));
 sky130_fd_sc_hd__mux2i_1 _206_ (.A0(net104),
    .A1(net40),
    .S(_071_),
    .Y(_085_));
 sky130_fd_sc_hd__nand2_1 _207_ (.A(_073_),
    .B(\main_reg[15] ),
    .Y(_086_));
 sky130_fd_sc_hd__o21ai_0 _208_ (.A1(_069_),
    .A2(_085_),
    .B1(_086_),
    .Y(_038_));
 sky130_fd_sc_hd__mux2i_1 _209_ (.A0(net105),
    .A1(net41),
    .S(_071_),
    .Y(_087_));
 sky130_fd_sc_hd__nand2_1 _210_ (.A(_073_),
    .B(\main_reg[16] ),
    .Y(_088_));
 sky130_fd_sc_hd__o21ai_0 _211_ (.A1(_069_),
    .A2(_087_),
    .B1(_088_),
    .Y(_039_));
 sky130_fd_sc_hd__buf_2 _212_ (.A(_068_),
    .X(_089_));
 sky130_fd_sc_hd__mux2i_1 _213_ (.A0(net106),
    .A1(net42),
    .S(_071_),
    .Y(_090_));
 sky130_fd_sc_hd__nand2_1 _214_ (.A(_073_),
    .B(\main_reg[17] ),
    .Y(_091_));
 sky130_fd_sc_hd__o21ai_0 _215_ (.A1(_089_),
    .A2(_090_),
    .B1(_091_),
    .Y(_040_));
 sky130_fd_sc_hd__mux2i_1 _216_ (.A0(net107),
    .A1(net43),
    .S(_071_),
    .Y(_092_));
 sky130_fd_sc_hd__nand2_1 _217_ (.A(_073_),
    .B(\main_reg[18] ),
    .Y(_093_));
 sky130_fd_sc_hd__o21ai_0 _218_ (.A1(_089_),
    .A2(_092_),
    .B1(_093_),
    .Y(_041_));
 sky130_fd_sc_hd__buf_8 _219_ (.A(_070_),
    .X(_094_));
 sky130_fd_sc_hd__mux2i_1 _220_ (.A0(net108),
    .A1(net44),
    .S(_094_),
    .Y(_095_));
 sky130_fd_sc_hd__clkbuf_4 _221_ (.A(_068_),
    .X(_096_));
 sky130_fd_sc_hd__nand2_1 _222_ (.A(_096_),
    .B(\main_reg[19] ),
    .Y(_097_));
 sky130_fd_sc_hd__o21ai_0 _223_ (.A1(_089_),
    .A2(_095_),
    .B1(_097_),
    .Y(_042_));
 sky130_fd_sc_hd__mux2i_1 _224_ (.A0(net109),
    .A1(net45),
    .S(_094_),
    .Y(_098_));
 sky130_fd_sc_hd__nand2_1 _225_ (.A(_096_),
    .B(\main_reg[1] ),
    .Y(_099_));
 sky130_fd_sc_hd__o21ai_0 _226_ (.A1(_089_),
    .A2(_098_),
    .B1(_099_),
    .Y(_043_));
 sky130_fd_sc_hd__mux2i_1 _227_ (.A0(net110),
    .A1(net46),
    .S(_094_),
    .Y(_100_));
 sky130_fd_sc_hd__nand2_1 _228_ (.A(_096_),
    .B(\main_reg[20] ),
    .Y(_101_));
 sky130_fd_sc_hd__o21ai_0 _229_ (.A1(_089_),
    .A2(_100_),
    .B1(_101_),
    .Y(_044_));
 sky130_fd_sc_hd__mux2i_1 _230_ (.A0(net111),
    .A1(net47),
    .S(_094_),
    .Y(_102_));
 sky130_fd_sc_hd__nand2_1 _231_ (.A(_096_),
    .B(\main_reg[21] ),
    .Y(_103_));
 sky130_fd_sc_hd__o21ai_0 _232_ (.A1(_089_),
    .A2(_102_),
    .B1(_103_),
    .Y(_045_));
 sky130_fd_sc_hd__mux2i_1 _233_ (.A0(net112),
    .A1(net48),
    .S(_094_),
    .Y(_104_));
 sky130_fd_sc_hd__nand2_1 _234_ (.A(_096_),
    .B(\main_reg[22] ),
    .Y(_105_));
 sky130_fd_sc_hd__o21ai_0 _235_ (.A1(_089_),
    .A2(_104_),
    .B1(_105_),
    .Y(_046_));
 sky130_fd_sc_hd__mux2i_1 _236_ (.A0(net113),
    .A1(net49),
    .S(_094_),
    .Y(_106_));
 sky130_fd_sc_hd__nand2_1 _237_ (.A(_096_),
    .B(\main_reg[23] ),
    .Y(_107_));
 sky130_fd_sc_hd__o21ai_0 _238_ (.A1(_089_),
    .A2(_106_),
    .B1(_107_),
    .Y(_047_));
 sky130_fd_sc_hd__mux2i_1 _239_ (.A0(net114),
    .A1(net50),
    .S(_094_),
    .Y(_108_));
 sky130_fd_sc_hd__nand2_1 _240_ (.A(_096_),
    .B(\main_reg[24] ),
    .Y(_109_));
 sky130_fd_sc_hd__o21ai_0 _241_ (.A1(_089_),
    .A2(_108_),
    .B1(_109_),
    .Y(_048_));
 sky130_fd_sc_hd__mux2i_1 _242_ (.A0(net115),
    .A1(net51),
    .S(_094_),
    .Y(_110_));
 sky130_fd_sc_hd__nand2_1 _243_ (.A(_096_),
    .B(\main_reg[25] ),
    .Y(_111_));
 sky130_fd_sc_hd__o21ai_0 _244_ (.A1(_089_),
    .A2(_110_),
    .B1(_111_),
    .Y(_049_));
 sky130_fd_sc_hd__buf_2 _245_ (.A(_068_),
    .X(_112_));
 sky130_fd_sc_hd__mux2i_1 _246_ (.A0(net116),
    .A1(net52),
    .S(_094_),
    .Y(_113_));
 sky130_fd_sc_hd__nand2_1 _247_ (.A(_096_),
    .B(\main_reg[26] ),
    .Y(_114_));
 sky130_fd_sc_hd__o21ai_0 _248_ (.A1(_112_),
    .A2(_113_),
    .B1(_114_),
    .Y(_050_));
 sky130_fd_sc_hd__mux2i_1 _249_ (.A0(net117),
    .A1(net53),
    .S(_094_),
    .Y(_115_));
 sky130_fd_sc_hd__nand2_1 _250_ (.A(_096_),
    .B(\main_reg[27] ),
    .Y(_116_));
 sky130_fd_sc_hd__o21ai_0 _251_ (.A1(_112_),
    .A2(_115_),
    .B1(_116_),
    .Y(_051_));
 sky130_fd_sc_hd__buf_8 _252_ (.A(_070_),
    .X(_117_));
 sky130_fd_sc_hd__mux2i_1 _253_ (.A0(net118),
    .A1(net54),
    .S(_117_),
    .Y(_118_));
 sky130_fd_sc_hd__clkbuf_4 _254_ (.A(_068_),
    .X(_119_));
 sky130_fd_sc_hd__nand2_1 _255_ (.A(_119_),
    .B(\main_reg[28] ),
    .Y(_120_));
 sky130_fd_sc_hd__o21ai_0 _256_ (.A1(_112_),
    .A2(_118_),
    .B1(_120_),
    .Y(_052_));
 sky130_fd_sc_hd__mux2i_1 _257_ (.A0(net119),
    .A1(net55),
    .S(_117_),
    .Y(_121_));
 sky130_fd_sc_hd__nand2_1 _258_ (.A(_119_),
    .B(\main_reg[29] ),
    .Y(_122_));
 sky130_fd_sc_hd__o21ai_0 _259_ (.A1(_112_),
    .A2(_121_),
    .B1(_122_),
    .Y(_053_));
 sky130_fd_sc_hd__mux2i_1 _260_ (.A0(net120),
    .A1(net56),
    .S(_117_),
    .Y(_123_));
 sky130_fd_sc_hd__nand2_1 _261_ (.A(_119_),
    .B(\main_reg[2] ),
    .Y(_124_));
 sky130_fd_sc_hd__o21ai_0 _262_ (.A1(_112_),
    .A2(_123_),
    .B1(_124_),
    .Y(_054_));
 sky130_fd_sc_hd__mux2i_1 _263_ (.A0(net121),
    .A1(net57),
    .S(_117_),
    .Y(_125_));
 sky130_fd_sc_hd__nand2_1 _264_ (.A(_119_),
    .B(\main_reg[30] ),
    .Y(_126_));
 sky130_fd_sc_hd__o21ai_0 _265_ (.A1(_112_),
    .A2(_125_),
    .B1(_126_),
    .Y(_055_));
 sky130_fd_sc_hd__mux2i_1 _266_ (.A0(net122),
    .A1(net58),
    .S(_117_),
    .Y(_127_));
 sky130_fd_sc_hd__nand2_1 _267_ (.A(_119_),
    .B(\main_reg[31] ),
    .Y(_128_));
 sky130_fd_sc_hd__o21ai_0 _268_ (.A1(_112_),
    .A2(_127_),
    .B1(_128_),
    .Y(_056_));
 sky130_fd_sc_hd__mux2i_1 _269_ (.A0(net123),
    .A1(net59),
    .S(_117_),
    .Y(_129_));
 sky130_fd_sc_hd__nand2_1 _270_ (.A(_119_),
    .B(\main_reg[3] ),
    .Y(_130_));
 sky130_fd_sc_hd__o21ai_0 _271_ (.A1(_112_),
    .A2(_129_),
    .B1(_130_),
    .Y(_057_));
 sky130_fd_sc_hd__mux2i_1 _272_ (.A0(net124),
    .A1(net60),
    .S(_117_),
    .Y(_131_));
 sky130_fd_sc_hd__nand2_1 _273_ (.A(_119_),
    .B(\main_reg[4] ),
    .Y(_132_));
 sky130_fd_sc_hd__o21ai_0 _274_ (.A1(_112_),
    .A2(_131_),
    .B1(_132_),
    .Y(_058_));
 sky130_fd_sc_hd__mux2i_1 _275_ (.A0(net125),
    .A1(net61),
    .S(_117_),
    .Y(_133_));
 sky130_fd_sc_hd__nand2_1 _276_ (.A(_119_),
    .B(\main_reg[5] ),
    .Y(_134_));
 sky130_fd_sc_hd__o21ai_0 _277_ (.A1(_112_),
    .A2(_133_),
    .B1(_134_),
    .Y(_059_));
 sky130_fd_sc_hd__mux2i_1 _278_ (.A0(net126),
    .A1(net62),
    .S(_117_),
    .Y(_135_));
 sky130_fd_sc_hd__nand2_1 _279_ (.A(_119_),
    .B(\main_reg[6] ),
    .Y(_136_));
 sky130_fd_sc_hd__o21ai_0 _280_ (.A1(_068_),
    .A2(_135_),
    .B1(_136_),
    .Y(_060_));
 sky130_fd_sc_hd__mux2i_1 _281_ (.A0(net127),
    .A1(net63),
    .S(_117_),
    .Y(_137_));
 sky130_fd_sc_hd__nand2_1 _282_ (.A(_119_),
    .B(\main_reg[7] ),
    .Y(_138_));
 sky130_fd_sc_hd__o21ai_0 _283_ (.A1(_068_),
    .A2(_137_),
    .B1(_138_),
    .Y(_061_));
 sky130_fd_sc_hd__mux2i_1 _284_ (.A0(net128),
    .A1(net64),
    .S(_070_),
    .Y(_139_));
 sky130_fd_sc_hd__nand2_1 _285_ (.A(_069_),
    .B(\main_reg[8] ),
    .Y(_140_));
 sky130_fd_sc_hd__o21ai_0 _286_ (.A1(_068_),
    .A2(_139_),
    .B1(_140_),
    .Y(_062_));
 sky130_fd_sc_hd__mux2i_1 _287_ (.A0(net129),
    .A1(net65),
    .S(_070_),
    .Y(_141_));
 sky130_fd_sc_hd__nand2_1 _288_ (.A(_069_),
    .B(\main_reg[9] ),
    .Y(_142_));
 sky130_fd_sc_hd__o21ai_0 _289_ (.A1(_068_),
    .A2(_141_),
    .B1(_142_),
    .Y(_063_));
 sky130_fd_sc_hd__buf_6 _290_ (.A(use_shadow_out),
    .X(_143_));
 sky130_fd_sc_hd__buf_6 _291_ (.A(_143_),
    .X(_144_));
 sky130_fd_sc_hd__mux2_1 _292_ (.A0(\main_reg[0] ),
    .A1(net98),
    .S(_144_),
    .X(net66));
 sky130_fd_sc_hd__mux2_1 _293_ (.A0(\main_reg[10] ),
    .A1(net99),
    .S(_144_),
    .X(net67));
 sky130_fd_sc_hd__mux2_1 _294_ (.A0(\main_reg[11] ),
    .A1(net100),
    .S(_144_),
    .X(net68));
 sky130_fd_sc_hd__mux2_1 _295_ (.A0(\main_reg[12] ),
    .A1(net101),
    .S(_144_),
    .X(net69));
 sky130_fd_sc_hd__mux2_1 _296_ (.A0(\main_reg[13] ),
    .A1(net102),
    .S(_144_),
    .X(net70));
 sky130_fd_sc_hd__mux2_1 _297_ (.A0(\main_reg[14] ),
    .A1(net103),
    .S(_144_),
    .X(net71));
 sky130_fd_sc_hd__mux2_1 _298_ (.A0(\main_reg[15] ),
    .A1(net104),
    .S(_144_),
    .X(net72));
 sky130_fd_sc_hd__mux2_1 _299_ (.A0(\main_reg[16] ),
    .A1(net105),
    .S(_144_),
    .X(net73));
 sky130_fd_sc_hd__mux2_1 _300_ (.A0(\main_reg[17] ),
    .A1(net106),
    .S(_144_),
    .X(net74));
 sky130_fd_sc_hd__mux2_1 _301_ (.A0(\main_reg[18] ),
    .A1(net107),
    .S(_144_),
    .X(net75));
 sky130_fd_sc_hd__buf_6 _302_ (.A(_143_),
    .X(_145_));
 sky130_fd_sc_hd__mux2_1 _303_ (.A0(\main_reg[19] ),
    .A1(net108),
    .S(_145_),
    .X(net76));
 sky130_fd_sc_hd__mux2_1 _304_ (.A0(\main_reg[1] ),
    .A1(net109),
    .S(_145_),
    .X(net77));
 sky130_fd_sc_hd__mux2_1 _305_ (.A0(\main_reg[20] ),
    .A1(net110),
    .S(_145_),
    .X(net78));
 sky130_fd_sc_hd__mux2_1 _306_ (.A0(\main_reg[21] ),
    .A1(net111),
    .S(_145_),
    .X(net79));
 sky130_fd_sc_hd__mux2_1 _307_ (.A0(\main_reg[22] ),
    .A1(net112),
    .S(_145_),
    .X(net80));
 sky130_fd_sc_hd__mux2_1 _308_ (.A0(\main_reg[23] ),
    .A1(net113),
    .S(_145_),
    .X(net81));
 sky130_fd_sc_hd__mux2_1 _309_ (.A0(\main_reg[24] ),
    .A1(net114),
    .S(_145_),
    .X(net82));
 sky130_fd_sc_hd__mux2_1 _310_ (.A0(\main_reg[25] ),
    .A1(net115),
    .S(_145_),
    .X(net83));
 sky130_fd_sc_hd__mux2_1 _311_ (.A0(\main_reg[26] ),
    .A1(net116),
    .S(_145_),
    .X(net84));
 sky130_fd_sc_hd__mux2_1 _312_ (.A0(\main_reg[27] ),
    .A1(net117),
    .S(_145_),
    .X(net85));
 sky130_fd_sc_hd__buf_8 _313_ (.A(_143_),
    .X(_146_));
 sky130_fd_sc_hd__mux2_1 _314_ (.A0(\main_reg[28] ),
    .A1(net118),
    .S(_146_),
    .X(net86));
 sky130_fd_sc_hd__mux2_1 _315_ (.A0(\main_reg[29] ),
    .A1(net119),
    .S(_146_),
    .X(net87));
 sky130_fd_sc_hd__mux2_1 _316_ (.A0(\main_reg[2] ),
    .A1(net120),
    .S(_146_),
    .X(net88));
 sky130_fd_sc_hd__mux2_1 _317_ (.A0(\main_reg[30] ),
    .A1(net121),
    .S(_146_),
    .X(net89));
 sky130_fd_sc_hd__mux2_1 _318_ (.A0(\main_reg[31] ),
    .A1(net122),
    .S(_146_),
    .X(net90));
 sky130_fd_sc_hd__mux2_1 _319_ (.A0(\main_reg[3] ),
    .A1(net123),
    .S(_146_),
    .X(net91));
 sky130_fd_sc_hd__mux2_1 _320_ (.A0(\main_reg[4] ),
    .A1(net124),
    .S(_146_),
    .X(net92));
 sky130_fd_sc_hd__mux2_1 _321_ (.A0(\main_reg[5] ),
    .A1(net125),
    .S(_146_),
    .X(net93));
 sky130_fd_sc_hd__mux2_1 _322_ (.A0(\main_reg[6] ),
    .A1(net126),
    .S(_146_),
    .X(net94));
 sky130_fd_sc_hd__mux2_1 _323_ (.A0(\main_reg[7] ),
    .A1(net127),
    .S(_146_),
    .X(net95));
 sky130_fd_sc_hd__mux2_1 _324_ (.A0(\main_reg[8] ),
    .A1(net128),
    .S(_143_),
    .X(net96));
 sky130_fd_sc_hd__mux2_1 _325_ (.A0(\main_reg[9] ),
    .A1(net129),
    .S(_143_),
    .X(net97));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[0]$_DFFE_PN0P_  (.D(_000_),
    .Q(\main_reg[0] ),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[10]$_DFFE_PN0P_  (.D(_001_),
    .Q(\main_reg[10] ),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[11]$_DFFE_PN0P_  (.D(_002_),
    .Q(\main_reg[11] ),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[12]$_DFFE_PN0P_  (.D(_003_),
    .Q(\main_reg[12] ),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[13]$_DFFE_PN0P_  (.D(_004_),
    .Q(\main_reg[13] ),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[14]$_DFFE_PN0P_  (.D(_005_),
    .Q(\main_reg[14] ),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[15]$_DFFE_PN0P_  (.D(_006_),
    .Q(\main_reg[15] ),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[16]$_DFFE_PN0P_  (.D(_007_),
    .Q(\main_reg[16] ),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[17]$_DFFE_PN0P_  (.D(_008_),
    .Q(\main_reg[17] ),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[18]$_DFFE_PN0P_  (.D(_009_),
    .Q(\main_reg[18] ),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[19]$_DFFE_PN0P_  (.D(_010_),
    .Q(\main_reg[19] ),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[1]$_DFFE_PN0P_  (.D(_011_),
    .Q(\main_reg[1] ),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[20]$_DFFE_PN0P_  (.D(_012_),
    .Q(\main_reg[20] ),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[21]$_DFFE_PN0P_  (.D(_013_),
    .Q(\main_reg[21] ),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[22]$_DFFE_PN0P_  (.D(_014_),
    .Q(\main_reg[22] ),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[23]$_DFFE_PN0P_  (.D(_015_),
    .Q(\main_reg[23] ),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[24]$_DFFE_PN0P_  (.D(_016_),
    .Q(\main_reg[24] ),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[25]$_DFFE_PN0P_  (.D(_017_),
    .Q(\main_reg[25] ),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[26]$_DFFE_PN0P_  (.D(_018_),
    .Q(\main_reg[26] ),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[27]$_DFFE_PN0P_  (.D(_019_),
    .Q(\main_reg[27] ),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[28]$_DFFE_PN0P_  (.D(_020_),
    .Q(\main_reg[28] ),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[29]$_DFFE_PN0P_  (.D(_021_),
    .Q(\main_reg[29] ),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[2]$_DFFE_PN0P_  (.D(_022_),
    .Q(\main_reg[2] ),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[30]$_DFFE_PN0P_  (.D(_023_),
    .Q(\main_reg[30] ),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[31]$_DFFE_PN0P_  (.D(_024_),
    .Q(\main_reg[31] ),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[3]$_DFFE_PN0P_  (.D(_025_),
    .Q(\main_reg[3] ),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[4]$_DFFE_PN0P_  (.D(_026_),
    .Q(\main_reg[4] ),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[5]$_DFFE_PN0P_  (.D(_027_),
    .Q(\main_reg[5] ),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[6]$_DFFE_PN0P_  (.D(_028_),
    .Q(\main_reg[6] ),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[7]$_DFFE_PN0P_  (.D(_029_),
    .Q(\main_reg[7] ),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[8]$_DFFE_PN0P_  (.D(_030_),
    .Q(\main_reg[8] ),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \main_reg[9]$_DFFE_PN0P_  (.D(_031_),
    .Q(\main_reg[9] ),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[0]$_DFFE_PN0P_  (.D(_032_),
    .Q(net98),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[10]$_DFFE_PN0P_  (.D(_033_),
    .Q(net99),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[11]$_DFFE_PN0P_  (.D(_034_),
    .Q(net100),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[12]$_DFFE_PN0P_  (.D(_035_),
    .Q(net101),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[13]$_DFFE_PN0P_  (.D(_036_),
    .Q(net102),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[14]$_DFFE_PN0P_  (.D(_037_),
    .Q(net103),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[15]$_DFFE_PN0P_  (.D(_038_),
    .Q(net104),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[16]$_DFFE_PN0P_  (.D(_039_),
    .Q(net105),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[17]$_DFFE_PN0P_  (.D(_040_),
    .Q(net106),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[18]$_DFFE_PN0P_  (.D(_041_),
    .Q(net107),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[19]$_DFFE_PN0P_  (.D(_042_),
    .Q(net108),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[1]$_DFFE_PN0P_  (.D(_043_),
    .Q(net109),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[20]$_DFFE_PN0P_  (.D(_044_),
    .Q(net110),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[21]$_DFFE_PN0P_  (.D(_045_),
    .Q(net111),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[22]$_DFFE_PN0P_  (.D(_046_),
    .Q(net112),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[23]$_DFFE_PN0P_  (.D(_047_),
    .Q(net113),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[24]$_DFFE_PN0P_  (.D(_048_),
    .Q(net114),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[25]$_DFFE_PN0P_  (.D(_049_),
    .Q(net115),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[26]$_DFFE_PN0P_  (.D(_050_),
    .Q(net116),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[27]$_DFFE_PN0P_  (.D(_051_),
    .Q(net117),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[28]$_DFFE_PN0P_  (.D(_052_),
    .Q(net118),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[29]$_DFFE_PN0P_  (.D(_053_),
    .Q(net119),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[2]$_DFFE_PN0P_  (.D(_054_),
    .Q(net120),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[30]$_DFFE_PN0P_  (.D(_055_),
    .Q(net121),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[31]$_DFFE_PN0P_  (.D(_056_),
    .Q(net122),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[3]$_DFFE_PN0P_  (.D(_057_),
    .Q(net123),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[4]$_DFFE_PN0P_  (.D(_058_),
    .Q(net124),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[5]$_DFFE_PN0P_  (.D(_059_),
    .Q(net125),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[6]$_DFFE_PN0P_  (.D(_060_),
    .Q(net126),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[7]$_DFFE_PN0P_  (.D(_061_),
    .Q(net127),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[8]$_DFFE_PN0P_  (.D(_062_),
    .Q(net128),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shadow_reg[9]$_DFFE_PN0P_  (.D(_063_),
    .Q(net129),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__buf_16 hold1 (.A(net130),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_74 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(main_data_in[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(main_data_in[10]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(main_data_in[11]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(main_data_in[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(main_data_in[13]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(main_data_in[14]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(main_data_in[15]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(main_data_in[16]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(main_data_in[17]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(main_data_in[18]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(main_data_in[19]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(main_data_in[1]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(main_data_in[20]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(main_data_in[21]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(main_data_in[22]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(main_data_in[23]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(main_data_in[24]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(main_data_in[25]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(main_data_in[26]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(main_data_in[27]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(main_data_in[28]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(main_data_in[29]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(main_data_in[2]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(main_data_in[30]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(main_data_in[31]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(main_data_in[3]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(main_data_in[4]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(main_data_in[5]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(main_data_in[6]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(main_data_in[7]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(main_data_in[8]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(main_data_in[9]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(shadow_data_in[0]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(shadow_data_in[10]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(shadow_data_in[11]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(shadow_data_in[12]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(shadow_data_in[13]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(shadow_data_in[14]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(shadow_data_in[15]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(shadow_data_in[16]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(shadow_data_in[17]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(shadow_data_in[18]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(shadow_data_in[19]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(shadow_data_in[1]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(shadow_data_in[20]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(shadow_data_in[21]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(shadow_data_in[22]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(shadow_data_in[23]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(shadow_data_in[24]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(shadow_data_in[25]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(shadow_data_in[26]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(shadow_data_in[27]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(shadow_data_in[28]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(shadow_data_in[29]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(shadow_data_in[2]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(shadow_data_in[30]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(shadow_data_in[31]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(shadow_data_in[3]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(shadow_data_in[4]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(shadow_data_in[5]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(shadow_data_in[6]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(shadow_data_in[7]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(shadow_data_in[8]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(shadow_data_in[9]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 output65 (.A(net66),
    .X(main_data_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output66 (.A(net67),
    .X(main_data_out[10]));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net68),
    .X(main_data_out[11]));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net69),
    .X(main_data_out[12]));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(net70),
    .X(main_data_out[13]));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net71),
    .X(main_data_out[14]));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(net72),
    .X(main_data_out[15]));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(net73),
    .X(main_data_out[16]));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(net74),
    .X(main_data_out[17]));
 sky130_fd_sc_hd__clkbuf_1 output74 (.A(net75),
    .X(main_data_out[18]));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(net76),
    .X(main_data_out[19]));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(net77),
    .X(main_data_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output77 (.A(net78),
    .X(main_data_out[20]));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(net79),
    .X(main_data_out[21]));
 sky130_fd_sc_hd__clkbuf_1 output79 (.A(net80),
    .X(main_data_out[22]));
 sky130_fd_sc_hd__clkbuf_1 output80 (.A(net81),
    .X(main_data_out[23]));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(net82),
    .X(main_data_out[24]));
 sky130_fd_sc_hd__clkbuf_1 output82 (.A(net83),
    .X(main_data_out[25]));
 sky130_fd_sc_hd__clkbuf_1 output83 (.A(net84),
    .X(main_data_out[26]));
 sky130_fd_sc_hd__clkbuf_1 output84 (.A(net85),
    .X(main_data_out[27]));
 sky130_fd_sc_hd__clkbuf_1 output85 (.A(net86),
    .X(main_data_out[28]));
 sky130_fd_sc_hd__clkbuf_1 output86 (.A(net87),
    .X(main_data_out[29]));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(net88),
    .X(main_data_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output88 (.A(net89),
    .X(main_data_out[30]));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(net90),
    .X(main_data_out[31]));
 sky130_fd_sc_hd__clkbuf_1 output90 (.A(net91),
    .X(main_data_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output91 (.A(net92),
    .X(main_data_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output92 (.A(net93),
    .X(main_data_out[5]));
 sky130_fd_sc_hd__clkbuf_1 output93 (.A(net94),
    .X(main_data_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output94 (.A(net95),
    .X(main_data_out[7]));
 sky130_fd_sc_hd__clkbuf_1 output95 (.A(net96),
    .X(main_data_out[8]));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(net97),
    .X(main_data_out[9]));
 sky130_fd_sc_hd__clkbuf_1 output97 (.A(net98),
    .X(shadow_data_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output98 (.A(net99),
    .X(shadow_data_out[10]));
 sky130_fd_sc_hd__clkbuf_1 output99 (.A(net100),
    .X(shadow_data_out[11]));
 sky130_fd_sc_hd__clkbuf_1 output100 (.A(net101),
    .X(shadow_data_out[12]));
 sky130_fd_sc_hd__clkbuf_1 output101 (.A(net102),
    .X(shadow_data_out[13]));
 sky130_fd_sc_hd__clkbuf_1 output102 (.A(net103),
    .X(shadow_data_out[14]));
 sky130_fd_sc_hd__clkbuf_1 output103 (.A(net104),
    .X(shadow_data_out[15]));
 sky130_fd_sc_hd__clkbuf_1 output104 (.A(net105),
    .X(shadow_data_out[16]));
 sky130_fd_sc_hd__clkbuf_1 output105 (.A(net106),
    .X(shadow_data_out[17]));
 sky130_fd_sc_hd__clkbuf_1 output106 (.A(net107),
    .X(shadow_data_out[18]));
 sky130_fd_sc_hd__clkbuf_1 output107 (.A(net108),
    .X(shadow_data_out[19]));
 sky130_fd_sc_hd__clkbuf_1 output108 (.A(net109),
    .X(shadow_data_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(net110),
    .X(shadow_data_out[20]));
 sky130_fd_sc_hd__clkbuf_1 output110 (.A(net111),
    .X(shadow_data_out[21]));
 sky130_fd_sc_hd__clkbuf_1 output111 (.A(net112),
    .X(shadow_data_out[22]));
 sky130_fd_sc_hd__clkbuf_1 output112 (.A(net113),
    .X(shadow_data_out[23]));
 sky130_fd_sc_hd__clkbuf_1 output113 (.A(net114),
    .X(shadow_data_out[24]));
 sky130_fd_sc_hd__clkbuf_1 output114 (.A(net115),
    .X(shadow_data_out[25]));
 sky130_fd_sc_hd__clkbuf_1 output115 (.A(net116),
    .X(shadow_data_out[26]));
 sky130_fd_sc_hd__clkbuf_1 output116 (.A(net117),
    .X(shadow_data_out[27]));
 sky130_fd_sc_hd__clkbuf_1 output117 (.A(net118),
    .X(shadow_data_out[28]));
 sky130_fd_sc_hd__clkbuf_1 output118 (.A(net119),
    .X(shadow_data_out[29]));
 sky130_fd_sc_hd__clkbuf_1 output119 (.A(net120),
    .X(shadow_data_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output120 (.A(net121),
    .X(shadow_data_out[30]));
 sky130_fd_sc_hd__clkbuf_1 output121 (.A(net122),
    .X(shadow_data_out[31]));
 sky130_fd_sc_hd__clkbuf_1 output122 (.A(net123),
    .X(shadow_data_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output123 (.A(net124),
    .X(shadow_data_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output124 (.A(net125),
    .X(shadow_data_out[5]));
 sky130_fd_sc_hd__clkbuf_1 output125 (.A(net126),
    .X(shadow_data_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output126 (.A(net127),
    .X(shadow_data_out[7]));
 sky130_fd_sc_hd__clkbuf_1 output127 (.A(net128),
    .X(shadow_data_out[8]));
 sky130_fd_sc_hd__clkbuf_1 output128 (.A(net129),
    .X(shadow_data_out[9]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload0 (.A(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload1 (.A(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload2 (.A(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload3 (.A(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload4 (.A(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net130));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_134 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_140 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_54 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_92 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_36 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_168 ();
endmodule
