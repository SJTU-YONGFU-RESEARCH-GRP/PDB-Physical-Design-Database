module configurable_param_fifo (almost_empty,
    almost_full,
    clk,
    empty,
    full,
    rd_en,
    rst_n,
    wr_en,
    rd_data,
    wr_data);
 output almost_empty;
 output almost_full;
 input clk;
 output empty;
 output full;
 input rd_en;
 input rst_n;
 input wr_en;
 output [7:0] rd_data;
 input [7:0] wr_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire \mem[0][0] ;
 wire \mem[0][1] ;
 wire \mem[0][2] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[10][0] ;
 wire \mem[10][1] ;
 wire \mem[10][2] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[11][0] ;
 wire \mem[11][1] ;
 wire \mem[11][2] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[12][0] ;
 wire \mem[12][1] ;
 wire \mem[12][2] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[13][0] ;
 wire \mem[13][1] ;
 wire \mem[13][2] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[14][0] ;
 wire \mem[14][1] ;
 wire \mem[14][2] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[15][0] ;
 wire \mem[15][1] ;
 wire \mem[15][2] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[1][0] ;
 wire \mem[1][1] ;
 wire \mem[1][2] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[2][0] ;
 wire \mem[2][1] ;
 wire \mem[2][2] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[3][0] ;
 wire \mem[3][1] ;
 wire \mem[3][2] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[4][0] ;
 wire \mem[4][1] ;
 wire \mem[4][2] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[5][0] ;
 wire \mem[5][1] ;
 wire \mem[5][2] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[6][0] ;
 wire \mem[6][1] ;
 wire \mem[6][2] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[7][0] ;
 wire \mem[7][1] ;
 wire \mem[7][2] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[8][0] ;
 wire \mem[8][1] ;
 wire \mem[8][2] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[9][0] ;
 wire \mem[9][1] ;
 wire \mem[9][2] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \rd_addr[0] ;
 wire \rd_addr[1] ;
 wire \rd_addr[2] ;
 wire \rd_addr[3] ;
 wire \rd_data_reg[0] ;
 wire \rd_data_reg[1] ;
 wire \rd_data_reg[2] ;
 wire \rd_data_reg[3] ;
 wire \rd_data_reg[4] ;
 wire \rd_data_reg[5] ;
 wire \rd_data_reg[6] ;
 wire \rd_data_reg[7] ;
 wire \rd_ptr[4] ;
 wire rd_valid;
 wire \wr_addr[0] ;
 wire \wr_addr[1] ;
 wire \wr_addr[2] ;
 wire \wr_addr[3] ;
 wire \wr_ptr[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;

 sky130_fd_sc_hd__xor2_1 _204_ (.A(\wr_ptr[4] ),
    .B(\rd_ptr[4] ),
    .X(_040_));
 sky130_fd_sc_hd__nand4_1 _205_ (.A(_194_),
    .B(_189_),
    .C(_192_),
    .D(_186_),
    .Y(_041_));
 sky130_fd_sc_hd__nor2_1 _206_ (.A(_040_),
    .B(_041_),
    .Y(net15));
 sky130_fd_sc_hd__and2b_1 _207_ (.A_N(_041_),
    .B(_040_),
    .X(net16));
 sky130_fd_sc_hd__nor2b_1 _208_ (.A(net15),
    .B_N(net2),
    .Y(_042_));
 sky130_fd_sc_hd__buf_2 _209_ (.A(_042_),
    .X(_000_));
 sky130_fd_sc_hd__clkbuf_8 _210_ (.A(\wr_addr[3] ),
    .X(_043_));
 sky130_fd_sc_hd__buf_6 _211_ (.A(\wr_addr[2] ),
    .X(_044_));
 sky130_fd_sc_hd__nor2b_1 _212_ (.A(net16),
    .B_N(net12),
    .Y(_045_));
 sky130_fd_sc_hd__buf_4 _213_ (.A(_045_),
    .X(_046_));
 sky130_fd_sc_hd__nand2_4 _214_ (.A(_197_),
    .B(_046_),
    .Y(_047_));
 sky130_fd_sc_hd__nor3_4 _215_ (.A(_043_),
    .B(_044_),
    .C(_047_),
    .Y(_001_));
 sky130_fd_sc_hd__nand2_4 _216_ (.A(_200_),
    .B(_046_),
    .Y(_048_));
 sky130_fd_sc_hd__nor3_4 _217_ (.A(_043_),
    .B(_044_),
    .C(_048_),
    .Y(_008_));
 sky130_fd_sc_hd__nand2_4 _218_ (.A(_198_),
    .B(_046_),
    .Y(_049_));
 sky130_fd_sc_hd__nor3_4 _219_ (.A(_043_),
    .B(_044_),
    .C(_049_),
    .Y(_009_));
 sky130_fd_sc_hd__nand2_4 _220_ (.A(_202_),
    .B(_046_),
    .Y(_050_));
 sky130_fd_sc_hd__nor3_4 _221_ (.A(_043_),
    .B(_044_),
    .C(_050_),
    .Y(_010_));
 sky130_fd_sc_hd__nand2b_4 _222_ (.A_N(_043_),
    .B(_044_),
    .Y(_051_));
 sky130_fd_sc_hd__nor2_4 _223_ (.A(_047_),
    .B(_051_),
    .Y(_011_));
 sky130_fd_sc_hd__nor2_4 _224_ (.A(_048_),
    .B(_051_),
    .Y(_012_));
 sky130_fd_sc_hd__nor2_4 _225_ (.A(_049_),
    .B(_051_),
    .Y(_013_));
 sky130_fd_sc_hd__nor2_4 _226_ (.A(_050_),
    .B(_051_),
    .Y(_014_));
 sky130_fd_sc_hd__nand2b_4 _227_ (.A_N(_044_),
    .B(_043_),
    .Y(_052_));
 sky130_fd_sc_hd__nor2_4 _228_ (.A(_047_),
    .B(_052_),
    .Y(_015_));
 sky130_fd_sc_hd__nor2_4 _229_ (.A(_048_),
    .B(_052_),
    .Y(_016_));
 sky130_fd_sc_hd__nor2_4 _230_ (.A(_049_),
    .B(_052_),
    .Y(_002_));
 sky130_fd_sc_hd__nor2_4 _231_ (.A(_050_),
    .B(_052_),
    .Y(_003_));
 sky130_fd_sc_hd__nand2_2 _232_ (.A(_043_),
    .B(_044_),
    .Y(_053_));
 sky130_fd_sc_hd__nor2_4 _233_ (.A(_047_),
    .B(_053_),
    .Y(_004_));
 sky130_fd_sc_hd__nor2_4 _234_ (.A(_048_),
    .B(_053_),
    .Y(_005_));
 sky130_fd_sc_hd__nor2_4 _235_ (.A(_049_),
    .B(_053_),
    .Y(_006_));
 sky130_fd_sc_hd__nand4_2 _236_ (.A(_043_),
    .B(_044_),
    .C(_202_),
    .D(_046_),
    .Y(_054_));
 sky130_fd_sc_hd__clkinv_4 _237_ (.A(_054_),
    .Y(_007_));
 sky130_fd_sc_hd__buf_6 _238_ (.A(\rd_addr[1] ),
    .X(_055_));
 sky130_fd_sc_hd__buf_6 _239_ (.A(_055_),
    .X(_056_));
 sky130_fd_sc_hd__buf_4 _240_ (.A(_056_),
    .X(_057_));
 sky130_fd_sc_hd__inv_1 _241_ (.A(_057_),
    .Y(_181_));
 sky130_fd_sc_hd__buf_4 _242_ (.A(\rd_addr[3] ),
    .X(_058_));
 sky130_fd_sc_hd__inv_2 _243_ (.A(_058_),
    .Y(_187_));
 sky130_fd_sc_hd__inv_2 _244_ (.A(\rd_addr[2] ),
    .Y(_190_));
 sky130_fd_sc_hd__inv_1 _245_ (.A(_193_),
    .Y(_182_));
 sky130_fd_sc_hd__clkinvlp_4 _246_ (.A(\wr_addr[0] ),
    .Y(_018_));
 sky130_fd_sc_hd__inv_1 _247_ (.A(\wr_addr[1] ),
    .Y(_196_));
 sky130_fd_sc_hd__xnor2_1 _248_ (.A(_192_),
    .B(_183_),
    .Y(_059_));
 sky130_fd_sc_hd__inv_1 _249_ (.A(_194_),
    .Y(_060_));
 sky130_fd_sc_hd__inv_1 _250_ (.A(net13),
    .Y(_061_));
 sky130_fd_sc_hd__nand3_1 _251_ (.A(_060_),
    .B(_184_),
    .C(_061_),
    .Y(_062_));
 sky130_fd_sc_hd__a21o_1 _252_ (.A1(_182_),
    .A2(_186_),
    .B1(_185_),
    .X(_063_));
 sky130_fd_sc_hd__a21oi_1 _253_ (.A1(_192_),
    .A2(_063_),
    .B1(_191_),
    .Y(_064_));
 sky130_fd_sc_hd__xor2_1 _254_ (.A(_189_),
    .B(_064_),
    .X(_065_));
 sky130_fd_sc_hd__a21o_1 _255_ (.A1(_192_),
    .A2(_183_),
    .B1(_191_),
    .X(_066_));
 sky130_fd_sc_hd__a21oi_1 _256_ (.A1(_189_),
    .A2(_066_),
    .B1(_188_),
    .Y(_067_));
 sky130_fd_sc_hd__xnor2_1 _257_ (.A(_040_),
    .B(_067_),
    .Y(_068_));
 sky130_fd_sc_hd__a41o_1 _258_ (.A1(_059_),
    .A2(_062_),
    .A3(_065_),
    .A4(_068_),
    .B1(net15),
    .X(_020_));
 sky130_fd_sc_hd__a21oi_1 _259_ (.A1(_060_),
    .A2(net14),
    .B1(_184_),
    .Y(_069_));
 sky130_fd_sc_hd__nor2b_1 _260_ (.A(net16),
    .B_N(_068_),
    .Y(_070_));
 sky130_fd_sc_hd__o31ai_1 _261_ (.A1(_059_),
    .A2(_065_),
    .A3(_069_),
    .B1(_070_),
    .Y(_021_));
 sky130_fd_sc_hd__buf_8 _262_ (.A(_055_),
    .X(_071_));
 sky130_fd_sc_hd__buf_4 _263_ (.A(\rd_addr[2] ),
    .X(_072_));
 sky130_fd_sc_hd__mux4_1 _264_ (.A0(\mem[1][0] ),
    .A1(\mem[3][0] ),
    .A2(\mem[5][0] ),
    .A3(\mem[7][0] ),
    .S0(_071_),
    .S1(_072_),
    .X(_073_));
 sky130_fd_sc_hd__buf_6 _265_ (.A(\rd_addr[0] ),
    .X(_074_));
 sky130_fd_sc_hd__nor2b_1 _266_ (.A(_058_),
    .B_N(_074_),
    .Y(_075_));
 sky130_fd_sc_hd__clkbuf_4 _267_ (.A(_075_),
    .X(_076_));
 sky130_fd_sc_hd__nor2_4 _268_ (.A(_074_),
    .B(_058_),
    .Y(_077_));
 sky130_fd_sc_hd__mux4_1 _269_ (.A0(\mem[0][0] ),
    .A1(\mem[2][0] ),
    .A2(\mem[4][0] ),
    .A3(\mem[6][0] ),
    .S0(_071_),
    .S1(_072_),
    .X(_078_));
 sky130_fd_sc_hd__a22oi_2 _270_ (.A1(_073_),
    .A2(_076_),
    .B1(_077_),
    .B2(_078_),
    .Y(_079_));
 sky130_fd_sc_hd__nand3_4 _271_ (.A(_074_),
    .B(_072_),
    .C(_058_),
    .Y(_080_));
 sky130_fd_sc_hd__buf_6 _272_ (.A(_056_),
    .X(_081_));
 sky130_fd_sc_hd__mux2i_1 _273_ (.A0(\mem[13][0] ),
    .A1(\mem[15][0] ),
    .S(_081_),
    .Y(_082_));
 sky130_fd_sc_hd__or3_1 _274_ (.A(_074_),
    .B(\rd_addr[2] ),
    .C(_187_),
    .X(_083_));
 sky130_fd_sc_hd__buf_2 _275_ (.A(_083_),
    .X(_084_));
 sky130_fd_sc_hd__mux2i_1 _276_ (.A0(\mem[8][0] ),
    .A1(\mem[10][0] ),
    .S(_057_),
    .Y(_085_));
 sky130_fd_sc_hd__o22ai_1 _277_ (.A1(_080_),
    .A2(_082_),
    .B1(_084_),
    .B2(_085_),
    .Y(_086_));
 sky130_fd_sc_hd__or3_1 _278_ (.A(_074_),
    .B(_190_),
    .C(_187_),
    .X(_087_));
 sky130_fd_sc_hd__clkbuf_4 _279_ (.A(_087_),
    .X(_088_));
 sky130_fd_sc_hd__buf_6 _280_ (.A(_056_),
    .X(_089_));
 sky130_fd_sc_hd__mux2i_1 _281_ (.A0(\mem[12][0] ),
    .A1(\mem[14][0] ),
    .S(_089_),
    .Y(_090_));
 sky130_fd_sc_hd__nand3_4 _282_ (.A(_074_),
    .B(_190_),
    .C(_058_),
    .Y(_091_));
 sky130_fd_sc_hd__mux2i_1 _283_ (.A0(\mem[9][0] ),
    .A1(\mem[11][0] ),
    .S(_057_),
    .Y(_092_));
 sky130_fd_sc_hd__o22ai_1 _284_ (.A1(_088_),
    .A2(_090_),
    .B1(_091_),
    .B2(_092_),
    .Y(_093_));
 sky130_fd_sc_hd__nor2_1 _285_ (.A(_086_),
    .B(_093_),
    .Y(_094_));
 sky130_fd_sc_hd__buf_4 _286_ (.A(_042_),
    .X(_095_));
 sky130_fd_sc_hd__nor2_1 _287_ (.A(\rd_data_reg[0] ),
    .B(_095_),
    .Y(_096_));
 sky130_fd_sc_hd__a31oi_1 _288_ (.A1(_000_),
    .A2(_079_),
    .A3(_094_),
    .B1(_096_),
    .Y(_022_));
 sky130_fd_sc_hd__mux4_1 _289_ (.A0(\mem[1][1] ),
    .A1(\mem[3][1] ),
    .A2(\mem[5][1] ),
    .A3(\mem[7][1] ),
    .S0(_071_),
    .S1(_072_),
    .X(_097_));
 sky130_fd_sc_hd__buf_4 _290_ (.A(\rd_addr[2] ),
    .X(_098_));
 sky130_fd_sc_hd__mux4_1 _291_ (.A0(\mem[0][1] ),
    .A1(\mem[2][1] ),
    .A2(\mem[4][1] ),
    .A3(\mem[6][1] ),
    .S0(_056_),
    .S1(_098_),
    .X(_099_));
 sky130_fd_sc_hd__a22oi_2 _292_ (.A1(_076_),
    .A2(_097_),
    .B1(_099_),
    .B2(_077_),
    .Y(_100_));
 sky130_fd_sc_hd__mux2i_1 _293_ (.A0(\mem[12][1] ),
    .A1(\mem[14][1] ),
    .S(_081_),
    .Y(_101_));
 sky130_fd_sc_hd__mux2i_1 _294_ (.A0(\mem[9][1] ),
    .A1(\mem[11][1] ),
    .S(_089_),
    .Y(_102_));
 sky130_fd_sc_hd__o22ai_2 _295_ (.A1(_088_),
    .A2(_101_),
    .B1(_102_),
    .B2(_091_),
    .Y(_103_));
 sky130_fd_sc_hd__mux2i_1 _296_ (.A0(\mem[8][1] ),
    .A1(\mem[10][1] ),
    .S(_089_),
    .Y(_104_));
 sky130_fd_sc_hd__mux2i_1 _297_ (.A0(\mem[13][1] ),
    .A1(\mem[15][1] ),
    .S(_057_),
    .Y(_105_));
 sky130_fd_sc_hd__o22ai_1 _298_ (.A1(_084_),
    .A2(_104_),
    .B1(_105_),
    .B2(_080_),
    .Y(_106_));
 sky130_fd_sc_hd__nor2_1 _299_ (.A(_103_),
    .B(_106_),
    .Y(_107_));
 sky130_fd_sc_hd__nor2_1 _300_ (.A(\rd_data_reg[1] ),
    .B(_095_),
    .Y(_108_));
 sky130_fd_sc_hd__a31oi_1 _301_ (.A1(_000_),
    .A2(_100_),
    .A3(_107_),
    .B1(_108_),
    .Y(_023_));
 sky130_fd_sc_hd__mux4_1 _302_ (.A0(\mem[1][2] ),
    .A1(\mem[3][2] ),
    .A2(\mem[5][2] ),
    .A3(\mem[7][2] ),
    .S0(_071_),
    .S1(_072_),
    .X(_109_));
 sky130_fd_sc_hd__mux4_1 _303_ (.A0(\mem[0][2] ),
    .A1(\mem[2][2] ),
    .A2(\mem[4][2] ),
    .A3(\mem[6][2] ),
    .S0(_056_),
    .S1(_098_),
    .X(_110_));
 sky130_fd_sc_hd__a22oi_2 _304_ (.A1(_076_),
    .A2(_109_),
    .B1(_110_),
    .B2(_077_),
    .Y(_111_));
 sky130_fd_sc_hd__mux2i_1 _305_ (.A0(\mem[12][2] ),
    .A1(\mem[14][2] ),
    .S(_081_),
    .Y(_112_));
 sky130_fd_sc_hd__mux2i_2 _306_ (.A0(\mem[9][2] ),
    .A1(\mem[11][2] ),
    .S(_081_),
    .Y(_113_));
 sky130_fd_sc_hd__o22ai_2 _307_ (.A1(_088_),
    .A2(_112_),
    .B1(_113_),
    .B2(_091_),
    .Y(_114_));
 sky130_fd_sc_hd__mux2i_1 _308_ (.A0(\mem[8][2] ),
    .A1(\mem[10][2] ),
    .S(_089_),
    .Y(_115_));
 sky130_fd_sc_hd__mux2i_1 _309_ (.A0(\mem[13][2] ),
    .A1(\mem[15][2] ),
    .S(_057_),
    .Y(_116_));
 sky130_fd_sc_hd__o22ai_1 _310_ (.A1(_084_),
    .A2(_115_),
    .B1(_116_),
    .B2(_080_),
    .Y(_117_));
 sky130_fd_sc_hd__nor2_1 _311_ (.A(_114_),
    .B(_117_),
    .Y(_118_));
 sky130_fd_sc_hd__nor2_1 _312_ (.A(\rd_data_reg[2] ),
    .B(_095_),
    .Y(_119_));
 sky130_fd_sc_hd__a31oi_1 _313_ (.A1(_000_),
    .A2(_111_),
    .A3(_118_),
    .B1(_119_),
    .Y(_024_));
 sky130_fd_sc_hd__mux4_1 _314_ (.A0(\mem[1][3] ),
    .A1(\mem[3][3] ),
    .A2(\mem[5][3] ),
    .A3(\mem[7][3] ),
    .S0(_071_),
    .S1(_072_),
    .X(_120_));
 sky130_fd_sc_hd__mux4_1 _315_ (.A0(\mem[0][3] ),
    .A1(\mem[2][3] ),
    .A2(\mem[4][3] ),
    .A3(\mem[6][3] ),
    .S0(_056_),
    .S1(_098_),
    .X(_121_));
 sky130_fd_sc_hd__a22oi_1 _316_ (.A1(_076_),
    .A2(_120_),
    .B1(_121_),
    .B2(_077_),
    .Y(_122_));
 sky130_fd_sc_hd__mux2i_1 _317_ (.A0(\mem[12][3] ),
    .A1(\mem[14][3] ),
    .S(_081_),
    .Y(_123_));
 sky130_fd_sc_hd__mux2i_1 _318_ (.A0(\mem[9][3] ),
    .A1(\mem[11][3] ),
    .S(_081_),
    .Y(_124_));
 sky130_fd_sc_hd__o22ai_2 _319_ (.A1(_088_),
    .A2(_123_),
    .B1(_124_),
    .B2(_091_),
    .Y(_125_));
 sky130_fd_sc_hd__mux2i_2 _320_ (.A0(\mem[8][3] ),
    .A1(\mem[10][3] ),
    .S(_089_),
    .Y(_126_));
 sky130_fd_sc_hd__mux2i_1 _321_ (.A0(\mem[13][3] ),
    .A1(\mem[15][3] ),
    .S(_057_),
    .Y(_127_));
 sky130_fd_sc_hd__o22ai_1 _322_ (.A1(_084_),
    .A2(_126_),
    .B1(_127_),
    .B2(_080_),
    .Y(_128_));
 sky130_fd_sc_hd__nor2_1 _323_ (.A(_125_),
    .B(_128_),
    .Y(_129_));
 sky130_fd_sc_hd__nor2_1 _324_ (.A(\rd_data_reg[3] ),
    .B(_095_),
    .Y(_130_));
 sky130_fd_sc_hd__a31oi_1 _325_ (.A1(_000_),
    .A2(_122_),
    .A3(_129_),
    .B1(_130_),
    .Y(_025_));
 sky130_fd_sc_hd__mux4_1 _326_ (.A0(\mem[1][4] ),
    .A1(\mem[3][4] ),
    .A2(\mem[5][4] ),
    .A3(\mem[7][4] ),
    .S0(_071_),
    .S1(_072_),
    .X(_131_));
 sky130_fd_sc_hd__mux4_1 _327_ (.A0(\mem[0][4] ),
    .A1(\mem[2][4] ),
    .A2(\mem[4][4] ),
    .A3(\mem[6][4] ),
    .S0(_071_),
    .S1(_098_),
    .X(_132_));
 sky130_fd_sc_hd__a22oi_2 _328_ (.A1(_076_),
    .A2(_131_),
    .B1(_132_),
    .B2(_077_),
    .Y(_133_));
 sky130_fd_sc_hd__mux2i_1 _329_ (.A0(\mem[12][4] ),
    .A1(\mem[14][4] ),
    .S(_056_),
    .Y(_134_));
 sky130_fd_sc_hd__mux2i_1 _330_ (.A0(\mem[9][4] ),
    .A1(\mem[11][4] ),
    .S(_081_),
    .Y(_135_));
 sky130_fd_sc_hd__o22ai_2 _331_ (.A1(_088_),
    .A2(_134_),
    .B1(_135_),
    .B2(_091_),
    .Y(_136_));
 sky130_fd_sc_hd__mux2i_1 _332_ (.A0(\mem[8][4] ),
    .A1(\mem[10][4] ),
    .S(_089_),
    .Y(_137_));
 sky130_fd_sc_hd__mux2i_1 _333_ (.A0(\mem[13][4] ),
    .A1(\mem[15][4] ),
    .S(_057_),
    .Y(_138_));
 sky130_fd_sc_hd__o22ai_1 _334_ (.A1(_084_),
    .A2(_137_),
    .B1(_138_),
    .B2(_080_),
    .Y(_139_));
 sky130_fd_sc_hd__nor2_1 _335_ (.A(_136_),
    .B(_139_),
    .Y(_140_));
 sky130_fd_sc_hd__nor2_1 _336_ (.A(\rd_data_reg[4] ),
    .B(_095_),
    .Y(_141_));
 sky130_fd_sc_hd__a31oi_1 _337_ (.A1(_000_),
    .A2(_133_),
    .A3(_140_),
    .B1(_141_),
    .Y(_026_));
 sky130_fd_sc_hd__mux4_1 _338_ (.A0(\mem[1][5] ),
    .A1(\mem[3][5] ),
    .A2(\mem[5][5] ),
    .A3(\mem[7][5] ),
    .S0(_055_),
    .S1(_072_),
    .X(_142_));
 sky130_fd_sc_hd__mux4_1 _339_ (.A0(\mem[0][5] ),
    .A1(\mem[2][5] ),
    .A2(\mem[4][5] ),
    .A3(\mem[6][5] ),
    .S0(_071_),
    .S1(_098_),
    .X(_143_));
 sky130_fd_sc_hd__a22oi_2 _340_ (.A1(_076_),
    .A2(_142_),
    .B1(_143_),
    .B2(_077_),
    .Y(_144_));
 sky130_fd_sc_hd__mux2i_2 _341_ (.A0(\mem[12][5] ),
    .A1(\mem[14][5] ),
    .S(_056_),
    .Y(_145_));
 sky130_fd_sc_hd__mux2i_1 _342_ (.A0(\mem[9][5] ),
    .A1(\mem[11][5] ),
    .S(_081_),
    .Y(_146_));
 sky130_fd_sc_hd__o22ai_2 _343_ (.A1(_088_),
    .A2(_145_),
    .B1(_146_),
    .B2(_091_),
    .Y(_147_));
 sky130_fd_sc_hd__mux2i_1 _344_ (.A0(\mem[8][5] ),
    .A1(\mem[10][5] ),
    .S(_089_),
    .Y(_148_));
 sky130_fd_sc_hd__mux2i_1 _345_ (.A0(\mem[13][5] ),
    .A1(\mem[15][5] ),
    .S(_057_),
    .Y(_149_));
 sky130_fd_sc_hd__o22ai_1 _346_ (.A1(_084_),
    .A2(_148_),
    .B1(_149_),
    .B2(_080_),
    .Y(_150_));
 sky130_fd_sc_hd__nor2_1 _347_ (.A(_147_),
    .B(_150_),
    .Y(_151_));
 sky130_fd_sc_hd__nor2_1 _348_ (.A(\rd_data_reg[5] ),
    .B(_095_),
    .Y(_152_));
 sky130_fd_sc_hd__a31oi_1 _349_ (.A1(_000_),
    .A2(_144_),
    .A3(_151_),
    .B1(_152_),
    .Y(_027_));
 sky130_fd_sc_hd__mux4_1 _350_ (.A0(\mem[1][6] ),
    .A1(\mem[3][6] ),
    .A2(\mem[5][6] ),
    .A3(\mem[7][6] ),
    .S0(_055_),
    .S1(_072_),
    .X(_153_));
 sky130_fd_sc_hd__mux4_2 _351_ (.A0(\mem[0][6] ),
    .A1(\mem[2][6] ),
    .A2(\mem[4][6] ),
    .A3(\mem[6][6] ),
    .S0(_071_),
    .S1(_098_),
    .X(_154_));
 sky130_fd_sc_hd__a22oi_2 _352_ (.A1(_076_),
    .A2(_153_),
    .B1(_154_),
    .B2(_077_),
    .Y(_155_));
 sky130_fd_sc_hd__mux2i_2 _353_ (.A0(\mem[12][6] ),
    .A1(\mem[14][6] ),
    .S(_056_),
    .Y(_156_));
 sky130_fd_sc_hd__mux2i_1 _354_ (.A0(\mem[9][6] ),
    .A1(\mem[11][6] ),
    .S(_081_),
    .Y(_157_));
 sky130_fd_sc_hd__o22ai_2 _355_ (.A1(_088_),
    .A2(_156_),
    .B1(_157_),
    .B2(_091_),
    .Y(_158_));
 sky130_fd_sc_hd__mux2i_2 _356_ (.A0(\mem[8][6] ),
    .A1(\mem[10][6] ),
    .S(_089_),
    .Y(_159_));
 sky130_fd_sc_hd__mux2i_1 _357_ (.A0(\mem[13][6] ),
    .A1(\mem[15][6] ),
    .S(_057_),
    .Y(_160_));
 sky130_fd_sc_hd__o22ai_1 _358_ (.A1(_084_),
    .A2(_159_),
    .B1(_160_),
    .B2(_080_),
    .Y(_161_));
 sky130_fd_sc_hd__nor2_1 _359_ (.A(_158_),
    .B(_161_),
    .Y(_162_));
 sky130_fd_sc_hd__nor2_1 _360_ (.A(\rd_data_reg[6] ),
    .B(_095_),
    .Y(_163_));
 sky130_fd_sc_hd__a31oi_1 _361_ (.A1(_000_),
    .A2(_155_),
    .A3(_162_),
    .B1(_163_),
    .Y(_028_));
 sky130_fd_sc_hd__mux4_1 _362_ (.A0(\mem[1][7] ),
    .A1(\mem[3][7] ),
    .A2(\mem[5][7] ),
    .A3(\mem[7][7] ),
    .S0(_055_),
    .S1(_072_),
    .X(_164_));
 sky130_fd_sc_hd__mux4_1 _363_ (.A0(\mem[0][7] ),
    .A1(\mem[2][7] ),
    .A2(\mem[4][7] ),
    .A3(\mem[6][7] ),
    .S0(_071_),
    .S1(_098_),
    .X(_165_));
 sky130_fd_sc_hd__a22oi_2 _364_ (.A1(_076_),
    .A2(_164_),
    .B1(_165_),
    .B2(_077_),
    .Y(_166_));
 sky130_fd_sc_hd__mux2i_1 _365_ (.A0(\mem[12][7] ),
    .A1(\mem[14][7] ),
    .S(_056_),
    .Y(_167_));
 sky130_fd_sc_hd__mux2i_1 _366_ (.A0(\mem[9][7] ),
    .A1(\mem[11][7] ),
    .S(_081_),
    .Y(_168_));
 sky130_fd_sc_hd__o22ai_2 _367_ (.A1(_088_),
    .A2(_167_),
    .B1(_168_),
    .B2(_091_),
    .Y(_169_));
 sky130_fd_sc_hd__mux2i_1 _368_ (.A0(\mem[8][7] ),
    .A1(\mem[10][7] ),
    .S(_089_),
    .Y(_170_));
 sky130_fd_sc_hd__mux2i_1 _369_ (.A0(\mem[13][7] ),
    .A1(\mem[15][7] ),
    .S(_089_),
    .Y(_171_));
 sky130_fd_sc_hd__o22ai_1 _370_ (.A1(_084_),
    .A2(_170_),
    .B1(_171_),
    .B2(_080_),
    .Y(_172_));
 sky130_fd_sc_hd__nor2_1 _371_ (.A(_169_),
    .B(_172_),
    .Y(_173_));
 sky130_fd_sc_hd__nor2_1 _372_ (.A(\rd_data_reg[7] ),
    .B(_095_),
    .Y(_174_));
 sky130_fd_sc_hd__a31oi_1 _373_ (.A1(_000_),
    .A2(_166_),
    .A3(_173_),
    .B1(_174_),
    .Y(_029_));
 sky130_fd_sc_hd__xor2_1 _374_ (.A(_074_),
    .B(_095_),
    .X(_030_));
 sky130_fd_sc_hd__nand2_1 _375_ (.A(_017_),
    .B(_095_),
    .Y(_175_));
 sky130_fd_sc_hd__o21ai_0 _376_ (.A1(_181_),
    .A2(_000_),
    .B1(_175_),
    .Y(_031_));
 sky130_fd_sc_hd__nand2_1 _377_ (.A(_195_),
    .B(_042_),
    .Y(_176_));
 sky130_fd_sc_hd__xnor2_1 _378_ (.A(_098_),
    .B(_176_),
    .Y(_032_));
 sky130_fd_sc_hd__nand4_1 _379_ (.A(_074_),
    .B(_057_),
    .C(_098_),
    .D(_042_),
    .Y(_177_));
 sky130_fd_sc_hd__xnor2_1 _380_ (.A(_058_),
    .B(_177_),
    .Y(_033_));
 sky130_fd_sc_hd__nand4_1 _381_ (.A(_098_),
    .B(_058_),
    .C(_195_),
    .D(_042_),
    .Y(_178_));
 sky130_fd_sc_hd__xnor2_1 _382_ (.A(\rd_ptr[4] ),
    .B(_178_),
    .Y(_034_));
 sky130_fd_sc_hd__xnor2_1 _383_ (.A(_018_),
    .B(_046_),
    .Y(_035_));
 sky130_fd_sc_hd__nand2_1 _384_ (.A(_019_),
    .B(_046_),
    .Y(_179_));
 sky130_fd_sc_hd__o21ai_0 _385_ (.A1(_196_),
    .A2(_046_),
    .B1(_179_),
    .Y(_036_));
 sky130_fd_sc_hd__xnor2_1 _386_ (.A(_044_),
    .B(_050_),
    .Y(_037_));
 sky130_fd_sc_hd__nand4_1 _387_ (.A(_044_),
    .B(\wr_addr[1] ),
    .C(\wr_addr[0] ),
    .D(_046_),
    .Y(_180_));
 sky130_fd_sc_hd__xnor2_1 _388_ (.A(_043_),
    .B(_180_),
    .Y(_038_));
 sky130_fd_sc_hd__xnor2_1 _389_ (.A(\wr_ptr[4] ),
    .B(_054_),
    .Y(_039_));
 sky130_fd_sc_hd__and2_0 _390_ (.A(\rd_data_reg[0] ),
    .B(rd_valid),
    .X(net17));
 sky130_fd_sc_hd__and2_0 _391_ (.A(\rd_data_reg[1] ),
    .B(rd_valid),
    .X(net18));
 sky130_fd_sc_hd__and2_0 _392_ (.A(\rd_data_reg[2] ),
    .B(rd_valid),
    .X(net19));
 sky130_fd_sc_hd__and2_0 _393_ (.A(\rd_data_reg[3] ),
    .B(rd_valid),
    .X(net20));
 sky130_fd_sc_hd__and2_0 _394_ (.A(\rd_data_reg[4] ),
    .B(rd_valid),
    .X(net21));
 sky130_fd_sc_hd__and2_0 _395_ (.A(\rd_data_reg[5] ),
    .B(rd_valid),
    .X(net22));
 sky130_fd_sc_hd__and2_0 _396_ (.A(\rd_data_reg[6] ),
    .B(rd_valid),
    .X(net23));
 sky130_fd_sc_hd__and2_0 _397_ (.A(\rd_data_reg[7] ),
    .B(rd_valid),
    .X(net24));
 sky130_fd_sc_hd__fa_1 _398_ (.A(_181_),
    .B(\wr_addr[1] ),
    .CIN(_182_),
    .COUT(_183_),
    .SUM(_184_));
 sky130_fd_sc_hd__ha_1 _399_ (.A(_181_),
    .B(\wr_addr[1] ),
    .COUT(_185_),
    .SUM(_186_));
 sky130_fd_sc_hd__ha_1 _400_ (.A(_187_),
    .B(\wr_addr[3] ),
    .COUT(_188_),
    .SUM(_189_));
 sky130_fd_sc_hd__ha_1 _401_ (.A(_190_),
    .B(\wr_addr[2] ),
    .COUT(_191_),
    .SUM(_192_));
 sky130_fd_sc_hd__ha_1 _402_ (.A(\rd_addr[0] ),
    .B(_018_),
    .COUT(_193_),
    .SUM(_194_));
 sky130_fd_sc_hd__ha_1 _403_ (.A(\rd_addr[0] ),
    .B(\rd_addr[1] ),
    .COUT(_195_),
    .SUM(_017_));
 sky130_fd_sc_hd__ha_1 _404_ (.A(_018_),
    .B(_196_),
    .COUT(_197_),
    .SUM(_019_));
 sky130_fd_sc_hd__ha_1 _405_ (.A(_018_),
    .B(\wr_addr[1] ),
    .COUT(_198_),
    .SUM(_199_));
 sky130_fd_sc_hd__ha_1 _406_ (.A(\wr_addr[0] ),
    .B(_196_),
    .COUT(_200_),
    .SUM(_201_));
 sky130_fd_sc_hd__ha_1 _407_ (.A(\wr_addr[0] ),
    .B(\wr_addr[1] ),
    .COUT(_202_),
    .SUM(_203_));
 sky130_fd_sc_hd__dfstp_1 \almost_empty_reg$_DFFE_PN1P_  (.D(_020_),
    .Q(net13),
    .SET_B(net3),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \almost_full_reg$_DFFE_PN0P_  (.D(_021_),
    .Q(net14),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][0]$_DFFE_PP_  (.D(net4),
    .DE(_001_),
    .Q(\mem[0][0] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][1]$_DFFE_PP_  (.D(net5),
    .DE(_001_),
    .Q(\mem[0][1] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][2]$_DFFE_PP_  (.D(net6),
    .DE(_001_),
    .Q(\mem[0][2] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][3]$_DFFE_PP_  (.D(net7),
    .DE(_001_),
    .Q(\mem[0][3] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][4]$_DFFE_PP_  (.D(net8),
    .DE(_001_),
    .Q(\mem[0][4] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][5]$_DFFE_PP_  (.D(net9),
    .DE(_001_),
    .Q(\mem[0][5] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][6]$_DFFE_PP_  (.D(net10),
    .DE(_001_),
    .Q(\mem[0][6] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][7]$_DFFE_PP_  (.D(net11),
    .DE(_001_),
    .Q(\mem[0][7] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][0]$_DFFE_PP_  (.D(net4),
    .DE(_002_),
    .Q(\mem[10][0] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][1]$_DFFE_PP_  (.D(net5),
    .DE(_002_),
    .Q(\mem[10][1] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][2]$_DFFE_PP_  (.D(net6),
    .DE(_002_),
    .Q(\mem[10][2] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][3]$_DFFE_PP_  (.D(net7),
    .DE(_002_),
    .Q(\mem[10][3] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][4]$_DFFE_PP_  (.D(net8),
    .DE(_002_),
    .Q(\mem[10][4] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][5]$_DFFE_PP_  (.D(net9),
    .DE(_002_),
    .Q(\mem[10][5] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][6]$_DFFE_PP_  (.D(net10),
    .DE(_002_),
    .Q(\mem[10][6] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][7]$_DFFE_PP_  (.D(net11),
    .DE(_002_),
    .Q(\mem[10][7] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][0]$_DFFE_PP_  (.D(net4),
    .DE(_003_),
    .Q(\mem[11][0] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][1]$_DFFE_PP_  (.D(net5),
    .DE(_003_),
    .Q(\mem[11][1] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][2]$_DFFE_PP_  (.D(net6),
    .DE(_003_),
    .Q(\mem[11][2] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][3]$_DFFE_PP_  (.D(net7),
    .DE(_003_),
    .Q(\mem[11][3] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][4]$_DFFE_PP_  (.D(net8),
    .DE(_003_),
    .Q(\mem[11][4] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][5]$_DFFE_PP_  (.D(net9),
    .DE(_003_),
    .Q(\mem[11][5] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][6]$_DFFE_PP_  (.D(net10),
    .DE(_003_),
    .Q(\mem[11][6] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][7]$_DFFE_PP_  (.D(net11),
    .DE(_003_),
    .Q(\mem[11][7] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][0]$_DFFE_PP_  (.D(net4),
    .DE(_004_),
    .Q(\mem[12][0] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][1]$_DFFE_PP_  (.D(net5),
    .DE(_004_),
    .Q(\mem[12][1] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][2]$_DFFE_PP_  (.D(net6),
    .DE(_004_),
    .Q(\mem[12][2] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][3]$_DFFE_PP_  (.D(net7),
    .DE(_004_),
    .Q(\mem[12][3] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][4]$_DFFE_PP_  (.D(net8),
    .DE(_004_),
    .Q(\mem[12][4] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][5]$_DFFE_PP_  (.D(net9),
    .DE(_004_),
    .Q(\mem[12][5] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][6]$_DFFE_PP_  (.D(net10),
    .DE(_004_),
    .Q(\mem[12][6] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][7]$_DFFE_PP_  (.D(net11),
    .DE(_004_),
    .Q(\mem[12][7] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][0]$_DFFE_PP_  (.D(net4),
    .DE(_005_),
    .Q(\mem[13][0] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][1]$_DFFE_PP_  (.D(net5),
    .DE(_005_),
    .Q(\mem[13][1] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][2]$_DFFE_PP_  (.D(net6),
    .DE(_005_),
    .Q(\mem[13][2] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][3]$_DFFE_PP_  (.D(net7),
    .DE(_005_),
    .Q(\mem[13][3] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][4]$_DFFE_PP_  (.D(net8),
    .DE(_005_),
    .Q(\mem[13][4] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][5]$_DFFE_PP_  (.D(net9),
    .DE(_005_),
    .Q(\mem[13][5] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][6]$_DFFE_PP_  (.D(net10),
    .DE(_005_),
    .Q(\mem[13][6] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][7]$_DFFE_PP_  (.D(net11),
    .DE(_005_),
    .Q(\mem[13][7] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][0]$_DFFE_PP_  (.D(net4),
    .DE(_006_),
    .Q(\mem[14][0] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][1]$_DFFE_PP_  (.D(net5),
    .DE(_006_),
    .Q(\mem[14][1] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][2]$_DFFE_PP_  (.D(net6),
    .DE(_006_),
    .Q(\mem[14][2] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][3]$_DFFE_PP_  (.D(net7),
    .DE(_006_),
    .Q(\mem[14][3] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][4]$_DFFE_PP_  (.D(net8),
    .DE(_006_),
    .Q(\mem[14][4] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][5]$_DFFE_PP_  (.D(net9),
    .DE(_006_),
    .Q(\mem[14][5] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][6]$_DFFE_PP_  (.D(net10),
    .DE(_006_),
    .Q(\mem[14][6] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][7]$_DFFE_PP_  (.D(net11),
    .DE(_006_),
    .Q(\mem[14][7] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][0]$_DFFE_PP_  (.D(net4),
    .DE(_007_),
    .Q(\mem[15][0] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][1]$_DFFE_PP_  (.D(net5),
    .DE(_007_),
    .Q(\mem[15][1] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][2]$_DFFE_PP_  (.D(net6),
    .DE(_007_),
    .Q(\mem[15][2] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][3]$_DFFE_PP_  (.D(net7),
    .DE(_007_),
    .Q(\mem[15][3] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][4]$_DFFE_PP_  (.D(net8),
    .DE(_007_),
    .Q(\mem[15][4] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][5]$_DFFE_PP_  (.D(net9),
    .DE(_007_),
    .Q(\mem[15][5] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][6]$_DFFE_PP_  (.D(net10),
    .DE(_007_),
    .Q(\mem[15][6] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][7]$_DFFE_PP_  (.D(net11),
    .DE(_007_),
    .Q(\mem[15][7] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][0]$_DFFE_PP_  (.D(net4),
    .DE(_008_),
    .Q(\mem[1][0] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][1]$_DFFE_PP_  (.D(net5),
    .DE(_008_),
    .Q(\mem[1][1] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][2]$_DFFE_PP_  (.D(net6),
    .DE(_008_),
    .Q(\mem[1][2] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][3]$_DFFE_PP_  (.D(net7),
    .DE(_008_),
    .Q(\mem[1][3] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][4]$_DFFE_PP_  (.D(net8),
    .DE(_008_),
    .Q(\mem[1][4] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][5]$_DFFE_PP_  (.D(net9),
    .DE(_008_),
    .Q(\mem[1][5] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][6]$_DFFE_PP_  (.D(net10),
    .DE(_008_),
    .Q(\mem[1][6] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][7]$_DFFE_PP_  (.D(net11),
    .DE(_008_),
    .Q(\mem[1][7] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][0]$_DFFE_PP_  (.D(net4),
    .DE(_009_),
    .Q(\mem[2][0] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][1]$_DFFE_PP_  (.D(net5),
    .DE(_009_),
    .Q(\mem[2][1] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][2]$_DFFE_PP_  (.D(net6),
    .DE(_009_),
    .Q(\mem[2][2] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][3]$_DFFE_PP_  (.D(net7),
    .DE(_009_),
    .Q(\mem[2][3] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][4]$_DFFE_PP_  (.D(net8),
    .DE(_009_),
    .Q(\mem[2][4] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][5]$_DFFE_PP_  (.D(net9),
    .DE(_009_),
    .Q(\mem[2][5] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][6]$_DFFE_PP_  (.D(net10),
    .DE(_009_),
    .Q(\mem[2][6] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][7]$_DFFE_PP_  (.D(net11),
    .DE(_009_),
    .Q(\mem[2][7] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][0]$_DFFE_PP_  (.D(net4),
    .DE(_010_),
    .Q(\mem[3][0] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][1]$_DFFE_PP_  (.D(net5),
    .DE(_010_),
    .Q(\mem[3][1] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][2]$_DFFE_PP_  (.D(net6),
    .DE(_010_),
    .Q(\mem[3][2] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][3]$_DFFE_PP_  (.D(net7),
    .DE(_010_),
    .Q(\mem[3][3] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][4]$_DFFE_PP_  (.D(net8),
    .DE(_010_),
    .Q(\mem[3][4] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][5]$_DFFE_PP_  (.D(net9),
    .DE(_010_),
    .Q(\mem[3][5] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][6]$_DFFE_PP_  (.D(net10),
    .DE(_010_),
    .Q(\mem[3][6] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][7]$_DFFE_PP_  (.D(net11),
    .DE(_010_),
    .Q(\mem[3][7] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][0]$_DFFE_PP_  (.D(net4),
    .DE(_011_),
    .Q(\mem[4][0] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][1]$_DFFE_PP_  (.D(net5),
    .DE(_011_),
    .Q(\mem[4][1] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][2]$_DFFE_PP_  (.D(net6),
    .DE(_011_),
    .Q(\mem[4][2] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][3]$_DFFE_PP_  (.D(net7),
    .DE(_011_),
    .Q(\mem[4][3] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][4]$_DFFE_PP_  (.D(net8),
    .DE(_011_),
    .Q(\mem[4][4] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][5]$_DFFE_PP_  (.D(net9),
    .DE(_011_),
    .Q(\mem[4][5] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][6]$_DFFE_PP_  (.D(net10),
    .DE(_011_),
    .Q(\mem[4][6] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][7]$_DFFE_PP_  (.D(net11),
    .DE(_011_),
    .Q(\mem[4][7] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][0]$_DFFE_PP_  (.D(net4),
    .DE(_012_),
    .Q(\mem[5][0] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][1]$_DFFE_PP_  (.D(net5),
    .DE(_012_),
    .Q(\mem[5][1] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][2]$_DFFE_PP_  (.D(net6),
    .DE(_012_),
    .Q(\mem[5][2] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][3]$_DFFE_PP_  (.D(net7),
    .DE(_012_),
    .Q(\mem[5][3] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][4]$_DFFE_PP_  (.D(net8),
    .DE(_012_),
    .Q(\mem[5][4] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][5]$_DFFE_PP_  (.D(net9),
    .DE(_012_),
    .Q(\mem[5][5] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][6]$_DFFE_PP_  (.D(net10),
    .DE(_012_),
    .Q(\mem[5][6] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][7]$_DFFE_PP_  (.D(net11),
    .DE(_012_),
    .Q(\mem[5][7] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][0]$_DFFE_PP_  (.D(net4),
    .DE(_013_),
    .Q(\mem[6][0] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][1]$_DFFE_PP_  (.D(net5),
    .DE(_013_),
    .Q(\mem[6][1] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][2]$_DFFE_PP_  (.D(net6),
    .DE(_013_),
    .Q(\mem[6][2] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][3]$_DFFE_PP_  (.D(net7),
    .DE(_013_),
    .Q(\mem[6][3] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][4]$_DFFE_PP_  (.D(net8),
    .DE(_013_),
    .Q(\mem[6][4] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][5]$_DFFE_PP_  (.D(net9),
    .DE(_013_),
    .Q(\mem[6][5] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][6]$_DFFE_PP_  (.D(net10),
    .DE(_013_),
    .Q(\mem[6][6] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][7]$_DFFE_PP_  (.D(net11),
    .DE(_013_),
    .Q(\mem[6][7] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][0]$_DFFE_PP_  (.D(net4),
    .DE(_014_),
    .Q(\mem[7][0] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][1]$_DFFE_PP_  (.D(net5),
    .DE(_014_),
    .Q(\mem[7][1] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][2]$_DFFE_PP_  (.D(net6),
    .DE(_014_),
    .Q(\mem[7][2] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][3]$_DFFE_PP_  (.D(net7),
    .DE(_014_),
    .Q(\mem[7][3] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][4]$_DFFE_PP_  (.D(net8),
    .DE(_014_),
    .Q(\mem[7][4] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][5]$_DFFE_PP_  (.D(net9),
    .DE(_014_),
    .Q(\mem[7][5] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][6]$_DFFE_PP_  (.D(net10),
    .DE(_014_),
    .Q(\mem[7][6] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][7]$_DFFE_PP_  (.D(net11),
    .DE(_014_),
    .Q(\mem[7][7] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][0]$_DFFE_PP_  (.D(net4),
    .DE(_015_),
    .Q(\mem[8][0] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][1]$_DFFE_PP_  (.D(net5),
    .DE(_015_),
    .Q(\mem[8][1] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][2]$_DFFE_PP_  (.D(net6),
    .DE(_015_),
    .Q(\mem[8][2] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][3]$_DFFE_PP_  (.D(net7),
    .DE(_015_),
    .Q(\mem[8][3] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][4]$_DFFE_PP_  (.D(net8),
    .DE(_015_),
    .Q(\mem[8][4] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][5]$_DFFE_PP_  (.D(net9),
    .DE(_015_),
    .Q(\mem[8][5] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][6]$_DFFE_PP_  (.D(net10),
    .DE(_015_),
    .Q(\mem[8][6] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][7]$_DFFE_PP_  (.D(net11),
    .DE(_015_),
    .Q(\mem[8][7] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][0]$_DFFE_PP_  (.D(net4),
    .DE(_016_),
    .Q(\mem[9][0] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][1]$_DFFE_PP_  (.D(net5),
    .DE(_016_),
    .Q(\mem[9][1] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][2]$_DFFE_PP_  (.D(net6),
    .DE(_016_),
    .Q(\mem[9][2] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][3]$_DFFE_PP_  (.D(net7),
    .DE(_016_),
    .Q(\mem[9][3] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][4]$_DFFE_PP_  (.D(net8),
    .DE(_016_),
    .Q(\mem[9][4] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][5]$_DFFE_PP_  (.D(net9),
    .DE(_016_),
    .Q(\mem[9][5] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][6]$_DFFE_PP_  (.D(net10),
    .DE(_016_),
    .Q(\mem[9][6] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][7]$_DFFE_PP_  (.D(net11),
    .DE(_016_),
    .Q(\mem[9][7] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_reg[0]$_DFFE_PN0P_  (.D(_022_),
    .Q(\rd_data_reg[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_reg[1]$_DFFE_PN0P_  (.D(_023_),
    .Q(\rd_data_reg[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_reg[2]$_DFFE_PN0P_  (.D(_024_),
    .Q(\rd_data_reg[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_reg[3]$_DFFE_PN0P_  (.D(_025_),
    .Q(\rd_data_reg[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_reg[4]$_DFFE_PN0P_  (.D(_026_),
    .Q(\rd_data_reg[4] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_reg[5]$_DFFE_PN0P_  (.D(_027_),
    .Q(\rd_data_reg[5] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_reg[6]$_DFFE_PN0P_  (.D(_028_),
    .Q(\rd_data_reg[6] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_reg[7]$_DFFE_PN0P_  (.D(_029_),
    .Q(\rd_data_reg[7] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[0]$_DFFE_PN0P_  (.D(_030_),
    .Q(\rd_addr[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[1]$_DFFE_PN0P_  (.D(_031_),
    .Q(\rd_addr[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[2]$_DFFE_PN0P_  (.D(_032_),
    .Q(\rd_addr[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[3]$_DFFE_PN0P_  (.D(_033_),
    .Q(\rd_addr[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[4]$_DFFE_PN0P_  (.D(_034_),
    .Q(\rd_ptr[4] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \rd_valid$_DFF_PN0_  (.D(_000_),
    .Q(rd_valid),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[0]$_DFFE_PN0P_  (.D(_035_),
    .Q(\wr_addr[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \wr_ptr[1]$_DFFE_PN0P_  (.D(_036_),
    .Q(\wr_addr[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[2]$_DFFE_PN0P_  (.D(_037_),
    .Q(\wr_addr[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[3]$_DFFE_PN0P_  (.D(_038_),
    .Q(\wr_addr[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[4]$_DFFE_PN0P_  (.D(_039_),
    .Q(\wr_ptr[4] ),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__buf_8 hold1 (.A(net3),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_135 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(rd_en),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(net25),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(wr_data[0]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_8 input4 (.A(net27),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input5 (.A(net30),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input6 (.A(wr_data[3]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input7 (.A(net29),
    .X(net8));
 sky130_fd_sc_hd__buf_6 input8 (.A(net26),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_8 input9 (.A(net28),
    .X(net10));
 sky130_fd_sc_hd__buf_4 input10 (.A(wr_data[7]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(wr_en),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 output12 (.A(net13),
    .X(almost_empty));
 sky130_fd_sc_hd__clkbuf_1 output13 (.A(net14),
    .X(almost_full));
 sky130_fd_sc_hd__clkbuf_1 output14 (.A(net15),
    .X(empty));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net16),
    .X(full));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net17),
    .X(rd_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net18),
    .X(rd_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net19),
    .X(rd_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net20),
    .X(rd_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net21),
    .X(rd_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net22),
    .X(rd_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net23),
    .X(rd_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net24),
    .X(rd_data[7]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload0 (.A(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload1 (.A(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload2 (.A(clknet_4_2_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload3 (.A(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload4 (.A(clknet_4_4_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload5 (.A(clknet_4_5_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload6 (.A(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload7 (.A(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkinv_1 clkload8 (.A(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkinv_1 clkload9 (.A(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload10 (.A(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload11 (.A(clknet_4_12_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload12 (.A(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload13 (.A(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload14 (.A(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net25));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(wr_data[5]),
    .X(net26));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(wr_data[1]),
    .X(net27));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(wr_data[6]),
    .X(net28));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(wr_data[4]),
    .X(net29));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(wr_data[2]),
    .X(net30));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_214 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_210 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_83 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_220 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_90 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_87 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_162 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_220 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_184 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_214 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_219 ();
endmodule
