module parameterized_i2c_master (ack_error,
    busy,
    clk,
    done,
    read,
    rst_n,
    scl,
    scl_internal_debug,
    sda,
    sda_internal_debug,
    start,
    stop,
    write,
    addr,
    bit_counter_debug,
    data_in,
    data_out,
    phase,
    shift_reg_debug,
    state);
 output ack_error;
 output busy;
 input clk;
 output done;
 input read;
 input rst_n;
 output scl;
 output scl_internal_debug;
 inout sda;
 output sda_internal_debug;
 input start;
 input stop;
 input write;
 input [6:0] addr;
 output [2:0] bit_counter_debug;
 input [7:0] data_in;
 output [7:0] data_out;
 output [1:0] phase;
 output [7:0] shift_reg_debug;
 output [3:0] state;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire clknet_0_clk;
 wire cmd_read;
 wire cmd_write;
 wire \divider_counter[0] ;
 wire \divider_counter[1] ;
 wire \divider_counter[2] ;
 wire \divider_counter[3] ;
 wire \divider_counter[4] ;
 wire \divider_counter[5] ;
 wire \divider_counter[6] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net54;

 sky130_fd_sc_hd__buf_2 _278_ (.A(net23),
    .X(_039_));
 sky130_fd_sc_hd__inv_1 _279_ (.A(_039_),
    .Y(_259_));
 sky130_fd_sc_hd__or4_2 _280_ (.A(\divider_counter[5] ),
    .B(\divider_counter[4] ),
    .C(\divider_counter[3] ),
    .D(\divider_counter[2] ),
    .X(_040_));
 sky130_fd_sc_hd__nor4_4 _281_ (.A(\divider_counter[6] ),
    .B(\divider_counter[1] ),
    .C(\divider_counter[0] ),
    .D(_040_),
    .Y(_041_));
 sky130_fd_sc_hd__buf_2 _282_ (.A(_041_),
    .X(_042_));
 sky130_fd_sc_hd__nor2_1 _283_ (.A(\divider_counter[0] ),
    .B(_042_),
    .Y(_000_));
 sky130_fd_sc_hd__nor2_1 _284_ (.A(_258_),
    .B(_042_),
    .Y(_001_));
 sky130_fd_sc_hd__or4_2 _285_ (.A(\divider_counter[6] ),
    .B(\divider_counter[1] ),
    .C(\divider_counter[0] ),
    .D(_040_),
    .X(_043_));
 sky130_fd_sc_hd__xnor2_1 _286_ (.A(\divider_counter[2] ),
    .B(_257_),
    .Y(_044_));
 sky130_fd_sc_hd__nand2_1 _287_ (.A(_043_),
    .B(_044_),
    .Y(_002_));
 sky130_fd_sc_hd__nor3_1 _288_ (.A(\divider_counter[1] ),
    .B(\divider_counter[2] ),
    .C(\divider_counter[0] ),
    .Y(_045_));
 sky130_fd_sc_hd__xor2_1 _289_ (.A(\divider_counter[3] ),
    .B(_045_),
    .X(_003_));
 sky130_fd_sc_hd__nor2_1 _290_ (.A(\divider_counter[3] ),
    .B(\divider_counter[2] ),
    .Y(_046_));
 sky130_fd_sc_hd__a21oi_1 _291_ (.A1(_257_),
    .A2(_046_),
    .B1(\divider_counter[4] ),
    .Y(_047_));
 sky130_fd_sc_hd__and3_1 _292_ (.A(\divider_counter[4] ),
    .B(_257_),
    .C(_046_),
    .X(_048_));
 sky130_fd_sc_hd__o21ai_0 _293_ (.A1(_047_),
    .A2(_048_),
    .B1(_043_),
    .Y(_004_));
 sky130_fd_sc_hd__nor2_1 _294_ (.A(\divider_counter[1] ),
    .B(\divider_counter[0] ),
    .Y(_049_));
 sky130_fd_sc_hd__nand3b_1 _295_ (.A_N(\divider_counter[4] ),
    .B(_046_),
    .C(_049_),
    .Y(_050_));
 sky130_fd_sc_hd__xnor2_1 _296_ (.A(\divider_counter[5] ),
    .B(_050_),
    .Y(_005_));
 sky130_fd_sc_hd__nor2_1 _297_ (.A(_257_),
    .B(_049_),
    .Y(_051_));
 sky130_fd_sc_hd__inv_1 _298_ (.A(_257_),
    .Y(_052_));
 sky130_fd_sc_hd__o21ai_0 _299_ (.A1(_052_),
    .A2(_040_),
    .B1(\divider_counter[6] ),
    .Y(_053_));
 sky130_fd_sc_hd__o31ai_1 _300_ (.A1(\divider_counter[6] ),
    .A2(_040_),
    .A3(_051_),
    .B1(_053_),
    .Y(_006_));
 sky130_fd_sc_hd__clkbuf_4 _301_ (.A(net51),
    .X(_054_));
 sky130_fd_sc_hd__buf_2 _302_ (.A(_054_),
    .X(_055_));
 sky130_fd_sc_hd__buf_2 _303_ (.A(net50),
    .X(_056_));
 sky130_fd_sc_hd__nor3_2 _304_ (.A(net49),
    .B(net48),
    .C(_056_),
    .Y(_057_));
 sky130_fd_sc_hd__nand2_1 _305_ (.A(_055_),
    .B(_057_),
    .Y(_058_));
 sky130_fd_sc_hd__buf_2 _306_ (.A(_275_),
    .X(_059_));
 sky130_fd_sc_hd__buf_2 _307_ (.A(_059_),
    .X(_060_));
 sky130_fd_sc_hd__nand2_1 _308_ (.A(_060_),
    .B(_041_),
    .Y(_061_));
 sky130_fd_sc_hd__nor2_1 _309_ (.A(_058_),
    .B(_061_),
    .Y(_007_));
 sky130_fd_sc_hd__inv_1 _310_ (.A(\divider_counter[0] ),
    .Y(_255_));
 sky130_fd_sc_hd__inv_1 _311_ (.A(net36),
    .Y(_267_));
 sky130_fd_sc_hd__inv_1 _312_ (.A(\divider_counter[1] ),
    .Y(_256_));
 sky130_fd_sc_hd__inv_1 _313_ (.A(net24),
    .Y(_260_));
 sky130_fd_sc_hd__inv_1 _314_ (.A(net37),
    .Y(_268_));
 sky130_fd_sc_hd__clkbuf_4 _315_ (.A(_054_),
    .X(_062_));
 sky130_fd_sc_hd__buf_2 _316_ (.A(net49),
    .X(_063_));
 sky130_fd_sc_hd__buf_2 _317_ (.A(_063_),
    .X(_064_));
 sky130_fd_sc_hd__buf_4 _318_ (.A(net48),
    .X(_065_));
 sky130_fd_sc_hd__clkbuf_4 _319_ (.A(_065_),
    .X(_066_));
 sky130_fd_sc_hd__buf_2 _320_ (.A(_271_),
    .X(_067_));
 sky130_fd_sc_hd__nor2b_1 _321_ (.A(_056_),
    .B_N(_067_),
    .Y(_068_));
 sky130_fd_sc_hd__clkbuf_4 _322_ (.A(net48),
    .X(_069_));
 sky130_fd_sc_hd__clkinvlp_4 _323_ (.A(_069_),
    .Y(_070_));
 sky130_fd_sc_hd__buf_2 _324_ (.A(_056_),
    .X(_071_));
 sky130_fd_sc_hd__inv_1 _325_ (.A(_071_),
    .Y(_072_));
 sky130_fd_sc_hd__nand2_1 _326_ (.A(_070_),
    .B(_072_),
    .Y(_073_));
 sky130_fd_sc_hd__buf_2 _327_ (.A(_071_),
    .X(_074_));
 sky130_fd_sc_hd__nand3_1 _328_ (.A(_066_),
    .B(_074_),
    .C(_067_),
    .Y(_075_));
 sky130_fd_sc_hd__a21oi_1 _329_ (.A1(_073_),
    .A2(_075_),
    .B1(_064_),
    .Y(_076_));
 sky130_fd_sc_hd__a31oi_1 _330_ (.A1(_064_),
    .A2(_066_),
    .A3(_068_),
    .B1(_076_),
    .Y(_077_));
 sky130_fd_sc_hd__inv_1 _331_ (.A(net19),
    .Y(_078_));
 sky130_fd_sc_hd__nor2_2 _332_ (.A(_063_),
    .B(_069_),
    .Y(_079_));
 sky130_fd_sc_hd__and3_1 _333_ (.A(_063_),
    .B(_065_),
    .C(_067_),
    .X(_080_));
 sky130_fd_sc_hd__a21oi_1 _334_ (.A1(_078_),
    .A2(_079_),
    .B1(_080_),
    .Y(_081_));
 sky130_fd_sc_hd__nor3_1 _335_ (.A(_054_),
    .B(_071_),
    .C(_081_),
    .Y(_082_));
 sky130_fd_sc_hd__o41a_1 _336_ (.A1(_062_),
    .A2(_043_),
    .A3(_077_),
    .A4(_082_),
    .B1(net22),
    .X(_008_));
 sky130_fd_sc_hd__inv_1 _337_ (.A(_063_),
    .Y(_083_));
 sky130_fd_sc_hd__nor2_1 _338_ (.A(_069_),
    .B(_054_),
    .Y(_084_));
 sky130_fd_sc_hd__a21boi_2 _339_ (.A1(_083_),
    .A2(_072_),
    .B1_N(_084_),
    .Y(_085_));
 sky130_fd_sc_hd__nand2_1 _340_ (.A(_039_),
    .B(_085_),
    .Y(_086_));
 sky130_fd_sc_hd__o21ai_0 _341_ (.A1(_063_),
    .A2(_071_),
    .B1(_084_),
    .Y(_087_));
 sky130_fd_sc_hd__buf_2 _342_ (.A(net25),
    .X(_088_));
 sky130_fd_sc_hd__inv_1 _343_ (.A(_088_),
    .Y(_089_));
 sky130_fd_sc_hd__nand3_2 _344_ (.A(_260_),
    .B(_089_),
    .C(_259_),
    .Y(_090_));
 sky130_fd_sc_hd__nor2b_2 _345_ (.A(net51),
    .B_N(_056_),
    .Y(_091_));
 sky130_fd_sc_hd__nand2b_1 _346_ (.A_N(net20),
    .B(cmd_read),
    .Y(_092_));
 sky130_fd_sc_hd__nand4_1 _347_ (.A(_064_),
    .B(_065_),
    .C(_091_),
    .D(_092_),
    .Y(_093_));
 sky130_fd_sc_hd__o21ai_0 _348_ (.A1(_087_),
    .A2(_090_),
    .B1(_093_),
    .Y(_094_));
 sky130_fd_sc_hd__o21ai_0 _349_ (.A1(_070_),
    .A2(_071_),
    .B1(_063_),
    .Y(_095_));
 sky130_fd_sc_hd__nand2_1 _350_ (.A(_070_),
    .B(_071_),
    .Y(_096_));
 sky130_fd_sc_hd__a211oi_1 _351_ (.A1(_095_),
    .A2(_096_),
    .B1(_054_),
    .C1(_059_),
    .Y(_097_));
 sky130_fd_sc_hd__nand2b_2 _352_ (.A_N(net51),
    .B(_069_),
    .Y(_098_));
 sky130_fd_sc_hd__nor2b_1 _353_ (.A(net20),
    .B_N(cmd_write),
    .Y(_099_));
 sky130_fd_sc_hd__nand2b_1 _354_ (.A_N(net49),
    .B(_056_),
    .Y(_100_));
 sky130_fd_sc_hd__nand2b_1 _355_ (.A_N(_056_),
    .B(net49),
    .Y(_101_));
 sky130_fd_sc_hd__o22a_1 _356_ (.A1(_099_),
    .A2(_100_),
    .B1(_101_),
    .B2(_059_),
    .X(_102_));
 sky130_fd_sc_hd__nor2_1 _357_ (.A(_054_),
    .B(_071_),
    .Y(_103_));
 sky130_fd_sc_hd__and3_1 _358_ (.A(_063_),
    .B(_069_),
    .C(_059_),
    .X(_104_));
 sky130_fd_sc_hd__nand3_1 _359_ (.A(net22),
    .B(_103_),
    .C(_104_),
    .Y(_105_));
 sky130_fd_sc_hd__nor2b_1 _360_ (.A(net49),
    .B_N(_069_),
    .Y(_106_));
 sky130_fd_sc_hd__mux2i_1 _361_ (.A0(_067_),
    .A1(_059_),
    .S(_056_),
    .Y(_107_));
 sky130_fd_sc_hd__a221oi_2 _362_ (.A1(_078_),
    .A2(_057_),
    .B1(_106_),
    .B2(_107_),
    .C1(_054_),
    .Y(_108_));
 sky130_fd_sc_hd__o2111ai_4 _363_ (.A1(_098_),
    .A2(_102_),
    .B1(_105_),
    .C1(_108_),
    .D1(_041_),
    .Y(_109_));
 sky130_fd_sc_hd__a211oi_2 _364_ (.A1(_060_),
    .A2(_094_),
    .B1(_097_),
    .C1(_109_),
    .Y(_110_));
 sky130_fd_sc_hd__mux2_1 _365_ (.A0(_039_),
    .A1(_086_),
    .S(_110_),
    .X(_009_));
 sky130_fd_sc_hd__nand2_1 _366_ (.A(_262_),
    .B(_085_),
    .Y(_111_));
 sky130_fd_sc_hd__nand2_1 _367_ (.A(_110_),
    .B(_111_),
    .Y(_112_));
 sky130_fd_sc_hd__o21ai_0 _368_ (.A1(_260_),
    .A2(_110_),
    .B1(_112_),
    .Y(_010_));
 sky130_fd_sc_hd__clkbuf_2 _369_ (.A(_261_),
    .X(_113_));
 sky130_fd_sc_hd__o21ai_0 _370_ (.A1(_113_),
    .A2(_087_),
    .B1(_110_),
    .Y(_114_));
 sky130_fd_sc_hd__and4_1 _371_ (.A(_088_),
    .B(_113_),
    .C(_085_),
    .D(_110_),
    .X(_115_));
 sky130_fd_sc_hd__a21oi_1 _372_ (.A1(_089_),
    .A2(_114_),
    .B1(_115_),
    .Y(_011_));
 sky130_fd_sc_hd__nor4_2 _373_ (.A(_063_),
    .B(_069_),
    .C(net51),
    .D(_056_),
    .Y(_116_));
 sky130_fd_sc_hd__nand3_2 _374_ (.A(net19),
    .B(_042_),
    .C(_116_),
    .Y(_117_));
 sky130_fd_sc_hd__mux2_1 _375_ (.A0(net17),
    .A1(cmd_read),
    .S(_117_),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _376_ (.A0(net21),
    .A1(cmd_write),
    .S(_117_),
    .X(_014_));
 sky130_fd_sc_hd__nor2b_2 _377_ (.A(net48),
    .B_N(net49),
    .Y(_118_));
 sky130_fd_sc_hd__nand2_2 _378_ (.A(_091_),
    .B(_118_),
    .Y(_119_));
 sky130_fd_sc_hd__nor3_4 _379_ (.A(_061_),
    .B(_090_),
    .C(_119_),
    .Y(_120_));
 sky130_fd_sc_hd__mux2_1 _380_ (.A0(net27),
    .A1(net40),
    .S(_120_),
    .X(_015_));
 sky130_fd_sc_hd__mux2_1 _381_ (.A0(net28),
    .A1(net41),
    .S(_120_),
    .X(_016_));
 sky130_fd_sc_hd__mux2_1 _382_ (.A0(net29),
    .A1(net42),
    .S(_120_),
    .X(_017_));
 sky130_fd_sc_hd__mux2_1 _383_ (.A0(net30),
    .A1(net43),
    .S(_120_),
    .X(_018_));
 sky130_fd_sc_hd__mux2_1 _384_ (.A0(net31),
    .A1(net44),
    .S(_120_),
    .X(_019_));
 sky130_fd_sc_hd__mux2_1 _385_ (.A0(net32),
    .A1(net45),
    .S(_120_),
    .X(_020_));
 sky130_fd_sc_hd__mux2_1 _386_ (.A0(net33),
    .A1(net46),
    .S(_120_),
    .X(_021_));
 sky130_fd_sc_hd__mux2_1 _387_ (.A0(net34),
    .A1(net47),
    .S(_120_),
    .X(_022_));
 sky130_fd_sc_hd__a21oi_1 _388_ (.A1(_095_),
    .A2(_096_),
    .B1(_062_),
    .Y(_121_));
 sky130_fd_sc_hd__nand2_1 _389_ (.A(_041_),
    .B(_105_),
    .Y(_122_));
 sky130_fd_sc_hd__nor3_1 _390_ (.A(_060_),
    .B(_269_),
    .C(_098_),
    .Y(_123_));
 sky130_fd_sc_hd__clkbuf_4 _391_ (.A(_101_),
    .X(_124_));
 sky130_fd_sc_hd__o21ai_0 _392_ (.A1(_273_),
    .A2(_124_),
    .B1(_100_),
    .Y(_125_));
 sky130_fd_sc_hd__inv_1 _393_ (.A(_059_),
    .Y(_126_));
 sky130_fd_sc_hd__nor3_1 _394_ (.A(net24),
    .B(_088_),
    .C(_039_),
    .Y(_127_));
 sky130_fd_sc_hd__nor2_2 _395_ (.A(_126_),
    .B(_127_),
    .Y(_128_));
 sky130_fd_sc_hd__and2_0 _396_ (.A(_091_),
    .B(_118_),
    .X(_129_));
 sky130_fd_sc_hd__buf_2 _397_ (.A(_129_),
    .X(_130_));
 sky130_fd_sc_hd__a22o_1 _398_ (.A1(_123_),
    .A2(_125_),
    .B1(_128_),
    .B2(_130_),
    .X(_131_));
 sky130_fd_sc_hd__a211oi_1 _399_ (.A1(_270_),
    .A2(_121_),
    .B1(_122_),
    .C1(_131_),
    .Y(_132_));
 sky130_fd_sc_hd__nor2_1 _400_ (.A(_065_),
    .B(_060_),
    .Y(_133_));
 sky130_fd_sc_hd__nor3_1 _401_ (.A(_070_),
    .B(_126_),
    .C(_092_),
    .Y(_134_));
 sky130_fd_sc_hd__o21ai_0 _402_ (.A1(_070_),
    .A2(_060_),
    .B1(_083_),
    .Y(_135_));
 sky130_fd_sc_hd__o311a_1 _403_ (.A1(_083_),
    .A2(_133_),
    .A3(_134_),
    .B1(_091_),
    .C1(_135_),
    .X(_136_));
 sky130_fd_sc_hd__a31oi_1 _404_ (.A1(_074_),
    .A2(_126_),
    .A3(net20),
    .B1(_062_),
    .Y(_137_));
 sky130_fd_sc_hd__o2111ai_1 _405_ (.A1(net39),
    .A2(_127_),
    .B1(_079_),
    .C1(_060_),
    .D1(_091_),
    .Y(_138_));
 sky130_fd_sc_hd__and3b_1 _406_ (.A_N(_063_),
    .B(_069_),
    .C(_071_),
    .X(_139_));
 sky130_fd_sc_hd__clkbuf_4 _407_ (.A(_139_),
    .X(_140_));
 sky130_fd_sc_hd__nand3_1 _408_ (.A(net16),
    .B(_099_),
    .C(_140_),
    .Y(_141_));
 sky130_fd_sc_hd__o21a_1 _409_ (.A1(_069_),
    .A2(_071_),
    .B1(_054_),
    .X(_142_));
 sky130_fd_sc_hd__a311oi_1 _410_ (.A1(_074_),
    .A2(net20),
    .A3(_118_),
    .B1(_142_),
    .C1(_116_),
    .Y(_143_));
 sky130_fd_sc_hd__o2111ai_1 _411_ (.A1(_083_),
    .A2(_137_),
    .B1(_138_),
    .C1(_141_),
    .D1(_143_),
    .Y(_144_));
 sky130_fd_sc_hd__nor2_1 _412_ (.A(_136_),
    .B(_144_),
    .Y(_145_));
 sky130_fd_sc_hd__clkinvlp_4 _413_ (.A(_054_),
    .Y(_146_));
 sky130_fd_sc_hd__o2111ai_1 _414_ (.A1(cmd_read),
    .A2(net47),
    .B1(_064_),
    .C1(_065_),
    .D1(_146_),
    .Y(_147_));
 sky130_fd_sc_hd__nand2_1 _415_ (.A(_062_),
    .B(_079_),
    .Y(_148_));
 sky130_fd_sc_hd__a21o_1 _416_ (.A1(_083_),
    .A2(_067_),
    .B1(_098_),
    .X(_149_));
 sky130_fd_sc_hd__nor2b_1 _417_ (.A(_067_),
    .B_N(_059_),
    .Y(_150_));
 sky130_fd_sc_hd__a31oi_1 _418_ (.A1(_054_),
    .A2(_067_),
    .A3(_079_),
    .B1(_150_),
    .Y(_151_));
 sky130_fd_sc_hd__a32oi_1 _419_ (.A1(_060_),
    .A2(_147_),
    .A3(_148_),
    .B1(_149_),
    .B2(_151_),
    .Y(_152_));
 sky130_fd_sc_hd__nand2b_1 _420_ (.A_N(_088_),
    .B(net24),
    .Y(_153_));
 sky130_fd_sc_hd__mux2_1 _421_ (.A0(net42),
    .A1(net43),
    .S(_039_),
    .X(_154_));
 sky130_fd_sc_hd__o2111ai_1 _422_ (.A1(_153_),
    .A2(_154_),
    .B1(_126_),
    .C1(_079_),
    .D1(_091_),
    .Y(_155_));
 sky130_fd_sc_hd__mux4_1 _423_ (.A0(net40),
    .A1(net41),
    .A2(net44),
    .A3(net45),
    .S0(_039_),
    .S1(_088_),
    .X(_156_));
 sky130_fd_sc_hd__nand2_1 _424_ (.A(net24),
    .B(_088_),
    .Y(_157_));
 sky130_fd_sc_hd__mux2_1 _425_ (.A0(net46),
    .A1(net47),
    .S(_039_),
    .X(_158_));
 sky130_fd_sc_hd__o22ai_1 _426_ (.A1(net24),
    .A2(_156_),
    .B1(_157_),
    .B2(_158_),
    .Y(_159_));
 sky130_fd_sc_hd__nor2_1 _427_ (.A(_155_),
    .B(_159_),
    .Y(_160_));
 sky130_fd_sc_hd__a21oi_1 _428_ (.A1(_072_),
    .A2(_152_),
    .B1(_160_),
    .Y(_161_));
 sky130_fd_sc_hd__o211ai_1 _429_ (.A1(_060_),
    .A2(net47),
    .B1(_103_),
    .C1(_118_),
    .Y(_162_));
 sky130_fd_sc_hd__nand4_1 _430_ (.A(_132_),
    .B(_145_),
    .C(_161_),
    .D(_162_),
    .Y(_163_));
 sky130_fd_sc_hd__nand4b_1 _431_ (.A_N(net39),
    .B(_128_),
    .C(_145_),
    .D(_161_),
    .Y(_164_));
 sky130_fd_sc_hd__o211a_1 _432_ (.A1(net39),
    .A2(_132_),
    .B1(_163_),
    .C1(_164_),
    .X(_026_));
 sky130_fd_sc_hd__nand4b_1 _433_ (.A_N(net22),
    .B(cmd_read),
    .C(_103_),
    .D(_104_),
    .Y(_165_));
 sky130_fd_sc_hd__a211o_1 _434_ (.A1(_067_),
    .A2(_118_),
    .B1(_106_),
    .C1(_072_),
    .X(_166_));
 sky130_fd_sc_hd__o311ai_4 _435_ (.A1(_065_),
    .A2(_124_),
    .A3(_128_),
    .B1(_165_),
    .C1(_166_),
    .Y(_167_));
 sky130_fd_sc_hd__nor2_4 _436_ (.A(_109_),
    .B(_167_),
    .Y(_168_));
 sky130_fd_sc_hd__inv_1 _437_ (.A(net9),
    .Y(_169_));
 sky130_fd_sc_hd__mux2i_1 _438_ (.A0(cmd_read),
    .A1(net9),
    .S(_074_),
    .Y(_170_));
 sky130_fd_sc_hd__o22ai_1 _439_ (.A1(_169_),
    .A2(_124_),
    .B1(_170_),
    .B2(_064_),
    .Y(_171_));
 sky130_fd_sc_hd__a32oi_1 _440_ (.A1(_064_),
    .A2(_074_),
    .A3(net17),
    .B1(_171_),
    .B2(_146_),
    .Y(_172_));
 sky130_fd_sc_hd__o21ai_0 _441_ (.A1(_062_),
    .A2(_079_),
    .B1(net17),
    .Y(_173_));
 sky130_fd_sc_hd__o21ai_0 _442_ (.A1(_070_),
    .A2(_172_),
    .B1(_173_),
    .Y(_174_));
 sky130_fd_sc_hd__xnor2_1 _443_ (.A(_088_),
    .B(_113_),
    .Y(_175_));
 sky130_fd_sc_hd__o31ai_1 _444_ (.A1(_262_),
    .A2(_090_),
    .A3(_175_),
    .B1(_130_),
    .Y(_176_));
 sky130_fd_sc_hd__a21boi_0 _445_ (.A1(_176_),
    .A2(_168_),
    .B1_N(net40),
    .Y(_177_));
 sky130_fd_sc_hd__a21o_1 _446_ (.A1(_168_),
    .A2(_174_),
    .B1(_177_),
    .X(_027_));
 sky130_fd_sc_hd__mux2i_1 _447_ (.A0(net40),
    .A1(net10),
    .S(_066_),
    .Y(_178_));
 sky130_fd_sc_hd__nor2_1 _448_ (.A(_124_),
    .B(_178_),
    .Y(_179_));
 sky130_fd_sc_hd__a21oi_1 _449_ (.A1(net10),
    .A2(_140_),
    .B1(_179_),
    .Y(_180_));
 sky130_fd_sc_hd__nand2_1 _450_ (.A(_263_),
    .B(_175_),
    .Y(_181_));
 sky130_fd_sc_hd__a21boi_1 _451_ (.A1(_065_),
    .A2(_071_),
    .B1_N(_064_),
    .Y(_182_));
 sky130_fd_sc_hd__o21ai_4 _452_ (.A1(_140_),
    .A2(_182_),
    .B1(_146_),
    .Y(_183_));
 sky130_fd_sc_hd__a32oi_1 _453_ (.A1(net41),
    .A2(_130_),
    .A3(_181_),
    .B1(_183_),
    .B2(net2),
    .Y(_184_));
 sky130_fd_sc_hd__o21ai_0 _454_ (.A1(_055_),
    .A2(_180_),
    .B1(_184_),
    .Y(_185_));
 sky130_fd_sc_hd__mux2_1 _455_ (.A0(net41),
    .A1(_185_),
    .S(_168_),
    .X(_028_));
 sky130_fd_sc_hd__nand2_1 _456_ (.A(_088_),
    .B(_113_),
    .Y(_186_));
 sky130_fd_sc_hd__o21ai_0 _457_ (.A1(_113_),
    .A2(_153_),
    .B1(_186_),
    .Y(_187_));
 sky130_fd_sc_hd__nand3_1 _458_ (.A(_262_),
    .B(_259_),
    .C(_187_),
    .Y(_188_));
 sky130_fd_sc_hd__nand3_1 _459_ (.A(net42),
    .B(_130_),
    .C(_188_),
    .Y(_189_));
 sky130_fd_sc_hd__mux2i_1 _460_ (.A0(net41),
    .A1(net11),
    .S(_066_),
    .Y(_190_));
 sky130_fd_sc_hd__nor2_1 _461_ (.A(_124_),
    .B(_190_),
    .Y(_191_));
 sky130_fd_sc_hd__a21oi_1 _462_ (.A1(net11),
    .A2(_140_),
    .B1(_191_),
    .Y(_192_));
 sky130_fd_sc_hd__nand2_1 _463_ (.A(net3),
    .B(_183_),
    .Y(_193_));
 sky130_fd_sc_hd__o21ai_0 _464_ (.A1(_055_),
    .A2(_192_),
    .B1(_193_),
    .Y(_194_));
 sky130_fd_sc_hd__mux2i_1 _465_ (.A0(net42),
    .A1(_194_),
    .S(_168_),
    .Y(_195_));
 sky130_fd_sc_hd__nand2_1 _466_ (.A(_189_),
    .B(_195_),
    .Y(_029_));
 sky130_fd_sc_hd__mux2i_1 _467_ (.A0(net42),
    .A1(net12),
    .S(_065_),
    .Y(_196_));
 sky130_fd_sc_hd__nor2_1 _468_ (.A(_124_),
    .B(_196_),
    .Y(_197_));
 sky130_fd_sc_hd__a21oi_1 _469_ (.A1(net12),
    .A2(_140_),
    .B1(_197_),
    .Y(_198_));
 sky130_fd_sc_hd__nand2_1 _470_ (.A(_265_),
    .B(_175_),
    .Y(_199_));
 sky130_fd_sc_hd__a32oi_1 _471_ (.A1(net43),
    .A2(_130_),
    .A3(_199_),
    .B1(_183_),
    .B2(net4),
    .Y(_200_));
 sky130_fd_sc_hd__o21ai_0 _472_ (.A1(_055_),
    .A2(_198_),
    .B1(_200_),
    .Y(_201_));
 sky130_fd_sc_hd__mux2_1 _473_ (.A0(net43),
    .A1(_201_),
    .S(_168_),
    .X(_030_));
 sky130_fd_sc_hd__nor2_1 _474_ (.A(_262_),
    .B(_039_),
    .Y(_202_));
 sky130_fd_sc_hd__a21oi_1 _475_ (.A1(_187_),
    .A2(_202_),
    .B1(_119_),
    .Y(_203_));
 sky130_fd_sc_hd__nand2_1 _476_ (.A(net44),
    .B(_203_),
    .Y(_204_));
 sky130_fd_sc_hd__mux2i_1 _477_ (.A0(net43),
    .A1(net13),
    .S(_066_),
    .Y(_205_));
 sky130_fd_sc_hd__nor2_1 _478_ (.A(_124_),
    .B(_205_),
    .Y(_206_));
 sky130_fd_sc_hd__a21oi_1 _479_ (.A1(net13),
    .A2(_140_),
    .B1(_206_),
    .Y(_207_));
 sky130_fd_sc_hd__nand2_1 _480_ (.A(net5),
    .B(_183_),
    .Y(_208_));
 sky130_fd_sc_hd__o21ai_0 _481_ (.A1(_055_),
    .A2(_207_),
    .B1(_208_),
    .Y(_209_));
 sky130_fd_sc_hd__mux2i_1 _482_ (.A0(net44),
    .A1(_209_),
    .S(_168_),
    .Y(_210_));
 sky130_fd_sc_hd__nand2_1 _483_ (.A(_204_),
    .B(_210_),
    .Y(_031_));
 sky130_fd_sc_hd__mux2i_1 _484_ (.A0(net44),
    .A1(net14),
    .S(_065_),
    .Y(_211_));
 sky130_fd_sc_hd__nor2_1 _485_ (.A(_124_),
    .B(_211_),
    .Y(_212_));
 sky130_fd_sc_hd__a21oi_1 _486_ (.A1(net14),
    .A2(_140_),
    .B1(_212_),
    .Y(_213_));
 sky130_fd_sc_hd__xor2_1 _487_ (.A(_088_),
    .B(_113_),
    .X(_214_));
 sky130_fd_sc_hd__nand2_1 _488_ (.A(_263_),
    .B(_214_),
    .Y(_215_));
 sky130_fd_sc_hd__a32oi_1 _489_ (.A1(net45),
    .A2(_130_),
    .A3(_215_),
    .B1(_183_),
    .B2(net6),
    .Y(_216_));
 sky130_fd_sc_hd__o21ai_0 _490_ (.A1(_062_),
    .A2(_213_),
    .B1(_216_),
    .Y(_217_));
 sky130_fd_sc_hd__mux2_1 _491_ (.A0(net45),
    .A1(_217_),
    .S(_168_),
    .X(_032_));
 sky130_fd_sc_hd__mux2i_1 _492_ (.A0(_089_),
    .A1(_153_),
    .S(_113_),
    .Y(_218_));
 sky130_fd_sc_hd__a31oi_1 _493_ (.A1(_262_),
    .A2(_259_),
    .A3(_218_),
    .B1(_119_),
    .Y(_219_));
 sky130_fd_sc_hd__o31ai_1 _494_ (.A1(_109_),
    .A2(_167_),
    .A3(_219_),
    .B1(net46),
    .Y(_220_));
 sky130_fd_sc_hd__mux2i_1 _495_ (.A0(net45),
    .A1(net15),
    .S(_066_),
    .Y(_221_));
 sky130_fd_sc_hd__nor2_1 _496_ (.A(_124_),
    .B(_221_),
    .Y(_222_));
 sky130_fd_sc_hd__a21oi_1 _497_ (.A1(net15),
    .A2(_140_),
    .B1(_222_),
    .Y(_223_));
 sky130_fd_sc_hd__nand2_1 _498_ (.A(net7),
    .B(_183_),
    .Y(_224_));
 sky130_fd_sc_hd__o21ai_0 _499_ (.A1(_055_),
    .A2(_223_),
    .B1(_224_),
    .Y(_225_));
 sky130_fd_sc_hd__nand2_1 _500_ (.A(_168_),
    .B(_225_),
    .Y(_226_));
 sky130_fd_sc_hd__nand2_1 _501_ (.A(_220_),
    .B(_226_),
    .Y(_033_));
 sky130_fd_sc_hd__mux2i_1 _502_ (.A0(net46),
    .A1(net16),
    .S(_065_),
    .Y(_227_));
 sky130_fd_sc_hd__nor2_1 _503_ (.A(_124_),
    .B(_227_),
    .Y(_228_));
 sky130_fd_sc_hd__a21oi_1 _504_ (.A1(net16),
    .A2(_140_),
    .B1(_228_),
    .Y(_229_));
 sky130_fd_sc_hd__nand2_1 _505_ (.A(_265_),
    .B(_214_),
    .Y(_230_));
 sky130_fd_sc_hd__a32oi_1 _506_ (.A1(net47),
    .A2(_130_),
    .A3(_230_),
    .B1(_183_),
    .B2(net8),
    .Y(_231_));
 sky130_fd_sc_hd__o21ai_0 _507_ (.A1(_062_),
    .A2(_229_),
    .B1(_231_),
    .Y(_232_));
 sky130_fd_sc_hd__mux2_1 _508_ (.A0(net47),
    .A1(_232_),
    .S(_168_),
    .X(_034_));
 sky130_fd_sc_hd__a21o_1 _509_ (.A1(_069_),
    .A2(_068_),
    .B1(net51),
    .X(_233_));
 sky130_fd_sc_hd__a2111oi_1 _510_ (.A1(_063_),
    .A2(_233_),
    .B1(_142_),
    .C1(_116_),
    .D1(_059_),
    .Y(_234_));
 sky130_fd_sc_hd__a2111o_2 _511_ (.A1(_085_),
    .A2(_128_),
    .B1(_234_),
    .C1(_122_),
    .D1(_082_),
    .X(_235_));
 sky130_fd_sc_hd__mux2_1 _512_ (.A0(_084_),
    .A1(_066_),
    .S(_235_),
    .X(_035_));
 sky130_fd_sc_hd__nand3_1 _513_ (.A(_064_),
    .B(_066_),
    .C(_060_),
    .Y(_236_));
 sky130_fd_sc_hd__nor3_1 _514_ (.A(_062_),
    .B(_074_),
    .C(_236_),
    .Y(_237_));
 sky130_fd_sc_hd__nand2_1 _515_ (.A(_064_),
    .B(_074_),
    .Y(_238_));
 sky130_fd_sc_hd__a211oi_1 _516_ (.A1(_066_),
    .A2(_092_),
    .B1(_238_),
    .C1(_062_),
    .Y(_239_));
 sky130_fd_sc_hd__a221oi_1 _517_ (.A1(cmd_read),
    .A2(_237_),
    .B1(_106_),
    .B2(_103_),
    .C1(_239_),
    .Y(_240_));
 sky130_fd_sc_hd__nor3_1 _518_ (.A(_066_),
    .B(_055_),
    .C(_074_),
    .Y(_241_));
 sky130_fd_sc_hd__o21ai_0 _519_ (.A1(_241_),
    .A2(_235_),
    .B1(_064_),
    .Y(_242_));
 sky130_fd_sc_hd__o21ai_0 _520_ (.A1(_235_),
    .A2(_240_),
    .B1(_242_),
    .Y(_036_));
 sky130_fd_sc_hd__nor2_1 _521_ (.A(_070_),
    .B(_099_),
    .Y(_243_));
 sky130_fd_sc_hd__o22ai_1 _522_ (.A1(_074_),
    .A2(_236_),
    .B1(_243_),
    .B2(_100_),
    .Y(_244_));
 sky130_fd_sc_hd__a21oi_1 _523_ (.A1(_146_),
    .A2(_244_),
    .B1(_239_),
    .Y(_245_));
 sky130_fd_sc_hd__nand2_1 _524_ (.A(_074_),
    .B(_235_),
    .Y(_246_));
 sky130_fd_sc_hd__o21ai_0 _525_ (.A1(_235_),
    .A2(_245_),
    .B1(_246_),
    .Y(_037_));
 sky130_fd_sc_hd__o21ai_0 _526_ (.A1(_098_),
    .A2(_102_),
    .B1(_093_),
    .Y(_247_));
 sky130_fd_sc_hd__mux2_1 _527_ (.A0(_247_),
    .A1(_055_),
    .S(_235_),
    .X(_038_));
 sky130_fd_sc_hd__a21o_1 _528_ (.A1(_078_),
    .A2(_057_),
    .B1(_062_),
    .X(_248_));
 sky130_fd_sc_hd__o211ai_1 _529_ (.A1(_060_),
    .A2(_058_),
    .B1(_248_),
    .C1(_042_),
    .Y(_249_));
 sky130_fd_sc_hd__o21a_1 _530_ (.A1(net26),
    .A2(_042_),
    .B1(_249_),
    .X(_012_));
 sky130_fd_sc_hd__o21ai_0 _531_ (.A1(_269_),
    .A2(_067_),
    .B1(_042_),
    .Y(_250_));
 sky130_fd_sc_hd__o21ai_0 _532_ (.A1(_267_),
    .A2(_042_),
    .B1(_250_),
    .Y(_023_));
 sky130_fd_sc_hd__nand2_1 _533_ (.A(_270_),
    .B(_042_),
    .Y(_251_));
 sky130_fd_sc_hd__o21ai_0 _534_ (.A1(_268_),
    .A2(_042_),
    .B1(_251_),
    .Y(_024_));
 sky130_fd_sc_hd__nand2_1 _535_ (.A(net38),
    .B(_043_),
    .Y(_252_));
 sky130_fd_sc_hd__nand3_1 _536_ (.A(_055_),
    .B(_269_),
    .C(_057_),
    .Y(_253_));
 sky130_fd_sc_hd__o311ai_0 _537_ (.A1(_055_),
    .A2(_270_),
    .A3(_057_),
    .B1(_253_),
    .C1(_042_),
    .Y(_254_));
 sky130_fd_sc_hd__nand2_1 _538_ (.A(_252_),
    .B(_254_),
    .Y(_025_));
 sky130_fd_sc_hd__ha_1 _539_ (.A(_255_),
    .B(_256_),
    .COUT(_257_),
    .SUM(_258_));
 sky130_fd_sc_hd__ha_1 _540_ (.A(_259_),
    .B(_260_),
    .COUT(_261_),
    .SUM(_262_));
 sky130_fd_sc_hd__ha_1 _541_ (.A(net23),
    .B(_260_),
    .COUT(_263_),
    .SUM(_264_));
 sky130_fd_sc_hd__ha_1 _542_ (.A(net23),
    .B(net24),
    .COUT(_265_),
    .SUM(_266_));
 sky130_fd_sc_hd__ha_1 _543_ (.A(_267_),
    .B(_268_),
    .COUT(_269_),
    .SUM(_270_));
 sky130_fd_sc_hd__ha_1 _544_ (.A(_267_),
    .B(net37),
    .COUT(_271_),
    .SUM(_272_));
 sky130_fd_sc_hd__ha_1 _545_ (.A(net36),
    .B(_268_),
    .COUT(_273_),
    .SUM(_274_));
 sky130_fd_sc_hd__ha_1 _546_ (.A(net36),
    .B(net37),
    .COUT(_275_),
    .SUM(_276_));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__buf_4 _548_ (.A(net52),
    .X(scl));
 sky130_fd_sc_hd__buf_4 _549_ (.A(net53),
    .X(sda));
 sky130_fd_sc_hd__dfrtp_1 \ack_error$_DFFE_PN0P_  (.D(_008_),
    .Q(net22),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfstp_1 \bit_counter_debug[0]$_DFFE_PN1P_  (.D(_009_),
    .Q(net23),
    .SET_B(net18),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfstp_2 \bit_counter_debug[1]$_DFFE_PN1P_  (.D(_010_),
    .Q(net24),
    .SET_B(net18),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfstp_1 \bit_counter_debug[2]$_DFFE_PN1P_  (.D(_011_),
    .Q(net25),
    .SET_B(net18),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \busy$_DFFE_PN0N_  (.D(_012_),
    .Q(net26),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \cmd_read$_DFFE_PN0P_  (.D(_013_),
    .Q(cmd_read),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \cmd_write$_DFFE_PN0P_  (.D(_014_),
    .Q(cmd_write),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out[0]$_DFFE_PN0P_  (.D(_015_),
    .Q(net27),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out[1]$_DFFE_PN0P_  (.D(_016_),
    .Q(net28),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out[2]$_DFFE_PN0P_  (.D(_017_),
    .Q(net29),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out[3]$_DFFE_PN0P_  (.D(_018_),
    .Q(net30),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out[4]$_DFFE_PN0P_  (.D(_019_),
    .Q(net31),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out[5]$_DFFE_PN0P_  (.D(_020_),
    .Q(net32),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out[6]$_DFFE_PN0P_  (.D(_021_),
    .Q(net33),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out[7]$_DFFE_PN0P_  (.D(_022_),
    .Q(net34),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \divider_counter[0]$_DFF_PN0_  (.D(_000_),
    .Q(\divider_counter[0] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \divider_counter[1]$_DFF_PN0_  (.D(_001_),
    .Q(\divider_counter[1] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfstp_1 \divider_counter[2]$_DFF_PN1_  (.D(_002_),
    .Q(\divider_counter[2] ),
    .SET_B(net18),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfstp_1 \divider_counter[3]$_DFF_PN1_  (.D(_003_),
    .Q(\divider_counter[3] ),
    .SET_B(net18),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfstp_1 \divider_counter[4]$_DFF_PN1_  (.D(_004_),
    .Q(\divider_counter[4] ),
    .SET_B(net18),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfstp_1 \divider_counter[5]$_DFF_PN1_  (.D(_005_),
    .Q(\divider_counter[5] ),
    .SET_B(net18),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfstp_1 \divider_counter[6]$_DFF_PN1_  (.D(_006_),
    .Q(\divider_counter[6] ),
    .SET_B(net18),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \done$_DFF_PN0_  (.D(_007_),
    .Q(net35),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \phase[0]$_DFFE_PN0N_  (.D(_023_),
    .Q(net36),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \phase[1]$_DFFE_PN0N_  (.D(_024_),
    .Q(net37),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfstp_1 \scl_internal$_DFFE_PN1N_  (.D(_025_),
    .Q(net38),
    .SET_B(net18),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfstp_1 \sda_internal$_DFFE_PN1P_  (.D(_026_),
    .Q(net39),
    .SET_B(net18),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shift_reg_debug[0]$_DFFE_PN0P_  (.D(_027_),
    .Q(net40),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shift_reg_debug[1]$_DFFE_PN0P_  (.D(_028_),
    .Q(net41),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \shift_reg_debug[2]$_DFFE_PN0P_  (.D(_029_),
    .Q(net42),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \shift_reg_debug[3]$_DFFE_PN0P_  (.D(_030_),
    .Q(net43),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \shift_reg_debug[4]$_DFFE_PN0P_  (.D(_031_),
    .Q(net44),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \shift_reg_debug[5]$_DFFE_PN0P_  (.D(_032_),
    .Q(net45),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \shift_reg_debug[6]$_DFFE_PN0P_  (.D(_033_),
    .Q(net46),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \shift_reg_debug[7]$_DFFE_PN0P_  (.D(_034_),
    .Q(net47),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \state[0]$_DFFE_PN0P_  (.D(_035_),
    .Q(net48),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \state[1]$_DFFE_PN0P_  (.D(_036_),
    .Q(net49),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \state[2]$_DFFE_PN0P_  (.D(_037_),
    .Q(net50),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \state[3]$_DFFE_PN0P_  (.D(_038_),
    .Q(net51),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__buf_12 hold1 (.A(net18),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_66 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(addr[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(addr[1]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(addr[2]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(addr[3]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(addr[4]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(addr[5]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(addr[6]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(data_in[0]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(data_in[1]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(data_in[2]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(data_in[3]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(data_in[4]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(data_in[5]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(data_in[6]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(data_in[7]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(read),
    .X(net17));
 sky130_fd_sc_hd__buf_4 input17 (.A(net54),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(start),
    .X(net19));
 sky130_fd_sc_hd__dlymetal6s2s_1 input19 (.A(stop),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(write),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net22),
    .X(ack_error));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net23),
    .X(bit_counter_debug[0]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net24),
    .X(bit_counter_debug[1]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net25),
    .X(bit_counter_debug[2]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net26),
    .X(busy));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net27),
    .X(data_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net28),
    .X(data_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net29),
    .X(data_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(net30),
    .X(data_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output30 (.A(net31),
    .X(data_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(net32),
    .X(data_out[5]));
 sky130_fd_sc_hd__clkbuf_1 output32 (.A(net33),
    .X(data_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output33 (.A(net34),
    .X(data_out[7]));
 sky130_fd_sc_hd__clkbuf_1 output34 (.A(net35),
    .X(done));
 sky130_fd_sc_hd__clkbuf_1 output35 (.A(net36),
    .X(phase[0]));
 sky130_fd_sc_hd__clkbuf_1 output36 (.A(net37),
    .X(phase[1]));
 sky130_fd_sc_hd__clkbuf_1 output37 (.A(net38),
    .X(scl_internal_debug));
 sky130_fd_sc_hd__clkbuf_1 output38 (.A(net39),
    .X(sda_internal_debug));
 sky130_fd_sc_hd__clkbuf_1 output39 (.A(net40),
    .X(shift_reg_debug[0]));
 sky130_fd_sc_hd__clkbuf_1 output40 (.A(net41),
    .X(shift_reg_debug[1]));
 sky130_fd_sc_hd__clkbuf_1 output41 (.A(net42),
    .X(shift_reg_debug[2]));
 sky130_fd_sc_hd__clkbuf_1 output42 (.A(net43),
    .X(shift_reg_debug[3]));
 sky130_fd_sc_hd__clkbuf_1 output43 (.A(net44),
    .X(shift_reg_debug[4]));
 sky130_fd_sc_hd__clkbuf_1 output44 (.A(net45),
    .X(shift_reg_debug[5]));
 sky130_fd_sc_hd__clkbuf_1 output45 (.A(net46),
    .X(shift_reg_debug[6]));
 sky130_fd_sc_hd__clkbuf_1 output46 (.A(net47),
    .X(shift_reg_debug[7]));
 sky130_fd_sc_hd__clkbuf_1 output47 (.A(net48),
    .X(state[0]));
 sky130_fd_sc_hd__clkbuf_1 output48 (.A(net49),
    .X(state[1]));
 sky130_fd_sc_hd__clkbuf_1 output49 (.A(net50),
    .X(state[2]));
 sky130_fd_sc_hd__clkbuf_1 output50 (.A(net51),
    .X(state[3]));
 sky130_fd_sc_hd__conb_1 _548__51 (.LO(net52));
 sky130_fd_sc_hd__conb_1 _549__52 (.LO(net53));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload0 (.A(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkinv_1 clkload1 (.A(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkinv_1 clkload2 (.A(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net54));
 sky130_fd_sc_hd__fill_1 FILLER_0_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_120 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_60 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_66 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_53 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_23 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_151 ();
endmodule
