
* cell bidirectional_fifo
* pin b_to_a_count[1]
* pin b_to_a_count[2]
* pin b_to_a_count[0]
* pin a_almost_empty
* pin b_to_a_count[3]
* pin a_almost_full
* pin a_rd_data[5]
* pin a_rd_data[6]
* pin a_rd_en
* pin b_wr_en
* pin a_rd_data[7]
* pin a_rd_data[2]
* pin a_rd_data[1]
* pin a_full
* pin a_empty
* pin PWELL
* pin NWELL
* pin clk
* pin b_rd_data[3]
* pin b_rd_data[5]
* pin b_rd_data[4]
* pin rst_n
* pin b_wr_data[2]
* pin b_to_a_count[4]
* pin b_rd_data[6]
* pin b_rd_data[0]
* pin b_rd_data[2]
* pin b_rd_data[7]
* pin a_rd_data[0]
* pin a_rd_data[4]
* pin b_rd_data[1]
* pin b_wr_data[1]
* pin a_rd_data[3]
* pin a_to_b_count[3]
* pin b_almost_empty
* pin b_almost_full
* pin a_to_b_count[2]
* pin b_wr_data[3]
* pin a_to_b_count[0]
* pin b_wr_data[0]
* pin b_wr_data[7]
* pin b_wr_data[6]
* pin b_wr_data[4]
* pin a_to_b_count[1]
* pin b_wr_data[5]
* pin a_wr_data[2]
* pin a_wr_data[1]
* pin b_rd_en
* pin a_wr_data[6]
* pin a_wr_data[7]
* pin a_wr_data[0]
* pin a_wr_en
* pin a_wr_data[3]
* pin a_wr_data[5]
* pin a_wr_data[4]
* pin b_empty
* pin b_full
* pin a_to_b_count[4]
.SUBCKT bidirectional_fifo 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 22 162 276
+ 277 278 279 293 328 329 381 382 427 515 551 552 587 588 757 794 795 796 840
+ 881 882 1004 1046 1085 1086 1087 1207 1208 1243 1313 1314 1359 1369 1381 1384
+ 1387 1388 1391 1392
* net 1 b_to_a_count[1]
* net 2 b_to_a_count[2]
* net 3 b_to_a_count[0]
* net 4 a_almost_empty
* net 5 b_to_a_count[3]
* net 6 a_almost_full
* net 7 a_rd_data[5]
* net 8 a_rd_data[6]
* net 9 a_rd_en
* net 10 b_wr_en
* net 11 a_rd_data[7]
* net 12 a_rd_data[2]
* net 13 a_rd_data[1]
* net 14 a_full
* net 15 a_empty
* net 16 PWELL
* net 22 NWELL
* net 162 clk
* net 276 b_rd_data[3]
* net 277 b_rd_data[5]
* net 278 b_rd_data[4]
* net 279 rst_n
* net 293 b_wr_data[2]
* net 328 b_to_a_count[4]
* net 329 b_rd_data[6]
* net 381 b_rd_data[0]
* net 382 b_rd_data[2]
* net 427 b_rd_data[7]
* net 515 a_rd_data[0]
* net 551 a_rd_data[4]
* net 552 b_rd_data[1]
* net 587 b_wr_data[1]
* net 588 a_rd_data[3]
* net 757 a_to_b_count[3]
* net 794 b_almost_empty
* net 795 b_almost_full
* net 796 a_to_b_count[2]
* net 840 b_wr_data[3]
* net 881 a_to_b_count[0]
* net 882 b_wr_data[0]
* net 1004 b_wr_data[7]
* net 1046 b_wr_data[6]
* net 1085 b_wr_data[4]
* net 1086 a_to_b_count[1]
* net 1087 b_wr_data[5]
* net 1207 a_wr_data[2]
* net 1208 a_wr_data[1]
* net 1243 b_rd_en
* net 1313 a_wr_data[6]
* net 1314 a_wr_data[7]
* net 1359 a_wr_data[0]
* net 1369 a_wr_en
* net 1381 a_wr_data[3]
* net 1384 a_wr_data[5]
* net 1387 a_wr_data[4]
* net 1388 b_empty
* net 1391 b_full
* net 1392 a_to_b_count[4]
* cell instance $3 r0 *1 357.96,1.4
X$3 28 16 22 1 BUF_X1
* cell instance $9 r0 *1 358.53,1.4
X$9 27 16 22 2 BUF_X1
* cell instance $15 r0 *1 359.1,1.4
X$15 34 16 22 3 BUF_X1
* cell instance $20 m0 *1 362.14,4.2
X$20 44 16 22 4 BUF_X1
* cell instance $26 m0 *1 361.57,4.2
X$26 24 16 22 5 BUF_X1
* cell instance $32 r0 *1 361.95,1.4
X$32 20 16 22 6 BUF_X1
* cell instance $39 r0 *1 363.09,1.4
X$39 19 16 22 7 BUF_X1
* cell instance $44 m0 *1 364.99,4.2
X$44 21 16 22 8 BUF_X1
* cell instance $54 r0 *1 365.18,231
X$54 9 16 22 23 CLKBUF_X3
* cell instance $60 r0 *1 366.32,298.2
X$60 10 16 22 25 BUF_X2
* cell instance $63 r0 *1 367.84,1.4
X$63 18 16 22 11 BUF_X1
* cell instance $68 m0 *1 371.83,4.2
X$68 322 16 22 12 BUF_X1
* cell instance $75 r0 *1 373.54,1.4
X$75 17 16 22 13 BUF_X1
* cell instance $80 r0 *1 374.87,1.4
X$80 40 16 22 14 BUF_X1
* cell instance $87 r0 *1 383.23,1.4
X$87 26 16 22 15 BUF_X1
* cell instance $91 m0 *1 359.67,345.8
X$91 261 199 271 16 22 272 MUX2_X1
* cell instance $93 m0 *1 361,345.8
X$93 255 150 22 16 271 AND2_X1
* cell instance $94 m0 *1 361.76,345.8
X$94 16 53 262 272 125 22 DFF_X1
* cell instance $95 m0 *1 364.99,345.8
X$95 16 143 246 275 125 22 DFF_X1
* cell instance $99 m0 *1 378.1,345.8
X$99 201 231 41 22 16 254 OAI21_X4
* cell instance $102 m0 *1 381.52,345.8
X$102 16 1404 264 273 307 22 DFF_X1
* cell instance $103 m0 *1 384.75,345.8
X$103 264 54 195 16 22 273 MUX2_X1
* cell instance $108 m0 *1 354.35,345.8
X$108 16 1453 260 258 104 22 DFF_X1
* cell instance $112 r0 *1 354.16,345.8
X$112 260 257 22 16 280 AND2_X1
* cell instance $113 r0 *1 354.92,345.8
X$113 280 274 281 16 22 258 MUX2_X1
* cell instance $114 r0 *1 356.25,345.8
X$114 259 260 16 22 281 NOR2_X1
* cell instance $117 r0 *1 359.1,345.8
X$117 300 257 22 16 261 AND2_X1
* cell instance $123 r0 *1 362.14,345.8
X$123 152 262 300 22 16 302 HA_X1
* cell instance $125 r0 *1 364.8,345.8
X$125 301 231 79 16 274 22 AOI21_X1
* cell instance $127 r0 *1 367.08,345.8
X$127 246 16 22 282 CLKBUF_X3
* cell instance $129 r0 *1 368.22,345.8
X$129 262 16 22 263 BUF_X2
* cell instance $133 r0 *1 371.07,345.8
X$133 221 231 41 22 16 304 OAI21_X4
* cell instance $135 r0 *1 373.73,345.8
X$135 222 231 41 22 16 332 OAI21_X4
* cell instance $136 r0 *1 376.2,345.8
X$136 156 231 41 22 16 637 OAI21_X4
* cell instance $137 r0 *1 378.67,345.8
X$137 203 231 41 22 16 514 OAI21_X4
* cell instance $141 r0 *1 383.23,345.8
X$141 263 22 286 16 BUF_X4
* cell instance $145 r0 *1 386.65,345.8
X$145 309 65 195 16 22 284 MUX2_X1
* cell instance $148 r0 *1 390.26,345.8
X$148 16 1623 265 310 307 22 DFF_X1
* cell instance $149 r0 *1 393.49,345.8
X$149 265 181 168 16 22 310 MUX2_X1
* cell instance $156 m0 *1 397.29,345.8
X$156 266 22 114 16 BUF_X4
* cell instance $162 r0 *1 397.48,345.8
X$162 265 114 267 16 22 324 MUX2_X1
* cell instance $168 r0 *1 404.7,345.8
X$168 285 54 183 16 22 305 MUX2_X1
* cell instance $172 r0 *1 407.36,345.8
X$172 287 65 183 16 22 288 MUX2_X1
* cell instance $176 m0 *1 417.24,345.8
X$176 239 286 250 16 22 292 MUX2_X1
* cell instance $181 m0 *1 423.51,345.8
X$181 16 1539 244 247 213 22 DFF_X1
* cell instance $186 r0 *1 425.79,345.8
X$186 244 114 240 16 22 268 MUX2_X1
* cell instance $188 m0 *1 429.59,345.8
X$188 211 114 241 16 22 366 MUX2_X1
* cell instance $192 m0 *1 431.87,345.8
X$192 16 1516 241 269 213 22 DFF_X1
* cell instance $859 m0 *1 2.85,348.6
X$859 294 16 22 278 BUF_X1
* cell instance $902 r0 *1 2.09,348.6
X$902 335 16 22 277 BUF_X1
* cell instance $976 m0 *1 305.33,348.6
X$976 16 314 104 1663 296 22 DFF_X2
* cell instance $983 m0 *1 345.42,348.6
X$983 279 16 22 174 BUF_X2
* cell instance $988 m0 *1 357.01,348.6
X$988 16 216 299 297 317 22 DFF_X1
* cell instance $990 m0 *1 361.76,348.6
X$990 299 16 22 319 CLKBUF_X3
* cell instance $1009 r0 *1 305.71,348.6
X$1009 311 296 312 16 22 342 NAND3_X1
* cell instance $1013 r0 *1 314.26,348.6
X$1013 16 336 315 1671 294 22 DFF_X2
* cell instance $1027 r0 *1 354.16,348.6
X$1027 174 16 22 311 CLKBUF_X3
* cell instance $1038 r0 *1 364.04,348.6
X$1038 259 319 16 22 318 NOR2_X1
* cell instance $1039 m0 *1 365.18,348.6
X$1039 302 319 282 23 16 22 301 NAND4_X1
* cell instance $1040 m0 *1 364.61,348.6
X$1040 259 282 16 22 303 NOR2_X1
* cell instance $1041 m0 *1 366.13,348.6
X$1041 302 23 16 22 337 NAND2_X1
* cell instance $1046 r0 *1 366.7,348.6
X$1046 337 231 200 16 338 22 AOI21_X1
* cell instance $1048 m0 *1 367.08,348.6
X$1048 283 338 303 16 22 275 MUX2_X1
* cell instance $1051 m0 *1 380.76,348.6
X$1051 263 22 308 16 BUF_X4
* cell instance $1054 m0 *1 383.04,348.6
X$1054 263 22 266 16 BUF_X4
* cell instance $1057 m0 *1 385.32,348.6
X$1057 264 308 309 16 22 499 MUX2_X1
* cell instance $1058 m0 *1 386.65,348.6
X$1058 16 1403 309 284 307 22 DFF_X1
* cell instance $1061 m0 *1 394.44,348.6
X$1061 16 1402 267 306 307 22 DFF_X1
* cell instance $1062 m0 *1 397.67,348.6
X$1062 267 212 168 16 22 306 MUX2_X1
* cell instance $1065 m0 *1 402.23,348.6
X$1065 16 1462 285 305 289 22 DFF_X1
* cell instance $1068 r0 *1 367.46,348.6
X$1068 109 379 16 22 283 NOR2_X1
* cell instance $1072 r0 *1 386.27,348.6
X$1072 159 16 22 307 CLKBUF_X3
* cell instance $1073 r0 *1 387.22,348.6
X$1073 307 16 22 1692 INV_X1
* cell instance $1081 m0 *1 407.93,348.6
X$1081 16 1452 287 288 289 22 DFF_X1
* cell instance $1082 m0 *1 406.6,348.6
X$1082 285 286 287 16 22 449 MUX2_X1
* cell instance $1084 m0 *1 412.87,348.6
X$1084 16 1427 290 298 289 22 DFF_X1
* cell instance $1085 m0 *1 411.54,348.6
X$1085 290 238 70 16 22 298 MUX2_X1
* cell instance $1086 m0 *1 416.1,348.6
X$1086 290 308 291 16 22 334 MUX2_X1
* cell instance $1087 m0 *1 417.43,348.6
X$1087 291 227 70 16 22 295 MUX2_X1
* cell instance $1088 m0 *1 418.76,348.6
X$1088 16 1397 291 295 289 22 DFF_X1
* cell instance $1105 r0 *1 421.61,348.6
X$1105 327 225 359 16 22 325 MUX2_X1
* cell instance $1110 r0 *1 431.49,348.6
X$1110 327 16 22 70 BUF_X2
* cell instance $1111 r0 *1 432.25,348.6
X$1111 70 332 326 16 22 331 MUX2_X1
* cell instance $1113 r0 *1 433.96,348.6
X$1113 16 1560 326 331 363 22 DFF_X1
* cell instance $1118 r0 *1 442.89,348.6
X$1118 293 16 22 327 CLKBUF_X2
* cell instance $1221 m0 *1 706.8,348.6
X$1221 39 16 22 328 BUF_X1
* cell instance $1233 m0 *1 294.5,354.2
X$1233 410 464 432 16 22 463 MUX2_X1
* cell instance $1234 m0 *1 296.02,354.2
X$1234 16 1482 410 463 339 22 DFF_X1
* cell instance $1236 m0 *1 299.44,354.2
X$1236 384 466 432 16 22 411 MUX2_X1
* cell instance $1242 m0 *1 288.04,354.2
X$1242 16 1534 383 406 339 22 DFF_X1
* cell instance $1244 m0 *1 291.27,354.2
X$1244 383 340 572 16 22 406 MUX2_X1
* cell instance $1248 r0 *1 288.04,354.2
X$1248 316 16 22 339 CLKBUF_X3
* cell instance $1249 r0 *1 288.99,354.2
X$1249 339 16 22 CLKBUF_X1
* cell instance $1254 r0 *1 298.3,354.2
X$1254 410 430 384 16 22 435 MUX2_X1
* cell instance $1259 r0 *1 302.48,354.2
X$1259 553 464 572 16 22 467 MUX2_X1
* cell instance $1261 r0 *1 305.33,354.2
X$1261 311 434 312 16 22 436 NAND3_X1
* cell instance $1262 r0 *1 306.09,354.2
X$1262 344 343 345 434 16 22 493 NAND4_X1
* cell instance $1266 r0 *1 309.13,354.2
X$1266 16 437 536 1669 456 22 DFF_X2
* cell instance $1270 r0 *1 314.07,354.2
X$1270 16 1618 438 470 315 22 DFF_X1
* cell instance $1271 m0 *1 315.78,354.2
X$1271 438 570 385 16 22 470 MUX2_X1
* cell instance $1273 m0 *1 317.11,354.2
X$1273 16 1530 472 473 315 22 DFF_X1
* cell instance $1276 m0 *1 323.57,354.2
X$1276 344 343 345 386 16 22 474 NAND4_X1
* cell instance $1277 m0 *1 324.52,354.2
X$1277 16 439 348 1661 386 22 DFF_X2
* cell instance $1278 m0 *1 328.13,354.2
X$1278 476 386 312 16 22 475 NAND3_X1
* cell instance $1282 m0 *1 341.24,354.2
X$1282 480 340 418 16 22 417 MUX2_X1
* cell instance $1283 m0 *1 342.57,354.2
X$1283 259 387 16 22 418 NOR2_X1
* cell instance $1285 m0 *1 343.33,354.2
X$1285 387 257 22 16 480 AND2_X1
* cell instance $1289 m0 *1 357.77,354.2
X$1289 349 16 22 109 CLKBUF_X3
* cell instance $1293 r0 *1 317.49,354.2
X$1293 438 430 472 16 22 471 MUX2_X1
* cell instance $1297 r0 *1 325.47,354.2
X$1297 475 474 620 16 22 439 NAND3_X1
* cell instance $1301 r0 *1 330.41,354.2
X$1301 150 16 22 476 CLKBUF_X3
* cell instance $1304 r0 *1 334.59,354.2
X$1304 349 312 440 16 22 NOR2_X4
* cell instance $1310 r0 *1 345.23,354.2
X$1310 387 442 16 22 825 XNOR2_X2
* cell instance $1312 r0 *1 347.32,354.2
X$1312 484 482 483 16 22 481 MUX2_X1
* cell instance $1318 m0 *1 362.33,354.2
X$1318 259 522 16 22 388 NOR2_X1
* cell instance $1324 m0 *1 364.8,354.2
X$1324 152 16 22 445 BUF_X2
* cell instance $1326 m0 *1 368.79,354.2
X$1326 16 425 317 1660 322 22 DFF_X2
* cell instance $1327 m0 *1 372.4,354.2
X$1327 476 322 443 16 22 444 NAND3_X1
* cell instance $1328 m0 *1 373.16,354.2
X$1328 444 389 421 16 22 425 NAND3_X1
* cell instance $1330 m0 *1 374.11,354.2
X$1330 476 17 443 16 22 424 NAND3_X1
* cell instance $1331 m0 *1 374.87,354.2
X$1331 16 491 307 1667 17 22 DFF_X2
* cell instance $1337 r0 *1 365.94,354.2
X$1337 200 29 345 19 16 22 531 NAND4_X1
* cell instance $1342 r0 *1 369.74,354.2
X$1342 349 443 392 16 22 NOR2_X4
* cell instance $1345 r0 *1 373.35,354.2
X$1345 445 16 22 402 CLKBUF_X3
* cell instance $1348 m0 *1 385.51,354.2
X$1348 16 1419 390 426 353 22 DFF_X1
* cell instance $1349 m0 *1 384.18,354.2
X$1349 323 286 390 16 22 446 MUX2_X1
* cell instance $1353 m0 *1 392.73,354.2
X$1353 159 16 22 353 CLKBUF_X3
* cell instance $1354 m0 *1 393.68,354.2
X$1354 16 1401 391 490 353 22 DFF_X1
* cell instance $1355 m0 *1 396.91,354.2
X$1355 375 114 391 16 22 487 MUX2_X1
* cell instance $1359 m0 *1 407.55,354.2
X$1359 39 41 397 478 392 421 16 22 OAI221_X2
* cell instance $1360 m0 *1 409.64,354.2
X$1360 39 41 413 479 392 419 16 22 OAI221_X2
* cell instance $1363 m0 *1 412.68,354.2
X$1363 394 452 477 451 395 396 16 22 479 OAI33_X1
* cell instance $1364 m0 *1 414.01,354.2
X$1364 394 525 453 451 416 358 16 22 478 OAI33_X1
* cell instance $1369 r0 *1 394.06,354.2
X$1369 353 16 22 1689 INV_X1
* cell instance $1372 r0 *1 396.72,354.2
X$1372 110 356 16 22 447 NOR2_X1
* cell instance $1374 r0 *1 398.05,354.2
X$1374 487 393 16 22 489 NOR2_X1
* cell instance $1376 r0 *1 398.81,354.2
X$1376 324 393 16 22 566 NOR2_X1
* cell instance $1379 r0 *1 401.28,354.2
X$1379 445 16 22 393 CLKBUF_X3
* cell instance $1383 r0 *1 404.89,354.2
X$1383 486 393 16 22 504 NOR2_X1
* cell instance $1386 r0 *1 406.6,354.2
X$1386 448 393 16 22 485 NOR2_X1
* cell instance $1390 r0 *1 408.5,354.2
X$1390 449 356 16 22 450 NOR2_X1
* cell instance $1396 r0 *1 414.96,354.2
X$1396 457 501 16 22 453 NOR2_X1
* cell instance $1400 m0 *1 418.76,354.2
X$1400 321 398 400 423 401 468 16 22 397 OAI33_X1
* cell instance $1401 m0 *1 420.28,354.2
X$1401 365 522 16 22 468 NOR2_X1
* cell instance $1402 m0 *1 420.85,354.2
X$1402 321 399 409 423 465 403 16 22 413 OAI33_X1
* cell instance $1404 m0 *1 422.37,354.2
X$1404 462 402 16 22 465 NOR2_X1
* cell instance $1405 m0 *1 422.94,354.2
X$1405 87 304 407 16 22 459 MUX2_X1
* cell instance $1406 m0 *1 424.27,354.2
X$1406 16 1480 407 459 289 22 DFF_X1
* cell instance $1410 r0 *1 419.71,354.2
X$1410 268 393 16 22 523 NOR2_X1
* cell instance $1413 r0 *1 421.42,354.2
X$1413 210 393 16 22 512 NOR2_X1
* cell instance $1415 r0 *1 423.51,354.2
X$1415 461 255 407 16 22 462 MUX2_X1
* cell instance $1417 m0 *1 431.11,354.2
X$1417 16 1535 404 458 363 22 DFF_X1
* cell instance $1422 m0 *1 438.33,354.2
X$1422 362 286 455 16 22 457 MUX2_X1
* cell instance $1433 r0 *1 437,354.2
X$1433 159 16 22 363 CLKBUF_X3
* cell instance $1548 m0 *1 1.33,351.4
X$1548 313 16 22 329 BUF_X1
* cell instance $1650 m0 *1 304.57,351.4
X$1650 333 368 367 16 22 330 NAND3_X1
* cell instance $1651 m0 *1 305.33,351.4
X$1651 311 313 312 16 22 333 NAND3_X1
* cell instance $1652 m0 *1 306.09,351.4
X$1652 344 343 150 313 16 22 368 NAND4_X1
* cell instance $1653 m0 *1 307.04,351.4
X$1653 344 343 345 296 16 22 369 NAND4_X1
* cell instance $1665 r0 *1 280.63,351.4
X$1665 16 1570 341 405 339 22 DFF_X1
* cell instance $1666 r0 *1 283.86,351.4
X$1666 341 340 432 16 22 405 MUX2_X1
* cell instance $1671 r0 *1 298.49,351.4
X$1671 16 1567 384 411 339 22 DFF_X1
* cell instance $1674 r0 *1 302.67,351.4
X$1674 16 330 315 1674 313 22 DFF_X2
* cell instance $1675 r0 *1 306.28,351.4
X$1675 342 369 412 16 22 314 NAND3_X1
* cell instance $1676 r0 *1 307.04,351.4
X$1676 16 414 315 1673 335 22 DFF_X2
* cell instance $1677 m0 *1 309.32,351.4
X$1677 311 335 312 16 22 370 NAND3_X1
* cell instance $1680 m0 *1 310.27,351.4
X$1680 344 343 345 335 16 22 415 NAND4_X1
* cell instance $1684 r0 *1 310.65,351.4
X$1684 370 415 346 16 22 414 NAND3_X1
* cell instance $1686 m0 *1 316.35,351.4
X$1686 372 347 373 16 22 336 NAND3_X1
* cell instance $1687 m0 *1 315.4,351.4
X$1687 344 343 345 294 16 22 347 NAND4_X1
* cell instance $1688 m0 *1 317.11,351.4
X$1688 311 294 312 16 22 372 NAND3_X1
* cell instance $1698 r0 *1 318.06,351.4
X$1698 472 340 385 16 22 473 MUX2_X1
* cell instance $1704 r0 *1 341.05,351.4
X$1704 16 1598 387 417 348 22 DFF_X1
* cell instance $1706 m0 *1 350.36,351.4
X$1706 174 16 22 349 INV_X2
* cell instance $1711 m0 *1 351.31,351.4
X$1711 174 16 22 257 BUF_X2
* cell instance $1715 m0 *1 353.97,351.4
X$1715 174 16 22 345 CLKBUF_X3
* cell instance $1720 r0 *1 354.73,351.4
X$1720 349 16 22 259 CLKBUF_X3
* cell instance $1723 r0 *1 356.63,351.4
X$1723 16 378 317 422 152 22 DFF_X2
* cell instance $1724 r0 *1 360.24,351.4
X$1724 422 150 22 16 420 AND2_X1
* cell instance $1726 r0 *1 361.19,351.4
X$1726 420 199 388 16 22 378 MUX2_X1
* cell instance $1728 m0 *1 363.09,351.4
X$1728 380 350 318 16 22 297 MUX2_X1
* cell instance $1732 m0 *1 366.13,351.4
X$1732 320 231 200 16 350 22 AOI21_X1
* cell instance $1733 m0 *1 365.56,351.4
X$1733 109 351 16 22 380 NOR2_X1
* cell instance $1735 m0 *1 367.65,351.4
X$1735 282 16 22 379 INV_X2
* cell instance $1736 m0 *1 368.22,351.4
X$1736 319 16 22 351 INV_X2
* cell instance $1737 m0 *1 368.79,351.4
X$1737 351 379 16 321 22 NAND2_X4
* cell instance $1738 m0 *1 370.5,351.4
X$1738 351 282 16 394 22 NAND2_X4
* cell instance $1744 r0 *1 365.75,351.4
X$1744 23 16 22 443 INV_X2
* cell instance $1745 r0 *1 366.32,351.4
X$1745 282 255 402 23 16 22 320 NAND4_X1
* cell instance $1747 r0 *1 368.79,351.4
X$1747 319 379 16 423 22 NAND2_X4
* cell instance $1748 r0 *1 370.5,351.4
X$1748 319 282 16 451 22 NAND2_X4
* cell instance $1750 r0 *1 372.4,351.4
X$1750 200 29 311 322 16 22 389 NAND4_X1
* cell instance $1754 r0 *1 375.82,351.4
X$1754 200 29 311 17 16 22 352 NAND4_X1
* cell instance $1755 r0 *1 376.77,351.4
X$1755 424 352 419 16 22 491 NAND3_X1
* cell instance $1759 r0 *1 380,351.4
X$1759 16 1651 323 377 307 22 DFF_X1
* cell instance $1760 m0 *1 382.66,351.4
X$1760 323 181 195 16 22 377 MUX2_X1
* cell instance $1768 r0 *1 385.89,351.4
X$1768 390 212 195 16 22 426 MUX2_X1
* cell instance $1771 r0 *1 390.45,351.4
X$1771 16 1624 375 376 353 22 DFF_X1
* cell instance $1773 m0 *1 391.21,351.4
X$1773 375 181 83 16 22 376 MUX2_X1
* cell instance $1775 m0 *1 401.66,351.4
X$1775 354 181 64 16 22 374 MUX2_X1
* cell instance $1779 r0 *1 393.87,351.4
X$1779 391 212 83 16 22 490 MUX2_X1
* cell instance $1781 r0 *1 395.96,351.4
X$1781 786 16 22 159 CLKBUF_X3
* cell instance $1785 r0 *1 400.52,351.4
X$1785 16 1550 354 374 353 22 DFF_X1
* cell instance $1786 r0 *1 403.75,351.4
X$1786 354 114 371 16 22 486 MUX2_X1
* cell instance $1787 m0 *1 405.08,351.4
X$1787 371 212 64 16 22 355 MUX2_X1
* cell instance $1794 r0 *1 405.27,351.4
X$1794 16 1643 371 355 353 22 DFF_X1
* cell instance $1797 r0 *1 413.06,351.4
X$1797 112 356 16 22 396 NOR2_X1
* cell instance $1800 r0 *1 414.2,351.4
X$1800 357 356 16 22 358 NOR2_X1
* cell instance $1803 r0 *1 416.67,351.4
X$1803 366 393 16 22 395 NOR2_X1
* cell instance $1805 m0 *1 417.62,351.4
X$1805 159 16 22 289 CLKBUF_X3
* cell instance $1807 m0 *1 418.57,351.4
X$1807 289 16 22 CLKBUF_X1
* cell instance $1809 m0 *1 420.66,351.4
X$1809 16 1423 359 325 289 22 DFF_X1
* cell instance $1810 m0 *1 423.89,351.4
X$1810 359 255 361 16 22 408 MUX2_X1
* cell instance $1813 r0 *1 418.19,351.4
X$1813 334 356 16 22 398 NOR2_X1
* cell instance $1814 r0 *1 418.76,351.4
X$1814 292 356 16 22 399 NOR2_X1
* cell instance $1815 r0 *1 419.33,351.4
X$1815 115 393 16 22 400 NOR2_X1
* cell instance $1818 r0 *1 420.47,351.4
X$1818 164 393 16 22 416 NOR2_X1
* cell instance $1819 r0 *1 421.04,351.4
X$1819 408 402 16 22 401 NOR2_X1
* cell instance $1820 r0 *1 421.61,351.4
X$1820 116 393 16 22 409 NOR2_X1
* cell instance $1886 m0 *1 280.44,354.2
X$1886 16 1536 428 429 339 22 DFF_X1
* cell instance $1889 r0 *1 280.44,354.2
X$1889 428 340 460 16 22 429 MUX2_X1
* cell instance $1893 r0 *1 283.86,354.2
X$1893 431 430 341 16 22 433 MUX2_X1
* cell instance $16987 m0 *1 306.85,410.2
X$16987 1298 1228 1377 16 22 1383 MUX2_X1
* cell instance $16988 m0 *1 308.18,410.2
X$16988 16 1406 1377 1383 1361 22 DFF_X1
* cell instance $16991 m0 *1 312.93,410.2
X$16991 16 1475 1378 1385 1299 22 DFF_X1
* cell instance $19365 m0 *1 277.02,404.6
X$19365 1334 1242 1354 16 22 1370 MUX2_X1
* cell instance $19368 m0 *1 278.54,404.6
X$19368 1334 1228 1371 16 22 1364 MUX2_X1
* cell instance $19370 r0 *1 278.73,404.6
X$19370 16 1631 1371 1364 1318 22 DFF_X1
* cell instance $19375 m0 *1 286.52,404.6
X$19375 16 1502 1352 1365 1361 22 DFF_X1
* cell instance $19378 r0 *1 289.18,404.6
X$19378 1351 1242 1366 16 22 1373 MUX2_X1
* cell instance $19380 r0 *1 290.51,404.6
X$19380 1366 930 1367 16 22 1095 MUX2_X1
* cell instance $19383 r0 *1 293.74,404.6
X$19383 1351 1228 1367 16 22 1368 MUX2_X1
* cell instance $19389 m0 *1 305.14,404.6
X$19389 16 1400 1363 1376 1361 22 DFF_X1
* cell instance $19392 m0 *1 309.89,404.6
X$19392 16 1524 1355 1375 1361 22 DFF_X1
* cell instance $19395 m0 *1 313.5,404.6
X$19395 16 1501 1356 1372 1325 22 DFF_X1
* cell instance $19398 m0 *1 318.44,404.6
X$19398 16 1474 1357 1374 1325 22 DFF_X1
* cell instance $19684 r0 *1 266.19,396.2
X$19684 1314 16 22 1292 CLKBUF_X2
* cell instance $19686 r0 *1 269.99,396.2
X$19686 16 1553 1346 1315 1318 22 DFF_X1
* cell instance $19692 r0 *1 277.97,396.2
X$19692 1292 1228 1316 16 22 1332 MUX2_X1
* cell instance $19697 r0 *1 282.15,396.2
X$19697 1292 1112 1319 16 22 1317 MUX2_X1
* cell instance $19700 r0 *1 284.24,396.2
X$19700 1334 16 22 432 BUF_X2
* cell instance $19702 r0 *1 285.76,396.2
X$19702 1334 1027 1321 16 22 1320 MUX2_X1
* cell instance $19705 m0 *1 288.42,396.2
X$19705 16 1510 1293 1336 1258 22 DFF_X1
* cell instance $19707 r0 *1 288.8,396.2
X$19707 432 1252 1293 16 22 1336 MUX2_X1
* cell instance $19709 m0 *1 291.65,396.2
X$19709 1321 1219 1293 16 22 1177 MUX2_X1
* cell instance $19715 r0 *1 300.01,396.2
X$19715 16 1634 1297 1295 1275 22 DFF_X1
* cell instance $19717 m0 *1 300.39,396.2
X$19717 432 1214 1297 16 22 1295 MUX2_X1
* cell instance $19718 m0 *1 301.72,396.2
X$19718 1352 1219 1297 16 22 1261 MUX2_X1
* cell instance $19722 r0 *1 304.38,396.2
X$19722 572 1214 1323 16 22 1324 MUX2_X1
* cell instance $19727 r0 *1 309.7,396.2
X$19727 1298 1027 1339 16 22 1340 MUX2_X1
* cell instance $19731 m0 *1 311.79,396.2
X$19731 1298 16 22 649 BUF_X2
* cell instance $19735 r0 *1 313.69,396.2
X$19735 1298 1112 1337 16 22 1338 MUX2_X1
* cell instance $19738 r0 *1 316.73,396.2
X$19738 1335 16 22 385 BUF_X2
* cell instance $19740 r0 *1 318.25,396.2
X$19740 1335 1027 1326 16 22 1333 MUX2_X1
* cell instance $19744 r0 *1 320.72,396.2
X$19744 385 1214 1330 16 22 1331 MUX2_X1
* cell instance $19745 r0 *1 322.05,396.2
X$19745 16 1576 1330 1331 1325 22 DFF_X1
* cell instance $19752 r0 *1 332.5,396.2
X$19752 16 1604 1300 1301 1299 22 DFF_X1
* cell instance $19753 m0 *1 332.5,396.2
X$19753 1280 1242 1300 16 22 1301 MUX2_X1
* cell instance $20062 r0 *1 358.91,320.6
X$20062 32 16 22 34 INV_X4
* cell instance $20065 m0 *1 360.05,320.6
X$20065 33 32 22 42 16 XOR2_X2
* cell instance $20070 m0 *1 361.95,320.6
X$20070 38 16 22 24 INV_X4
* cell instance $20079 m0 *1 383.42,320.6
X$20079 16 39 22 37 BUF_X8
* cell instance $20370 r0 *1 358.15,323.4
X$20370 46 16 22 31 INV_X4
* cell instance $20373 m0 *1 358.91,323.4
X$20373 33 16 22 45 INV_X1
* cell instance $20374 r0 *1 359.1,323.4
X$20374 36 32 45 46 22 16 50 AND4_X1
* cell instance $20375 m0 *1 359.29,323.4
X$20375 31 33 34 36 16 22 43 NOR4_X1
* cell instance $20377 m0 *1 360.24,323.4
X$20377 36 34 33 31 16 22 47 OR4_X1
* cell instance $20380 m0 *1 361.38,323.4
X$20380 48 36 22 38 16 XOR2_X2
* cell instance $20381 r0 *1 361.38,323.4
X$20381 51 48 47 16 22 49 MUX2_X1
* cell instance $20382 r0 *1 362.71,323.4
X$20382 50 43 48 22 16 96 MUX2_X2
* cell instance $20385 r0 *1 365.18,323.4
X$20385 16 41 22 49 BUF_X8
* cell instance $20680 r0 *1 357.77,326.2
X$20680 52 60 16 22 46 XNOR2_X2
* cell instance $20683 m0 *1 359.48,326.2
X$20683 46 45 32 36 16 22 51 NAND4_X1
* cell instance $20705 r0 *1 400.52,326.2
X$20705 16 1555 57 58 55 22 DFF_X1
* cell instance $23399 m0 *1 316.92,413
X$23399 1384 16 22 1298 CLKBUF_X2
* cell instance $23404 m0 *1 322.62,413
X$23404 1387 16 22 1335 CLKBUF_X2
* cell instance $68077 r0 *1 270.75,379.4
X$68077 1057 1141 1129 16 22 1167 MUX2_X1
* cell instance $68079 r0 *1 273.6,379.4
X$68079 16 1543 1116 1169 864 22 DFF_X1
* cell instance $68080 m0 *1 275.12,379.4
X$68080 1121 16 22 864 CLKBUF_X3
* cell instance $68081 m0 *1 274.36,379.4
X$68081 1057 16 22 740 BUF_X2
* cell instance $68082 m0 *1 276.07,379.4
X$68082 864 16 22 1685 INV_X1
* cell instance $68085 r0 *1 276.83,379.4
X$68085 1116 653 1142 16 22 1170 MUX2_X1
* cell instance $68086 r0 *1 278.16,379.4
X$68086 1170 1037 16 22 1059 NOR2_X1
* cell instance $68087 m0 *1 278.54,379.4
X$68087 1060 1037 16 22 1030 NOR2_X1
* cell instance $68095 r0 *1 279.68,379.4
X$68095 1131 1054 16 22 1061 NOR2_X1
* cell instance $68096 r0 *1 280.25,379.4
X$68096 1286 1117 16 22 1031 NOR2_X1
* cell instance $68099 r0 *1 281.77,379.4
X$68099 1171 1117 16 22 1010 NOR2_X1
* cell instance $68102 r0 *1 284.05,379.4
X$68102 1117 16 22 949 CLKBUF_X3
* cell instance $68103 m0 *1 286.14,379.4
X$68103 16 1476 1062 1093 864 22 DFF_X1
* cell instance $68104 m0 *1 284.81,379.4
X$68104 1057 1112 1062 16 22 1093 MUX2_X1
* cell instance $68111 r0 *1 289.37,379.4
X$68111 1054 16 22 1117 INV_X2
* cell instance $68113 m0 *1 291.46,379.4
X$68113 1095 1037 16 22 1096 NOR2_X1
* cell instance $68117 m0 *1 295.83,379.4
X$68117 1062 947 1063 16 22 1097 MUX2_X1
* cell instance $68120 m0 *1 298.87,379.4
X$68120 435 1029 16 22 1135 NOR2_X1
* cell instance $68123 r0 *1 294.5,379.4
X$68123 740 1214 1063 16 22 1145 MUX2_X1
* cell instance $68126 m0 *1 300.01,379.4
X$68126 1097 1069 16 22 1064 NOR2_X1
* cell instance $68128 m0 *1 300.58,379.4
X$68128 1134 1065 16 22 1099 NOR2_X1
* cell instance $68129 m0 *1 301.15,379.4
X$68129 1133 1065 16 22 1067 NOR2_X1
* cell instance $68134 r0 *1 300.58,379.4
X$68134 1176 949 16 22 1180 NOR2_X1
* cell instance $68135 r0 *1 301.15,379.4
X$68135 1178 1069 16 22 1066 NOR2_X1
* cell instance $68136 r0 *1 301.72,379.4
X$68136 1098 1146 1135 1034 1147 1181 16 22 1137 OAI33_X1
* cell instance $68137 r0 *1 303.05,379.4
X$68137 1098 1180 1014 1034 1179 1184 16 22 1101 OAI33_X1
* cell instance $68138 r0 *1 304.38,379.4
X$68138 1118 1069 16 22 1179 NOR2_X1
* cell instance $68140 r0 *1 305.14,379.4
X$68140 1183 1065 16 22 1120 NOR2_X1
* cell instance $68144 m0 *1 306.66,379.4
X$68144 1102 1029 16 22 1119 NOR2_X1
* cell instance $68147 r0 *1 306.66,379.4
X$68147 1098 1186 1119 1034 1148 1120 16 22 1103 OAI33_X1
* cell instance $68150 r0 *1 309.13,379.4
X$68150 1241 1037 16 22 1035 NOR2_X1
* cell instance $68153 m0 *1 309.89,379.4
X$68153 1068 1029 16 22 987 NOR2_X1
* cell instance $68156 m0 *1 315.78,379.4
X$68156 1139 1037 16 22 1105 NOR2_X1
* cell instance $68159 r0 *1 310.65,379.4
X$68159 894 16 22 1394 INV_X2
* cell instance $68160 r0 *1 311.22,379.4
X$68160 1121 16 22 894 CLKBUF_X3
* cell instance $68161 r0 *1 312.17,379.4
X$68161 1098 1190 1140 1034 1122 1192 16 22 990 OAI33_X1
* cell instance $68162 r0 *1 313.5,379.4
X$68162 1151 1037 16 22 1190 NOR2_X1
* cell instance $68165 m0 *1 316.73,379.4
X$68165 1106 1029 16 22 1104 NOR2_X1
* cell instance $68169 r0 *1 320.34,379.4
X$68169 1098 1198 1199 1034 1200 1197 16 22 1138 OAI33_X1
* cell instance $68172 r0 *1 322.62,379.4
X$68172 1117 16 22 1065 CLKBUF_X3
* cell instance $68173 r0 *1 323.57,379.4
X$68173 1117 16 22 1037 CLKBUF_X3
* cell instance $68174 m0 *1 325.47,379.4
X$68174 993 1069 16 22 1123 NOR2_X1
* cell instance $68175 m0 *1 324.52,379.4
X$68175 1054 16 22 1069 CLKBUF_X3
* cell instance $68179 r0 *1 324.9,379.4
X$68179 1245 1117 16 22 1202 NOR2_X1
* cell instance $68181 r0 *1 325.66,379.4
X$68181 1202 1136 1034 1123 1154 1098 16 22 1053 OAI33_X1
* cell instance $68185 m0 *1 327.94,379.4
X$68185 1110 1065 16 22 1109 NOR2_X1
* cell instance $68186 r0 *1 328.13,379.4
X$68186 1203 1054 16 22 1136 NOR2_X1
* cell instance $68187 r0 *1 328.7,379.4
X$68187 1038 1124 16 22 1034 NAND2_X2
* cell instance $68188 m0 *1 329.08,379.4
X$68188 1075 1072 16 981 22 NAND2_X4
* cell instance $68194 m0 *1 342.19,379.4
X$68194 1132 1073 743 16 482 22 AOI21_X1
* cell instance $68197 r0 *1 329.65,379.4
X$68197 1075 1124 16 22 1098 NAND2_X2
* cell instance $68201 r0 *1 331.93,379.4
X$68201 1204 1073 946 22 16 1141 OAI21_X4
* cell instance $68204 r0 *1 338.96,379.4
X$68204 1072 947 1069 770 16 22 1206 NAND4_X1
* cell instance $68205 r0 *1 339.91,379.4
X$68205 1206 1073 743 16 1126 22 AOI21_X1
* cell instance $68207 r0 *1 342.19,379.4
X$68207 1074 1038 1072 770 16 22 1132 NAND4_X1
* cell instance $68208 r0 *1 343.14,379.4
X$68208 1074 770 16 22 1205 NAND2_X1
* cell instance $68209 r0 *1 343.71,379.4
X$68209 1072 16 22 1124 INV_X1
* cell instance $68210 r0 *1 344.09,379.4
X$68210 109 1124 16 22 1156 NOR2_X1
* cell instance $68211 m0 *1 344.28,379.4
X$68211 1038 16 22 1075 INV_X2
* cell instance $68215 m0 *1 347.13,379.4
X$68215 259 1038 16 22 1076 NOR2_X1
* cell instance $68216 m0 *1 347.7,379.4
X$68216 16 1020 1115 1077 1078 22 DFF_X1
* cell instance $68217 m0 *1 350.93,379.4
X$68217 1115 16 22 1038 CLKBUF_X3
* cell instance $68225 r0 *1 345.04,379.4
X$68225 259 1072 16 22 1196 NOR2_X1
* cell instance $68227 r0 *1 346.37,379.4
X$68227 109 1075 16 22 1157 NOR2_X1
* cell instance $68228 r0 *1 346.94,379.4
X$68228 1157 1126 1076 16 22 1077 MUX2_X1
* cell instance $68235 r0 *1 361.95,379.4
X$68235 749 16 22 1078 CLKBUF_X3
* cell instance $68236 r0 *1 362.9,379.4
X$68236 1078 16 22 1396 INV_X2
* cell instance $68241 r0 *1 376.58,379.4
X$68241 16 1566 1079 1130 1078 22 DFF_X1
* cell instance $68243 m0 *1 377.34,379.4
X$68243 876 637 1079 16 22 1130 MUX2_X1
* cell instance $68248 m0 *1 383.61,379.4
X$68248 1018 255 1188 16 22 660 MUX2_X1
* cell instance $68250 m0 *1 387.22,379.4
X$68250 16 1513 1113 1114 1041 22 DFF_X1
* cell instance $68251 m0 *1 390.45,379.4
X$68251 960 225 1080 16 22 1128 MUX2_X1
* cell instance $68252 m0 *1 391.78,379.4
X$68252 749 16 22 1041 CLKBUF_X3
* cell instance $68253 m0 *1 392.73,379.4
X$68253 1041 16 22 CLKBUF_X1
* cell instance $68257 m0 *1 402.61,379.4
X$68257 16 1439 1107 1081 1162 22 DFF_X1
* cell instance $68264 r0 *1 388.36,379.4
X$68264 16 1565 1080 1128 1041 22 DFF_X1
* cell instance $68269 m0 *1 408.5,379.4
X$68269 16 1441 1082 1083 1162 22 DFF_X1
* cell instance $68271 m0 *1 419.33,379.4
X$68271 16 1470 1045 1044 838 22 DFF_X1
* cell instance $68273 m0 *1 422.75,379.4
X$68273 879 225 1084 16 22 1127 MUX2_X1
* cell instance $68276 m0 *1 427.31,379.4
X$68276 960 637 1094 16 22 1166 MUX2_X1
* cell instance $68285 r0 *1 420.28,379.4
X$68285 16 1596 1084 1127 1002 22 DFF_X1
* cell instance $68287 r0 *1 429.59,379.4
X$68287 749 16 22 1002 CLKBUF_X3
* cell instance $68288 r0 *1 430.54,379.4
X$68288 1002 16 22 CLKBUF_X1
* cell instance $68290 m0 *1 431.49,379.4
X$68290 16 1465 1090 1091 1002 22 DFF_X1
* cell instance $68296 m0 *1 437.57,379.4
X$68296 1085 16 22 939 BUF_X2
* cell instance $68538 m0 *1 269.61,393.4
X$68538 1292 1141 1304 16 22 1271 MUX2_X1
* cell instance $68547 r0 *1 269.42,393.4
X$68547 1292 976 1303 16 22 1302 MUX2_X1
* cell instance $68548 r0 *1 270.75,393.4
X$68548 16 1545 1303 1302 1258 22 DFF_X1
* cell instance $68549 m0 *1 272.27,393.4
X$68549 1304 906 1303 16 22 1131 MUX2_X1
* cell instance $68555 r0 *1 276.26,393.4
X$68555 16 1547 1305 1306 1258 22 DFF_X1
* cell instance $68556 m0 *1 277.21,393.4
X$68556 1292 1242 1305 16 22 1306 MUX2_X1
* cell instance $68559 m0 *1 279.11,393.4
X$68559 1305 930 1316 16 22 1286 MUX2_X1
* cell instance $68565 m0 *1 281.58,393.4
X$68565 1121 16 22 1258 CLKBUF_X3
* cell instance $68567 m0 *1 286.33,393.4
X$68567 16 1431 1273 1308 1258 22 DFF_X1
* cell instance $68578 r0 *1 296.78,393.4
X$68578 16 1653 1294 1310 1258 22 DFF_X1
* cell instance $68579 r0 *1 300.01,393.4
X$68579 572 1252 1294 16 22 1310 MUX2_X1
* cell instance $68580 r0 *1 301.34,393.4
X$68580 1296 1219 1294 16 22 1182 MUX2_X1
* cell instance $68582 m0 *1 303.81,393.4
X$68582 1319 1219 1289 16 22 1185 MUX2_X1
* cell instance $68587 m0 *1 307.61,393.4
X$68587 16 1479 1276 1311 1275 22 DFF_X1
* cell instance $68589 m0 *1 313.88,393.4
X$68589 649 1214 1278 16 22 1312 MUX2_X1
* cell instance $68590 m0 *1 315.21,393.4
X$68590 1337 947 1278 16 22 1277 MUX2_X1
* cell instance $68593 m0 *1 318.82,393.4
X$68593 385 1252 1279 16 22 1287 MUX2_X1
* cell instance $68594 m0 *1 320.15,393.4
X$68594 1326 1219 1279 16 22 1285 MUX2_X1
* cell instance $68598 m0 *1 325.47,393.4
X$68598 1307 930 1283 16 22 1245 MUX2_X1
* cell instance $68605 r0 *1 308.37,393.4
X$68605 649 1252 1276 16 22 1311 MUX2_X1
* cell instance $68608 r0 *1 310.27,393.4
X$68608 1339 1219 1276 16 22 1253 MUX2_X1
* cell instance $68612 r0 *1 314.26,393.4
X$68612 16 1582 1278 1312 1325 22 DFF_X1
* cell instance $68615 r0 *1 319.39,393.4
X$68615 930 22 1219 16 BUF_X4
* cell instance $68619 r0 *1 324.9,393.4
X$68619 16 1578 1307 1309 1299 22 DFF_X1
* cell instance $68620 r0 *1 328.13,393.4
X$68620 1280 1027 1307 16 22 1309 MUX2_X1
* cell instance $68622 m0 *1 331.93,393.4
X$68622 1300 947 1281 16 22 1110 MUX2_X1
* cell instance $68948 m0 *1 264.67,399
X$68948 1313 16 22 1334 CLKBUF_X2
* cell instance $68954 m0 *1 269.8,399
X$68954 1334 1141 1346 16 22 1315 MUX2_X1
* cell instance $68959 r0 *1 270.18,399
X$68959 1334 976 1347 16 22 1345 MUX2_X1
* cell instance $68960 r0 *1 271.51,399
X$68960 16 1628 1347 1345 1318 22 DFF_X1
* cell instance $68962 m0 *1 273.79,399
X$68962 1346 906 1347 16 22 1089 MUX2_X1
* cell instance $68966 m0 *1 277.02,399
X$68966 16 1509 1316 1332 1318 22 DFF_X1
* cell instance $68968 m0 *1 281.96,399
X$68968 16 1525 1319 1317 1318 22 DFF_X1
* cell instance $68970 m0 *1 285.95,399
X$68970 16 1414 1321 1320 1318 22 DFF_X1
* cell instance $68974 m0 *1 296.97,399
X$68974 1351 16 22 572 BUF_X2
* cell instance $68984 r0 *1 299.06,399
X$68984 16 1630 1296 1350 1275 22 DFF_X1
* cell instance $68985 m0 *1 300.58,399
X$68985 1351 1027 1296 16 22 1350 MUX2_X1
* cell instance $68989 m0 *1 303.62,399
X$68989 1322 947 1323 16 22 1118 MUX2_X1
* cell instance $68990 m0 *1 304.95,399
X$68990 16 1503 1323 1324 1275 22 DFF_X1
* cell instance $68992 m0 *1 308.94,399
X$68992 16 1483 1339 1340 1275 22 DFF_X1
* cell instance $68995 m0 *1 313.12,399
X$68995 16 1512 1337 1338 1325 22 DFF_X1
* cell instance $68999 r0 *1 303.81,399
X$68999 1121 16 22 1275 CLKBUF_X3
* cell instance $69000 r0 *1 304.76,399
X$69000 1275 16 22 1688 INV_X1
* cell instance $69005 m0 *1 317.49,399
X$69005 16 1505 1326 1333 1325 22 DFF_X1
* cell instance $69008 m0 *1 323.19,399
X$69008 1343 947 1330 16 22 1327 MUX2_X1
* cell instance $69009 m0 *1 324.52,399
X$69009 930 22 947 16 BUF_X4
* cell instance $69012 m0 *1 327.56,399
X$69012 1328 947 1329 16 22 1155 MUX2_X1
* cell instance $69015 r0 *1 320.34,399
X$69015 1121 16 22 1325 CLKBUF_X3
* cell instance $69016 r0 *1 321.29,399
X$69016 1325 16 22 CLKBUF_X1
* cell instance $69019 r0 *1 329.46,399
X$69019 16 1627 1329 1344 1325 22 DFF_X1
* cell instance $69020 m0 *1 330.22,399
X$69020 1280 976 1329 16 22 1344 MUX2_X1
* cell instance $69292 m0 *1 271.7,390.6
X$69292 16 1491 1246 1266 1258 22 DFF_X1
* cell instance $69301 r0 *1 268.85,390.6
X$69301 16 1556 1304 1271 1258 22 DFF_X1
* cell instance $69304 m0 *1 276.83,390.6
X$69304 16 1511 1259 1267 1258 22 DFF_X1
* cell instance $69308 m0 *1 293.93,390.6
X$69308 16 1493 1260 1269 1239 22 DFF_X1
* cell instance $69313 r0 *1 280.63,390.6
X$69313 1292 16 22 813 BUF_X2
* cell instance $69316 r0 *1 282.34,390.6
X$69316 1292 1027 1272 16 22 1288 MUX2_X1
* cell instance $69322 r0 *1 284.24,390.6
X$69322 16 1542 1272 1288 1258 22 DFF_X1
* cell instance $69323 r0 *1 287.47,390.6
X$69323 813 1252 1273 16 22 1308 MUX2_X1
* cell instance $69324 r0 *1 288.8,390.6
X$69324 1272 1219 1273 16 22 1183 MUX2_X1
* cell instance $69326 r0 *1 296.21,390.6
X$69326 16 1656 1290 1291 1239 22 DFF_X1
* cell instance $69327 m0 *1 297.73,390.6
X$69327 1290 871 572 16 22 1291 MUX2_X1
* cell instance $69331 m0 *1 302.86,390.6
X$69331 813 1214 1289 16 22 1274 MUX2_X1
* cell instance $69337 m0 *1 324.71,390.6
X$69337 619 1252 1283 16 22 1284 MUX2_X1
* cell instance $69343 r0 *1 302.29,390.6
X$69343 16 1654 1289 1274 1239 22 DFF_X1
* cell instance $69349 r0 *1 316.73,390.6
X$69349 16 1581 1279 1287 1249 22 DFF_X1
* cell instance $69353 r0 *1 323.95,390.6
X$69353 16 1580 1283 1284 1249 22 DFF_X1
* cell instance $69355 m0 *1 326.42,390.6
X$69355 1280 1112 1263 16 22 1268 MUX2_X1
* cell instance $69356 m0 *1 327.94,390.6
X$69356 1280 16 22 619 BUF_X2
* cell instance $69386 r0 *1 330.79,390.6
X$69386 1280 1228 1281 16 22 1282 MUX2_X1
* cell instance $69387 r0 *1 332.12,390.6
X$69387 16 1617 1281 1282 1299 22 DFF_X1
* cell instance $69618 m0 *1 269.61,382.2
X$69618 16 1436 1129 1167 864 22 DFF_X1
* cell instance $69622 m0 *1 275.31,382.2
X$69622 1057 1242 1116 16 22 1169 MUX2_X1
* cell instance $69634 r0 *1 275.69,382.2
X$69634 16 1541 1142 1227 864 22 DFF_X1
* cell instance $69637 m0 *1 284.62,382.2
X$69637 1057 1027 1143 16 22 1173 MUX2_X1
* cell instance $69638 m0 *1 286.14,382.2
X$69638 16 1486 1143 1173 1211 22 DFF_X1
* cell instance $69645 r0 *1 290.13,382.2
X$69645 16 1648 1144 1174 1211 22 DFF_X1
* cell instance $69647 m0 *1 290.51,382.2
X$69647 740 1252 1144 16 22 1174 MUX2_X1
* cell instance $69648 m0 *1 292.6,382.2
X$69648 1143 1219 1144 16 22 1134 MUX2_X1
* cell instance $69651 m0 *1 294.5,382.2
X$69651 16 1490 1063 1145 1239 22 DFF_X1
* cell instance $69655 m0 *1 300.96,382.2
X$69655 1177 1065 16 22 1181 NOR2_X1
* cell instance $69659 m0 *1 301.91,382.2
X$69659 1216 1037 16 22 1146 NOR2_X1
* cell instance $69661 m0 *1 302.86,382.2
X$69661 1261 1069 16 22 1147 NOR2_X1
* cell instance $69663 m0 *1 303.81,382.2
X$69663 1182 1065 16 22 1184 NOR2_X1
* cell instance $69668 m0 *1 307.04,382.2
X$69668 1185 1069 16 22 1148 NOR2_X1
* cell instance $69671 m0 *1 310.08,382.2
X$69671 16 1523 1150 1189 894 22 DFF_X1
* cell instance $69672 m0 *1 309.51,382.2
X$69672 1149 1037 16 22 1186 NOR2_X1
* cell instance $69673 m0 *1 313.31,382.2
X$69673 786 16 22 1121 CLKBUF_X3
* cell instance $69674 m0 *1 314.26,382.2
X$69674 1253 1065 16 22 1192 NOR2_X1
* cell instance $69678 r0 *1 311.22,382.2
X$69678 1150 855 649 16 22 1189 MUX2_X1
* cell instance $69679 r0 *1 312.55,382.2
X$69679 1150 653 1218 16 22 1151 MUX2_X1
* cell instance $69681 m0 *1 315.4,382.2
X$69681 1277 1069 16 22 1122 NOR2_X1
* cell instance $69686 r0 *1 316.16,382.2
X$69686 16 1584 1152 1233 894 22 DFF_X1
* cell instance $69688 m0 *1 317.11,382.2
X$69688 1152 855 385 16 22 1233 MUX2_X1
* cell instance $69689 m0 *1 320.15,382.2
X$69689 1194 1037 16 22 1198 NOR2_X1
* cell instance $69690 m0 *1 318.82,382.2
X$69690 1152 653 1247 16 22 1194 MUX2_X1
* cell instance $69693 m0 *1 321.29,382.2
X$69693 1285 1065 16 22 1197 NOR2_X1
* cell instance $69697 m0 *1 322.24,382.2
X$69697 1327 1069 16 22 1200 NOR2_X1
* cell instance $69698 m0 *1 325.85,382.2
X$69698 1153 1065 16 22 1154 NOR2_X1
* cell instance $69701 m0 *1 328.13,382.2
X$69701 1155 1069 16 22 1071 NOR2_X1
* cell instance $69704 m0 *1 331.93,382.2
X$69704 911 1073 946 22 16 1242 OAI21_X4
* cell instance $69705 m0 *1 334.4,382.2
X$69705 953 1073 946 22 16 1214 OAI21_X4
* cell instance $69708 m0 *1 343.14,382.2
X$69708 1205 1073 743 16 1201 22 AOI21_X1
* cell instance $69710 m0 *1 344.66,382.2
X$69710 1156 1201 1196 16 22 1195 MUX2_X1
* cell instance $69711 m0 *1 345.99,382.2
X$69711 16 957 1193 1195 1078 22 DFF_X1
* cell instance $69712 m0 *1 349.22,382.2
X$69712 1193 16 22 1072 CLKBUF_X3
* cell instance $69721 m0 *1 383.04,382.2
X$69721 876 253 1188 16 22 1191 MUX2_X1
* cell instance $69729 r0 *1 332.31,382.2
X$69729 1232 1073 946 22 16 1252 OAI21_X4
* cell instance $69730 r0 *1 334.78,382.2
X$69730 16 991 22 946 BUF_X8
* cell instance $69732 r0 *1 338.77,382.2
X$69732 1125 1073 946 22 16 1228 OAI21_X4
* cell instance $69735 r0 *1 343.52,382.2
X$69735 16 343 22 1073 BUF_X8
* cell instance $69748 r0 *1 381.71,382.2
X$69748 16 1563 1188 1191 1078 22 DFF_X1
* cell instance $69751 r0 *1 385.89,382.2
X$69751 16 1564 1158 1187 1041 22 DFF_X1
* cell instance $69752 r0 *1 389.12,382.2
X$69752 960 254 1158 16 22 1187 MUX2_X1
* cell instance $69755 r0 *1 392.16,382.2
X$69755 1158 266 1159 16 22 545 MUX2_X1
* cell instance $69896 m0 *1 287.85,407.4
X$69896 16 1504 1366 1373 1361 22 DFF_X1
* cell instance $69900 m0 *1 293.55,407.4
X$69900 16 1429 1367 1368 1361 22 DFF_X1
* cell instance $69917 m0 *1 299.63,407.4
X$69917 1121 16 22 1361 CLKBUF_X3
* cell instance $69919 m0 *1 300.58,407.4
X$69919 1361 16 22 CLKBUF_X1
* cell instance $69922 m0 *1 302.1,407.4
X$69922 1381 16 22 1351 CLKBUF_X2
* cell instance $69929 m0 *1 305.52,407.4
X$69929 16 1405 1382 1380 1361 22 DFF_X1
* cell instance $69930 m0 *1 314.83,407.4
X$69930 1335 1228 1379 16 22 1386 MUX2_X1
* cell instance $69931 m0 *1 316.16,407.4
X$69931 16 1478 1379 1386 1299 22 DFF_X1
* cell instance $69937 m0 *1 342.19,407.4
X$69937 1369 16 22 745 BUF_X2
* cell instance $69963 r0 *1 305.9,407.4
X$69963 1298 1242 1382 16 22 1380 MUX2_X1
* cell instance $69966 r0 *1 308.37,407.4
X$69966 1382 930 1377 16 22 1241 MUX2_X1
* cell instance $69971 r0 *1 314.07,407.4
X$69971 1335 1242 1378 16 22 1385 MUX2_X1
* cell instance $69974 r0 *1 315.97,407.4
X$69974 1378 930 1379 16 22 1139 MUX2_X1
* cell instance $70208 m0 *1 270.94,368.2
X$70208 16 1448 814 843 663 22 DFF_X1
* cell instance $70210 m0 *1 275.69,368.2
X$70210 761 666 814 16 22 928 MUX2_X1
* cell instance $70218 r0 *1 273.22,368.2
X$70218 883 664 813 16 22 885 MUX2_X1
* cell instance $70221 r0 *1 277.97,368.2
X$70221 865 570 813 16 22 887 MUX2_X1
* cell instance $70222 m0 *1 279.11,368.2
X$70222 16 1445 845 847 663 22 DFF_X1
* cell instance $70226 m0 *1 282.91,368.2
X$70226 16 1447 815 774 663 22 DFF_X1
* cell instance $70232 r0 *1 288.42,368.2
X$70232 16 1646 816 849 889 22 DFF_X1
* cell instance $70234 m0 *1 291.08,368.2
X$70234 763 666 816 16 22 933 MUX2_X1
* cell instance $70239 m0 *1 309.32,368.2
X$70239 742 666 776 16 22 777 MUX2_X1
* cell instance $70242 r0 *1 291.65,368.2
X$70242 816 664 572 16 22 849 MUX2_X1
* cell instance $70244 r0 *1 293.17,368.2
X$70244 16 1599 817 848 889 22 DFF_X1
* cell instance $70245 r0 *1 296.4,368.2
X$70245 817 855 740 16 22 848 MUX2_X1
* cell instance $70246 r0 *1 297.73,368.2
X$70246 817 653 818 16 22 819 MUX2_X1
* cell instance $70252 r0 *1 304.95,368.2
X$70252 895 466 813 16 22 893 MUX2_X1
* cell instance $70255 m0 *1 315.4,368.2
X$70255 16 1443 779 853 709 22 DFF_X1
* cell instance $70256 m0 *1 314.07,368.2
X$70256 766 666 779 16 22 778 MUX2_X1
* cell instance $70261 m0 *1 324.52,368.2
X$70261 821 611 619 16 22 809 MUX2_X1
* cell instance $70262 m0 *1 321.29,368.2
X$70262 16 1440 821 809 709 22 DFF_X1
* cell instance $70269 r0 *1 324.14,368.2
X$70269 821 906 696 16 22 822 MUX2_X1
* cell instance $70273 m0 *1 332.5,368.2
X$70273 823 812 782 16 22 811 NAND3_X2
* cell instance $70274 m0 *1 330.03,368.2
X$70274 16 466 811 780 743 22 AOI21_X4
* cell instance $70276 r0 *1 330.22,368.2
X$70276 16 855 856 737 743 22 AOI21_X4
* cell instance $70277 r0 *1 332.69,368.2
X$70277 823 700 782 16 22 856 NAND3_X1
* cell instance $70280 r0 *1 334.02,368.2
X$70280 824 16 22 901 BUF_X1
* cell instance $70281 m0 *1 334.4,368.2
X$70281 823 739 782 16 22 857 NAND3_X1
* cell instance $70283 m0 *1 335.16,368.2
X$70283 824 16 22 737 INV_X8
* cell instance $70287 r0 *1 334.59,368.2
X$70287 16 871 857 780 710 22 AOI21_X4
* cell instance $70288 r0 *1 337.06,368.2
X$70288 824 16 22 995 BUF_X1
* cell instance $70291 r0 *1 338.58,368.2
X$70291 812 16 22 872 INV_X1
* cell instance $70294 m0 *1 344.09,368.2
X$70294 783 16 22 782 INV_X4
* cell instance $70296 m0 *1 349.6,368.2
X$70296 783 957 826 22 16 860 HA_X1
* cell instance $70298 m0 *1 353.02,368.2
X$70298 784 829 860 826 861 835 22 16 AOI221_X2
* cell instance $70302 m0 *1 359.1,368.2
X$70302 832 863 835 22 16 710 MUX2_X2
* cell instance $70303 m0 *1 360.81,368.2
X$70303 835 830 22 804 16 XOR2_X2
* cell instance $70304 m0 *1 362.52,368.2
X$70304 16 836 758 737 787 841 22 NOR4_X4
* cell instance $70310 r0 *1 345.42,368.2
X$70310 825 905 22 824 16 XOR2_X2
* cell instance $70312 r0 *1 347.32,368.2
X$70312 607 915 831 22 16 859 HA_X1
* cell instance $70316 r0 *1 351.69,368.2
X$70316 859 16 22 829 INV_X1
* cell instance $70318 r0 *1 352.26,368.2
X$70318 830 826 22 16 827 AND2_X1
* cell instance $70319 r0 *1 353.02,368.2
X$70319 16 623 828 874 785 829 22 FA_X1
* cell instance $70320 r0 *1 356.06,368.2
X$70320 162 16 22 786 CLKBUF_X3
* cell instance $70323 r0 *1 358.72,368.2
X$70323 830 831 833 834 22 16 832 AND4_X1
* cell instance $70325 r0 *1 360.24,368.2
X$70325 862 16 22 833 INV_X1
* cell instance $70328 r0 *1 361.19,368.2
X$70328 836 862 842 830 16 22 863 NOR4_X1
* cell instance $70330 r0 *1 362.9,368.2
X$70330 831 16 22 842 INV_X4
* cell instance $70332 r0 *1 364.23,368.2
X$70332 862 831 22 787 16 XOR2_X2
* cell instance $70334 r0 *1 366.13,368.2
X$70334 836 16 22 839 BUF_X1
* cell instance $70335 r0 *1 366.7,368.2
X$70335 836 862 16 22 788 NAND2_X1
* cell instance $70340 r0 *1 375.44,368.2
X$70340 876 225 858 16 22 899 MUX2_X1
* cell instance $70343 r0 *1 377.34,368.2
X$70343 195 332 877 16 22 898 MUX2_X1
* cell instance $70346 r0 *1 379.81,368.2
X$70346 876 16 22 195 BUF_X2
* cell instance $70348 m0 *1 380,368.2
X$70348 789 227 195 16 22 790 MUX2_X1
* cell instance $70354 r0 *1 387.79,368.2
X$70354 16 1569 837 854 875 22 DFF_X1
* cell instance $70356 m0 *1 388.55,368.2
X$70356 83 332 837 16 22 854 MUX2_X1
* cell instance $70358 r0 *1 391.02,368.2
X$70358 917 520 837 16 22 717 MUX2_X1
* cell instance $70362 r0 *1 395.01,368.2
X$70362 719 227 168 16 22 896 MUX2_X1
* cell instance $70364 m0 *1 396.53,368.2
X$70364 749 16 22 1694 CLKBUF_X3
* cell instance $70366 m0 *1 397.48,368.2
X$70366 168 332 851 16 22 852 MUX2_X1
* cell instance $70367 m0 *1 398.81,368.2
X$70367 786 16 22 749 CLKBUF_X3
* cell instance $70369 m0 *1 399.95,368.2
X$70369 16 1500 799 800 510 22 DFF_X1
* cell instance $70373 m0 *1 413.06,368.2
X$70373 548 254 791 16 22 850 MUX2_X1
* cell instance $70375 m0 *1 415.15,368.2
X$70375 791 308 792 16 22 584 MUX2_X1
* cell instance $70378 r0 *1 396.91,368.2
X$70378 16 1583 851 852 875 22 DFF_X1
* cell instance $70383 r0 *1 408.31,368.2
X$70383 748 227 183 16 22 890 MUX2_X1
* cell instance $70388 r0 *1 412.49,368.2
X$70388 16 1586 791 850 838 22 DFF_X1
* cell instance $70390 m0 *1 418.19,368.2
X$70390 16 1515 792 846 510 22 DFF_X1
* cell instance $70391 m0 *1 416.86,368.2
X$70391 548 253 792 16 22 846 MUX2_X1
* cell instance $70392 m0 *1 421.42,368.2
X$70392 16 1487 752 793 586 22 DFF_X1
* cell instance $70397 m0 *1 430.16,368.2
X$70397 753 228 754 16 22 844 MUX2_X1
* cell instance $70448 m0 *1 707.18,368.2
X$70448 841 16 22 794 BUF_X1
* cell instance $70454 r0 *1 429.59,368.2
X$70454 16 1612 754 844 923 22 DFF_X1
* cell instance $70458 r0 *1 439.85,368.2
X$70458 840 16 22 753 CLKBUF_X2
* cell instance $70507 m0 *1 709.65,368.2
X$70507 839 16 22 796 BUF_X1
* cell instance $70647 m0 *1 271.13,373.8
X$70647 16 1437 927 926 864 22 DFF_X1
* cell instance $70650 m0 *1 280.63,373.8
X$70650 866 949 16 22 967 NOR2_X1
* cell instance $70662 r0 *1 278.92,373.8
X$70662 928 948 16 22 978 NOR2_X1
* cell instance $70663 r0 *1 279.49,373.8
X$70663 886 948 16 22 979 NOR2_X1
* cell instance $70664 r0 *1 280.06,373.8
X$70664 929 948 16 22 980 NOR2_X1
* cell instance $70665 r0 *1 280.63,373.8
X$70665 706 949 16 22 1009 NOR2_X1
* cell instance $70669 r0 *1 282.53,373.8
X$70669 950 949 16 22 1008 NOR2_X1
* cell instance $70671 r0 *1 283.48,373.8
X$70671 762 948 16 22 982 NOR2_X1
* cell instance $70674 m0 *1 284.62,373.8
X$70674 433 949 16 22 951 NOR2_X1
* cell instance $70678 m0 *1 296.02,373.8
X$70678 908 906 952 16 22 969 MUX2_X1
* cell instance $70682 m0 *1 311.03,373.8
X$70682 692 949 16 22 988 NOR2_X1
* cell instance $70691 r0 *1 286.14,373.8
X$70691 1054 16 22 948 CLKBUF_X3
* cell instance $70695 r0 *1 290.7,373.8
X$70695 614 949 16 22 983 NOR2_X1
* cell instance $70696 r0 *1 291.27,373.8
X$70696 933 948 16 22 1011 NOR2_X1
* cell instance $70699 r0 *1 293.74,373.8
X$70699 16 1600 952 1012 889 22 DFF_X1
* cell instance $70700 r0 *1 296.97,373.8
X$70700 952 871 460 16 22 1012 MUX2_X1
* cell instance $70703 r0 *1 298.87,373.8
X$70703 819 949 16 22 985 NOR2_X1
* cell instance $70706 r0 *1 300.01,373.8
X$70706 820 948 16 22 1033 NOR2_X1
* cell instance $70707 r0 *1 300.58,373.8
X$70707 969 949 16 22 986 NOR2_X1
* cell instance $70708 r0 *1 301.15,373.8
X$70708 690 948 16 22 1100 NOR2_X1
* cell instance $70713 r0 *1 315.02,373.8
X$70713 778 948 16 22 1022 NOR2_X1
* cell instance $70716 r0 *1 316.54,373.8
X$70716 471 949 16 22 1036 NOR2_X1
* cell instance $70718 r0 *1 323.19,373.8
X$70718 992 464 619 16 22 1025 MUX2_X1
* cell instance $70721 r0 *1 326.23,373.8
X$70721 822 1054 16 22 1108 NOR2_X1
* cell instance $70723 m0 *1 329.65,373.8
X$70723 16 464 945 737 743 22 AOI21_X4
* cell instance $70725 m0 *1 332.12,373.8
X$70725 782 700 698 22 16 1028 AND3_X1
* cell instance $70726 m0 *1 333.07,373.8
X$70726 782 711 698 22 16 1111 AND3_X1
* cell instance $70730 r0 *1 331.55,373.8
X$70730 669 711 823 22 16 1204 AND3_X1
* cell instance $70734 m0 *1 334.4,373.8
X$70734 912 781 823 16 22 NOR2_X4
* cell instance $70737 r0 *1 335.16,373.8
X$70737 1026 975 669 22 1232 16 NOR3_X2
* cell instance $70738 r0 *1 336.49,373.8
X$70738 1026 872 669 22 953 16 NOR3_X2
* cell instance $70739 m0 *1 337.82,373.8
X$70739 16 781 912 782 975 1125 22 NOR4_X4
* cell instance $70740 m0 *1 337.25,373.8
X$70740 912 745 16 22 1026 NAND2_X1
* cell instance $70744 r0 *1 340.1,373.8
X$70744 915 16 22 1054 CLKBUF_X3
* cell instance $70745 r0 *1 341.05,373.8
X$70745 946 780 770 22 954 16 OAI21_X1
* cell instance $70747 m0 *1 341.62,373.8
X$70747 16 955 870 1023 915 22 DFF_X2
* cell instance $70750 m0 *1 347.7,373.8
X$70750 912 257 22 16 1021 AND2_X1
* cell instance $70751 m0 *1 348.46,373.8
X$70751 259 912 16 22 956 NOR2_X1
* cell instance $70752 m0 *1 349.03,373.8
X$70752 972 22 912 16 BUF_X4
* cell instance $70757 r0 *1 342.95,373.8
X$70757 1023 257 22 16 1024 AND2_X1
* cell instance $70762 r0 *1 348.08,373.8
X$70762 1021 807 956 16 22 996 MUX2_X1
* cell instance $70764 m0 *1 351.69,373.8
X$70764 972 1020 973 22 16 944 HA_X1
* cell instance $70770 m0 *1 359.1,373.8
X$70770 16 946 22 958 BUF_X8
* cell instance $70786 r0 *1 378.29,373.8
X$70786 876 514 959 16 22 1019 MUX2_X1
* cell instance $70788 m0 *1 381.14,373.8
X$70788 16 1418 916 941 875 22 DFF_X1
* cell instance $70793 m0 *1 389.69,373.8
X$70793 960 228 917 16 22 940 MUX2_X1
* cell instance $70802 r0 *1 391.59,373.8
X$70802 16 1588 997 971 1041 22 DFF_X1
* cell instance $70803 m0 *1 393.87,373.8
X$70803 168 304 997 16 22 971 MUX2_X1
* cell instance $70806 m0 *1 395.96,373.8
X$70806 939 16 22 168 BUF_X2
* cell instance $70807 m0 *1 396.72,373.8
X$70807 16 1473 918 937 1041 22 DFF_X1
* cell instance $70812 m0 *1 402.04,373.8
X$70812 16 1494 919 936 838 22 DFF_X1
* cell instance $70816 m0 *1 406.6,373.8
X$70816 999 228 961 16 22 970 MUX2_X1
* cell instance $70818 m0 *1 407.93,373.8
X$70818 16 1495 961 970 838 22 DFF_X1
* cell instance $70822 m0 *1 412.87,373.8
X$70822 753 253 963 16 22 968 MUX2_X1
* cell instance $70823 m0 *1 411.54,373.8
X$70823 962 266 963 16 22 750 MUX2_X1
* cell instance $70829 r0 *1 412.68,373.8
X$70829 16 1587 963 968 923 22 DFF_X1
* cell instance $70832 m0 *1 418.38,373.8
X$70832 16 1514 920 934 923 22 DFF_X1
* cell instance $70834 m0 *1 423.89,373.8
X$70834 16 1421 921 922 923 22 DFF_X1
* cell instance $70841 r0 *1 426.36,373.8
X$70841 960 514 1001 16 22 1000 MUX2_X1
* cell instance $70842 r0 *1 427.69,373.8
X$70842 1001 286 1094 16 22 555 MUX2_X1
* cell instance $70843 m0 *1 429.97,373.8
X$70843 923 16 22 CLKBUF_X1
* cell instance $70844 m0 *1 429.02,373.8
X$70844 749 16 22 923 CLKBUF_X3
* cell instance $70846 m0 *1 430.73,373.8
X$70846 16 1420 964 966 923 22 DFF_X1
* cell instance $70900 r0 *1 431.49,373.8
X$70900 939 514 964 16 22 966 MUX2_X1
* cell instance $70901 r0 *1 432.82,373.8
X$70901 964 286 1090 16 22 645 MUX2_X1
* cell instance $70905 r0 *1 436.62,373.8
X$70905 999 514 1003 16 22 1047 MUX2_X1
* cell instance $70906 r0 *1 437.95,373.8
X$70906 1003 286 965 16 22 547 MUX2_X1
* cell instance $70907 r0 *1 439.28,373.8
X$70907 999 637 965 16 22 1005 MUX2_X1
* cell instance $70911 r0 *1 447.64,373.8
X$70911 1004 16 22 879 CLKBUF_X2
* cell instance $71096 m0 *1 270.37,371
X$71096 16 1438 883 885 864 22 DFF_X1
* cell instance $71108 r0 *1 272.65,371
X$71108 927 611 813 16 22 926 MUX2_X1
* cell instance $71109 r0 *1 273.98,371
X$71109 927 666 883 16 22 929 MUX2_X1
* cell instance $71111 m0 *1 276.45,371
X$71111 16 1446 865 887 889 22 DFF_X1
* cell instance $71113 m0 *1 279.68,371
X$71113 865 906 845 16 22 866 MUX2_X1
* cell instance $71118 r0 *1 280.25,371
X$71118 930 22 666 16 BUF_X4
* cell instance $71120 r0 *1 281.77,371
X$71120 907 430 815 16 22 950 MUX2_X1
* cell instance $71121 m0 *1 282.34,371
X$71121 907 570 740 16 22 867 MUX2_X1
* cell instance $71127 r0 *1 283.1,371
X$71127 16 1592 907 867 889 22 DFF_X1
* cell instance $71131 r0 *1 291.08,371
X$71131 316 16 22 889 CLKBUF_X3
* cell instance $71132 r0 *1 292.03,371
X$71132 889 16 22 CLKBUF_X1
* cell instance $71134 r0 *1 292.79,371
X$71134 16 1601 908 932 889 22 DFF_X1
* cell instance $71135 r0 *1 296.02,371
X$71135 908 855 460 16 22 932 MUX2_X1
* cell instance $71137 m0 *1 299.06,371
X$71137 16 1468 818 892 889 22 DFF_X1
* cell instance $71138 m0 *1 297.73,371
X$71138 818 871 740 16 22 892 MUX2_X1
* cell instance $71141 m0 *1 304,371
X$71141 16 1464 895 893 894 22 DFF_X1
* cell instance $71145 m0 *1 309.7,371
X$71145 897 464 649 16 22 935 MUX2_X1
* cell instance $71151 r0 *1 304.76,371
X$71151 775 430 895 16 22 1102 MUX2_X1
* cell instance $71156 r0 *1 308.94,371
X$71156 16 1626 897 935 894 22 DFF_X1
* cell instance $71157 m0 *1 312.36,371
X$71157 897 430 909 16 22 868 MUX2_X1
* cell instance $71163 m0 *1 322.24,371
X$71163 16 1457 900 869 870 22 DFF_X1
* cell instance $71167 m0 *1 333.26,371
X$71167 316 16 22 870 CLKBUF_X3
* cell instance $71169 m0 *1 334.4,371
X$71169 901 16 22 780 INV_X4
* cell instance $71171 m0 *1 338.39,371
X$71171 745 16 22 781 INV_X4
* cell instance $71172 m0 *1 339.34,371
X$71172 947 150 22 16 903 AND2_X1
* cell instance $71177 r0 *1 313.31,371
X$71177 909 466 649 16 22 938 MUX2_X1
* cell instance $71178 r0 *1 314.64,371
X$71178 16 1574 909 938 870 22 DFF_X1
* cell instance $71179 r0 *1 317.87,371
X$71179 930 22 430 16 BUF_X4
* cell instance $71183 r0 *1 322.81,371
X$71183 900 466 619 16 22 869 MUX2_X1
* cell instance $71185 r0 *1 324.33,371
X$71185 910 22 906 16 BUF_X4
* cell instance $71186 r0 *1 325.66,371
X$71186 910 22 930 16 BUF_X4
* cell instance $71189 r0 *1 327.56,371
X$71189 910 22 653 16 BUF_X4
* cell instance $71193 r0 *1 330.22,371
X$71193 914 16 22 910 CLKBUF_X2
* cell instance $71195 r0 *1 331.74,371
X$71195 669 700 823 22 16 911 AND3_X1
* cell instance $71196 r0 *1 332.69,371
X$71196 823 711 782 16 22 945 NAND3_X2
* cell instance $71197 r0 *1 334.02,371
X$71197 870 16 22 1690 INV_X1
* cell instance $71199 r0 *1 334.78,371
X$71199 745 912 22 16 698 AND2_X2
* cell instance $71201 r0 *1 336.49,371
X$71201 16 781 912 782 872 913 22 NOR4_X4
* cell instance $71202 r0 *1 339.91,371
X$71202 739 16 22 975 INV_X1
* cell instance $71205 m0 *1 342,371
X$71205 902 954 903 16 22 904 MUX2_X1
* cell instance $71206 m0 *1 341.24,371
X$71206 873 257 22 16 902 AND2_X1
* cell instance $71207 m0 *1 343.33,371
X$71207 16 785 914 904 870 22 DFF_X1
* cell instance $71211 m0 *1 351.31,371
X$71211 860 830 944 827 828 905 22 16 AOI221_X2
* cell instance $71212 m0 *1 353.4,371
X$71212 828 826 16 22 834 XNOR2_X2
* cell instance $71215 m0 *1 359.1,371
X$71215 834 833 831 830 16 22 943 NAND4_X1
* cell instance $71217 m0 *1 360.81,371
X$71217 834 16 22 836 INV_X4
* cell instance $71218 m0 *1 361.76,371
X$71218 830 842 862 836 16 22 942 OR4_X1
* cell instance $71220 m0 *1 364.42,371
X$71220 874 16 22 862 CLKBUF_X2
* cell instance $71224 m0 *1 373.54,371
X$71224 16 1459 858 899 875 22 DFF_X1
* cell instance $71225 m0 *1 376.77,371
X$71225 16 1538 877 898 875 22 DFF_X1
* cell instance $71229 r0 *1 341.62,371
X$71229 915 914 873 22 16 1074 HA_X1
* cell instance $71234 r0 *1 351.69,371
X$71234 973 16 22 830 BUF_X2
* cell instance $71238 r0 *1 359.48,371
X$71238 943 835 942 16 22 958 MUX2_X1
* cell instance $71243 r0 *1 364.61,371
X$71243 874 16 22 924 BUF_X1
* cell instance $71250 r0 *1 383.04,371
X$71250 876 228 916 16 22 941 MUX2_X1
* cell instance $71251 m0 *1 383.61,371
X$71251 916 266 877 16 22 715 MUX2_X1
* cell instance $71253 m0 *1 384.94,371
X$71253 882 16 22 876 CLKBUF_X2
* cell instance $71259 r0 *1 385.7,371
X$71259 749 16 22 875 CLKBUF_X3
* cell instance $71262 r0 *1 388.93,371
X$71262 16 1568 917 940 875 22 DFF_X1
* cell instance $71263 m0 *1 392.35,371
X$71263 16 1507 719 896 875 22 DFF_X1
* cell instance $71272 r0 *1 397.67,371
X$71272 939 228 918 16 22 937 MUX2_X1
* cell instance $71274 m0 *1 398.24,371
X$71274 918 520 851 16 22 878 MUX2_X1
* cell instance $71277 m0 *1 407.36,371
X$71277 16 1499 748 890 838 22 DFF_X1
* cell instance $71286 r0 *1 402.8,371
X$71286 64 332 919 16 22 936 MUX2_X1
* cell instance $71287 r0 *1 404.13,371
X$71287 961 520 919 16 22 676 MUX2_X1
* cell instance $71293 r0 *1 418.95,371
X$71293 183 332 920 16 22 934 MUX2_X1
* cell instance $71294 r0 *1 420.28,371
X$71294 921 520 920 16 22 730 MUX2_X1
* cell instance $71298 r0 *1 423.7,371
X$71298 879 228 921 16 22 922 MUX2_X1
* cell instance $71304 r0 *1 435.48,371
X$71304 16 1561 888 925 923 22 DFF_X1
* cell instance $71305 m0 *1 436.24,371
X$71305 879 514 888 16 22 925 MUX2_X1
* cell instance $71308 m0 *1 438.14,371
X$71308 888 286 880 16 22 639 MUX2_X1
* cell instance $71312 m0 *1 441.18,371
X$71312 16 1415 880 884 923 22 DFF_X1
* cell instance $71313 m0 *1 439.85,371
X$71313 879 637 880 16 22 884 MUX2_X1
* cell instance $71361 m0 *1 704.14,371
X$71361 842 16 22 881 BUF_X1
* cell instance $71559 r0 *1 271.89,359.8
X$71559 16 1593 612 640 663 22 DFF_X1
* cell instance $71560 r0 *1 275.12,359.8
X$71560 612 611 460 16 22 640 MUX2_X1
* cell instance $71564 r0 *1 279.11,359.8
X$71564 16 1594 613 642 663 22 DFF_X1
* cell instance $71565 r0 *1 282.34,359.8
X$71565 613 611 432 16 22 642 MUX2_X1
* cell instance $71567 m0 *1 289.75,359.8
X$71567 571 570 572 16 22 591 MUX2_X1
* cell instance $71568 m0 *1 286.52,359.8
X$71568 16 1425 571 591 668 22 DFF_X1
* cell instance $71571 m0 *1 295.64,359.8
X$71571 615 464 460 16 22 594 MUX2_X1
* cell instance $71575 m0 *1 300.96,359.8
X$71575 646 466 572 16 22 616 MUX2_X1
* cell instance $71579 m0 *1 307.61,359.8
X$71579 617 570 649 16 22 648 MUX2_X1
* cell instance $71582 m0 *1 311.22,359.8
X$71582 652 340 649 16 22 650 MUX2_X1
* cell instance $71585 m0 *1 317.11,359.8
X$71585 16 1442 538 537 315 22 DFF_X1
* cell instance $71590 r0 *1 293.55,359.8
X$71590 16 1605 615 594 668 22 DFF_X1
* cell instance $71591 r0 *1 296.78,359.8
X$71591 615 666 535 16 22 690 MUX2_X1
* cell instance $71595 r0 *1 300.77,359.8
X$71595 16 1595 646 616 536 22 DFF_X1
* cell instance $71598 r0 *1 305.14,359.8
X$71598 316 16 22 536 CLKBUF_X3
* cell instance $71599 r0 *1 306.09,359.8
X$71599 16 1609 617 648 536 22 DFF_X1
* cell instance $71602 r0 *1 310.27,359.8
X$71602 617 430 652 16 22 692 MUX2_X1
* cell instance $71603 r0 *1 311.6,359.8
X$71603 16 1632 652 650 709 22 DFF_X1
* cell instance $71606 m0 *1 321.67,359.8
X$71606 16 1409 574 601 315 22 DFF_X1
* cell instance $71608 m0 *1 324.9,359.8
X$71608 574 570 619 16 22 601 MUX2_X1
* cell instance $71612 m0 *1 328.7,359.8
X$71612 575 340 619 16 22 602 MUX2_X1
* cell instance $71614 m0 *1 330.22,359.8
X$71614 16 1407 575 602 709 22 DFF_X1
* cell instance $71615 m0 *1 333.45,359.8
X$71615 654 576 573 16 22 604 NAND3_X1
* cell instance $71618 m0 *1 341.81,359.8
X$71618 441 577 621 16 22 560 MUX2_X1
* cell instance $71619 m0 *1 343.14,359.8
X$71619 607 150 22 16 621 AND2_X1
* cell instance $71626 r0 *1 325.28,359.8
X$71626 574 653 575 16 22 974 MUX2_X1
* cell instance $71631 r0 *1 338.01,359.8
X$71631 770 16 22 312 INV_X4
* cell instance $71633 r0 *1 342,359.8
X$71633 497 622 1681 22 16 700 HA_X1
* cell instance $71636 r0 *1 345.61,359.8
X$71636 607 622 609 22 16 711 HA_X1
* cell instance $71638 m0 *1 346.56,359.8
X$71638 609 150 22 16 656 AND2_X1
* cell instance $71643 m0 *1 361.95,359.8
X$71643 16 610 317 1666 21 22 DFF_X2
* cell instance $71644 m0 *1 365.56,359.8
X$71644 476 21 443 16 22 578 NAND3_X1
* cell instance $71645 m0 *1 366.32,359.8
X$71645 578 579 598 16 22 610 NAND3_X1
* cell instance $71648 m0 *1 368.03,359.8
X$71648 476 18 443 16 22 608 NAND3_X1
* cell instance $71650 r0 *1 347.51,359.8
X$71650 623 257 22 16 624 AND2_X1
* cell instance $71651 r0 *1 348.27,359.8
X$71651 624 577 656 16 22 657 MUX2_X1
* cell instance $71652 r0 *1 349.6,359.8
X$71652 16 657 348 622 623 22 DFF_X2
* cell instance $71662 r0 *1 367.08,359.8
X$71662 16 658 317 1668 18 22 DFF_X2
* cell instance $71663 m0 *1 369.36,359.8
X$71663 608 539 596 16 22 658 NAND3_X1
* cell instance $71670 m0 *1 372.78,359.8
X$71670 541 625 600 16 22 563 NAND3_X1
* cell instance $71672 m0 *1 376.77,359.8
X$71672 200 29 311 550 16 22 606 NAND4_X1
* cell instance $71673 m0 *1 377.72,359.8
X$71673 476 550 443 16 22 605 NAND3_X1
* cell instance $71674 m0 *1 378.48,359.8
X$71674 605 606 603 16 22 626 NAND3_X1
* cell instance $71677 m0 *1 383.8,359.8
X$71677 627 498 392 41 39 22 16 603 OAI221_X1
* cell instance $71679 m0 *1 385.13,359.8
X$71679 233 402 16 22 629 NOR2_X1
* cell instance $71684 r0 *1 377.91,359.8
X$71684 16 626 580 1672 550 22 DFF_X2
* cell instance $71688 r0 *1 383.99,359.8
X$71688 659 402 16 22 543 NOR2_X1
* cell instance $71689 r0 *1 384.56,359.8
X$71689 660 522 16 22 628 NOR2_X1
* cell instance $71694 r0 *1 387.98,359.8
X$71694 633 16 22 544 CLKBUF_X3
* cell instance $71696 m0 *1 389.31,359.8
X$71696 16 1477 661 569 580 22 DFF_X1
* cell instance $71700 m0 *1 395.77,359.8
X$71700 39 41 581 503 392 600 16 22 OAI221_X2
* cell instance $71703 r0 *1 389.31,359.8
X$71703 702 308 661 16 22 630 MUX2_X1
* cell instance $71704 r0 *1 390.64,359.8
X$71704 630 544 16 22 631 NOR2_X1
* cell instance $71705 r0 *1 391.21,359.8
X$71705 321 631 500 423 701 672 16 22 662 OAI33_X1
* cell instance $71709 m0 *1 399.76,359.8
X$71709 721 544 16 22 582 NOR2_X1
* cell instance $71712 m0 *1 400.71,359.8
X$71712 645 501 16 22 599 NOR2_X1
* cell instance $71714 m0 *1 403.56,359.8
X$71714 167 501 16 22 634 NOR2_X1
* cell instance $71715 m0 *1 404.13,359.8
X$71715 39 41 635 597 392 598 16 22 OAI221_X2
* cell instance $71717 m0 *1 406.41,359.8
X$71717 39 41 595 506 392 596 16 22 OAI221_X2
* cell instance $71720 m0 *1 413.06,359.8
X$71720 584 544 16 22 452 NOR2_X1
* cell instance $71723 m0 *1 414.58,359.8
X$71723 638 501 16 22 477 NOR2_X1
* cell instance $71724 m0 *1 415.15,359.8
X$71724 641 501 16 22 593 NOR2_X1
* cell instance $71728 r0 *1 400.9,359.8
X$71728 445 16 22 633 INV_X2
* cell instance $71730 r0 *1 402.99,359.8
X$71730 633 16 22 356 CLKBUF_X3
* cell instance $71731 r0 *1 403.94,359.8
X$71731 321 693 634 423 675 677 16 22 635 OAI33_X1
* cell instance $71735 r0 *1 406.6,359.8
X$71735 724 633 16 22 655 NOR2_X1
* cell instance $71737 r0 *1 407.93,359.8
X$71737 639 445 16 22 583 NOR2_X1
* cell instance $71740 r0 *1 412.3,359.8
X$71740 750 544 16 22 636 NOR2_X1
* cell instance $71745 m0 *1 418.57,359.8
X$71745 16 1521 585 511 586 22 DFF_X1
* cell instance $71747 m0 *1 421.8,359.8
X$71747 16 1466 461 556 586 22 DFF_X1
* cell instance $71749 m0 *1 431.11,359.8
X$71749 16 1519 549 644 363 22 DFF_X1
* cell instance $71752 r0 *1 418.76,359.8
X$71752 651 356 16 22 647 NOR2_X1
* cell instance $71754 r0 *1 420.85,359.8
X$71754 321 647 512 423 680 683 16 22 592 OAI33_X1
* cell instance $71758 m0 *1 434.91,359.8
X$71758 16 1399 590 589 363 22 DFF_X1
* cell instance $71760 m0 *1 438.14,359.8
X$71760 548 637 590 16 22 589 MUX2_X1
* cell instance $71761 m0 *1 439.47,359.8
X$71761 587 16 22 548 CLKBUF_X2
* cell instance $71772 r0 *1 436.05,359.8
X$71772 548 514 643 16 22 681 MUX2_X1
* cell instance $71774 r0 *1 437.57,359.8
X$71774 643 286 590 16 22 638 MUX2_X1
* cell instance $71864 m0 *1 707.56,359.8
X$71864 542 16 22 588 BUF_X1
* cell instance $72021 m0 *1 274.17,362.6
X$72021 16 1435 665 684 663 22 DFF_X1
* cell instance $72022 m0 *1 277.4,362.6
X$72022 665 664 460 16 22 684 MUX2_X1
* cell instance $72026 m0 *1 281.2,362.6
X$72026 613 666 667 16 22 762 MUX2_X1
* cell instance $72027 m0 *1 282.53,362.6
X$72027 667 664 432 16 22 686 MUX2_X1
* cell instance $72028 m0 *1 283.86,362.6
X$72028 16 1433 667 686 668 22 DFF_X1
* cell instance $72033 m0 *1 301.53,362.6
X$72033 553 666 646 16 22 1013 MUX2_X1
* cell instance $72040 m0 *1 325.09,362.6
X$72040 696 664 619 16 22 695 MUX2_X1
* cell instance $72044 m0 *1 330.41,362.6
X$72044 698 700 669 16 22 697 NAND3_X2
* cell instance $72055 r0 *1 276.64,362.6
X$72055 612 666 665 16 22 886 MUX2_X1
* cell instance $72065 r0 *1 289.94,362.6
X$72065 763 611 572 16 22 687 MUX2_X1
* cell instance $72070 r0 *1 294.12,362.6
X$72070 316 16 22 668 CLKBUF_X3
* cell instance $72071 r0 *1 295.07,362.6
X$72071 668 16 22 CLKBUF_X1
* cell instance $72073 r0 *1 296.4,362.6
X$72073 16 1607 707 731 668 22 DFF_X1
* cell instance $72077 r0 *1 309.51,362.6
X$72077 742 611 649 16 22 734 MUX2_X1
* cell instance $72080 r0 *1 315.4,362.6
X$72080 766 611 385 16 22 735 MUX2_X1
* cell instance $72084 r0 *1 324.71,362.6
X$72084 16 1590 696 695 709 22 DFF_X1
* cell instance $72087 r0 *1 328.89,362.6
X$72087 16 570 697 737 743 22 AOI21_X4
* cell instance $72090 m0 *1 334.59,362.6
X$72090 698 739 669 16 22 670 NAND3_X1
* cell instance $72102 r0 *1 334.59,362.6
X$72102 16 340 670 737 710 22 AOI21_X4
* cell instance $72105 r0 *1 338.96,362.6
X$72105 710 16 22 344 CLKBUF_X3
* cell instance $72111 r0 *1 341.05,362.6
X$72111 497 623 1678 22 16 739 HA_X1
* cell instance $72124 m0 *1 380.76,362.6
X$72124 713 445 16 22 704 NOR2_X1
* cell instance $72128 m0 *1 383.61,362.6
X$72128 705 704 423 629 671 321 16 22 627 OAI33_X1
* cell instance $72129 m0 *1 384.94,362.6
X$72129 715 633 16 22 705 NOR2_X1
* cell instance $72135 r0 *1 384.18,362.6
X$72135 714 522 16 22 671 NOR2_X1
* cell instance $72139 r0 *1 386.84,362.6
X$72139 16 1573 702 703 580 22 DFF_X1
* cell instance $72141 m0 *1 388.17,362.6
X$72141 702 238 83 16 22 703 MUX2_X1
* cell instance $72143 m0 *1 391.78,362.6
X$72143 716 402 16 22 701 NOR2_X1
* cell instance $72144 m0 *1 392.35,362.6
X$72144 717 522 16 22 672 NOR2_X1
* cell instance $72147 r0 *1 393.11,362.6
X$72147 718 238 168 16 22 738 MUX2_X1
* cell instance $72148 m0 *1 393.49,362.6
X$72148 633 16 22 522 CLKBUF_X3
* cell instance $72154 r0 *1 395.01,362.6
X$72154 718 308 719 16 22 673 MUX2_X1
* cell instance $72158 m0 *1 396.53,362.6
X$72158 673 544 16 22 674 NOR2_X1
* cell instance $72160 m0 *1 397.1,362.6
X$72160 321 674 632 423 699 694 16 22 581 OAI33_X1
* cell instance $72165 m0 *1 403.94,362.6
X$72165 723 544 16 22 693 NOR2_X1
* cell instance $72168 r0 *1 397.86,362.6
X$72168 720 402 16 22 699 NOR2_X1
* cell instance $72171 r0 *1 399,362.6
X$72171 878 522 16 22 694 NOR2_X1
* cell instance $72174 r0 *1 401.85,362.6
X$72174 722 238 64 16 22 736 MUX2_X1
* cell instance $72177 r0 *1 404.89,362.6
X$72177 891 402 16 22 675 NOR2_X1
* cell instance $72178 m0 *1 405.08,362.6
X$72178 676 522 16 22 677 NOR2_X1
* cell instance $72182 m0 *1 407.93,362.6
X$72182 688 633 16 22 507 NOR2_X1
* cell instance $72187 m0 *1 414.01,362.6
X$72187 689 544 16 22 678 NOR2_X1
* cell instance $72193 r0 *1 410.97,362.6
X$72193 725 238 208 16 22 733 MUX2_X1
* cell instance $72194 r0 *1 412.3,362.6
X$72194 16 1572 725 733 510 22 DFF_X1
* cell instance $72196 m0 *1 414.96,362.6
X$72196 321 678 691 423 679 685 16 22 595 OAI33_X1
* cell instance $72199 m0 *1 418.76,362.6
X$72199 730 522 16 22 685 NOR2_X1
* cell instance $72202 r0 *1 415.53,362.6
X$72202 732 227 208 16 22 751 MUX2_X1
* cell instance $72203 r0 *1 416.86,362.6
X$72203 725 308 732 16 22 651 MUX2_X1
* cell instance $72205 m0 *1 420.66,362.6
X$72205 931 402 16 22 679 NOR2_X1
* cell instance $72213 r0 *1 421.8,362.6
X$72213 682 522 16 22 683 NOR2_X1
* cell instance $72214 r0 *1 422.37,362.6
X$72214 729 402 16 22 680 NOR2_X1
* cell instance $72218 r0 *1 425.03,362.6
X$72218 208 304 765 16 22 726 MUX2_X1
* cell instance $72221 r0 *1 428.07,362.6
X$72221 208 332 727 16 22 728 MUX2_X1
* cell instance $72222 r0 *1 429.4,362.6
X$72222 16 1611 727 728 586 22 DFF_X1
* cell instance $72225 m0 *1 435.29,362.6
X$72225 16 1428 643 681 586 22 DFF_X1
* cell instance $72435 m0 *1 269.61,376.6
X$72435 1057 976 977 16 22 1006 MUX2_X1
* cell instance $72444 r0 *1 267.52,376.6
X$72444 16 1640 977 1006 864 22 DFF_X1
* cell instance $72447 r0 *1 272.65,376.6
X$72447 1129 906 977 16 22 1088 MUX2_X1
* cell instance $72450 r0 *1 275.88,376.6
X$72450 1088 1029 16 22 1007 NOR2_X1
* cell instance $72451 r0 *1 276.45,376.6
X$72451 1058 1029 16 22 1048 NOR2_X1
* cell instance $72453 m0 *1 278.35,376.6
X$72453 981 1059 1007 1032 978 1008 16 22 1016 OAI33_X1
* cell instance $72455 m0 *1 279.68,376.6
X$72455 981 1030 1048 1032 979 1009 16 22 1049 OAI33_X1
* cell instance $72459 m0 *1 283.48,376.6
X$72459 981 1010 1092 1032 982 951 16 22 1051 OAI33_X1
* cell instance $72466 r0 *1 279.11,376.6
X$72466 1089 1029 16 22 1092 NOR2_X1
* cell instance $72467 r0 *1 279.68,376.6
X$72467 981 1031 1061 1032 980 967 16 22 1050 OAI33_X1
* cell instance $72471 m0 *1 290.7,376.6
X$72471 981 1096 984 1032 1011 983 16 22 1052 OAI33_X1
* cell instance $72476 m0 *1 302.67,376.6
X$72476 1013 948 16 22 1014 NOR2_X1
* cell instance $72477 m0 *1 303.24,376.6
X$72477 737 991 1015 1016 440 554 16 22 OAI221_X2
* cell instance $72478 m0 *1 305.33,376.6
X$72478 737 991 1017 1049 440 573 16 22 OAI221_X2
* cell instance $72482 r0 *1 291.08,376.6
X$72482 1348 1029 16 22 984 NOR2_X1
* cell instance $72487 r0 *1 299.82,376.6
X$72487 1098 985 1033 1034 1064 1099 16 22 1015 OAI33_X1
* cell instance $72488 r0 *1 301.15,376.6
X$72488 1098 986 1100 1034 1066 1067 16 22 1017 OAI33_X1
* cell instance $72489 r0 *1 302.48,376.6
X$72489 737 991 1137 1051 440 367 16 22 OAI221_X2
* cell instance $72491 r0 *1 304.76,376.6
X$72491 737 991 1101 1052 440 412 16 22 OAI221_X2
* cell instance $72494 r0 *1 307.8,376.6
X$72494 780 991 1103 1050 440 618 16 22 OAI221_X2
* cell instance $72495 m0 *1 310.65,376.6
X$72495 777 948 16 22 989 NOR2_X1
* cell instance $72496 m0 *1 309.32,376.6
X$72496 981 1035 987 1032 989 988 16 22 1056 OAI33_X1
* cell instance $72500 m0 *1 311.6,376.6
X$72500 737 991 990 1056 440 346 16 22 OAI221_X2
* cell instance $72503 m0 *1 320.72,376.6
X$72503 16 1410 992 1025 870 22 DFF_X1
* cell instance $72504 m0 *1 323.95,376.6
X$72504 992 947 900 16 22 993 MUX2_X1
* cell instance $72506 m0 *1 325.47,376.6
X$72506 991 737 994 1053 440 620 16 22 OAI221_X2
* cell instance $72511 r0 *1 313.31,376.6
X$72511 868 1029 16 22 1140 NOR2_X1
* cell instance $72514 r0 *1 315.78,376.6
X$72514 981 1105 1104 1032 1022 1036 16 22 1055 OAI33_X1
* cell instance $72515 r0 *1 317.11,376.6
X$72515 737 991 1138 1055 440 373 16 22 OAI221_X2
* cell instance $72516 r0 *1 319.2,376.6
X$72516 1054 16 22 1029 CLKBUF_X3
* cell instance $72518 r0 *1 320.34,376.6
X$72518 708 1029 16 22 1199 NOR2_X1
* cell instance $72522 r0 *1 325.66,376.6
X$72522 974 1037 16 22 1070 NOR2_X1
* cell instance $72523 r0 *1 326.23,376.6
X$72523 1070 1108 1032 1071 1109 981 16 22 994 OAI33_X1
* cell instance $72525 r0 *1 329.08,376.6
X$72525 1038 1072 16 1032 22 NAND2_X4
* cell instance $72528 r0 *1 332.5,376.6
X$72528 1111 995 946 22 16 1112 OAI21_X4
* cell instance $72530 m0 *1 332.5,376.6
X$72530 1028 995 946 22 16 1027 OAI21_X4
* cell instance $72535 r0 *1 336.87,376.6
X$72535 913 1073 946 22 16 976 OAI21_X4
* cell instance $72537 r0 *1 339.72,376.6
X$72537 16 1073 22 995 BUF_X8
* cell instance $72539 m0 *1 342.38,376.6
X$72539 1024 954 1039 16 22 955 MUX2_X1
* cell instance $72545 r0 *1 342.57,376.6
X$72545 259 1065 16 22 1039 NOR2_X1
* cell instance $72549 m0 *1 349.41,376.6
X$72549 16 1485 972 996 1078 22 DFF_X1
* cell instance $72555 m0 *1 375.63,376.6
X$72555 16 1537 959 1019 875 22 DFF_X1
* cell instance $72556 m0 *1 378.86,376.6
X$72556 959 255 1079 16 22 659 MUX2_X1
* cell instance $72569 r0 *1 381.71,376.6
X$72569 16 1614 1018 1040 1041 22 DFF_X1
* cell instance $72570 m0 *1 382.28,376.6
X$72570 876 254 1018 16 22 1040 MUX2_X1
* cell instance $72574 m0 *1 391.21,376.6
X$72574 960 16 22 83 BUF_X2
* cell instance $72580 r0 *1 387.03,376.6
X$72580 266 22 520 16 BUF_X4
* cell instance $72581 r0 *1 388.36,376.6
X$72581 83 304 1113 16 22 1114 MUX2_X1
* cell instance $72584 r0 *1 390.64,376.6
X$72584 1080 255 1113 16 22 716 MUX2_X1
* cell instance $72586 r0 *1 395.01,376.6
X$72586 16 1577 998 1042 1041 22 DFF_X1
* cell instance $72587 m0 *1 396.72,376.6
X$72587 998 255 997 16 22 720 MUX2_X1
* cell instance $72588 m0 *1 395.39,376.6
X$72588 939 225 998 16 22 1042 MUX2_X1
* cell instance $72594 r0 *1 403.56,376.6
X$72594 64 304 1107 16 22 1081 MUX2_X1
* cell instance $72596 m0 *1 404.51,376.6
X$72596 999 16 22 64 BUF_X2
* cell instance $72598 r0 *1 404.89,376.6
X$72598 1082 520 1107 16 22 891 MUX2_X1
* cell instance $72600 r0 *1 407.74,376.6
X$72600 999 225 1082 16 22 1083 MUX2_X1
* cell instance $72602 r0 *1 409.83,376.6
X$72602 266 22 255 16 BUF_X4
* cell instance $72604 m0 *1 412.3,376.6
X$72604 753 254 962 16 22 1043 MUX2_X1
* cell instance $72605 m0 *1 411.73,376.6
X$72605 838 16 22 CLKBUF_X1
* cell instance $72606 m0 *1 413.63,376.6
X$72606 749 16 22 838 CLKBUF_X3
* cell instance $72610 r0 *1 412.49,376.6
X$72610 16 1575 962 1043 838 22 DFF_X1
* cell instance $72611 m0 *1 415.15,376.6
X$72611 879 16 22 183 BUF_X2
* cell instance $72616 m0 *1 425.79,376.6
X$72616 16 1416 1001 1000 1002 22 DFF_X1
* cell instance $72619 m0 *1 435.86,376.6
X$72619 16 1522 1003 1047 1002 22 DFF_X1
* cell instance $72624 r0 *1 419.71,376.6
X$72624 183 304 1045 16 22 1044 MUX2_X1
* cell instance $72626 r0 *1 421.8,376.6
X$72626 1084 520 1045 16 22 931 MUX2_X1
* cell instance $72632 r0 *1 432.06,376.6
X$72632 939 637 1090 16 22 1091 MUX2_X1
* cell instance $72636 r0 *1 437.38,376.6
X$72636 1087 16 22 960 BUF_X2
* cell instance $72638 m0 *1 439.66,376.6
X$72638 16 1520 965 1005 1002 22 DFF_X1
* cell instance $72691 r0 *1 446.5,376.6
X$72691 1046 16 22 999 BUF_X2
* cell instance $72738 r0 *1 704.71,376.6
X$72738 924 16 22 1086 BUF_X1
* cell instance $72896 m0 *1 272.27,387.8
X$72896 1210 1141 1235 16 22 1244 MUX2_X1
* cell instance $72897 m0 *1 269.04,387.8
X$72897 16 1469 1235 1244 1211 22 DFF_X1
* cell instance $72900 m0 *1 277.4,387.8
X$72900 1246 653 1259 16 22 1060 MUX2_X1
* cell instance $72905 r0 *1 274.17,387.8
X$72905 1210 1242 1246 16 22 1266 MUX2_X1
* cell instance $72908 r0 *1 277.4,387.8
X$72908 1210 1228 1259 16 22 1267 MUX2_X1
* cell instance $72911 r0 *1 281.96,387.8
X$72911 16 1554 1250 1236 1211 22 DFF_X1
* cell instance $72913 m0 *1 282.15,387.8
X$72913 1210 1027 1250 16 22 1236 MUX2_X1
* cell instance $72916 m0 *1 285.95,387.8
X$72916 16 1451 1237 1251 1211 22 DFF_X1
* cell instance $72917 m0 *1 289.18,387.8
X$72917 1250 1219 1237 16 22 1133 MUX2_X1
* cell instance $72921 m0 *1 292.98,387.8
X$72921 16 1532 1215 1238 1239 22 DFF_X1
* cell instance $72931 r0 *1 295.26,387.8
X$72931 1260 855 572 16 22 1269 MUX2_X1
* cell instance $72933 m0 *1 300.58,387.8
X$72933 1257 871 432 16 22 1256 MUX2_X1
* cell instance $72934 m0 *1 297.35,387.8
X$72934 16 1528 1255 1240 1239 22 DFF_X1
* cell instance $72935 m0 *1 301.91,387.8
X$72935 16 1417 1257 1256 1239 22 DFF_X1
* cell instance $72938 r0 *1 297.35,387.8
X$72938 1260 653 1290 16 22 1176 MUX2_X1
* cell instance $72941 r0 *1 299.63,387.8
X$72941 1121 16 22 1239 CLKBUF_X3
* cell instance $72942 r0 *1 300.58,387.8
X$72942 1239 16 22 CLKBUF_X1
* cell instance $72945 r0 *1 304.57,387.8
X$72945 16 1657 1262 1270 1239 22 DFF_X1
* cell instance $72946 r0 *1 307.8,387.8
X$72946 1262 855 813 16 22 1270 MUX2_X1
* cell instance $72948 m0 *1 308.56,387.8
X$72948 1262 653 1231 16 22 1149 MUX2_X1
* cell instance $72952 m0 *1 312.74,387.8
X$72952 16 1496 1218 1254 894 22 DFF_X1
* cell instance $72957 m0 *1 318.06,387.8
X$72957 16 1497 1247 1248 1249 22 DFF_X1
* cell instance $72964 r0 *1 324.52,387.8
X$72964 1249 16 22 1693 INV_X1
* cell instance $72965 r0 *1 324.9,387.8
X$72965 16 1589 1263 1268 1249 22 DFF_X1
* cell instance $72966 m0 *1 325.66,387.8
X$72966 1121 16 22 1249 CLKBUF_X3
* cell instance $72972 m0 *1 342,387.8
X$72972 1243 16 22 770 BUF_X2
* cell instance $73038 r0 *1 328.13,387.8
X$73038 1263 653 1264 16 22 1203 MUX2_X1
* cell instance $73042 r0 *1 332.12,387.8
X$73042 619 1214 1264 16 22 1265 MUX2_X1
* cell instance $73043 r0 *1 333.45,387.8
X$73043 16 1616 1264 1265 1249 22 DFF_X1
* cell instance $73243 m0 *1 261.82,385
X$73243 1208 16 22 1210 CLKBUF_X2
* cell instance $73250 m0 *1 266.19,385
X$73250 1207 16 22 1057 CLKBUF_X2
* cell instance $73257 r0 *1 269.61,385
X$73257 16 1557 1212 1209 1211 22 DFF_X1
* cell instance $73258 m0 *1 271.7,385
X$73258 1235 906 1212 16 22 1058 MUX2_X1
* cell instance $73259 m0 *1 270.37,385
X$73259 1210 976 1212 16 22 1209 MUX2_X1
* cell instance $73261 m0 *1 276.07,385
X$73261 1210 16 22 460 BUF_X2
* cell instance $73262 m0 *1 276.83,385
X$73262 1057 1228 1142 16 22 1227 MUX2_X1
* cell instance $73266 m0 *1 283.48,385
X$73266 1210 1112 1213 16 22 1229 MUX2_X1
* cell instance $73267 m0 *1 284.81,385
X$73267 16 1450 1213 1229 1211 22 DFF_X1
* cell instance $73270 m0 *1 295.64,385
X$73270 1213 947 1215 16 22 1178 MUX2_X1
* cell instance $73275 m0 *1 307.04,385
X$73275 1231 871 813 16 22 1217 MUX2_X1
* cell instance $73284 r0 *1 282.72,385
X$73284 1121 16 22 1211 CLKBUF_X3
* cell instance $73288 r0 *1 283.67,385
X$73288 1211 16 22 1691 INV_X1
* cell instance $73291 r0 *1 287.28,385
X$73291 460 1252 1237 16 22 1251 MUX2_X1
* cell instance $73297 r0 *1 294.5,385
X$73297 460 1214 1215 16 22 1238 MUX2_X1
* cell instance $73301 r0 *1 297.92,385
X$73301 1255 855 432 16 22 1240 MUX2_X1
* cell instance $73304 r0 *1 300.2,385
X$73304 1255 653 1257 16 22 1216 MUX2_X1
* cell instance $73308 r0 *1 306.47,385
X$73308 16 1655 1231 1217 894 22 DFF_X1
* cell instance $73311 r0 *1 313.12,385
X$73311 1218 871 649 16 22 1254 MUX2_X1
* cell instance $73315 r0 *1 318.44,385
X$73315 1247 871 385 16 22 1248 MUX2_X1
* cell instance $73318 m0 *1 324.52,385
X$73318 1234 1219 1221 16 22 1153 MUX2_X1
* cell instance $73319 m0 *1 323.19,385
X$73319 1234 855 619 16 22 1220 MUX2_X1
* cell instance $73322 m0 *1 327.56,385
X$73322 1221 871 619 16 22 1222 MUX2_X1
* cell instance $73333 m0 *1 389.69,385
X$73333 16 1518 1159 1230 1162 22 DFF_X1
* cell instance $73334 m0 *1 392.92,385
X$73334 960 253 1159 16 22 1230 MUX2_X1
* cell instance $73338 m0 *1 398.24,385
X$73338 939 253 1161 16 22 1223 MUX2_X1
* cell instance $73342 r0 *1 323.76,385
X$73342 16 1615 1234 1220 1249 22 DFF_X1
* cell instance $73344 r0 *1 327.37,385
X$73344 16 1571 1221 1222 1249 22 DFF_X1
* cell instance $73364 r0 *1 398.43,385
X$73364 16 1585 1161 1223 1162 22 DFF_X1
* cell instance $73367 m0 *1 402.99,385
X$73367 16 1411 1224 1226 1162 22 DFF_X1
* cell instance $73589 m0 *1 272.65,365.4
X$73589 761 611 740 16 22 760 MUX2_X1
* cell instance $73590 m0 *1 273.98,365.4
X$73590 16 1434 761 760 663 22 DFF_X1
* cell instance $73601 r0 *1 273.03,365.4
X$73601 814 664 740 16 22 843 MUX2_X1
* cell instance $73603 m0 *1 278.54,365.4
X$73603 663 16 22 CLKBUF_X1
* cell instance $73604 m0 *1 277.59,365.4
X$73604 316 16 22 663 CLKBUF_X3
* cell instance $73608 m0 *1 288.99,365.4
X$73608 16 1492 763 687 668 22 DFF_X1
* cell instance $73611 m0 *1 295.45,365.4
X$73611 741 464 740 16 22 764 MUX2_X1
* cell instance $73614 r0 *1 280.82,365.4
X$73614 845 340 813 16 22 847 MUX2_X1
* cell instance $73616 r0 *1 282.34,365.4
X$73616 815 340 740 16 22 774 MUX2_X1
* cell instance $73621 r0 *1 294.69,365.4
X$73621 16 1606 741 764 668 22 DFF_X1
* cell instance $73622 m0 *1 298.49,365.4
X$73622 741 666 707 16 22 820 MUX2_X1
* cell instance $73623 m0 *1 297.16,365.4
X$73623 707 466 740 16 22 731 MUX2_X1
* cell instance $73628 m0 *1 308.37,365.4
X$73628 16 1424 742 734 536 22 DFF_X1
* cell instance $73630 m0 *1 314.64,365.4
X$73630 16 1488 766 735 709 22 DFF_X1
* cell instance $73635 r0 *1 301.72,365.4
X$73635 775 464 813 16 22 801 MUX2_X1
* cell instance $73636 r0 *1 303.05,365.4
X$73636 16 1613 775 801 668 22 DFF_X1
* cell instance $73639 r0 *1 307.23,365.4
X$73639 16 1610 776 803 536 22 DFF_X1
* cell instance $73640 r0 *1 310.46,365.4
X$73640 776 664 649 16 22 803 MUX2_X1
* cell instance $73643 r0 *1 314.07,365.4
X$73643 316 16 22 1695 CLKBUF_X3
* cell instance $73644 r0 *1 315.02,365.4
X$73644 779 664 385 16 22 853 MUX2_X1
* cell instance $73645 r0 *1 316.35,365.4
X$73645 786 16 22 316 CLKBUF_X3
* cell instance $73647 m0 *1 322.24,365.4
X$73647 709 16 22 1687 INV_X1
* cell instance $73648 m0 *1 321.29,365.4
X$73648 316 16 22 709 CLKBUF_X3
* cell instance $73652 m0 *1 327.94,365.4
X$73652 16 611 769 737 743 22 AOI21_X4
* cell instance $73653 m0 *1 330.41,365.4
X$73653 698 711 669 16 22 769 NAND3_X2
* cell instance $73661 r0 *1 328.13,365.4
X$73661 16 664 810 737 743 22 AOI21_X4
* cell instance $73663 r0 *1 330.79,365.4
X$73663 698 812 669 16 22 810 NAND3_X2
* cell instance $73665 m0 *1 339.91,365.4
X$73665 739 745 16 22 771 NAND2_X1
* cell instance $73666 m0 *1 337.44,365.4
X$73666 16 743 22 710 BUF_X8
* cell instance $73667 m0 *1 340.48,365.4
X$73667 771 780 344 16 744 22 AOI21_X1
* cell instance $73669 m0 *1 341.43,365.4
X$73669 497 623 669 745 16 22 808 NAND4_X1
* cell instance $73672 m0 *1 344.09,365.4
X$73672 109 782 16 22 712 NOR2_X1
* cell instance $73673 m0 *1 344.66,365.4
X$73673 712 744 773 16 22 806 MUX2_X1
* cell instance $73674 m0 *1 345.99,365.4
X$73674 259 669 16 22 773 NOR2_X1
* cell instance $73678 r0 *1 339.15,365.4
X$73678 781 743 780 16 577 22 AOI21_X2
* cell instance $73680 r0 *1 340.67,365.4
X$73680 808 780 344 16 807 22 AOI21_X1
* cell instance $73682 r0 *1 341.62,365.4
X$73682 607 623 1682 22 16 812 HA_X1
* cell instance $73687 r0 *1 346.37,365.4
X$73687 16 806 870 1676 783 22 DFF_X2
* cell instance $73689 m0 *1 346.94,365.4
X$73689 783 22 669 16 BUF_X4
* cell instance $73695 m0 *1 375.82,365.4
X$73695 195 304 746 16 22 802 MUX2_X1
* cell instance $73700 r0 *1 353.4,365.4
X$73700 826 805 22 16 784 AND2_X1
* cell instance $73701 r0 *1 354.16,365.4
X$73701 623 785 805 22 16 861 HA_X1
* cell instance $73709 r0 *1 363.28,365.4
X$73709 804 16 22 758 INV_X4
* cell instance $73710 r0 *1 364.23,365.4
X$73710 343 804 788 22 16 797 OAI21_X4
* cell instance $73715 r0 *1 374.87,365.4
X$73715 16 1644 746 802 580 22 DFF_X1
* cell instance $73717 m0 *1 379.24,365.4
X$73717 858 308 746 16 22 713 MUX2_X1
* cell instance $73719 m0 *1 380.57,365.4
X$73719 747 238 195 16 22 772 MUX2_X1
* cell instance $73720 m0 *1 381.9,365.4
X$73720 16 1408 747 772 580 22 DFF_X1
* cell instance $73721 m0 *1 385.13,365.4
X$73721 749 16 22 580 CLKBUF_X3
* cell instance $73722 m0 *1 386.08,365.4
X$73722 580 16 22 CLKBUF_X1
* cell instance $73726 m0 *1 391.97,365.4
X$73726 16 1484 718 738 580 22 DFF_X1
* cell instance $73730 m0 *1 399.95,365.4
X$73730 16 1498 722 736 510 22 DFF_X1
* cell instance $73731 m0 *1 403.18,365.4
X$73731 722 308 799 16 22 723 MUX2_X1
* cell instance $73736 r0 *1 380.19,365.4
X$73736 16 1552 789 790 580 22 DFF_X1
* cell instance $73737 r0 *1 383.42,365.4
X$73737 747 520 789 16 22 714 MUX2_X1
* cell instance $73743 r0 *1 401.85,365.4
X$73743 799 227 64 16 22 800 MUX2_X1
* cell instance $73747 r0 *1 407.17,365.4
X$73747 16 1579 767 768 510 22 DFF_X1
* cell instance $73748 m0 *1 408.12,365.4
X$73748 767 238 183 16 22 768 MUX2_X1
* cell instance $73751 m0 *1 410.02,365.4
X$73751 767 308 748 16 22 689 MUX2_X1
* cell instance $73754 m0 *1 411.54,365.4
X$73754 749 16 22 510 CLKBUF_X3
* cell instance $73755 m0 *1 412.49,365.4
X$73755 510 16 22 CLKBUF_X1
* cell instance $73759 m0 *1 415.53,365.4
X$73759 16 1481 732 751 510 22 DFF_X1
* cell instance $73766 r0 *1 423.32,365.4
X$73766 753 225 752 16 22 793 MUX2_X1
* cell instance $73767 m0 *1 423.89,365.4
X$73767 752 255 765 16 22 729 MUX2_X1
* cell instance $73769 m0 *1 425.22,365.4
X$73769 16 1426 765 726 586 22 DFF_X1
* cell instance $73770 m0 *1 428.45,365.4
X$73770 753 16 22 208 BUF_X2
* cell instance $73773 m0 *1 430.54,365.4
X$73773 754 520 727 16 22 682 MUX2_X1
* cell instance $73774 m0 *1 429.59,365.4
X$73774 749 16 22 586 CLKBUF_X3
* cell instance $73777 m0 *1 435.67,365.4
X$73777 753 514 755 16 22 798 MUX2_X1
* cell instance $73782 r0 *1 434.72,365.4
X$73782 16 1608 755 798 586 22 DFF_X1
* cell instance $73784 m0 *1 437.38,365.4
X$73784 755 286 756 16 22 641 MUX2_X1
* cell instance $73786 m0 *1 439.28,365.4
X$73786 753 637 756 16 22 759 MUX2_X1
* cell instance $73788 m0 *1 440.61,365.4
X$73788 16 1430 756 759 586 22 DFF_X1
* cell instance $73837 m0 *1 708.7,365.4
X$73837 758 16 22 757 BUF_X1
* cell instance $73888 r0 *1 709.08,365.4
X$73888 797 16 22 795 BUF_X1
* cell instance $74050 r0 *1 276.26,401.8
X$74050 16 1620 1354 1370 1318 22 DFF_X1
* cell instance $74051 m0 *1 279.87,401.8
X$74051 1318 16 22 1686 INV_X1
* cell instance $74052 m0 *1 278.92,401.8
X$74052 1121 16 22 1318 CLKBUF_X3
* cell instance $74057 r0 *1 279.49,401.8
X$74057 1354 930 1371 16 22 1171 MUX2_X1
* cell instance $74063 r0 *1 284.62,401.8
X$74063 1334 1112 1352 16 22 1365 MUX2_X1
* cell instance $74067 r0 *1 288.04,401.8
X$74067 16 1621 1341 1362 1361 22 DFF_X1
* cell instance $74068 m0 *1 289.18,401.8
X$74068 1351 1141 1341 16 22 1362 MUX2_X1
* cell instance $74071 m0 *1 290.7,401.8
X$74071 1341 906 1342 16 22 1348 MUX2_X1
* cell instance $74073 m0 *1 292.22,401.8
X$74073 1351 976 1342 16 22 1349 MUX2_X1
* cell instance $74074 m0 *1 293.55,401.8
X$74074 16 1531 1342 1349 1275 22 DFF_X1
* cell instance $74082 r0 *1 301.34,401.8
X$74082 16 1649 1322 1353 1275 22 DFF_X1
* cell instance $74083 m0 *1 301.91,401.8
X$74083 1351 1112 1322 16 22 1353 MUX2_X1
* cell instance $74090 m0 *1 322.43,401.8
X$74090 1335 1112 1343 16 22 1360 MUX2_X1
* cell instance $74092 m0 *1 325.28,401.8
X$74092 1299 16 22 1393 INV_X2
* cell instance $74093 m0 *1 325.85,401.8
X$74093 1121 16 22 1299 CLKBUF_X3
* cell instance $74098 r0 *1 305.9,401.8
X$74098 1298 1141 1363 16 22 1376 MUX2_X1
* cell instance $74101 r0 *1 308.94,401.8
X$74101 1363 906 1355 16 22 1068 MUX2_X1
* cell instance $74102 r0 *1 310.27,401.8
X$74102 1298 976 1355 16 22 1375 MUX2_X1
* cell instance $74104 r0 *1 314.64,401.8
X$74104 1335 1141 1356 16 22 1372 MUX2_X1
* cell instance $74106 r0 *1 316.35,401.8
X$74106 1356 906 1357 16 22 1106 MUX2_X1
* cell instance $74108 r0 *1 318.06,401.8
X$74108 1335 976 1357 16 22 1374 MUX2_X1
* cell instance $74113 r0 *1 322.24,401.8
X$74113 16 1625 1343 1360 1325 22 DFF_X1
* cell instance $74115 r0 *1 326.99,401.8
X$74115 16 1622 1328 1358 1299 22 DFF_X1
* cell instance $74117 m0 *1 327.18,401.8
X$74117 1280 1141 1328 16 22 1358 MUX2_X1
* cell instance $74143 r0 *1 330.22,401.8
X$74143 1359 16 22 1280 BUF_X1
* cell instance $75300 m0 *1 355.49,331.8
X$75300 93 16 22 36 BUF_X2
* cell instance $75301 m0 *1 356.25,331.8
X$75301 95 36 94 77 78 76 22 16 AOI221_X2
* cell instance $75331 r0 *1 355.49,331.8
X$75331 216 105 93 22 16 94 HA_X1
* cell instance $75337 m0 *1 361,331.8
X$75337 106 16 22 61 INV_X1
* cell instance $75342 m0 *1 367.08,331.8
X$75342 16 79 22 96 BUF_X8
* cell instance $75343 m0 *1 369.55,331.8
X$75343 81 22 80 16 BUF_X4
* cell instance $75344 m0 *1 370.88,331.8
X$75344 81 16 22 121 INV_X4
* cell instance $75350 m0 *1 389.31,331.8
X$75350 101 88 83 16 22 82 MUX2_X1
* cell instance $75353 m0 *1 392.92,331.8
X$75353 84 65 83 16 22 103 MUX2_X1
* cell instance $75354 m0 *1 394.25,331.8
X$75354 102 54 83 16 22 100 MUX2_X1
* cell instance $75361 m0 *1 423.13,331.8
X$75361 90 88 87 16 22 91 MUX2_X1
* cell instance $75362 m0 *1 424.46,331.8
X$75362 16 1460 90 91 71 22 DFF_X1
* cell instance $75416 r0 *1 368.03,331.8
X$75416 109 80 16 22 119 NOR2_X1
* cell instance $75417 r0 *1 368.6,331.8
X$75417 98 108 119 16 22 97 MUX2_X1
* cell instance $75418 r0 *1 369.93,331.8
X$75418 109 121 16 22 98 NOR2_X1
* cell instance $75422 r0 *1 378.86,331.8
X$75422 16 37 22 130 BUF_X8
* cell instance $75426 r0 *1 389.12,331.8
X$75426 16 1650 101 82 63 22 DFF_X1
* cell instance $75427 r0 *1 392.35,331.8
X$75427 16 1658 84 103 63 22 DFF_X1
* cell instance $75432 r0 *1 395.77,331.8
X$75432 102 86 84 16 22 110 MUX2_X1
* cell instance $75435 r0 *1 398.05,331.8
X$75435 16 1559 85 99 63 22 DFF_X1
* cell instance $75436 r0 *1 401.28,331.8
X$75436 85 88 64 16 22 99 MUX2_X1
* cell instance $75439 r0 *1 408.88,331.8
X$75439 159 16 22 55 CLKBUF_X3
* cell instance $75440 r0 *1 409.83,331.8
X$75440 55 16 22 CLKBUF_X1
* cell instance $75441 r0 *1 410.4,331.8
X$75441 111 54 87 16 22 117 MUX2_X1
* cell instance $75444 r0 *1 413.44,331.8
X$75444 136 65 87 16 22 113 MUX2_X1
* cell instance $75448 r0 *1 418.95,331.8
X$75448 72 114 142 16 22 115 MUX2_X1
* cell instance $75451 r0 *1 421.99,331.8
X$75451 16 1548 138 89 71 22 DFF_X1
* cell instance $75647 m0 *1 360.81,317.8
X$75647 31 33 16 22 30 NAND2_X1
* cell instance $75648 m0 *1 361.38,317.8
X$75648 31 16 22 27 BUF_X1
* cell instance $75677 r0 *1 359.29,317.8
X$75677 35 16 22 28 BUF_X1
* cell instance $75678 r0 *1 359.86,317.8
X$75678 35 16 22 33 CLKBUF_X2
* cell instance $75681 r0 *1 361.19,317.8
X$75681 16 37 24 31 42 44 22 NOR4_X4
* cell instance $75683 m0 *1 362.33,317.8
X$75683 29 38 30 22 16 20 OAI21_X4
* cell instance $75748 r0 *1 376.01,317.8
X$75748 41 29 40 16 22 NOR2_X4
* cell instance $75753 r0 *1 383.23,317.8
X$75753 39 41 26 16 22 NOR2_X4
* cell instance $75962 r0 *1 357.2,329
X$75962 36 60 22 16 77 AND2_X1
* cell instance $75963 m0 *1 357.96,329
X$75963 52 16 22 78 BUF_X2
* cell instance $75964 m0 *1 358.72,329
X$75964 16 61 52 35 59 53 22 FA_X1
* cell instance $75965 m0 *1 361.76,329
X$75965 60 74 22 16 62 AND2_X1
* cell instance $75966 m0 *1 362.52,329
X$75966 53 59 74 22 16 75 HA_X1
* cell instance $75969 m0 *1 367.65,329
X$75969 16 97 125 1659 81 22 DFF_X2
* cell instance $75975 m0 *1 401.66,329
X$75975 57 54 64 16 22 58 MUX2_X1
* cell instance $75982 r0 *1 361.76,329
X$75982 62 61 95 60 75 48 22 16 AOI221_X2
* cell instance $75984 r0 *1 365.37,329
X$75984 143 81 60 22 16 95 HA_X1
* cell instance $75991 r0 *1 392.16,329
X$75991 16 1652 102 100 63 22 DFF_X1
* cell instance $75997 r0 *1 404.32,329
X$75997 57 86 67 16 22 206 MUX2_X1
* cell instance $75999 m0 *1 404.89,329
X$75999 16 1461 67 66 55 22 DFF_X1
* cell instance $76001 m0 *1 411.92,329
X$76001 56 54 70 16 22 73 MUX2_X1
* cell instance $76002 m0 *1 413.25,329
X$76002 16 1471 69 68 71 22 DFF_X1
* cell instance $76056 r0 *1 405.65,329
X$76056 67 65 64 16 22 66 MUX2_X1
* cell instance $76060 r0 *1 409.45,329
X$76060 16 1635 56 73 55 22 DFF_X1
* cell instance $76061 r0 *1 412.68,329
X$76061 56 86 69 16 22 357 MUX2_X1
* cell instance $76062 r0 *1 414.01,329
X$76062 69 65 70 16 22 68 MUX2_X1
* cell instance $76063 r0 *1 415.34,329
X$76063 16 1633 72 92 71 22 DFF_X1
* cell instance $76064 r0 *1 418.57,329
X$76064 72 88 70 16 22 92 MUX2_X1
* cell instance $76284 m0 *1 351.31,337.4
X$76284 122 174 22 16 149 AND2_X1
* cell instance $76288 m0 *1 358.34,337.4
X$76288 124 150 22 16 151 AND2_X1
* cell instance $76295 r0 *1 356.25,337.4
X$76295 174 16 22 150 CLKBUF_X3
* cell instance $76298 r0 *1 357.77,337.4
X$76298 187 153 151 16 22 123 MUX2_X1
* cell instance $76299 r0 *1 359.1,337.4
X$76299 127 257 22 16 187 AND2_X1
* cell instance $76301 r0 *1 360.24,337.4
X$76301 59 174 22 16 189 AND2_X1
* cell instance $76303 r0 *1 361.19,337.4
X$76303 189 153 175 16 22 198 MUX2_X1
* cell instance $76305 m0 *1 361.76,337.4
X$76305 166 150 22 16 175 AND2_X1
* cell instance $76309 m0 *1 363.66,337.4
X$76309 124 154 166 22 16 147 HA_X1
* cell instance $76313 r0 *1 365.37,337.4
X$76313 176 79 37 16 153 22 AOI21_X2
* cell instance $76315 m0 *1 365.94,337.4
X$76315 127 154 1677 22 16 157 HA_X1
* cell instance $76316 m0 *1 368.6,337.4
X$76316 25 16 22 176 INV_X4
* cell instance $76323 r0 *1 369.55,337.4
X$76323 122 25 16 22 177 NAND2_X1
* cell instance $76325 m0 *1 370.88,337.4
X$76325 144 16 22 155 INV_X1
* cell instance $76327 m0 *1 371.26,337.4
X$76327 16 176 122 121 173 249 22 NOR4_X4
* cell instance $76328 m0 *1 374.68,337.4
X$76328 107 16 22 173 INV_X1
* cell instance $76330 m0 *1 376.58,337.4
X$76330 129 147 80 16 22 172 NAND3_X2
* cell instance $76331 m0 *1 377.91,337.4
X$76331 129 144 80 16 22 170 NAND3_X2
* cell instance $76334 m0 *1 381.52,337.4
X$76334 16 212 170 37 79 22 AOI21_X4
* cell instance $76339 r0 *1 370.88,337.4
X$76339 16 176 122 121 155 156 22 NOR4_X4
* cell instance $76340 r0 *1 374.3,337.4
X$76340 131 107 121 16 22 223 NAND3_X2
* cell instance $76341 r0 *1 375.63,337.4
X$76341 121 147 129 22 16 194 AND3_X1
* cell instance $76342 r0 *1 376.58,337.4
X$76342 131 157 121 16 22 226 NAND3_X2
* cell instance $76343 r0 *1 377.91,337.4
X$76343 121 157 129 22 16 202 AND3_X1
* cell instance $76345 r0 *1 380.38,337.4
X$76345 16 181 172 37 79 22 AOI21_X4
* cell instance $76348 r0 *1 385.13,337.4
X$76348 178 134 195 16 22 179 MUX2_X1
* cell instance $76353 r0 *1 392.16,337.4
X$76353 16 1647 158 169 63 22 DFF_X1
* cell instance $76355 m0 *1 394.25,337.4
X$76355 158 88 168 16 22 169 MUX2_X1
* cell instance $76363 m0 *1 428.45,337.4
X$76363 160 181 70 16 22 165 MUX2_X1
* cell instance $76364 m0 *1 429.78,337.4
X$76364 160 114 161 16 22 164 MUX2_X1
* cell instance $76367 r0 *1 395.58,337.4
X$76367 158 86 180 16 22 270 MUX2_X1
* cell instance $76368 r0 *1 396.91,337.4
X$76368 180 134 168 16 22 193 MUX2_X1
* cell instance $76369 r0 *1 398.24,337.4
X$76369 16 1546 180 193 205 22 DFF_X1
* cell instance $76375 r0 *1 410.4,337.4
X$76375 192 54 208 16 22 191 MUX2_X1
* cell instance $76378 r0 *1 414.01,337.4
X$76378 182 88 183 16 22 190 MUX2_X1
* cell instance $76379 r0 *1 415.34,337.4
X$76379 16 1639 184 188 55 22 DFF_X1
* cell instance $76380 r0 *1 418.57,337.4
X$76380 184 134 183 16 22 188 MUX2_X1
* cell instance $76385 r0 *1 422.75,337.4
X$76385 16 1540 209 186 213 22 DFF_X1
* cell instance $76388 r0 *1 426.55,337.4
X$76388 215 134 208 16 22 185 MUX2_X1
* cell instance $76390 m0 *1 431.68,337.4
X$76390 161 212 70 16 22 163 MUX2_X1
* cell instance $76395 m0 *1 434.34,337.4
X$76395 16 1533 161 163 71 22 DFF_X1
* cell instance $76673 r0 *1 342.57,343
X$76673 316 16 22 104 CLKBUF_X3
* cell instance $76674 r0 *1 343.52,343
X$76674 104 16 22 1395 INV_X2
* cell instance $76678 r0 *1 351.88,343
X$76678 16 1602 196 243 104 22 DFF_X1
* cell instance $76679 m0 *1 354.35,343
X$76679 196 174 22 16 242 AND2_X1
* cell instance $76681 m0 *1 355.11,343
X$76681 109 196 16 22 230 NOR2_X1
* cell instance $76682 m0 *1 355.68,343
X$76682 196 260 22 16 197 XNOR2_X1
* cell instance $76687 m0 *1 365.37,343
X$76687 16 231 22 232 BUF_X8
* cell instance $76691 r0 *1 355.11,343
X$76691 242 65 230 16 22 243 MUX2_X1
* cell instance $76698 r0 *1 369.17,343
X$76698 231 22 29 16 BUF_X4
* cell instance $76701 r0 *1 373.73,343
X$76701 249 231 41 22 16 253 OAI21_X4
* cell instance $76703 m0 *1 375.06,343
X$76703 194 251 41 22 16 225 OAI21_X4
* cell instance $76704 r0 *1 376.2,343
X$76704 232 16 22 251 BUF_X1
* cell instance $76706 m0 *1 378.1,343
X$76706 202 251 41 22 16 228 OAI21_X4
* cell instance $76710 m0 *1 382.66,343
X$76710 16 1529 229 256 125 22 DFF_X1
* cell instance $76717 r0 *1 384.37,343
X$76717 229 255 178 16 22 233 MUX2_X1
* cell instance $76721 r0 *1 392.92,343
X$76721 266 22 86 16 BUF_X4
* cell instance $76722 r0 *1 394.25,343
X$76722 16 1645 235 234 205 22 DFF_X1
* cell instance $76723 m0 *1 394.82,343
X$76723 235 65 168 16 22 234 MUX2_X1
* cell instance $76728 m0 *1 396.53,343
X$76728 16 1517 204 224 205 22 DFF_X1
* cell instance $76734 r0 *1 398.81,343
X$76734 204 86 235 16 22 527 MUX2_X1
* cell instance $76737 r0 *1 402.04,343
X$76737 16 1641 236 219 205 22 DFF_X1
* cell instance $76738 m0 *1 406.03,343
X$76738 159 16 22 205 CLKBUF_X3
* cell instance $76739 m0 *1 404.7,343
X$76739 236 212 183 16 22 219 MUX2_X1
* cell instance $76742 m0 *1 407.93,343
X$76742 16 1449 237 217 205 22 DFF_X1
* cell instance $76743 m0 *1 411.16,343
X$76743 192 86 237 16 22 207 MUX2_X1
* cell instance $76747 m0 *1 426.17,343
X$76747 159 16 22 213 CLKBUF_X3
* cell instance $76800 r0 *1 405.27,343
X$76800 220 114 236 16 22 448 MUX2_X1
* cell instance $76804 r0 *1 411.92,343
X$76804 239 238 87 16 22 252 MUX2_X1
* cell instance $76805 r0 *1 413.25,343
X$76805 16 1637 239 252 213 22 DFF_X1
* cell instance $76807 r0 *1 417.24,343
X$76807 250 227 87 16 22 248 MUX2_X1
* cell instance $76808 r0 *1 418.57,343
X$76808 16 1638 250 248 213 22 DFF_X1
* cell instance $76812 r0 *1 424.46,343
X$76812 244 181 208 16 22 247 MUX2_X1
* cell instance $76814 r0 *1 426.17,343
X$76814 240 212 208 16 22 245 MUX2_X1
* cell instance $76815 r0 *1 427.5,343
X$76815 16 1544 240 245 213 22 DFF_X1
* cell instance $76819 r0 *1 432.06,343
X$76819 241 212 87 16 22 269 MUX2_X1
* cell instance $77054 r0 *1 356.06,340.2
X$77054 76 197 22 232 16 XOR2_X2
* cell instance $77059 m0 *1 361,340.2
X$77059 16 198 125 154 59 22 DFF_X2
* cell instance $77063 m0 *1 366.51,340.2
X$77063 41 37 23 22 199 16 OAI21_X1
* cell instance $77064 r0 *1 367.27,340.2
X$77064 96 16 22 200 CLKBUF_X3
* cell instance $77065 m0 *1 368.6,340.2
X$77065 125 16 22 1684 INV_X1
* cell instance $77066 m0 *1 367.65,340.2
X$77066 159 16 22 125 CLKBUF_X3
* cell instance $77068 m0 *1 369.74,340.2
X$77068 177 155 80 22 221 16 NOR3_X2
* cell instance $77069 m0 *1 371.07,340.2
X$77069 122 176 131 16 22 NOR2_X4
* cell instance $77071 m0 *1 372.97,340.2
X$77071 177 173 80 22 222 16 NOR3_X2
* cell instance $77073 m0 *1 374.49,340.2
X$77073 16 227 223 130 96 22 AOI21_X4
* cell instance $77075 m0 *1 377.15,340.2
X$77075 80 157 131 22 16 201 AND3_X1
* cell instance $77076 m0 *1 378.1,340.2
X$77076 80 147 131 22 16 203 AND3_X1
* cell instance $77084 r0 *1 374.87,340.2
X$77084 232 16 22 130 INV_X4
* cell instance $77086 r0 *1 377.34,340.2
X$77086 16 238 226 130 79 22 AOI21_X4
* cell instance $77091 r0 *1 384.18,340.2
X$77091 229 88 195 16 22 256 MUX2_X1
* cell instance $77093 m0 *1 384.75,340.2
X$77093 16 1526 178 179 63 22 DFF_X1
* cell instance $77106 r0 *1 397.1,340.2
X$77106 204 54 168 16 22 224 MUX2_X1
* cell instance $77108 m0 *1 404.51,340.2
X$77108 220 181 183 16 22 218 MUX2_X1
* cell instance $77114 r0 *1 404.89,340.2
X$77114 16 1642 220 218 205 22 DFF_X1
* cell instance $77117 m0 *1 413.25,340.2
X$77117 16 1444 182 190 205 22 DFF_X1
* cell instance $77118 m0 *1 410.02,340.2
X$77118 16 1506 192 191 205 22 DFF_X1
* cell instance $77121 r0 *1 410.4,340.2
X$77121 237 65 208 16 22 217 MUX2_X1
* cell instance $77125 r0 *1 414.2,340.2
X$77125 182 86 184 16 22 454 MUX2_X1
* cell instance $77129 m0 *1 422.94,340.2
X$77129 209 88 208 16 22 186 MUX2_X1
* cell instance $77131 m0 *1 425.22,340.2
X$77131 209 114 215 16 22 210 MUX2_X1
* cell instance $77133 m0 *1 427.12,340.2
X$77133 16 1508 215 185 213 22 DFF_X1
* cell instance $77148 r0 *1 430.35,340.2
X$77148 211 181 87 16 22 214 MUX2_X1
* cell instance $77149 r0 *1 431.68,340.2
X$77149 16 1549 211 214 213 22 DFF_X1
* cell instance $77706 r0 *1 351.12,334.6
X$77706 149 139 141 16 22 140 MUX2_X1
* cell instance $77707 m0 *1 352.07,334.6
X$77707 16 1467 105 140 104 22 DFF_X1
* cell instance $77710 r0 *1 352.45,334.6
X$77710 109 122 16 22 141 NOR2_X1
* cell instance $77713 m0 *1 355.68,334.6
X$77713 105 22 122 16 BUF_X4
* cell instance $77716 m0 *1 359.48,334.6
X$77716 152 124 32 22 16 106 HA_X1
* cell instance $77722 r0 *1 357.39,334.6
X$77722 16 123 125 124 127 22 DFF_X2
* cell instance $77726 r0 *1 362.9,334.6
X$77726 124 59 1680 22 16 144 HA_X1
* cell instance $77727 r0 *1 364.8,334.6
X$77727 126 37 79 16 139 22 AOI21_X1
* cell instance $77728 r0 *1 365.56,334.6
X$77728 127 59 80 25 16 22 126 NAND4_X1
* cell instance $77729 r0 *1 366.51,334.6
X$77729 127 59 1679 22 16 107 HA_X1
* cell instance $77730 m0 *1 368.6,334.6
X$77730 107 25 16 22 128 NAND2_X1
* cell instance $77731 m0 *1 367.84,334.6
X$77731 128 37 79 16 108 22 AOI21_X1
* cell instance $77735 m0 *1 373.92,334.6
X$77735 129 107 80 16 22 145 NAND3_X1
* cell instance $77736 m0 *1 374.68,334.6
X$77736 16 65 145 130 96 22 AOI21_X4
* cell instance $77739 m0 *1 378.1,334.6
X$77739 129 157 80 16 22 120 NAND3_X2
* cell instance $77743 r0 *1 370.69,334.6
X$77743 25 122 22 16 129 AND2_X2
* cell instance $77748 r0 *1 377.15,334.6
X$77748 131 144 121 16 22 146 NAND3_X1
* cell instance $77749 r0 *1 377.91,334.6
X$77749 131 147 121 16 22 171 NAND3_X2
* cell instance $77750 r0 *1 379.24,334.6
X$77750 16 134 146 130 79 22 AOI21_X4
* cell instance $77752 m0 *1 379.81,334.6
X$77752 16 54 120 37 79 22 AOI21_X4
* cell instance $77758 r0 *1 382.28,334.6
X$77758 16 88 171 37 79 22 AOI21_X4
* cell instance $77762 r0 *1 386.84,334.6
X$77762 16 1629 132 148 63 22 DFF_X1
* cell instance $77764 m0 *1 387.98,334.6
X$77764 132 134 83 16 22 148 MUX2_X1
* cell instance $77768 m0 *1 400.14,334.6
X$77768 16 1398 135 118 55 22 DFF_X1
* cell instance $77769 m0 *1 403.37,334.6
X$77769 135 134 64 16 22 118 MUX2_X1
* cell instance $77771 m0 *1 407.74,334.6
X$77771 16 1432 111 117 55 22 DFF_X1
* cell instance $77774 m0 *1 411.92,334.6
X$77774 111 86 136 16 22 112 MUX2_X1
* cell instance $77775 m0 *1 413.25,334.6
X$77775 16 1527 136 113 55 22 DFF_X1
* cell instance $77778 m0 *1 418.19,334.6
X$77778 142 134 70 16 22 137 MUX2_X1
* cell instance $77783 r0 *1 390.26,334.6
X$77783 101 86 132 16 22 133 MUX2_X1
* cell instance $77785 r0 *1 392.35,334.6
X$77785 159 16 22 63 CLKBUF_X3
* cell instance $77786 r0 *1 393.3,334.6
X$77786 63 16 22 CLKBUF_X1
* cell instance $77792 r0 *1 401.47,334.6
X$77792 85 86 135 16 22 167 MUX2_X1
* cell instance $77797 r0 *1 418.19,334.6
X$77797 16 1636 142 137 71 22 DFF_X1
* cell instance $77799 m0 *1 423.51,334.6
X$77799 90 114 138 16 22 116 MUX2_X1
* cell instance $77800 m0 *1 422.18,334.6
X$77800 138 134 87 16 22 89 MUX2_X1
* cell instance $77801 m0 *1 424.84,334.6
X$77801 159 16 22 71 CLKBUF_X3
* cell instance $77813 r0 *1 423.7,334.6
X$77813 71 16 22 CLKBUF_X1
* cell instance $77818 r0 *1 427.12,334.6
X$77818 16 1558 160 165 71 22 DFF_X1
* cell instance $77929 m0 *1 5.32,354.2
X$77929 434 16 22 382 BUF_X1
* cell instance $77973 m0 *1 3.61,354.2
X$77973 386 16 22 381 BUF_X1
* cell instance $77979 r0 *1 3.23,354.2
X$77979 456 16 22 427 BUF_X1
* cell instance $78100 r0 *1 2.85,345.8
X$78100 296 16 22 276 BUF_X1
* cell instance $78318 m0 *1 319.77,709.8
X$78318 991 737 16 22 1389 NOR2_X1
* cell instance $78323 m0 *1 336.3,709.8
X$78323 991 343 16 22 1390 NOR2_X1
* cell instance $78367 r0 *1 319.77,709.8
X$78367 1389 16 22 1388 BUF_X1
* cell instance $78372 r0 *1 337.06,709.8
X$78372 1390 16 22 1391 BUF_X1
* cell instance $78379 r0 *1 359.67,709.8
X$78379 737 16 22 1392 BUF_X1
* cell instance $78567 m0 *1 438.14,351.4
X$78567 327 514 362 16 22 364 MUX2_X1
* cell instance $78569 m0 *1 439.47,351.4
X$78569 16 1489 362 364 363 22 DFF_X1
* cell instance $78579 m0 *1 425.6,351.4
X$78579 70 304 361 16 22 360 MUX2_X1
* cell instance $78583 r0 *1 425.6,351.4
X$78583 16 1551 361 360 289 22 DFF_X1
* cell instance $78586 r0 *1 430.73,351.4
X$78586 327 228 404 16 22 458 MUX2_X1
* cell instance $78587 r0 *1 432.06,351.4
X$78587 404 520 326 16 22 365 MUX2_X1
* cell instance $78749 m0 *1 277.78,357
X$78749 492 570 460 16 22 534 MUX2_X1
* cell instance $78751 m0 *1 279.87,357
X$78751 492 430 428 16 22 706 MUX2_X1
* cell instance $78761 r0 *1 277.78,357
X$78761 16 1591 492 534 339 22 DFF_X1
* cell instance $78763 m0 *1 282.53,357
X$78763 431 570 432 16 22 517 MUX2_X1
* cell instance $78765 m0 *1 283.86,357
X$78765 16 1412 431 517 339 22 DFF_X1
* cell instance $78773 r0 *1 289.56,357
X$78773 571 430 383 16 22 614 MUX2_X1
* cell instance $78776 r0 *1 295.45,357
X$78776 16 1619 535 521 536 22 DFF_X1
* cell instance $78778 m0 *1 297.35,357
X$78778 535 466 460 16 22 521 MUX2_X1
* cell instance $78781 m0 *1 300.77,357
X$78781 16 1413 553 467 536 22 DFF_X1
* cell instance $78783 m0 *1 304,357
X$78783 16 524 536 1662 434 22 DFF_X2
* cell instance $78786 r0 *1 304.76,357
X$78786 436 493 554 16 22 524 NAND3_X1
* cell instance $78790 m0 *1 308.75,357
X$78790 311 456 312 16 22 494 NAND3_X1
* cell instance $78792 r0 *1 309.13,357
X$78792 494 469 618 16 22 437 NAND3_X1
* cell instance $78793 m0 *1 310.08,357
X$78793 344 343 150 456 16 22 469 NAND4_X1
* cell instance $78799 m0 *1 316.16,357
X$78799 316 16 22 315 CLKBUF_X3
* cell instance $78801 m0 *1 317.11,357
X$78801 315 16 22 CLKBUF_X1
* cell instance $78804 m0 *1 319.39,357
X$78804 495 466 385 16 22 526 MUX2_X1
* cell instance $78805 m0 *1 320.72,357
X$78805 16 1422 495 526 315 22 DFF_X1
* cell instance $78811 m0 *1 340.86,357
X$78811 316 16 22 348 CLKBUF_X3
* cell instance $78812 m0 *1 341.81,357
X$78812 497 257 22 16 441 AND2_X1
* cell instance $78813 m0 *1 342.57,357
X$78813 348 16 22 1683 INV_X1
* cell instance $78815 m0 *1 343.71,357
X$78815 16 1458 442 481 348 22 DFF_X1
* cell instance $78816 m0 *1 346.94,357
X$78816 442 257 22 16 484 AND2_X1
* cell instance $78817 m0 *1 347.7,357
X$78817 109 442 16 22 483 NOR2_X1
* cell instance $78824 r0 *1 317.11,357
X$78824 538 464 385 16 22 537 MUX2_X1
* cell instance $78826 r0 *1 318.82,357
X$78826 538 430 495 16 22 708 MUX2_X1
* cell instance $78831 r0 *1 332.88,357
X$78831 344 343 345 496 16 22 576 NAND4_X1
* cell instance $78832 r0 *1 333.83,357
X$78832 476 496 312 16 22 654 NAND3_X1
* cell instance $78834 r0 *1 335.35,357
X$78834 16 604 348 1675 496 22 DFF_X2
* cell instance $78837 r0 *1 340.86,357
X$78837 16 560 348 607 497 22 DFF_X2
* cell instance $78846 m0 *1 365.94,357
X$78846 159 16 22 317 CLKBUF_X3
* cell instance $78847 m0 *1 362.33,357
X$78847 16 488 317 1665 19 22 DFF_X2
* cell instance $78848 m0 *1 366.89,357
X$78848 476 19 443 16 22 532 NAND3_X1
* cell instance $78849 m0 *1 367.65,357
X$78849 532 531 529 16 22 488 NAND3_X1
* cell instance $78854 m0 *1 379.81,357
X$78854 16 533 353 1664 542 22 DFF_X2
* cell instance $78857 m0 *1 385.13,357
X$78857 446 445 16 22 530 NOR2_X1
* cell instance $78863 r0 *1 365.75,357
X$78863 200 29 345 21 16 22 579 NAND4_X1
* cell instance $78864 r0 *1 366.7,357
X$78864 317 16 22 CLKBUF_X1
* cell instance $78867 r0 *1 368.98,357
X$78867 200 29 345 18 16 22 539 NAND4_X1
* cell instance $78869 r0 *1 371.45,357
X$78869 200 29 345 540 16 22 625 NAND4_X1
* cell instance $78870 r0 *1 372.4,357
X$78870 476 540 443 16 22 541 NAND3_X1
* cell instance $78871 r0 *1 373.16,357
X$78871 16 563 317 1670 540 22 DFF_X2
* cell instance $78872 r0 *1 376.77,357
X$78872 200 29 311 542 16 22 564 NAND4_X1
* cell instance $78873 r0 *1 377.72,357
X$78873 476 542 443 16 22 565 NAND3_X1
* cell instance $78874 r0 *1 378.48,357
X$78874 565 564 562 16 22 533 NAND3_X1
* cell instance $78878 r0 *1 383.99,357
X$78878 567 530 451 543 628 394 16 22 498 OAI33_X1
* cell instance $78880 r0 *1 386.08,357
X$78880 499 544 16 22 567 NOR2_X1
* cell instance $78885 r0 *1 391.02,357
X$78885 661 227 83 16 22 569 MUX2_X1
* cell instance $78886 m0 *1 391.59,357
X$78886 133 501 16 22 500 NOR2_X1
* cell instance $78890 m0 *1 392.73,357
X$78890 445 16 22 501 CLKBUF_X3
* cell instance $78894 m0 *1 399.95,357
X$78894 527 356 16 22 502 NOR2_X1
* cell instance $78898 r0 *1 392.54,357
X$78898 39 41 662 568 392 529 16 22 OAI221_X2
* cell instance $78900 r0 *1 394.82,357
X$78900 545 544 16 22 546 NOR2_X1
* cell instance $78901 r0 *1 395.39,357
X$78901 394 546 528 451 489 447 16 22 568 OAI33_X1
* cell instance $78903 r0 *1 397.1,357
X$78903 270 501 16 22 632 NOR2_X1
* cell instance $78906 r0 *1 399.38,357
X$78906 394 582 599 451 566 502 16 22 503 OAI33_X1
* cell instance $78907 r0 *1 400.71,357
X$78907 555 501 16 22 528 NOR2_X1
* cell instance $78911 r0 *1 404.89,357
X$78911 394 655 561 451 504 505 16 22 597 OAI33_X1
* cell instance $78913 m0 *1 405.46,357
X$78913 206 356 16 22 505 NOR2_X1
* cell instance $78915 m0 *1 412.3,357
X$78915 207 356 16 22 508 NOR2_X1
* cell instance $78917 m0 *1 415.91,357
X$78917 16 1455 557 509 510 22 DFF_X1
* cell instance $78922 r0 *1 407.74,357
X$78922 394 507 583 451 485 450 16 22 506 OAI33_X1
* cell instance $78924 r0 *1 409.45,357
X$78924 39 41 592 559 392 562 16 22 OAI221_X2
* cell instance $78925 r0 *1 411.54,357
X$78925 547 501 16 22 561 NOR2_X1
* cell instance $78926 r0 *1 412.11,357
X$78926 394 636 593 451 523 508 16 22 559 OAI33_X1
* cell instance $78929 r0 *1 414.01,357
X$78929 558 544 16 22 525 NOR2_X1
* cell instance $78932 r0 *1 415.15,357
X$78932 454 501 16 22 691 NOR2_X1
* cell instance $78934 r0 *1 415.91,357
X$78934 327 254 557 16 22 509 MUX2_X1
* cell instance $78935 r0 *1 417.24,357
X$78935 557 308 585 16 22 558 MUX2_X1
* cell instance $78937 r0 *1 418.76,357
X$78937 327 253 585 16 22 511 MUX2_X1
* cell instance $78940 m0 *1 421.8,357
X$78940 519 522 16 22 403 NOR2_X1
* cell instance $78946 r0 *1 424.08,357
X$78946 548 225 461 16 22 556 MUX2_X1
* cell instance $78949 r0 *1 431.87,357
X$78949 548 228 549 16 22 644 MUX2_X1
* cell instance $78950 r0 *1 433.2,357
X$78950 548 16 22 87 BUF_X2
* cell instance $78951 m0 *1 434.72,357
X$78951 87 332 513 16 22 518 MUX2_X1
* cell instance $78952 m0 *1 433.39,357
X$78952 549 520 513 16 22 519 MUX2_X1
* cell instance $78953 m0 *1 436.05,357
X$78953 16 1454 513 518 363 22 DFF_X1
* cell instance $78957 r0 *1 437,357
X$78957 363 16 22 CLKBUF_X1
* cell instance $78959 m0 *1 441.75,357
X$78959 16 1456 455 516 363 22 DFF_X1
* cell instance $78960 m0 *1 440.42,357
X$78960 327 637 455 16 22 516 MUX2_X1
* cell instance $79059 r0 *1 705.09,357
X$79059 540 16 22 551 BUF_X1
* cell instance $79064 r0 *1 710.03,357
X$79064 496 16 22 552 BUF_X1
* cell instance $79066 r0 *1 710.79,357
X$79066 550 16 22 515 BUF_X1
* cell instance $79110 m0 *1 416.29,382.2
X$79110 879 253 1165 16 22 1168 MUX2_X1
* cell instance $79114 m0 *1 427.69,382.2
X$79114 16 1463 1094 1166 1002 22 DFF_X1
* cell instance $79166 m0 *1 396.15,382.2
X$79166 939 254 1175 16 22 1160 MUX2_X1
* cell instance $79168 m0 *1 399.19,382.2
X$79168 1175 266 1161 16 22 721 MUX2_X1
* cell instance $79173 m0 *1 410.59,382.2
X$79173 16 1472 1164 1172 838 22 DFF_X1
* cell instance $79174 m0 *1 413.82,382.2
X$79174 1164 266 1165 16 22 688 MUX2_X1
* cell instance $79178 r0 *1 396.34,382.2
X$79178 16 1562 1175 1160 1162 22 DFF_X1
* cell instance $79180 r0 *1 402.61,382.2
X$79180 749 16 22 1162 CLKBUF_X3
* cell instance $79181 r0 *1 403.56,382.2
X$79181 1162 16 22 CLKBUF_X1
* cell instance $79183 r0 *1 404.51,382.2
X$79183 999 254 1224 16 22 1226 MUX2_X1
* cell instance $79184 r0 *1 405.84,382.2
X$79184 1224 266 1163 16 22 724 MUX2_X1
* cell instance $79185 r0 *1 407.17,382.2
X$79185 999 253 1163 16 22 1225 MUX2_X1
* cell instance $79186 r0 *1 408.5,382.2
X$79186 16 1597 1163 1225 1162 22 DFF_X1
* cell instance $79190 r0 *1 413.06,382.2
X$79190 879 254 1164 16 22 1172 MUX2_X1
* cell instance $79193 r0 *1 414.96,382.2
X$79193 16 1603 1165 1168 1002 22 DFF_X1
.ENDS bidirectional_fifo

* cell AOI21_X2
* pin A
* pin B2
* pin B1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT AOI21_X2 1 2 3 4 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 4 PWELL,VSS
* net 6 ZN
* net 7 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 7 1 5 7 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 6 2 5 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 5 3 6 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $7 r0 *1 0.21,0.2975 NMOS_VTL
M$7 6 1 4 4 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $9 r0 *1 0.59,0.2975 NMOS_VTL
M$9 9 2 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.78,0.2975 NMOS_VTL
M$10 6 3 9 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.97,0.2975 NMOS_VTL
M$11 8 3 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 1.16,0.2975 NMOS_VTL
M$12 4 2 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI21_X2

* cell NOR2_X4
* pin A2
* pin A1
* pin ZN
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT NOR2_X4 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 ZN
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 9 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 3 2 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 8 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 5 1 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 7 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 3 2 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.35,0.995 PMOS_VTL
M$7 6 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.54,0.995 PMOS_VTL
M$8 5 1 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 0.21,0.2975 NMOS_VTL
M$9 3 1 4 4 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.130725P PS=2.705U
+ PD=2.705U
* device instance $10 r0 *1 0.4,0.2975 NMOS_VTL
M$10 4 2 3 4 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.1162P PS=2.22U PD=2.22U
.ENDS NOR2_X4

* cell AND2_X2
* pin A1
* pin A2
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND2_X2 1 2 4 5 6
* net 1 A1
* net 2 A2
* net 4 NWELL,VDD
* net 5 PWELL,VSS
* net 6 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 3 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 4 2 3 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 7 1 3 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.36,0.2975 NMOS_VTL
M$6 5 2 7 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.55,0.2975 NMOS_VTL
M$7 6 3 5 5 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS AND2_X2

* cell NOR3_X2
* pin A3
* pin A2
* pin A1
* pin NWELL,VDD
* pin ZN
* pin PWELL,VSS
.SUBCKT NOR3_X2 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 NWELL,VDD
* net 5 ZN
* net 6 PWELL,VSS
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 10 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 9 2 10 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 5 3 9 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 8 3 5 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 7 2 8 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 4 1 7 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.21,0.2975 NMOS_VTL
M$7 5 1 6 6 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.072625P PS=1.595U
+ PD=1.595U
* device instance $8 r0 *1 0.4,0.2975 NMOS_VTL
M$8 6 2 5 6 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $9 r0 *1 0.59,0.2975 NMOS_VTL
M$9 5 3 6 6 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
.ENDS NOR3_X2

* cell OAI21_X1
* pin B2
* pin B1
* pin A
* pin NWELL,VDD
* pin ZN
* pin PWELL,VSS
.SUBCKT OAI21_X1 1 2 3 5 6 7
* net 1 B2
* net 2 B1
* net 3 A
* net 5 NWELL,VDD
* net 6 ZN
* net 7 PWELL,VSS
* device instance $1 r0 *1 0.195,0.995 PMOS_VTL
M$1 8 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.385,0.995 PMOS_VTL
M$2 6 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.575,0.995 PMOS_VTL
M$3 5 3 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.195,0.2975 NMOS_VTL
M$4 6 1 4 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.385,0.2975 NMOS_VTL
M$5 4 2 6 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.575,0.2975 NMOS_VTL
M$6 7 3 4 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI21_X1

* cell XNOR2_X2
* pin A
* pin B
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT XNOR2_X2 2 3 4 5 7
* net 2 A
* net 3 B
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 1.135,0.995 PMOS_VTL
M$1 7 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 1.325,0.995 PMOS_VTL
M$2 9 2 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 1.515,0.995 PMOS_VTL
M$3 5 3 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 1.705,0.995 PMOS_VTL
M$4 8 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.18,0.995 PMOS_VTL
M$5 7 1 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $7 r0 *1 0.56,0.995 PMOS_VTL
M$7 1 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 0.75,0.995 PMOS_VTL
M$8 5 2 1 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 1.135,0.2975 NMOS_VTL
M$9 6 2 7 4 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $11 r0 *1 1.515,0.2975 NMOS_VTL
M$11 6 3 7 4 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $13 r0 *1 0.18,0.2975 NMOS_VTL
M$13 6 1 4 4 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $15 r0 *1 0.56,0.2975 NMOS_VTL
M$15 10 3 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 0.75,0.2975 NMOS_VTL
M$16 1 2 10 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS XNOR2_X2

* cell FA_X1
* pin PWELL,VSS
* pin B
* pin CO
* pin S
* pin CI
* pin A
* pin NWELL,VDD
.SUBCKT FA_X1 1 2 3 8 11 12 14
* net 1 PWELL,VSS
* net 2 B
* net 3 CO
* net 8 S
* net 11 CI
* net 12 A
* net 14 NWELL,VDD
* device instance $1 r0 *1 0.385,1.0275 PMOS_VTL
M$1 17 2 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $2 r0 *1 0.575,1.0275 PMOS_VTL
M$2 4 12 17 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.765,1.0275 PMOS_VTL
M$3 15 11 4 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02265P PS=0.455U
+ PD=0.535U
* device instance $4 r0 *1 0.96,1.1025 PMOS_VTL
M$4 14 12 15 14 PMOS_VTL L=0.05U W=0.315U AS=0.02265P AD=0.02205P PS=0.535U
+ PD=0.455U
* device instance $5 r0 *1 1.15,1.1025 PMOS_VTL
M$5 15 2 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.033075P PS=0.455U
+ PD=0.84U
* device instance $6 r0 *1 0.195,0.995 PMOS_VTL
M$6 14 4 3 14 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.033075P PS=1.47U
+ PD=0.77U
* device instance $7 r0 *1 1.49,1.1525 PMOS_VTL
M$7 16 2 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $8 r0 *1 1.68,1.1525 PMOS_VTL
M$8 14 11 16 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $9 r0 *1 1.87,1.1525 PMOS_VTL
M$9 16 12 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $10 r0 *1 2.06,1.1525 PMOS_VTL
M$10 7 4 16 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.023625P PS=0.455U
+ PD=0.465U
* device instance $11 r0 *1 2.26,1.1525 PMOS_VTL
M$11 18 11 7 14 PMOS_VTL L=0.05U W=0.315U AS=0.023625P AD=0.02205P PS=0.465U
+ PD=0.455U
* device instance $12 r0 *1 2.45,1.1525 PMOS_VTL
M$12 19 2 18 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $13 r0 *1 2.64,1.1525 PMOS_VTL
M$13 19 12 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $14 r0 *1 2.83,0.995 PMOS_VTL
M$14 8 7 14 14 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U
+ PD=1.47U
* device instance $15 r0 *1 0.385,0.32 NMOS_VTL
M$15 13 2 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.021875P AD=0.0147P PS=0.555U
+ PD=0.35U
* device instance $16 r0 *1 0.575,0.32 NMOS_VTL
M$16 4 12 13 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $17 r0 *1 0.765,0.32 NMOS_VTL
M$17 5 11 4 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.015225P PS=0.35U
+ PD=0.355U
* device instance $18 r0 *1 0.96,0.32 NMOS_VTL
M$18 1 12 5 1 NMOS_VTL L=0.05U W=0.21U AS=0.015225P AD=0.0147P PS=0.355U
+ PD=0.35U
* device instance $19 r0 *1 1.15,0.32 NMOS_VTL
M$19 5 2 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.02205P PS=0.35U PD=0.63U
* device instance $20 r0 *1 0.195,0.2975 NMOS_VTL
M$20 1 4 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.021875P PS=1.04U
+ PD=0.555U
* device instance $21 r0 *1 1.49,0.195 NMOS_VTL
M$21 6 2 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $22 r0 *1 1.68,0.195 NMOS_VTL
M$22 1 11 6 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $23 r0 *1 1.87,0.195 NMOS_VTL
M$23 6 12 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $24 r0 *1 2.06,0.195 NMOS_VTL
M$24 7 4 6 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.01575P PS=0.35U PD=0.36U
* device instance $25 r0 *1 2.26,0.195 NMOS_VTL
M$25 9 11 7 1 NMOS_VTL L=0.05U W=0.21U AS=0.01575P AD=0.0147P PS=0.36U PD=0.35U
* device instance $26 r0 *1 2.45,0.195 NMOS_VTL
M$26 10 2 9 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $27 r0 *1 2.64,0.195 NMOS_VTL
M$27 1 12 10 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
* device instance $28 r0 *1 2.83,0.2975 NMOS_VTL
M$28 8 7 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS FA_X1

* cell INV_X8
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT INV_X8 1 2 3 4
* net 1 A
* net 2 PWELL,VSS
* net 3 NWELL,VDD
* net 4 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 3 3 PMOS_VTL L=0.05U W=5.04U AS=0.37485P AD=0.37485P PS=6.86U PD=6.86U
* device instance $9 r0 *1 0.17,0.2975 NMOS_VTL
M$9 4 1 2 2 NMOS_VTL L=0.05U W=3.32U AS=0.246925P AD=0.246925P PS=4.925U
+ PD=4.925U
.ENDS INV_X8

* cell AND3_X1
* pin A1
* pin A2
* pin A3
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND3_X1 1 2 3 5 6 7
* net 1 A1
* net 2 A2
* net 3 A3
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 5 1 4 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 4 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 4 3 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 4 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.195 NMOS_VTL
M$5 8 1 4 6 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $6 r0 *1 0.36,0.195 NMOS_VTL
M$6 9 2 8 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $7 r0 *1 0.55,0.195 NMOS_VTL
M$7 6 3 9 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $8 r0 *1 0.74,0.2975 NMOS_VTL
M$8 7 4 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AND3_X1

* cell NAND3_X2
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND3_X2 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 6 1 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.11025P PS=2.24U PD=2.24U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 5 2 6 5 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 6 3 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $7 r0 *1 0.21,0.2975 NMOS_VTL
M$7 10 1 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $8 r0 *1 0.4,0.2975 NMOS_VTL
M$8 9 2 10 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.59,0.2975 NMOS_VTL
M$9 6 3 9 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.78,0.2975 NMOS_VTL
M$10 8 3 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.97,0.2975 NMOS_VTL
M$11 7 2 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 1.16,0.2975 NMOS_VTL
M$12 4 1 7 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND3_X2

* cell AOI21_X4
* pin PWELL,VSS
* pin ZN
* pin A
* pin B2
* pin B1
* pin NWELL,VDD
.SUBCKT AOI21_X4 1 2 3 4 5 11
* net 1 PWELL,VSS
* net 2 ZN
* net 3 A
* net 4 B2
* net 5 B1
* net 11 NWELL,VDD
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 11 3 10 11 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.945,0.995 PMOS_VTL
M$5 2 4 10 11 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $6 r0 *1 1.135,0.995 PMOS_VTL
M$6 10 5 2 11 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.1764P PS=3.08U PD=3.08U
* device instance $13 r0 *1 0.185,0.2975 NMOS_VTL
M$13 2 3 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $17 r0 *1 0.945,0.2975 NMOS_VTL
M$17 8 4 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $18 r0 *1 1.135,0.2975 NMOS_VTL
M$18 2 5 8 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 1.325,0.2975 NMOS_VTL
M$19 9 5 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $20 r0 *1 1.515,0.2975 NMOS_VTL
M$20 1 4 9 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $21 r0 *1 1.705,0.2975 NMOS_VTL
M$21 6 4 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $22 r0 *1 1.895,0.2975 NMOS_VTL
M$22 2 5 6 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $23 r0 *1 2.085,0.2975 NMOS_VTL
M$23 7 5 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $24 r0 *1 2.275,0.2975 NMOS_VTL
M$24 1 4 7 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI21_X4

* cell NAND2_X2
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND2_X2 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.195,0.995 PMOS_VTL
M$1 5 1 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.11025P PS=2.24U PD=2.24U
* device instance $2 r0 *1 0.385,0.995 PMOS_VTL
M$2 4 2 5 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $5 r0 *1 0.195,0.2975 NMOS_VTL
M$5 7 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.385,0.2975 NMOS_VTL
M$6 5 2 7 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.575,0.2975 NMOS_VTL
M$7 6 2 5 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.765,0.2975 NMOS_VTL
M$8 3 1 6 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND2_X2

* cell AOI21_X1
* pin A
* pin B2
* pin B1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT AOI21_X1 1 2 3 4 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 4 PWELL,VSS
* net 6 ZN
* net 7 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 6 2 5 7 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 5 3 6 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 7 1 5 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.21,0.2975 NMOS_VTL
M$4 8 2 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.4,0.2975 NMOS_VTL
M$5 6 3 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.59,0.2975 NMOS_VTL
M$6 4 1 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI21_X1

* cell NAND2_X4
* pin A2
* pin A1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT NAND2_X4 1 2 4 5 6
* net 1 A2
* net 2 A1
* net 4 PWELL,VSS
* net 5 ZN
* net 6 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 5 1 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 5 2 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $9 r0 *1 0.21,0.2975 NMOS_VTL
M$9 4 1 3 4 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $13 r0 *1 0.97,0.2975 NMOS_VTL
M$13 5 2 3 4 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS NAND2_X4

* cell OAI221_X2
* pin C2
* pin C1
* pin B1
* pin B2
* pin A
* pin ZN
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT OAI221_X2 1 2 3 4 5 7 9 10
* net 1 C2
* net 2 C1
* net 3 B1
* net 4 B2
* net 5 A
* net 7 ZN
* net 9 PWELL,VSS
* net 10 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 12 1 10 10 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 7 2 12 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 11 2 7 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 10 1 11 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 7 5 10 10 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 14 3 7 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.35,0.995 PMOS_VTL
M$7 10 4 14 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.54,0.995 PMOS_VTL
M$8 13 4 10 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $9 r0 *1 1.73,0.995 PMOS_VTL
M$9 7 3 13 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $11 r0 *1 0.21,0.2975 NMOS_VTL
M$11 7 1 6 9 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $12 r0 *1 0.4,0.2975 NMOS_VTL
M$12 6 2 7 9 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $15 r0 *1 0.97,0.2975 NMOS_VTL
M$15 8 5 6 9 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $16 r0 *1 1.16,0.2975 NMOS_VTL
M$16 9 3 8 9 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $17 r0 *1 1.35,0.2975 NMOS_VTL
M$17 8 4 9 9 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
.ENDS OAI221_X2

* cell OAI221_X1
* pin B2
* pin B1
* pin A
* pin C2
* pin C1
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT OAI221_X1 1 2 3 4 5 7 8 9
* net 1 B2
* net 2 B1
* net 3 A
* net 4 C2
* net 5 C1
* net 7 NWELL,VDD
* net 8 PWELL,VSS
* net 9 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 12 1 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 9 2 12 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 7 3 9 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 11 4 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 9 5 11 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.17,0.2975 NMOS_VTL
M$6 8 1 6 8 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $7 r0 *1 0.36,0.2975 NMOS_VTL
M$7 6 2 8 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.55,0.2975 NMOS_VTL
M$8 10 3 6 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.74,0.2975 NMOS_VTL
M$9 9 4 10 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.93,0.2975 NMOS_VTL
M$10 10 5 9 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI221_X1

* cell OAI21_X4
* pin A
* pin B2
* pin B1
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT OAI21_X4 1 2 3 5 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 1 5 5 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 11 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 7 3 11 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.31,0.995 PMOS_VTL
M$7 10 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.5,0.995 PMOS_VTL
M$8 5 2 10 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $9 r0 *1 1.69,0.995 PMOS_VTL
M$9 9 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $10 r0 *1 1.88,0.995 PMOS_VTL
M$10 7 3 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $11 r0 *1 2.07,0.995 PMOS_VTL
M$11 8 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $12 r0 *1 2.26,0.995 PMOS_VTL
M$12 5 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $13 r0 *1 0.17,0.2975 NMOS_VTL
M$13 6 1 4 6 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $17 r0 *1 0.93,0.2975 NMOS_VTL
M$17 7 2 4 6 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
* device instance $18 r0 *1 1.12,0.2975 NMOS_VTL
M$18 4 3 7 6 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.1162P PS=2.22U PD=2.22U
.ENDS OAI21_X4

* cell NAND2_X1
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND2_X1 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 5 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 4 2 5 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.185,0.2975 NMOS_VTL
M$3 6 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $4 r0 *1 0.375,0.2975 NMOS_VTL
M$4 5 2 6 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND2_X1

* cell NOR4_X1
* pin A4
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NOR4_X1 1 2 3 4 5 6 7
* net 1 A4
* net 2 A3
* net 3 A2
* net 4 A1
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 10 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 9 2 10 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 8 3 9 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 4 8 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 7 1 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.36,0.2975 NMOS_VTL
M$6 5 2 7 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.55,0.2975 NMOS_VTL
M$7 7 3 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.74,0.2975 NMOS_VTL
M$8 5 4 7 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NOR4_X1

* cell AND4_X1
* pin A1
* pin A2
* pin A3
* pin A4
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND4_X1 1 2 3 4 6 7 8
* net 1 A1
* net 2 A2
* net 3 A3
* net 4 A4
* net 6 NWELL,VDD
* net 7 PWELL,VSS
* net 8 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 5 1 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 6 2 5 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 5 3 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $4 r0 *1 0.74,1.1525 PMOS_VTL
M$4 5 4 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 8 5 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.17,0.195 NMOS_VTL
M$6 10 1 5 7 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $7 r0 *1 0.36,0.195 NMOS_VTL
M$7 11 2 10 7 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $8 r0 *1 0.55,0.195 NMOS_VTL
M$8 9 3 11 7 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $9 r0 *1 0.74,0.195 NMOS_VTL
M$9 7 4 9 7 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $10 r0 *1 0.93,0.2975 NMOS_VTL
M$10 8 5 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AND4_X1

* cell OR4_X1
* pin A1
* pin A2
* pin A3
* pin A4
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR4_X1 1 2 3 4 5 7 8
* net 1 A1
* net 2 A2
* net 3 A3
* net 4 A4
* net 5 PWELL,VSS
* net 7 NWELL,VDD
* net 8 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 10 1 6 7 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 9 2 10 7 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 11 3 9 7 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $4 r0 *1 0.74,1.1525 PMOS_VTL
M$4 11 4 7 7 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 8 6 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.17,0.195 NMOS_VTL
M$6 6 1 5 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $7 r0 *1 0.36,0.195 NMOS_VTL
M$7 5 2 6 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $8 r0 *1 0.55,0.195 NMOS_VTL
M$8 6 3 5 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $9 r0 *1 0.74,0.195 NMOS_VTL
M$9 5 4 6 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $10 r0 *1 0.93,0.2975 NMOS_VTL
M$10 8 6 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OR4_X1

* cell CLKBUF_X2
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT CLKBUF_X2 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.17,0.1875 NMOS_VTL
M$4 3 1 2 3 NMOS_VTL L=0.05U W=0.195U AS=0.020475P AD=0.01365P PS=0.6U PD=0.335U
* device instance $5 r0 *1 0.36,0.1875 NMOS_VTL
M$5 5 2 3 3 NMOS_VTL L=0.05U W=0.39U AS=0.0273P AD=0.034125P PS=0.67U PD=0.935U
.ENDS CLKBUF_X2

* cell BUF_X8
* pin PWELL,VSS
* pin Z
* pin NWELL,VDD
* pin A
.SUBCKT BUF_X8 1 3 4 5
* net 1 PWELL,VSS
* net 3 Z
* net 4 NWELL,VDD
* net 5 A
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 2 5 4 4 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 3 2 4 4 PMOS_VTL L=0.05U W=5.04U AS=0.3528P AD=0.37485P PS=6.16U PD=6.86U
* device instance $13 r0 *1 0.17,0.2975 NMOS_VTL
M$13 2 5 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $17 r0 *1 0.93,0.2975 NMOS_VTL
M$17 3 2 1 1 NMOS_VTL L=0.05U W=3.32U AS=0.2324P AD=0.246925P PS=4.44U PD=4.925U
.ENDS BUF_X8

* cell INV_X4
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT INV_X4 1 2 3 4
* net 1 A
* net 2 PWELL,VSS
* net 3 NWELL,VDD
* net 4 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 3 3 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.19845P PS=3.78U PD=3.78U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 4 1 2 2 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.130725P PS=2.705U
+ PD=2.705U
.ENDS INV_X4

* cell NOR4_X4
* pin PWELL,VSS
* pin A1
* pin A2
* pin A3
* pin A4
* pin ZN
* pin NWELL,VDD
.SUBCKT NOR4_X4 1 2 3 4 5 6 10
* net 1 PWELL,VSS
* net 2 A1
* net 3 A2
* net 4 A3
* net 5 A4
* net 6 ZN
* net 10 NWELL,VDD
* device instance $1 r0 *1 1.92,0.995 PMOS_VTL
M$1 8 4 9 10 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 2.68,0.995 PMOS_VTL
M$5 10 5 9 10 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $9 r0 *1 0.17,0.995 PMOS_VTL
M$9 6 2 7 10 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $13 r0 *1 0.93,0.995 PMOS_VTL
M$13 8 3 7 10 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $17 r0 *1 1.92,0.2975 NMOS_VTL
M$17 1 4 6 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $21 r0 *1 2.68,0.2975 NMOS_VTL
M$21 1 5 6 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
* device instance $25 r0 *1 0.17,0.2975 NMOS_VTL
M$25 6 2 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $29 r0 *1 0.93,0.2975 NMOS_VTL
M$29 6 3 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS NOR4_X4

* cell MUX2_X2
* pin A
* pin B
* pin S
* pin NWELL,VDD
* pin PWELL,VSS
* pin Z
.SUBCKT MUX2_X2 1 2 3 6 7 8
* net 1 A
* net 2 B
* net 3 S
* net 6 NWELL,VDD
* net 7 PWELL,VSS
* net 8 Z
* device instance $1 r0 *1 1.16,0.995 PMOS_VTL
M$1 8 4 6 6 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.077175P PS=2.24U PD=1.54U
* device instance $3 r0 *1 1.54,1.1525 PMOS_VTL
M$3 9 3 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.033075P PS=0.77U
+ PD=0.84U
* device instance $4 r0 *1 0.215,0.995 PMOS_VTL
M$4 6 1 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $5 r0 *1 0.405,0.995 PMOS_VTL
M$5 5 9 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 0.595,0.995 PMOS_VTL
M$6 4 2 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.045675P PS=0.77U PD=0.775U
* device instance $7 r0 *1 0.79,0.995 PMOS_VTL
M$7 5 3 4 6 PMOS_VTL L=0.05U W=0.63U AS=0.045675P AD=0.0693P PS=0.775U PD=1.48U
* device instance $8 r0 *1 1.54,0.195 NMOS_VTL
M$8 9 3 7 7 NMOS_VTL L=0.05U W=0.21U AS=0.021875P AD=0.02205P PS=0.555U PD=0.63U
* device instance $9 r0 *1 1.16,0.2975 NMOS_VTL
M$9 8 4 7 7 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.050925P PS=1.595U
+ PD=1.11U
* device instance $11 r0 *1 0.215,0.2975 NMOS_VTL
M$11 11 1 4 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $12 r0 *1 0.405,0.2975 NMOS_VTL
M$12 7 9 11 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.595,0.2975 NMOS_VTL
M$13 10 2 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.0300875P PS=0.555U
+ PD=0.56U
* device instance $14 r0 *1 0.79,0.2975 NMOS_VTL
M$14 4 3 10 7 NMOS_VTL L=0.05U W=0.415U AS=0.0300875P AD=0.043575P PS=0.56U
+ PD=1.04U
.ENDS MUX2_X2

* cell INV_X2
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT INV_X2 1 2 3 4
* net 1 A
* net 2 PWELL,VSS
* net 3 NWELL,VDD
* net 4 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 4 1 3 3 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.11025P PS=2.24U PD=2.24U
* device instance $3 r0 *1 0.185,0.2975 NMOS_VTL
M$3 4 1 2 2 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.072625P PS=1.595U
+ PD=1.595U
.ENDS INV_X2

* cell OAI33_X1
* pin B3
* pin B2
* pin B1
* pin A1
* pin A2
* pin A3
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OAI33_X1 1 2 3 4 5 6 7 8 10
* net 1 B3
* net 2 B2
* net 3 B1
* net 4 A1
* net 5 A2
* net 6 A3
* net 7 PWELL,VSS
* net 8 NWELL,VDD
* net 10 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 14 1 8 8 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 13 2 14 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.565,0.995 PMOS_VTL
M$3 10 3 13 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.755,0.995 PMOS_VTL
M$4 12 4 10 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.945,0.995 PMOS_VTL
M$5 11 5 12 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.135,0.995 PMOS_VTL
M$6 8 6 11 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.185,0.2975 NMOS_VTL
M$7 9 1 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $8 r0 *1 0.375,0.2975 NMOS_VTL
M$8 7 2 9 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.565,0.2975 NMOS_VTL
M$9 9 3 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.755,0.2975 NMOS_VTL
M$10 10 4 9 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.945,0.2975 NMOS_VTL
M$11 9 5 10 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 1.135,0.2975 NMOS_VTL
M$12 10 6 9 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI33_X1

* cell BUF_X1
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT BUF_X1 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 2 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.033075P PS=0.77U
+ PD=0.84U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.17,0.195 NMOS_VTL
M$3 3 1 2 3 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.021875P PS=0.63U PD=0.555U
* device instance $4 r0 *1 0.36,0.2975 NMOS_VTL
M$4 5 2 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS BUF_X1

* cell CLKBUF_X1
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT CLKBUF_X1 1 3 4
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.19,1.1525 PMOS_VTL
M$1 2 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.033075P PS=0.77U
+ PD=0.84U
* device instance $2 r0 *1 0.38,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.19,0.2075 NMOS_VTL
M$3 3 1 2 3 NMOS_VTL L=0.05U W=0.095U AS=0.009975P AD=0.01015P PS=0.4U PD=0.335U
* device instance $4 r0 *1 0.38,0.2575 NMOS_VTL
M$4 5 2 3 3 NMOS_VTL L=0.05U W=0.195U AS=0.01015P AD=0.020475P PS=0.335U PD=0.6U
.ENDS CLKBUF_X1

* cell DFF_X1
* pin PWELL,VSS
* pin QN
* pin Q
* pin D
* pin CK
* pin NWELL,VDD
.SUBCKT DFF_X1 1 8 9 14 15 16
* net 1 PWELL,VSS
* net 8 QN
* net 9 Q
* net 14 D
* net 15 CK
* net 16 NWELL,VDD
* device instance $1 r0 *1 2.85,0.995 PMOS_VTL
M$1 16 6 8 16 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 3.04,0.995 PMOS_VTL
M$2 9 7 16 16 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.185,0.9425 PMOS_VTL
M$3 16 5 2 16 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.014175P PS=0.84U
+ PD=0.455U
* device instance $4 r0 *1 0.375,1.055 PMOS_VTL
M$4 17 3 16 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.0063P PS=0.455U
+ PD=0.23U
* device instance $5 r0 *1 0.565,1.055 PMOS_VTL
M$5 17 5 4 16 PMOS_VTL L=0.05U W=0.09U AS=0.018075P AD=0.0063P PS=0.565U
+ PD=0.23U
* device instance $6 r0 *1 0.76,0.975 PMOS_VTL
M$6 18 2 4 16 PMOS_VTL L=0.05U W=0.42U AS=0.018075P AD=0.0294P PS=0.565U
+ PD=0.56U
* device instance $7 r0 *1 0.95,0.975 PMOS_VTL
M$7 16 14 18 16 PMOS_VTL L=0.05U W=0.42U AS=0.0294P AD=0.025725P PS=0.56U
+ PD=0.56U
* device instance $8 r0 *1 1.14,1.0275 PMOS_VTL
M$8 3 4 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.025725P AD=0.0567P PS=0.56U
+ PD=0.99U
* device instance $9 r0 *1 1.555,1.0275 PMOS_VTL
M$9 16 15 5 16 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $10 r0 *1 1.745,1.0275 PMOS_VTL
M$10 19 4 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $11 r0 *1 1.935,1.0275 PMOS_VTL
M$11 6 5 19 16 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.014175P PS=0.455U
+ PD=0.455U
* device instance $12 r0 *1 2.125,1.14 PMOS_VTL
M$12 20 2 6 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.006525P PS=0.455U
+ PD=0.235U
* device instance $13 r0 *1 2.32,1.14 PMOS_VTL
M$13 20 7 16 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.006525P PS=0.455U
+ PD=0.235U
* device instance $14 r0 *1 2.51,1.0275 PMOS_VTL
M$14 7 6 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.014175P AD=0.033075P PS=0.455U
+ PD=0.84U
* device instance $15 r0 *1 2.85,0.2975 NMOS_VTL
M$15 1 6 8 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $16 r0 *1 3.04,0.2975 NMOS_VTL
M$16 9 7 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
* device instance $17 r0 *1 2.125,0.345 NMOS_VTL
M$17 12 5 6 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.006525P PS=0.35U
+ PD=0.235U
* device instance $18 r0 *1 2.32,0.345 NMOS_VTL
M$18 12 7 1 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.006525P PS=0.35U
+ PD=0.235U
* device instance $19 r0 *1 1.555,0.36 NMOS_VTL
M$19 1 15 5 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $20 r0 *1 1.745,0.36 NMOS_VTL
M$20 13 4 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $21 r0 *1 1.935,0.36 NMOS_VTL
M$21 6 2 13 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0105P PS=0.35U PD=0.35U
* device instance $22 r0 *1 2.51,0.36 NMOS_VTL
M$22 7 6 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0105P AD=0.02205P PS=0.35U PD=0.63U
* device instance $23 r0 *1 0.185,0.285 NMOS_VTL
M$23 1 5 2 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0105P PS=0.63U PD=0.35U
* device instance $24 r0 *1 0.375,0.345 NMOS_VTL
M$24 10 3 1 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.0063P PS=0.35U PD=0.23U
* device instance $25 r0 *1 0.565,0.345 NMOS_VTL
M$25 10 2 4 1 NMOS_VTL L=0.05U W=0.09U AS=0.013P AD=0.0063P PS=0.42U PD=0.23U
* device instance $26 r0 *1 1.14,0.285 NMOS_VTL
M$26 3 4 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.016975P AD=0.02205P PS=0.415U
+ PD=0.63U
* device instance $27 r0 *1 0.76,0.3175 NMOS_VTL
M$27 11 5 4 1 NMOS_VTL L=0.05U W=0.275U AS=0.013P AD=0.01925P PS=0.42U PD=0.415U
* device instance $28 r0 *1 0.95,0.3175 NMOS_VTL
M$28 1 14 11 1 NMOS_VTL L=0.05U W=0.275U AS=0.01925P AD=0.016975P PS=0.415U
+ PD=0.415U
.ENDS DFF_X1

* cell DFF_X2
* pin PWELL,VSS
* pin D
* pin CK
* pin QN
* pin Q
* pin NWELL,VDD
.SUBCKT DFF_X2 1 6 8 10 11 16
* net 1 PWELL,VSS
* net 6 D
* net 8 CK
* net 10 QN
* net 11 Q
* net 16 NWELL,VDD
* device instance $1 r0 *1 2.855,0.995 PMOS_VTL
M$1 10 9 16 16 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $3 r0 *1 3.235,0.995 PMOS_VTL
M$3 11 2 16 16 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $5 r0 *1 0.2,0.9275 PMOS_VTL
M$5 16 7 3 16 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.014175P PS=0.84U
+ PD=0.455U
* device instance $6 r0 *1 0.39,1.04 PMOS_VTL
M$6 17 4 16 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.0063P PS=0.455U
+ PD=0.23U
* device instance $7 r0 *1 0.58,1.04 PMOS_VTL
M$7 17 7 5 16 PMOS_VTL L=0.05U W=0.09U AS=0.01785P AD=0.0063P PS=0.56U PD=0.23U
* device instance $8 r0 *1 0.77,0.975 PMOS_VTL
M$8 18 3 5 16 PMOS_VTL L=0.05U W=0.42U AS=0.01785P AD=0.0294P PS=0.56U PD=0.56U
* device instance $9 r0 *1 0.96,0.975 PMOS_VTL
M$9 16 6 18 16 PMOS_VTL L=0.05U W=0.42U AS=0.0294P AD=0.025725P PS=0.56U
+ PD=0.56U
* device instance $10 r0 *1 1.15,1.0275 PMOS_VTL
M$10 4 5 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.025725P AD=0.0567P PS=0.56U
+ PD=0.99U
* device instance $11 r0 *1 2.135,0.915 PMOS_VTL
M$11 20 3 9 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.0063P PS=0.455U
+ PD=0.23U
* device instance $12 r0 *1 2.325,0.915 PMOS_VTL
M$12 20 2 16 16 PMOS_VTL L=0.05U W=0.09U AS=0.0252P AD=0.0063P PS=0.77U PD=0.23U
* device instance $13 r0 *1 1.565,1.0275 PMOS_VTL
M$13 16 8 7 16 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $14 r0 *1 1.755,1.0275 PMOS_VTL
M$14 19 5 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $15 r0 *1 1.945,1.0275 PMOS_VTL
M$15 9 7 19 16 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.014175P PS=0.455U
+ PD=0.455U
* device instance $16 r0 *1 2.515,0.995 PMOS_VTL
M$16 2 9 16 16 PMOS_VTL L=0.05U W=0.63U AS=0.0252P AD=0.06615P PS=0.77U PD=1.47U
* device instance $17 r0 *1 2.855,0.2975 NMOS_VTL
M$17 10 9 1 1 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U
+ PD=1.11U
* device instance $19 r0 *1 3.235,0.2975 NMOS_VTL
M$19 11 2 1 1 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U
+ PD=1.595U
* device instance $21 r0 *1 0.39,0.31 NMOS_VTL
M$21 12 4 1 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.0063P PS=0.35U PD=0.23U
* device instance $22 r0 *1 0.58,0.31 NMOS_VTL
M$22 12 3 5 1 NMOS_VTL L=0.05U W=0.09U AS=0.012775P AD=0.0063P PS=0.415U
+ PD=0.23U
* device instance $23 r0 *1 1.15,0.25 NMOS_VTL
M$23 4 5 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.016975P AD=0.02205P PS=0.415U
+ PD=0.63U
* device instance $24 r0 *1 0.77,0.2825 NMOS_VTL
M$24 13 7 5 1 NMOS_VTL L=0.05U W=0.275U AS=0.012775P AD=0.01925P PS=0.415U
+ PD=0.415U
* device instance $25 r0 *1 0.96,0.2825 NMOS_VTL
M$25 1 6 13 1 NMOS_VTL L=0.05U W=0.275U AS=0.01925P AD=0.016975P PS=0.415U
+ PD=0.415U
* device instance $26 r0 *1 0.2,0.37 NMOS_VTL
M$26 1 7 3 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0105P PS=0.63U PD=0.35U
* device instance $27 r0 *1 1.565,0.35 NMOS_VTL
M$27 1 8 7 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $28 r0 *1 1.755,0.35 NMOS_VTL
M$28 14 5 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $29 r0 *1 1.945,0.35 NMOS_VTL
M$29 9 3 14 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0105P PS=0.35U PD=0.35U
* device instance $30 r0 *1 2.135,0.41 NMOS_VTL
M$30 15 7 9 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.0063P PS=0.35U PD=0.23U
* device instance $31 r0 *1 2.325,0.41 NMOS_VTL
M$31 15 2 1 1 NMOS_VTL L=0.05U W=0.09U AS=0.017675P AD=0.0063P PS=0.555U
+ PD=0.23U
* device instance $32 r0 *1 2.515,0.2975 NMOS_VTL
M$32 2 9 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.017675P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS DFF_X2

* cell HA_X1
* pin A
* pin B
* pin S
* pin NWELL,VDD
* pin PWELL,VSS
* pin CO
.SUBCKT HA_X1 1 2 4 5 6 9
* net 1 A
* net 2 B
* net 4 S
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 9 CO
* device instance $1 r0 *1 0.785,1.0275 PMOS_VTL
M$1 10 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.0338625P AD=0.02205P PS=0.775U
+ PD=0.455U
* device instance $2 r0 *1 0.975,1.0275 PMOS_VTL
M$2 7 1 10 5 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.033075P PS=0.455U
+ PD=0.84U
* device instance $3 r0 *1 0.21,0.995 PMOS_VTL
M$3 4 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $4 r0 *1 0.4,0.995 PMOS_VTL
M$4 3 1 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.59,0.995 PMOS_VTL
M$5 5 7 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0338625P PS=0.77U PD=0.775U
* device instance $6 r0 *1 1.345,1.0275 PMOS_VTL
M$6 8 1 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $7 r0 *1 1.535,1.0275 PMOS_VTL
M$7 8 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $8 r0 *1 1.725,0.995 PMOS_VTL
M$8 9 8 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 1.345,0.195 NMOS_VTL
M$9 12 1 8 6 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $10 r0 *1 1.535,0.195 NMOS_VTL
M$10 6 2 12 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
* device instance $11 r0 *1 1.725,0.2975 NMOS_VTL
M$11 9 8 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
* device instance $12 r0 *1 0.785,0.195 NMOS_VTL
M$12 7 2 6 6 NMOS_VTL L=0.05U W=0.21U AS=0.0224P AD=0.0147P PS=0.56U PD=0.35U
* device instance $13 r0 *1 0.975,0.195 NMOS_VTL
M$13 6 1 7 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.02205P PS=0.35U PD=0.63U
* device instance $14 r0 *1 0.21,0.2975 NMOS_VTL
M$14 11 2 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $15 r0 *1 0.4,0.2975 NMOS_VTL
M$15 4 1 11 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 0.59,0.2975 NMOS_VTL
M$16 6 7 4 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.0224P PS=0.555U PD=0.56U
.ENDS HA_X1

* cell CLKBUF_X3
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT CLKBUF_X3 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=1.89U AS=0.1323P AD=0.15435P PS=2.31U PD=3.01U
* device instance $5 r0 *1 0.17,0.1875 NMOS_VTL
M$5 3 1 2 3 NMOS_VTL L=0.05U W=0.195U AS=0.020475P AD=0.01365P PS=0.6U PD=0.335U
* device instance $6 r0 *1 0.36,0.1875 NMOS_VTL
M$6 5 2 3 3 NMOS_VTL L=0.05U W=0.585U AS=0.04095P AD=0.047775P PS=1.005U
+ PD=1.27U
.ENDS CLKBUF_X3

* cell NAND3_X1
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND3_X1 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 6 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.2975 NMOS_VTL
M$4 8 1 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.36,0.2975 NMOS_VTL
M$5 7 2 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 3 7 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND3_X1

* cell BUF_X4
* pin A
* pin NWELL,VDD
* pin Z
* pin PWELL,VSS
.SUBCKT BUF_X4 1 3 4 5
* net 1 A
* net 3 NWELL,VDD
* net 4 Z
* net 5 PWELL,VSS
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 2 1 3 3 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 4 2 3 3 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $7 r0 *1 0.17,0.2975 NMOS_VTL
M$7 2 1 5 5 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $9 r0 *1 0.55,0.2975 NMOS_VTL
M$9 4 2 5 5 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS BUF_X4

* cell NOR2_X1
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NOR2_X1 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 6 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 5 2 6 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.185,0.2975 NMOS_VTL
M$3 5 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $4 r0 *1 0.375,0.2975 NMOS_VTL
M$4 3 2 5 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NOR2_X1

* cell MUX2_X1
* pin A
* pin S
* pin B
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT MUX2_X1 1 2 3 5 6 8
* net 1 A
* net 2 S
* net 3 B
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 8 Z
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 6 2 4 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 9 1 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 7 2 9 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $4 r0 *1 0.74,1.1525 PMOS_VTL
M$4 10 4 7 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $5 r0 *1 0.93,1.1525 PMOS_VTL
M$5 10 3 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 8 7 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.17,0.195 NMOS_VTL
M$7 5 2 4 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $8 r0 *1 0.36,0.195 NMOS_VTL
M$8 12 1 5 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $9 r0 *1 0.55,0.195 NMOS_VTL
M$9 7 4 12 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $10 r0 *1 0.74,0.195 NMOS_VTL
M$10 11 2 7 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $11 r0 *1 0.93,0.195 NMOS_VTL
M$11 5 3 11 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
* device instance $12 r0 *1 1.12,0.2975 NMOS_VTL
M$12 8 7 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS MUX2_X1

* cell NAND4_X1
* pin A4
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND4_X1 1 2 3 4 5 6 7
* net 1 A4
* net 2 A3
* net 3 A2
* net 4 A1
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 6 2 7 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 7 3 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 6 4 7 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 10 1 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.36,0.2975 NMOS_VTL
M$6 9 2 10 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.55,0.2975 NMOS_VTL
M$7 8 3 9 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.74,0.2975 NMOS_VTL
M$8 7 4 8 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND4_X1

* cell XNOR2_X1
* pin A
* pin B
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT XNOR2_X1 1 2 4 5 7
* net 1 A
* net 2 B
* net 4 NWELL,VDD
* net 5 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.18,1.1525 PMOS_VTL
M$1 3 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.37,1.1525 PMOS_VTL
M$2 3 2 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.0338625P AD=0.02205P PS=0.775U
+ PD=0.455U
* device instance $3 r0 *1 0.565,0.995 PMOS_VTL
M$3 7 3 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.0338625P AD=0.0441P PS=0.775U PD=0.77U
* device instance $4 r0 *1 0.755,0.995 PMOS_VTL
M$4 8 1 7 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.945,0.995 PMOS_VTL
M$5 4 2 8 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.18,0.195 NMOS_VTL
M$6 9 1 3 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $7 r0 *1 0.37,0.195 NMOS_VTL
M$7 5 2 9 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0224P PS=0.35U PD=0.56U
* device instance $8 r0 *1 0.565,0.2975 NMOS_VTL
M$8 6 3 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.0224P AD=0.02905P PS=0.56U PD=0.555U
* device instance $9 r0 *1 0.755,0.2975 NMOS_VTL
M$9 7 1 6 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.945,0.2975 NMOS_VTL
M$10 6 2 7 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS XNOR2_X1

* cell XOR2_X2
* pin B
* pin A
* pin NWELL,VDD
* pin Z
* pin PWELL,VSS
.SUBCKT XOR2_X2 1 2 4 5 7
* net 1 B
* net 2 A
* net 4 NWELL,VDD
* net 5 Z
* net 7 PWELL,VSS
* device instance $1 r0 *1 0.2,0.995 PMOS_VTL
M$1 8 2 3 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.39,0.995 PMOS_VTL
M$2 4 1 8 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.58,0.995 PMOS_VTL
M$3 6 3 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.77,0.995 PMOS_VTL
M$4 5 2 6 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $5 r0 *1 0.96,0.995 PMOS_VTL
M$5 6 1 5 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $9 r0 *1 0.2,0.2975 NMOS_VTL
M$9 3 2 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $10 r0 *1 0.39,0.2975 NMOS_VTL
M$10 7 1 3 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.58,0.2975 NMOS_VTL
M$11 5 3 7 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $12 r0 *1 0.77,0.2975 NMOS_VTL
M$12 10 2 5 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.96,0.2975 NMOS_VTL
M$13 7 1 10 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 1.15,0.2975 NMOS_VTL
M$14 9 1 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 1.34,0.2975 NMOS_VTL
M$15 5 2 9 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
.ENDS XOR2_X2

* cell AOI221_X2
* pin B1
* pin B2
* pin A
* pin C2
* pin C1
* pin ZN
* pin NWELL,VDD
* pin PWELL,VSS
.SUBCKT AOI221_X2 1 2 3 4 5 6 8 9
* net 1 B1
* net 2 B2
* net 3 A
* net 4 C2
* net 5 C1
* net 6 ZN
* net 8 NWELL,VDD
* net 9 PWELL,VSS
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 3 10 8 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.09135P PS=2.24U PD=1.55U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 8 1 7 8 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 7 2 8 8 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $7 r0 *1 1.32,0.995 PMOS_VTL
M$7 6 4 10 8 PMOS_VTL L=0.05U W=1.26U AS=0.09135P AD=0.11025P PS=1.55U PD=2.24U
* device instance $8 r0 *1 1.51,0.995 PMOS_VTL
M$8 10 5 6 8 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $11 r0 *1 0.17,0.2975 NMOS_VTL
M$11 6 3 9 9 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.060175P PS=1.595U
+ PD=1.12U
* device instance $12 r0 *1 0.36,0.2975 NMOS_VTL
M$12 14 1 6 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.55,0.2975 NMOS_VTL
M$13 9 2 14 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 0.74,0.2975 NMOS_VTL
M$14 13 2 9 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 0.93,0.2975 NMOS_VTL
M$15 6 1 13 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $17 r0 *1 1.32,0.2975 NMOS_VTL
M$17 12 4 9 9 NMOS_VTL L=0.05U W=0.415U AS=0.031125P AD=0.02905P PS=0.565U
+ PD=0.555U
* device instance $18 r0 *1 1.51,0.2975 NMOS_VTL
M$18 6 5 12 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 1.7,0.2975 NMOS_VTL
M$19 11 5 6 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $20 r0 *1 1.89,0.2975 NMOS_VTL
M$20 9 4 11 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI221_X2

* cell INV_X1
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT INV_X1 1 2 3 4
* net 1 A
* net 2 PWELL,VSS
* net 3 NWELL,VDD
* net 4 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 3 3 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.06615P PS=1.47U PD=1.47U
* device instance $2 r0 *1 0.17,0.2975 NMOS_VTL
M$2 4 1 2 2 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.043575P PS=1.04U
+ PD=1.04U
.ENDS INV_X1

* cell AND2_X1
* pin A1
* pin A2
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND2_X1 1 2 4 5 6
* net 1 A1
* net 2 A2
* net 4 NWELL,VDD
* net 5 PWELL,VSS
* net 6 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 3 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 3 2 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.195 NMOS_VTL
M$4 7 1 3 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $5 r0 *1 0.36,0.195 NMOS_VTL
M$5 5 2 7 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 3 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AND2_X1

* cell BUF_X2
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT BUF_X2 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 4 1 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.21,0.2975 NMOS_VTL
M$4 3 1 2 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.4,0.2975 NMOS_VTL
M$5 5 2 3 3 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS BUF_X2
