module parameterized_barrel_rotator (direction,
    data_in,
    data_out,
    rotate_amount);
 input direction;
 input [31:0] data_in;
 output [31:0] data_out;
 input [4:0] rotate_amount;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;

 sky130_fd_sc_hd__inv_2 _396_ (.A(net34),
    .Y(_369_));
 sky130_fd_sc_hd__clkbuf_4 _397_ (.A(_369_),
    .X(_370_));
 sky130_fd_sc_hd__clkbuf_4 _398_ (.A(_370_),
    .X(_392_));
 sky130_fd_sc_hd__inv_1 _399_ (.A(net35),
    .Y(_393_));
 sky130_fd_sc_hd__inv_1 _400_ (.A(net33),
    .Y(_371_));
 sky130_fd_sc_hd__clkbuf_4 _401_ (.A(_394_),
    .X(_372_));
 sky130_fd_sc_hd__buf_4 _402_ (.A(_395_),
    .X(_373_));
 sky130_fd_sc_hd__nor2_1 _403_ (.A(net35),
    .B(_373_),
    .Y(_374_));
 sky130_fd_sc_hd__o22ai_2 _404_ (.A1(_372_),
    .A2(_373_),
    .B1(_374_),
    .B2(net36),
    .Y(_375_));
 sky130_fd_sc_hd__nor2_1 _405_ (.A(net36),
    .B(_394_),
    .Y(_376_));
 sky130_fd_sc_hd__o21ai_1 _406_ (.A1(_373_),
    .A2(_376_),
    .B1(net35),
    .Y(_377_));
 sky130_fd_sc_hd__inv_2 _407_ (.A(net36),
    .Y(_378_));
 sky130_fd_sc_hd__a31oi_2 _408_ (.A1(_378_),
    .A2(_393_),
    .A3(_369_),
    .B1(_371_),
    .Y(_379_));
 sky130_fd_sc_hd__a41oi_4 _409_ (.A1(_371_),
    .A2(_369_),
    .A3(_375_),
    .A4(_377_),
    .B1(_379_),
    .Y(_380_));
 sky130_fd_sc_hd__xnor2_2 _410_ (.A(net37),
    .B(_380_),
    .Y(_381_));
 sky130_fd_sc_hd__buf_2 _411_ (.A(_381_),
    .X(_382_));
 sky130_fd_sc_hd__nand2b_1 _412_ (.A_N(_394_),
    .B(net33),
    .Y(_383_));
 sky130_fd_sc_hd__clkbuf_4 _413_ (.A(_383_),
    .X(_384_));
 sky130_fd_sc_hd__xnor2_4 _414_ (.A(net36),
    .B(_384_),
    .Y(_385_));
 sky130_fd_sc_hd__buf_4 _415_ (.A(_385_),
    .X(_386_));
 sky130_fd_sc_hd__buf_4 _416_ (.A(net33),
    .X(_387_));
 sky130_fd_sc_hd__or2_2 _417_ (.A(net35),
    .B(net34),
    .X(_388_));
 sky130_fd_sc_hd__clkbuf_4 _418_ (.A(_373_),
    .X(_389_));
 sky130_fd_sc_hd__nor2b_1 _419_ (.A(_389_),
    .B_N(_372_),
    .Y(_390_));
 sky130_fd_sc_hd__or3_1 _420_ (.A(net38),
    .B(net37),
    .C(net36),
    .X(_391_));
 sky130_fd_sc_hd__nor4_4 _421_ (.A(_387_),
    .B(_388_),
    .C(_390_),
    .D(_391_),
    .Y(_000_));
 sky130_fd_sc_hd__nor2_2 _422_ (.A(_386_),
    .B(_000_),
    .Y(_001_));
 sky130_fd_sc_hd__and2b_2 _423_ (.A_N(net33),
    .B(net34),
    .X(_002_));
 sky130_fd_sc_hd__xnor2_4 _424_ (.A(_373_),
    .B(_002_),
    .Y(_003_));
 sky130_fd_sc_hd__buf_4 _425_ (.A(net34),
    .X(_004_));
 sky130_fd_sc_hd__buf_4 _426_ (.A(_004_),
    .X(_005_));
 sky130_fd_sc_hd__mux2i_2 _427_ (.A0(net17),
    .A1(net18),
    .S(_005_),
    .Y(_006_));
 sky130_fd_sc_hd__nand2_1 _428_ (.A(_003_),
    .B(_006_),
    .Y(_007_));
 sky130_fd_sc_hd__nand2b_2 _429_ (.A_N(net33),
    .B(net34),
    .Y(_008_));
 sky130_fd_sc_hd__xnor2_4 _430_ (.A(_373_),
    .B(_008_),
    .Y(_009_));
 sky130_fd_sc_hd__buf_6 _431_ (.A(_009_),
    .X(_010_));
 sky130_fd_sc_hd__buf_4 _432_ (.A(_010_),
    .X(_011_));
 sky130_fd_sc_hd__mux2i_2 _433_ (.A0(net19),
    .A1(net20),
    .S(_004_),
    .Y(_012_));
 sky130_fd_sc_hd__nand2_1 _434_ (.A(_011_),
    .B(_012_),
    .Y(_013_));
 sky130_fd_sc_hd__buf_4 _435_ (.A(_005_),
    .X(_014_));
 sky130_fd_sc_hd__xor2_4 _436_ (.A(net33),
    .B(_373_),
    .X(_015_));
 sky130_fd_sc_hd__nand2_1 _437_ (.A(net22),
    .B(_015_),
    .Y(_016_));
 sky130_fd_sc_hd__xnor2_2 _438_ (.A(_387_),
    .B(_389_),
    .Y(_017_));
 sky130_fd_sc_hd__buf_6 _439_ (.A(_017_),
    .X(_018_));
 sky130_fd_sc_hd__nand2_1 _440_ (.A(net25),
    .B(_018_),
    .Y(_019_));
 sky130_fd_sc_hd__buf_4 _441_ (.A(_389_),
    .X(_020_));
 sky130_fd_sc_hd__buf_4 _442_ (.A(_389_),
    .X(_021_));
 sky130_fd_sc_hd__nor2b_1 _443_ (.A(_021_),
    .B_N(net21),
    .Y(_022_));
 sky130_fd_sc_hd__buf_4 _444_ (.A(_004_),
    .X(_023_));
 sky130_fd_sc_hd__a211oi_2 _445_ (.A1(_020_),
    .A2(net24),
    .B1(_022_),
    .C1(_023_),
    .Y(_024_));
 sky130_fd_sc_hd__a31oi_4 _446_ (.A1(_014_),
    .A2(_016_),
    .A3(_019_),
    .B1(_024_),
    .Y(_025_));
 sky130_fd_sc_hd__buf_4 _447_ (.A(_386_),
    .X(_026_));
 sky130_fd_sc_hd__a32oi_4 _448_ (.A1(_001_),
    .A2(_007_),
    .A3(_013_),
    .B1(_025_),
    .B2(_026_),
    .Y(_027_));
 sky130_fd_sc_hd__mux2i_2 _449_ (.A0(net8),
    .A1(net10),
    .S(_010_),
    .Y(_028_));
 sky130_fd_sc_hd__xnor2_4 _450_ (.A(_378_),
    .B(_384_),
    .Y(_029_));
 sky130_fd_sc_hd__clkbuf_4 _451_ (.A(_029_),
    .X(_030_));
 sky130_fd_sc_hd__clkbuf_4 _452_ (.A(_030_),
    .X(_031_));
 sky130_fd_sc_hd__nand2_1 _453_ (.A(_370_),
    .B(_031_),
    .Y(_032_));
 sky130_fd_sc_hd__nand2_4 _454_ (.A(_023_),
    .B(_030_),
    .Y(_033_));
 sky130_fd_sc_hd__mux2i_4 _455_ (.A0(net9),
    .A1(net11),
    .S(_009_),
    .Y(_034_));
 sky130_fd_sc_hd__o22ai_4 _456_ (.A1(_028_),
    .A2(_032_),
    .B1(_033_),
    .B2(_034_),
    .Y(_035_));
 sky130_fd_sc_hd__mux2i_4 _457_ (.A0(net15),
    .A1(net16),
    .S(_004_),
    .Y(_036_));
 sky130_fd_sc_hd__mux2_1 _458_ (.A0(net13),
    .A1(net14),
    .S(_004_),
    .X(_037_));
 sky130_fd_sc_hd__nor2_1 _459_ (.A(_011_),
    .B(_037_),
    .Y(_038_));
 sky130_fd_sc_hd__a211oi_4 _460_ (.A1(_011_),
    .A2(_036_),
    .B1(_038_),
    .C1(_031_),
    .Y(_039_));
 sky130_fd_sc_hd__nor3_1 _461_ (.A(_382_),
    .B(_035_),
    .C(_039_),
    .Y(_040_));
 sky130_fd_sc_hd__a21oi_1 _462_ (.A1(_382_),
    .A2(_027_),
    .B1(_040_),
    .Y(_041_));
 sky130_fd_sc_hd__buf_2 _463_ (.A(net36),
    .X(_042_));
 sky130_fd_sc_hd__nor2_1 _464_ (.A(net37),
    .B(_042_),
    .Y(_043_));
 sky130_fd_sc_hd__a31oi_2 _465_ (.A1(_378_),
    .A2(_372_),
    .A3(_388_),
    .B1(_387_),
    .Y(_044_));
 sky130_fd_sc_hd__a31oi_4 _466_ (.A1(_387_),
    .A2(_372_),
    .A3(_043_),
    .B1(_044_),
    .Y(_045_));
 sky130_fd_sc_hd__xor2_4 _467_ (.A(net38),
    .B(_045_),
    .X(_046_));
 sky130_fd_sc_hd__mux2i_2 _468_ (.A0(net32),
    .A1(net3),
    .S(_010_),
    .Y(_047_));
 sky130_fd_sc_hd__mux2i_2 _469_ (.A0(net5),
    .A1(net7),
    .S(_009_),
    .Y(_048_));
 sky130_fd_sc_hd__clkbuf_4 _470_ (.A(_385_),
    .X(_049_));
 sky130_fd_sc_hd__mux2i_2 _471_ (.A0(_047_),
    .A1(_048_),
    .S(_049_),
    .Y(_050_));
 sky130_fd_sc_hd__nor2_1 _472_ (.A(_005_),
    .B(_386_),
    .Y(_051_));
 sky130_fd_sc_hd__mux2i_2 _473_ (.A0(net31),
    .A1(net2),
    .S(_009_),
    .Y(_052_));
 sky130_fd_sc_hd__mux2i_1 _474_ (.A0(net4),
    .A1(net6),
    .S(_010_),
    .Y(_053_));
 sky130_fd_sc_hd__nor2_1 _475_ (.A(_023_),
    .B(_030_),
    .Y(_054_));
 sky130_fd_sc_hd__a22oi_1 _476_ (.A1(_051_),
    .A2(_052_),
    .B1(_053_),
    .B2(_054_),
    .Y(_055_));
 sky130_fd_sc_hd__o21ai_2 _477_ (.A1(_392_),
    .A2(_050_),
    .B1(_055_),
    .Y(_056_));
 sky130_fd_sc_hd__mux2i_4 _478_ (.A0(net12),
    .A1(net26),
    .S(_009_),
    .Y(_057_));
 sky130_fd_sc_hd__mux2i_4 _479_ (.A0(net28),
    .A1(net30),
    .S(_009_),
    .Y(_058_));
 sky130_fd_sc_hd__mux2i_1 _480_ (.A0(_057_),
    .A1(_058_),
    .S(_049_),
    .Y(_059_));
 sky130_fd_sc_hd__mux2i_4 _481_ (.A0(net27),
    .A1(net29),
    .S(_009_),
    .Y(_060_));
 sky130_fd_sc_hd__mux2_1 _482_ (.A0(net1),
    .A1(net23),
    .S(_021_),
    .X(_061_));
 sky130_fd_sc_hd__nor2_1 _483_ (.A(_049_),
    .B(_061_),
    .Y(_062_));
 sky130_fd_sc_hd__a21oi_1 _484_ (.A1(_026_),
    .A2(_060_),
    .B1(_062_),
    .Y(_063_));
 sky130_fd_sc_hd__mux2i_1 _485_ (.A0(_059_),
    .A1(_063_),
    .S(_392_),
    .Y(_064_));
 sky130_fd_sc_hd__xor2_4 _486_ (.A(net37),
    .B(_380_),
    .X(_065_));
 sky130_fd_sc_hd__clkbuf_4 _487_ (.A(_065_),
    .X(_066_));
 sky130_fd_sc_hd__mux2i_1 _488_ (.A0(_056_),
    .A1(_064_),
    .S(_066_),
    .Y(_067_));
 sky130_fd_sc_hd__nor2_1 _489_ (.A(_000_),
    .B(_046_),
    .Y(_068_));
 sky130_fd_sc_hd__a22o_1 _490_ (.A1(_041_),
    .A2(_046_),
    .B1(_067_),
    .B2(_068_),
    .X(net39));
 sky130_fd_sc_hd__xnor2_1 _491_ (.A(net38),
    .B(_045_),
    .Y(_069_));
 sky130_fd_sc_hd__clkbuf_4 _492_ (.A(_069_),
    .X(_070_));
 sky130_fd_sc_hd__buf_2 _493_ (.A(_070_),
    .X(_071_));
 sky130_fd_sc_hd__mux2i_2 _494_ (.A0(net23),
    .A1(net27),
    .S(_009_),
    .Y(_072_));
 sky130_fd_sc_hd__nand2_1 _495_ (.A(_389_),
    .B(net31),
    .Y(_073_));
 sky130_fd_sc_hd__nand2b_1 _496_ (.A_N(_373_),
    .B(net29),
    .Y(_074_));
 sky130_fd_sc_hd__a21oi_1 _497_ (.A1(_073_),
    .A2(_074_),
    .B1(_002_),
    .Y(_075_));
 sky130_fd_sc_hd__nand2b_1 _498_ (.A_N(_373_),
    .B(net31),
    .Y(_076_));
 sky130_fd_sc_hd__nand2_1 _499_ (.A(_389_),
    .B(net29),
    .Y(_077_));
 sky130_fd_sc_hd__a21oi_1 _500_ (.A1(_076_),
    .A2(_077_),
    .B1(_008_),
    .Y(_078_));
 sky130_fd_sc_hd__nor2_1 _501_ (.A(_075_),
    .B(_078_),
    .Y(_079_));
 sky130_fd_sc_hd__mux2i_4 _502_ (.A0(net26),
    .A1(net28),
    .S(_009_),
    .Y(_080_));
 sky130_fd_sc_hd__mux2i_4 _503_ (.A0(net30),
    .A1(net32),
    .S(_009_),
    .Y(_081_));
 sky130_fd_sc_hd__clkbuf_4 _504_ (.A(_023_),
    .X(_082_));
 sky130_fd_sc_hd__mux4_1 _505_ (.A0(_072_),
    .A1(_079_),
    .A2(_080_),
    .A3(_081_),
    .S0(_386_),
    .S1(_082_),
    .X(_083_));
 sky130_fd_sc_hd__or2_0 _506_ (.A(_388_),
    .B(_391_),
    .X(_084_));
 sky130_fd_sc_hd__or3_1 _507_ (.A(_387_),
    .B(_390_),
    .C(_084_),
    .X(_085_));
 sky130_fd_sc_hd__clkbuf_4 _508_ (.A(_085_),
    .X(_086_));
 sky130_fd_sc_hd__nand2_1 _509_ (.A(_381_),
    .B(_086_),
    .Y(_087_));
 sky130_fd_sc_hd__mux2i_1 _510_ (.A0(net21),
    .A1(net22),
    .S(_005_),
    .Y(_088_));
 sky130_fd_sc_hd__mux2i_2 _511_ (.A0(_012_),
    .A1(_088_),
    .S(_010_),
    .Y(_089_));
 sky130_fd_sc_hd__or2_0 _512_ (.A(_049_),
    .B(_089_),
    .X(_090_));
 sky130_fd_sc_hd__nor2_1 _513_ (.A(_388_),
    .B(_391_),
    .Y(_091_));
 sky130_fd_sc_hd__or3_1 _514_ (.A(_387_),
    .B(net34),
    .C(_389_),
    .X(_092_));
 sky130_fd_sc_hd__nand3b_1 _515_ (.A_N(_092_),
    .B(_393_),
    .C(_372_),
    .Y(_093_));
 sky130_fd_sc_hd__nand3b_1 _516_ (.A_N(_042_),
    .B(net35),
    .C(_372_),
    .Y(_094_));
 sky130_fd_sc_hd__nand2b_1 _517_ (.A_N(_372_),
    .B(_042_),
    .Y(_095_));
 sky130_fd_sc_hd__nand2_1 _518_ (.A(net38),
    .B(net37),
    .Y(_096_));
 sky130_fd_sc_hd__a211oi_2 _519_ (.A1(_094_),
    .A2(_095_),
    .B1(_096_),
    .C1(_092_),
    .Y(_097_));
 sky130_fd_sc_hd__a21oi_2 _520_ (.A1(_091_),
    .A2(_093_),
    .B1(_097_),
    .Y(_098_));
 sky130_fd_sc_hd__clkbuf_4 _521_ (.A(_098_),
    .X(_099_));
 sky130_fd_sc_hd__buf_4 _522_ (.A(_030_),
    .X(_100_));
 sky130_fd_sc_hd__inv_1 _523_ (.A(net24),
    .Y(_101_));
 sky130_fd_sc_hd__nand2_1 _524_ (.A(_023_),
    .B(net25),
    .Y(_102_));
 sky130_fd_sc_hd__o32ai_1 _525_ (.A1(_023_),
    .A2(_020_),
    .A3(_101_),
    .B1(_018_),
    .B2(_102_),
    .Y(_103_));
 sky130_fd_sc_hd__o21ai_0 _526_ (.A1(_100_),
    .A2(_103_),
    .B1(_086_),
    .Y(_104_));
 sky130_fd_sc_hd__mux2i_1 _527_ (.A0(net12),
    .A1(net25),
    .S(_015_),
    .Y(_105_));
 sky130_fd_sc_hd__mux2_1 _528_ (.A0(net24),
    .A1(net1),
    .S(_389_),
    .X(_106_));
 sky130_fd_sc_hd__nor2_1 _529_ (.A(_023_),
    .B(_106_),
    .Y(_107_));
 sky130_fd_sc_hd__a21oi_1 _530_ (.A1(_082_),
    .A2(_105_),
    .B1(_107_),
    .Y(_108_));
 sky130_fd_sc_hd__o21ai_0 _531_ (.A1(_100_),
    .A2(_108_),
    .B1(_098_),
    .Y(_109_));
 sky130_fd_sc_hd__o22ai_1 _532_ (.A1(_099_),
    .A2(_104_),
    .B1(_109_),
    .B2(_382_),
    .Y(_110_));
 sky130_fd_sc_hd__a2bb2oi_1 _533_ (.A1_N(_083_),
    .A2_N(_087_),
    .B1(_090_),
    .B2(_110_),
    .Y(_111_));
 sky130_fd_sc_hd__buf_2 _534_ (.A(_065_),
    .X(_112_));
 sky130_fd_sc_hd__mux2i_4 _535_ (.A0(net11),
    .A1(net14),
    .S(_018_),
    .Y(_113_));
 sky130_fd_sc_hd__mux2i_1 _536_ (.A0(net10),
    .A1(net13),
    .S(_020_),
    .Y(_114_));
 sky130_fd_sc_hd__mux2i_1 _537_ (.A0(_113_),
    .A1(_114_),
    .S(_370_),
    .Y(_115_));
 sky130_fd_sc_hd__nor3_1 _538_ (.A(_030_),
    .B(_011_),
    .C(_036_),
    .Y(_116_));
 sky130_fd_sc_hd__a21oi_1 _539_ (.A1(_100_),
    .A2(_115_),
    .B1(_116_),
    .Y(_117_));
 sky130_fd_sc_hd__nor2_1 _540_ (.A(_031_),
    .B(_006_),
    .Y(_118_));
 sky130_fd_sc_hd__nand2_1 _541_ (.A(_011_),
    .B(_118_),
    .Y(_119_));
 sky130_fd_sc_hd__o21ai_1 _542_ (.A1(_000_),
    .A2(_117_),
    .B1(_119_),
    .Y(_120_));
 sky130_fd_sc_hd__nand2b_1 _543_ (.A_N(_021_),
    .B(net2),
    .Y(_121_));
 sky130_fd_sc_hd__nand2_1 _544_ (.A(_020_),
    .B(net4),
    .Y(_122_));
 sky130_fd_sc_hd__and2_0 _545_ (.A(_121_),
    .B(_122_),
    .X(_123_));
 sky130_fd_sc_hd__mux2i_1 _546_ (.A0(net6),
    .A1(net8),
    .S(_020_),
    .Y(_124_));
 sky130_fd_sc_hd__mux2i_1 _547_ (.A0(_123_),
    .A1(_124_),
    .S(_049_),
    .Y(_125_));
 sky130_fd_sc_hd__mux2_1 _548_ (.A0(net7),
    .A1(net9),
    .S(_018_),
    .X(_126_));
 sky130_fd_sc_hd__nor2_2 _549_ (.A(_369_),
    .B(_029_),
    .Y(_127_));
 sky130_fd_sc_hd__mux2i_4 _550_ (.A0(net3),
    .A1(net5),
    .S(_018_),
    .Y(_128_));
 sky130_fd_sc_hd__nor3_1 _551_ (.A(_392_),
    .B(_026_),
    .C(_128_),
    .Y(_129_));
 sky130_fd_sc_hd__a221oi_2 _552_ (.A1(_392_),
    .A2(_125_),
    .B1(_126_),
    .B2(_127_),
    .C1(_129_),
    .Y(_130_));
 sky130_fd_sc_hd__o21ai_0 _553_ (.A1(_000_),
    .A2(_130_),
    .B1(_112_),
    .Y(_131_));
 sky130_fd_sc_hd__o211ai_1 _554_ (.A1(_112_),
    .A2(_120_),
    .B1(_131_),
    .C1(_071_),
    .Y(_132_));
 sky130_fd_sc_hd__o21ai_0 _555_ (.A1(_071_),
    .A2(_111_),
    .B1(_132_),
    .Y(net40));
 sky130_fd_sc_hd__clkbuf_4 _556_ (.A(_381_),
    .X(_133_));
 sky130_fd_sc_hd__nand3_1 _557_ (.A(_082_),
    .B(_031_),
    .C(_060_),
    .Y(_134_));
 sky130_fd_sc_hd__nand2_1 _558_ (.A(_127_),
    .B(_052_),
    .Y(_135_));
 sky130_fd_sc_hd__a22oi_1 _559_ (.A1(_051_),
    .A2(_080_),
    .B1(_081_),
    .B2(_054_),
    .Y(_136_));
 sky130_fd_sc_hd__and3_1 _560_ (.A(_134_),
    .B(_135_),
    .C(_136_),
    .X(_137_));
 sky130_fd_sc_hd__mux2_1 _561_ (.A0(net20),
    .A1(net22),
    .S(_021_),
    .X(_138_));
 sky130_fd_sc_hd__nand2_1 _562_ (.A(_030_),
    .B(_138_),
    .Y(_139_));
 sky130_fd_sc_hd__nor2b_1 _563_ (.A(_389_),
    .B_N(net25),
    .Y(_140_));
 sky130_fd_sc_hd__a21o_1 _564_ (.A1(_020_),
    .A2(net12),
    .B1(_140_),
    .X(_141_));
 sky130_fd_sc_hd__nand2_1 _565_ (.A(_049_),
    .B(_141_),
    .Y(_142_));
 sky130_fd_sc_hd__a21oi_1 _566_ (.A1(_139_),
    .A2(_142_),
    .B1(_082_),
    .Y(_143_));
 sky130_fd_sc_hd__mux2i_1 _567_ (.A0(net21),
    .A1(net24),
    .S(_010_),
    .Y(_144_));
 sky130_fd_sc_hd__mux2i_2 _568_ (.A0(net1),
    .A1(net23),
    .S(_018_),
    .Y(_145_));
 sky130_fd_sc_hd__nand2_4 _569_ (.A(_023_),
    .B(_386_),
    .Y(_146_));
 sky130_fd_sc_hd__o22ai_1 _570_ (.A1(_033_),
    .A2(_144_),
    .B1(_145_),
    .B2(_146_),
    .Y(_147_));
 sky130_fd_sc_hd__clkbuf_4 _571_ (.A(_065_),
    .X(_148_));
 sky130_fd_sc_hd__o21a_1 _572_ (.A1(_143_),
    .A2(_147_),
    .B1(_148_),
    .X(_149_));
 sky130_fd_sc_hd__a21o_1 _573_ (.A1(_091_),
    .A2(_093_),
    .B1(_097_),
    .X(_150_));
 sky130_fd_sc_hd__clkbuf_4 _574_ (.A(_150_),
    .X(_151_));
 sky130_fd_sc_hd__a211oi_1 _575_ (.A1(_133_),
    .A2(_137_),
    .B1(_149_),
    .C1(_151_),
    .Y(_152_));
 sky130_fd_sc_hd__clkbuf_4 _576_ (.A(_046_),
    .X(_153_));
 sky130_fd_sc_hd__mux2i_1 _577_ (.A0(_138_),
    .A1(_140_),
    .S(_386_),
    .Y(_154_));
 sky130_fd_sc_hd__o22ai_1 _578_ (.A1(_033_),
    .A2(_144_),
    .B1(_154_),
    .B2(_082_),
    .Y(_155_));
 sky130_fd_sc_hd__nor3_2 _579_ (.A(_387_),
    .B(_372_),
    .C(_084_),
    .Y(_156_));
 sky130_fd_sc_hd__a211o_1 _580_ (.A1(_148_),
    .A2(_155_),
    .B1(_156_),
    .C1(_099_),
    .X(_157_));
 sky130_fd_sc_hd__nand2_1 _581_ (.A(_153_),
    .B(_157_),
    .Y(_158_));
 sky130_fd_sc_hd__mux2i_2 _582_ (.A0(net4),
    .A1(net8),
    .S(_385_),
    .Y(_159_));
 sky130_fd_sc_hd__mux2i_1 _583_ (.A0(net5),
    .A1(net9),
    .S(_386_),
    .Y(_160_));
 sky130_fd_sc_hd__nor2b_1 _584_ (.A(_004_),
    .B_N(_021_),
    .Y(_161_));
 sky130_fd_sc_hd__a32oi_1 _585_ (.A1(_014_),
    .A2(_003_),
    .A3(_159_),
    .B1(_160_),
    .B2(_161_),
    .Y(_162_));
 sky130_fd_sc_hd__nand3_1 _586_ (.A(_387_),
    .B(_372_),
    .C(_020_),
    .Y(_163_));
 sky130_fd_sc_hd__o21ai_0 _587_ (.A1(_387_),
    .A2(_020_),
    .B1(_163_),
    .Y(_164_));
 sky130_fd_sc_hd__mux2i_1 _588_ (.A0(net6),
    .A1(net10),
    .S(_042_),
    .Y(_165_));
 sky130_fd_sc_hd__and2_0 _589_ (.A(_042_),
    .B(net6),
    .X(_166_));
 sky130_fd_sc_hd__nand2_1 _590_ (.A(_005_),
    .B(_020_),
    .Y(_167_));
 sky130_fd_sc_hd__a2111oi_0 _591_ (.A1(_378_),
    .A2(net10),
    .B1(_384_),
    .C1(_166_),
    .D1(_167_),
    .Y(_168_));
 sky130_fd_sc_hd__a31oi_1 _592_ (.A1(_014_),
    .A2(_164_),
    .A3(_165_),
    .B1(_168_),
    .Y(_169_));
 sky130_fd_sc_hd__nor2_2 _593_ (.A(_004_),
    .B(_021_),
    .Y(_170_));
 sky130_fd_sc_hd__nand2_1 _594_ (.A(net3),
    .B(_030_),
    .Y(_171_));
 sky130_fd_sc_hd__nand2_1 _595_ (.A(net7),
    .B(_049_),
    .Y(_172_));
 sky130_fd_sc_hd__nand3_1 _596_ (.A(_170_),
    .B(_171_),
    .C(_172_),
    .Y(_173_));
 sky130_fd_sc_hd__and3_1 _597_ (.A(_162_),
    .B(_169_),
    .C(_173_),
    .X(_174_));
 sky130_fd_sc_hd__mux2i_4 _598_ (.A0(net16),
    .A1(net17),
    .S(_005_),
    .Y(_175_));
 sky130_fd_sc_hd__mux2i_2 _599_ (.A0(net18),
    .A1(net19),
    .S(_005_),
    .Y(_176_));
 sky130_fd_sc_hd__mux2i_4 _600_ (.A0(_175_),
    .A1(_176_),
    .S(_010_),
    .Y(_177_));
 sky130_fd_sc_hd__mux2i_2 _601_ (.A0(net11),
    .A1(net13),
    .S(_004_),
    .Y(_178_));
 sky130_fd_sc_hd__mux2i_2 _602_ (.A0(net14),
    .A1(net15),
    .S(_004_),
    .Y(_179_));
 sky130_fd_sc_hd__mux2i_1 _603_ (.A0(_178_),
    .A1(_179_),
    .S(_010_),
    .Y(_180_));
 sky130_fd_sc_hd__mux2i_2 _604_ (.A0(_177_),
    .A1(_180_),
    .S(_031_),
    .Y(_181_));
 sky130_fd_sc_hd__nor3_1 _605_ (.A(_148_),
    .B(_000_),
    .C(_181_),
    .Y(_182_));
 sky130_fd_sc_hd__a21oi_1 _606_ (.A1(_112_),
    .A2(_174_),
    .B1(_182_),
    .Y(_183_));
 sky130_fd_sc_hd__o22ai_1 _607_ (.A1(_152_),
    .A2(_158_),
    .B1(_183_),
    .B2(_153_),
    .Y(net41));
 sky130_fd_sc_hd__a21oi_1 _608_ (.A1(_001_),
    .A2(_037_),
    .B1(_118_),
    .Y(_184_));
 sky130_fd_sc_hd__nand2_1 _609_ (.A(_031_),
    .B(_036_),
    .Y(_185_));
 sky130_fd_sc_hd__nand2_1 _610_ (.A(_026_),
    .B(_012_),
    .Y(_186_));
 sky130_fd_sc_hd__a31oi_1 _611_ (.A1(_086_),
    .A2(_185_),
    .A3(_186_),
    .B1(_003_),
    .Y(_187_));
 sky130_fd_sc_hd__a21oi_1 _612_ (.A1(_003_),
    .A2(_184_),
    .B1(_187_),
    .Y(_188_));
 sky130_fd_sc_hd__mux4_2 _613_ (.A0(_034_),
    .A1(_028_),
    .A2(_048_),
    .A3(_053_),
    .S0(_369_),
    .S1(_031_),
    .X(_189_));
 sky130_fd_sc_hd__nand2_1 _614_ (.A(_066_),
    .B(_189_),
    .Y(_190_));
 sky130_fd_sc_hd__o21ai_0 _615_ (.A1(_066_),
    .A2(_188_),
    .B1(_190_),
    .Y(_191_));
 sky130_fd_sc_hd__nand2_4 _616_ (.A(_046_),
    .B(_099_),
    .Y(_192_));
 sky130_fd_sc_hd__mux4_1 _617_ (.A0(_047_),
    .A1(_052_),
    .A2(_058_),
    .A3(_060_),
    .S0(_370_),
    .S1(_031_),
    .X(_193_));
 sky130_fd_sc_hd__o21ai_0 _618_ (.A1(_014_),
    .A2(_061_),
    .B1(_026_),
    .Y(_194_));
 sky130_fd_sc_hd__a21o_1 _619_ (.A1(_082_),
    .A2(_057_),
    .B1(_194_),
    .X(_195_));
 sky130_fd_sc_hd__nand2_1 _620_ (.A(_001_),
    .B(_025_),
    .Y(_196_));
 sky130_fd_sc_hd__nand2_1 _621_ (.A(_195_),
    .B(_196_),
    .Y(_197_));
 sky130_fd_sc_hd__a2bb2oi_1 _622_ (.A1_N(_087_),
    .A2_N(_193_),
    .B1(_197_),
    .B2(_112_),
    .Y(_198_));
 sky130_fd_sc_hd__o22ai_1 _623_ (.A1(_153_),
    .A2(_191_),
    .B1(_192_),
    .B2(_198_),
    .Y(net42));
 sky130_fd_sc_hd__mux2i_4 _624_ (.A0(_175_),
    .A1(_179_),
    .S(_003_),
    .Y(_199_));
 sky130_fd_sc_hd__mux2i_4 _625_ (.A0(net18),
    .A1(net20),
    .S(_021_),
    .Y(_200_));
 sky130_fd_sc_hd__mux2i_2 _626_ (.A0(net19),
    .A1(net21),
    .S(_017_),
    .Y(_201_));
 sky130_fd_sc_hd__mux2i_4 _627_ (.A0(_200_),
    .A1(_201_),
    .S(_023_),
    .Y(_202_));
 sky130_fd_sc_hd__mux2i_2 _628_ (.A0(_199_),
    .A1(_202_),
    .S(_026_),
    .Y(_203_));
 sky130_fd_sc_hd__mux2i_1 _629_ (.A0(net10),
    .A1(net13),
    .S(_010_),
    .Y(_204_));
 sky130_fd_sc_hd__mux2i_1 _630_ (.A0(net6),
    .A1(net8),
    .S(_010_),
    .Y(_205_));
 sky130_fd_sc_hd__mux4_2 _631_ (.A0(_034_),
    .A1(_048_),
    .A2(_204_),
    .A3(_205_),
    .S0(_029_),
    .S1(_082_),
    .X(_206_));
 sky130_fd_sc_hd__mux2i_2 _632_ (.A0(_203_),
    .A1(_206_),
    .S(_148_),
    .Y(_207_));
 sky130_fd_sc_hd__nand2_1 _633_ (.A(net32),
    .B(_170_),
    .Y(_208_));
 sky130_fd_sc_hd__nand2_1 _634_ (.A(net28),
    .B(_170_),
    .Y(_209_));
 sky130_fd_sc_hd__mux2_1 _635_ (.A0(_208_),
    .A1(_209_),
    .S(_029_),
    .X(_210_));
 sky130_fd_sc_hd__o211ai_1 _636_ (.A1(_075_),
    .A2(_078_),
    .B1(_014_),
    .C1(_031_),
    .Y(_211_));
 sky130_fd_sc_hd__nand2_1 _637_ (.A(_042_),
    .B(net3),
    .Y(_212_));
 sky130_fd_sc_hd__nand2b_1 _638_ (.A_N(_042_),
    .B(net30),
    .Y(_213_));
 sky130_fd_sc_hd__a21boi_0 _639_ (.A1(_212_),
    .A2(_213_),
    .B1_N(_384_),
    .Y(_214_));
 sky130_fd_sc_hd__nand2b_1 _640_ (.A_N(_042_),
    .B(net3),
    .Y(_215_));
 sky130_fd_sc_hd__nand2_1 _641_ (.A(_042_),
    .B(net30),
    .Y(_216_));
 sky130_fd_sc_hd__a21oi_1 _642_ (.A1(_215_),
    .A2(_216_),
    .B1(_384_),
    .Y(_217_));
 sky130_fd_sc_hd__o21ai_0 _643_ (.A1(_214_),
    .A2(_217_),
    .B1(_161_),
    .Y(_218_));
 sky130_fd_sc_hd__a21oi_1 _644_ (.A1(_121_),
    .A2(_122_),
    .B1(_002_),
    .Y(_219_));
 sky130_fd_sc_hd__nand2_1 _645_ (.A(_020_),
    .B(net2),
    .Y(_220_));
 sky130_fd_sc_hd__nand2b_1 _646_ (.A_N(_021_),
    .B(net4),
    .Y(_221_));
 sky130_fd_sc_hd__a21oi_1 _647_ (.A1(_220_),
    .A2(_221_),
    .B1(_008_),
    .Y(_222_));
 sky130_fd_sc_hd__o211ai_1 _648_ (.A1(_219_),
    .A2(_222_),
    .B1(_023_),
    .C1(_049_),
    .Y(_223_));
 sky130_fd_sc_hd__nand4_2 _649_ (.A(_210_),
    .B(_211_),
    .C(_218_),
    .D(_223_),
    .Y(_224_));
 sky130_fd_sc_hd__mux2i_4 _650_ (.A0(net23),
    .A1(net27),
    .S(_018_),
    .Y(_225_));
 sky130_fd_sc_hd__mux2i_4 _651_ (.A0(net22),
    .A1(net25),
    .S(_021_),
    .Y(_226_));
 sky130_fd_sc_hd__mux2i_1 _652_ (.A0(net12),
    .A1(net26),
    .S(_021_),
    .Y(_227_));
 sky130_fd_sc_hd__mux2_1 _653_ (.A0(_226_),
    .A1(_227_),
    .S(_385_),
    .X(_228_));
 sky130_fd_sc_hd__mux2_1 _654_ (.A0(net1),
    .A1(net24),
    .S(_015_),
    .X(_229_));
 sky130_fd_sc_hd__nand3_1 _655_ (.A(_014_),
    .B(_030_),
    .C(_229_),
    .Y(_230_));
 sky130_fd_sc_hd__o221ai_4 _656_ (.A1(_146_),
    .A2(_225_),
    .B1(_228_),
    .B2(_014_),
    .C1(_230_),
    .Y(_231_));
 sky130_fd_sc_hd__mux2_1 _657_ (.A0(_224_),
    .A1(_231_),
    .S(_065_),
    .X(_232_));
 sky130_fd_sc_hd__nor2_4 _658_ (.A(_070_),
    .B(_151_),
    .Y(_233_));
 sky130_fd_sc_hd__a22oi_1 _659_ (.A1(_070_),
    .A2(_207_),
    .B1(_232_),
    .B2(_233_),
    .Y(_234_));
 sky130_fd_sc_hd__nor2_1 _660_ (.A(_000_),
    .B(_234_),
    .Y(net43));
 sky130_fd_sc_hd__nand2_1 _661_ (.A(_003_),
    .B(_036_),
    .Y(_235_));
 sky130_fd_sc_hd__nand2_1 _662_ (.A(_011_),
    .B(_006_),
    .Y(_236_));
 sky130_fd_sc_hd__a32o_1 _663_ (.A1(_001_),
    .A2(_235_),
    .A3(_236_),
    .B1(_089_),
    .B2(_026_),
    .X(_237_));
 sky130_fd_sc_hd__mux2_1 _664_ (.A0(_124_),
    .A1(_114_),
    .S(_386_),
    .X(_238_));
 sky130_fd_sc_hd__nand3_1 _665_ (.A(_082_),
    .B(_031_),
    .C(_126_),
    .Y(_239_));
 sky130_fd_sc_hd__o221ai_4 _666_ (.A1(_146_),
    .A2(_113_),
    .B1(_238_),
    .B2(_082_),
    .C1(_239_),
    .Y(_240_));
 sky130_fd_sc_hd__mux2i_2 _667_ (.A0(_237_),
    .A1(_240_),
    .S(_148_),
    .Y(_241_));
 sky130_fd_sc_hd__nand2_1 _668_ (.A(_026_),
    .B(_123_),
    .Y(_242_));
 sky130_fd_sc_hd__nand3_1 _669_ (.A(_100_),
    .B(_073_),
    .C(_074_),
    .Y(_243_));
 sky130_fd_sc_hd__nand3_1 _670_ (.A(_392_),
    .B(_242_),
    .C(_243_),
    .Y(_244_));
 sky130_fd_sc_hd__o221ai_4 _671_ (.A1(_033_),
    .A2(_081_),
    .B1(_128_),
    .B2(_146_),
    .C1(_244_),
    .Y(_245_));
 sky130_fd_sc_hd__nand2_1 _672_ (.A(net28),
    .B(_018_),
    .Y(_246_));
 sky130_fd_sc_hd__nand2_1 _673_ (.A(net26),
    .B(_015_),
    .Y(_247_));
 sky130_fd_sc_hd__nand2_1 _674_ (.A(_246_),
    .B(_247_),
    .Y(_248_));
 sky130_fd_sc_hd__mux2_1 _675_ (.A0(net23),
    .A1(net27),
    .S(_389_),
    .X(_249_));
 sky130_fd_sc_hd__mux2_1 _676_ (.A0(_106_),
    .A1(_249_),
    .S(_385_),
    .X(_250_));
 sky130_fd_sc_hd__nor3_1 _677_ (.A(_370_),
    .B(_049_),
    .C(_105_),
    .Y(_251_));
 sky130_fd_sc_hd__a221oi_2 _678_ (.A1(_127_),
    .A2(_248_),
    .B1(_250_),
    .B2(_392_),
    .C1(_251_),
    .Y(_252_));
 sky130_fd_sc_hd__nand2_1 _679_ (.A(_112_),
    .B(_252_),
    .Y(_253_));
 sky130_fd_sc_hd__o21ai_1 _680_ (.A1(_112_),
    .A2(_245_),
    .B1(_253_),
    .Y(_254_));
 sky130_fd_sc_hd__o22ai_1 _681_ (.A1(_153_),
    .A2(_241_),
    .B1(_254_),
    .B2(_192_),
    .Y(net44));
 sky130_fd_sc_hd__o21ai_0 _682_ (.A1(_214_),
    .A2(_217_),
    .B1(_170_),
    .Y(_255_));
 sky130_fd_sc_hd__nand2_1 _683_ (.A(net5),
    .B(_161_),
    .Y(_256_));
 sky130_fd_sc_hd__nand2_1 _684_ (.A(net32),
    .B(_161_),
    .Y(_257_));
 sky130_fd_sc_hd__mux2_1 _685_ (.A0(_256_),
    .A1(_257_),
    .S(_030_),
    .X(_258_));
 sky130_fd_sc_hd__a21o_1 _686_ (.A1(_378_),
    .A2(net2),
    .B1(_166_),
    .X(_259_));
 sky130_fd_sc_hd__mux2i_1 _687_ (.A0(net6),
    .A1(net2),
    .S(_042_),
    .Y(_260_));
 sky130_fd_sc_hd__nor3_1 _688_ (.A(_384_),
    .B(_167_),
    .C(_260_),
    .Y(_261_));
 sky130_fd_sc_hd__a31oi_1 _689_ (.A1(_014_),
    .A2(_164_),
    .A3(_259_),
    .B1(_261_),
    .Y(_262_));
 sky130_fd_sc_hd__nand3_1 _690_ (.A(_005_),
    .B(net4),
    .C(_015_),
    .Y(_263_));
 sky130_fd_sc_hd__nand3_1 _691_ (.A(_005_),
    .B(net31),
    .C(_015_),
    .Y(_264_));
 sky130_fd_sc_hd__mux2_1 _692_ (.A0(_263_),
    .A1(_264_),
    .S(_029_),
    .X(_265_));
 sky130_fd_sc_hd__nand4_2 _693_ (.A(_255_),
    .B(_258_),
    .C(_262_),
    .D(_265_),
    .Y(_266_));
 sky130_fd_sc_hd__o21ai_0 _694_ (.A1(_049_),
    .A2(_141_),
    .B1(_392_),
    .Y(_267_));
 sky130_fd_sc_hd__a21o_1 _695_ (.A1(_026_),
    .A2(_080_),
    .B1(_267_),
    .X(_268_));
 sky130_fd_sc_hd__o221ai_2 _696_ (.A1(_146_),
    .A2(_060_),
    .B1(_145_),
    .B2(_033_),
    .C1(_268_),
    .Y(_269_));
 sky130_fd_sc_hd__mux2i_1 _697_ (.A0(_266_),
    .A1(_269_),
    .S(_066_),
    .Y(_270_));
 sky130_fd_sc_hd__mux2_1 _698_ (.A0(net9),
    .A1(net10),
    .S(net34),
    .X(_271_));
 sky130_fd_sc_hd__mux2_1 _699_ (.A0(net7),
    .A1(net8),
    .S(_004_),
    .X(_272_));
 sky130_fd_sc_hd__mux2_1 _700_ (.A0(_271_),
    .A1(_272_),
    .S(_003_),
    .X(_273_));
 sky130_fd_sc_hd__mux2_1 _701_ (.A0(_180_),
    .A1(_273_),
    .S(_030_),
    .X(_274_));
 sky130_fd_sc_hd__and2_0 _702_ (.A(_066_),
    .B(_274_),
    .X(_275_));
 sky130_fd_sc_hd__nand2_1 _703_ (.A(net21),
    .B(_015_),
    .Y(_276_));
 sky130_fd_sc_hd__nand2_1 _704_ (.A(net24),
    .B(_018_),
    .Y(_277_));
 sky130_fd_sc_hd__nor2_1 _705_ (.A(_014_),
    .B(_138_),
    .Y(_278_));
 sky130_fd_sc_hd__a311oi_1 _706_ (.A1(_082_),
    .A2(_276_),
    .A3(_277_),
    .B1(_278_),
    .C1(_100_),
    .Y(_279_));
 sky130_fd_sc_hd__a21oi_2 _707_ (.A1(_100_),
    .A2(_177_),
    .B1(_279_),
    .Y(_280_));
 sky130_fd_sc_hd__nor3_1 _708_ (.A(_066_),
    .B(_000_),
    .C(_280_),
    .Y(_281_));
 sky130_fd_sc_hd__o21ai_0 _709_ (.A1(_275_),
    .A2(_281_),
    .B1(_071_),
    .Y(_282_));
 sky130_fd_sc_hd__o21ai_0 _710_ (.A1(_192_),
    .A2(_270_),
    .B1(_282_),
    .Y(net45));
 sky130_fd_sc_hd__a22o_1 _711_ (.A1(_041_),
    .A2(_070_),
    .B1(_067_),
    .B2(_233_),
    .X(net46));
 sky130_fd_sc_hd__mux2i_1 _712_ (.A0(net2),
    .A1(net6),
    .S(_386_),
    .Y(_283_));
 sky130_fd_sc_hd__nand2_1 _713_ (.A(_014_),
    .B(_011_),
    .Y(_284_));
 sky130_fd_sc_hd__o32ai_1 _714_ (.A1(_370_),
    .A2(_018_),
    .A3(_283_),
    .B1(_284_),
    .B2(_159_),
    .Y(_285_));
 sky130_fd_sc_hd__a21oi_2 _715_ (.A1(_392_),
    .A2(_050_),
    .B1(_285_),
    .Y(_286_));
 sky130_fd_sc_hd__mux4_1 _716_ (.A0(_057_),
    .A1(_058_),
    .A2(_072_),
    .A3(_079_),
    .S0(_385_),
    .S1(_005_),
    .X(_287_));
 sky130_fd_sc_hd__mux2_1 _717_ (.A0(_286_),
    .A1(_287_),
    .S(_148_),
    .X(_288_));
 sky130_fd_sc_hd__mux2i_2 _718_ (.A0(_200_),
    .A1(_226_),
    .S(_385_),
    .Y(_289_));
 sky130_fd_sc_hd__nor3_1 _719_ (.A(_370_),
    .B(_386_),
    .C(_201_),
    .Y(_290_));
 sky130_fd_sc_hd__a221oi_4 _720_ (.A1(_127_),
    .A2(_229_),
    .B1(_289_),
    .B2(_370_),
    .C1(_290_),
    .Y(_291_));
 sky130_fd_sc_hd__nand2_1 _721_ (.A(_003_),
    .B(_271_),
    .Y(_292_));
 sky130_fd_sc_hd__o21ai_2 _722_ (.A1(_003_),
    .A2(_178_),
    .B1(_292_),
    .Y(_293_));
 sky130_fd_sc_hd__mux2i_2 _723_ (.A0(_199_),
    .A1(_293_),
    .S(_100_),
    .Y(_294_));
 sky130_fd_sc_hd__mux2_1 _724_ (.A0(_291_),
    .A1(_294_),
    .S(_148_),
    .X(_295_));
 sky130_fd_sc_hd__nand2_2 _725_ (.A(_086_),
    .B(_070_),
    .Y(_296_));
 sky130_fd_sc_hd__o22ai_1 _726_ (.A1(_192_),
    .A2(_288_),
    .B1(_295_),
    .B2(_296_),
    .Y(net47));
 sky130_fd_sc_hd__o2111ai_1 _727_ (.A1(_100_),
    .A2(_108_),
    .B1(_090_),
    .C1(_382_),
    .D1(_099_),
    .Y(_297_));
 sky130_fd_sc_hd__a21boi_0 _728_ (.A1(_112_),
    .A2(_120_),
    .B1_N(_297_),
    .Y(_298_));
 sky130_fd_sc_hd__mux2i_1 _729_ (.A0(_083_),
    .A1(_130_),
    .S(_382_),
    .Y(_299_));
 sky130_fd_sc_hd__nand3_1 _730_ (.A(_086_),
    .B(_233_),
    .C(_299_),
    .Y(_300_));
 sky130_fd_sc_hd__o21ai_0 _731_ (.A1(_153_),
    .A2(_298_),
    .B1(_300_),
    .Y(net48));
 sky130_fd_sc_hd__mux2i_1 _732_ (.A0(_137_),
    .A1(_174_),
    .S(_133_),
    .Y(_301_));
 sky130_fd_sc_hd__nor3_1 _733_ (.A(_148_),
    .B(_143_),
    .C(_147_),
    .Y(_302_));
 sky130_fd_sc_hd__a211o_1 _734_ (.A1(_066_),
    .A2(_181_),
    .B1(_302_),
    .C1(_000_),
    .X(_303_));
 sky130_fd_sc_hd__o22ai_1 _735_ (.A1(_192_),
    .A2(_301_),
    .B1(_303_),
    .B2(_153_),
    .Y(net49));
 sky130_fd_sc_hd__o22ai_1 _736_ (.A1(_296_),
    .A2(_288_),
    .B1(_295_),
    .B2(_071_),
    .Y(net50));
 sky130_fd_sc_hd__o211ai_1 _737_ (.A1(_151_),
    .A2(_195_),
    .B1(_196_),
    .C1(_133_),
    .Y(_304_));
 sky130_fd_sc_hd__o21ai_0 _738_ (.A1(_133_),
    .A2(_188_),
    .B1(_304_),
    .Y(_305_));
 sky130_fd_sc_hd__mux2i_1 _739_ (.A0(_189_),
    .A1(_193_),
    .S(_066_),
    .Y(_306_));
 sky130_fd_sc_hd__nand2_1 _740_ (.A(_233_),
    .B(_306_),
    .Y(_307_));
 sky130_fd_sc_hd__o21ai_0 _741_ (.A1(_153_),
    .A2(_305_),
    .B1(_307_),
    .Y(net51));
 sky130_fd_sc_hd__nand2_1 _742_ (.A(_099_),
    .B(_231_),
    .Y(_308_));
 sky130_fd_sc_hd__a21oi_1 _743_ (.A1(net24),
    .A2(_015_),
    .B1(_370_),
    .Y(_309_));
 sky130_fd_sc_hd__a21oi_2 _744_ (.A1(_370_),
    .A2(_226_),
    .B1(_309_),
    .Y(_310_));
 sky130_fd_sc_hd__a31oi_1 _745_ (.A1(_100_),
    .A2(_151_),
    .A3(_310_),
    .B1(_148_),
    .Y(_311_));
 sky130_fd_sc_hd__a22o_1 _746_ (.A1(_066_),
    .A2(_203_),
    .B1(_308_),
    .B2(_311_),
    .X(_312_));
 sky130_fd_sc_hd__nand2_1 _747_ (.A(_133_),
    .B(_206_),
    .Y(_313_));
 sky130_fd_sc_hd__o21ai_0 _748_ (.A1(_133_),
    .A2(_224_),
    .B1(_313_),
    .Y(_314_));
 sky130_fd_sc_hd__o22ai_1 _749_ (.A1(_296_),
    .A2(_312_),
    .B1(_314_),
    .B2(_192_),
    .Y(net52));
 sky130_fd_sc_hd__nor3_1 _750_ (.A(_148_),
    .B(_151_),
    .C(_252_),
    .Y(_315_));
 sky130_fd_sc_hd__a21oi_1 _751_ (.A1(_112_),
    .A2(_237_),
    .B1(_315_),
    .Y(_316_));
 sky130_fd_sc_hd__mux2i_1 _752_ (.A0(_240_),
    .A1(_245_),
    .S(_066_),
    .Y(_317_));
 sky130_fd_sc_hd__nand3_1 _753_ (.A(net1),
    .B(_011_),
    .C(_156_),
    .Y(_318_));
 sky130_fd_sc_hd__o221ai_1 _754_ (.A1(_153_),
    .A2(_316_),
    .B1(_317_),
    .B2(_192_),
    .C1(_318_),
    .Y(net53));
 sky130_fd_sc_hd__nand3_1 _755_ (.A(net25),
    .B(_100_),
    .C(_170_),
    .Y(_319_));
 sky130_fd_sc_hd__o21ai_0 _756_ (.A1(_099_),
    .A2(_319_),
    .B1(_382_),
    .Y(_320_));
 sky130_fd_sc_hd__a21oi_1 _757_ (.A1(_099_),
    .A2(_269_),
    .B1(_320_),
    .Y(_321_));
 sky130_fd_sc_hd__nand2_1 _758_ (.A(_112_),
    .B(_280_),
    .Y(_322_));
 sky130_fd_sc_hd__nand2_1 _759_ (.A(_068_),
    .B(_322_),
    .Y(_323_));
 sky130_fd_sc_hd__mux2_1 _760_ (.A0(_266_),
    .A1(_274_),
    .S(_381_),
    .X(_324_));
 sky130_fd_sc_hd__a32oi_1 _761_ (.A1(net12),
    .A2(_011_),
    .A3(_156_),
    .B1(_233_),
    .B2(_324_),
    .Y(_325_));
 sky130_fd_sc_hd__o21ai_0 _762_ (.A1(_321_),
    .A2(_323_),
    .B1(_325_),
    .Y(net54));
 sky130_fd_sc_hd__o21ai_0 _763_ (.A1(_035_),
    .A2(_039_),
    .B1(_382_),
    .Y(_326_));
 sky130_fd_sc_hd__o21a_1 _764_ (.A1(_382_),
    .A2(_056_),
    .B1(_326_),
    .X(_327_));
 sky130_fd_sc_hd__mux2_1 _765_ (.A0(_059_),
    .A1(_063_),
    .S(_392_),
    .X(_328_));
 sky130_fd_sc_hd__nor2_1 _766_ (.A(_382_),
    .B(_027_),
    .Y(_329_));
 sky130_fd_sc_hd__a31oi_1 _767_ (.A1(_133_),
    .A2(_086_),
    .A3(_328_),
    .B1(_329_),
    .Y(_330_));
 sky130_fd_sc_hd__nand2_1 _768_ (.A(net1),
    .B(_003_),
    .Y(_331_));
 sky130_fd_sc_hd__nand2_1 _769_ (.A(net23),
    .B(_011_),
    .Y(_332_));
 sky130_fd_sc_hd__nand2_1 _770_ (.A(_331_),
    .B(_332_),
    .Y(_333_));
 sky130_fd_sc_hd__nand2_1 _771_ (.A(_156_),
    .B(_333_),
    .Y(_334_));
 sky130_fd_sc_hd__o221ai_1 _772_ (.A1(_192_),
    .A2(_327_),
    .B1(_330_),
    .B2(_153_),
    .C1(_334_),
    .Y(net55));
 sky130_fd_sc_hd__mux2i_1 _773_ (.A0(_286_),
    .A1(_294_),
    .S(_381_),
    .Y(_335_));
 sky130_fd_sc_hd__or3_1 _774_ (.A(_387_),
    .B(_372_),
    .C(_084_),
    .X(_336_));
 sky130_fd_sc_hd__buf_2 _775_ (.A(_336_),
    .X(_337_));
 sky130_fd_sc_hd__nor2_1 _776_ (.A(_057_),
    .B(_337_),
    .Y(_338_));
 sky130_fd_sc_hd__a22oi_2 _777_ (.A1(_001_),
    .A2(_202_),
    .B1(_310_),
    .B2(_026_),
    .Y(_339_));
 sky130_fd_sc_hd__nand3_1 _778_ (.A(_086_),
    .B(_070_),
    .C(_151_),
    .Y(_340_));
 sky130_fd_sc_hd__mux2_1 _779_ (.A0(_287_),
    .A1(_291_),
    .S(_065_),
    .X(_341_));
 sky130_fd_sc_hd__nand2_1 _780_ (.A(_070_),
    .B(_099_),
    .Y(_342_));
 sky130_fd_sc_hd__o22ai_1 _781_ (.A1(_339_),
    .A2(_340_),
    .B1(_341_),
    .B2(_342_),
    .Y(_343_));
 sky130_fd_sc_hd__a211o_1 _782_ (.A1(_233_),
    .A2(_335_),
    .B1(_338_),
    .C1(_343_),
    .X(net56));
 sky130_fd_sc_hd__nand3_1 _783_ (.A(_133_),
    .B(_119_),
    .C(_117_),
    .Y(_344_));
 sky130_fd_sc_hd__nand3_1 _784_ (.A(_131_),
    .B(_233_),
    .C(_344_),
    .Y(_345_));
 sky130_fd_sc_hd__o221ai_1 _785_ (.A1(_153_),
    .A2(_111_),
    .B1(_337_),
    .B2(_072_),
    .C1(_345_),
    .Y(net57));
 sky130_fd_sc_hd__a211oi_1 _786_ (.A1(_112_),
    .A2(_174_),
    .B1(_182_),
    .C1(_070_),
    .Y(_346_));
 sky130_fd_sc_hd__a311oi_1 _787_ (.A1(_133_),
    .A2(_086_),
    .A3(_137_),
    .B1(_149_),
    .C1(_046_),
    .Y(_347_));
 sky130_fd_sc_hd__nor3_2 _788_ (.A(_000_),
    .B(_046_),
    .C(_098_),
    .Y(_348_));
 sky130_fd_sc_hd__nor2_1 _789_ (.A(_080_),
    .B(_337_),
    .Y(_349_));
 sky130_fd_sc_hd__a21oi_1 _790_ (.A1(_155_),
    .A2(_348_),
    .B1(_349_),
    .Y(_350_));
 sky130_fd_sc_hd__o31ai_1 _791_ (.A1(_151_),
    .A2(_346_),
    .A3(_347_),
    .B1(_350_),
    .Y(net58));
 sky130_fd_sc_hd__nor2_1 _792_ (.A(_060_),
    .B(_337_),
    .Y(_351_));
 sky130_fd_sc_hd__a21oi_1 _793_ (.A1(_025_),
    .A2(_348_),
    .B1(_351_),
    .Y(_352_));
 sky130_fd_sc_hd__o221ai_1 _794_ (.A1(_191_),
    .A2(_192_),
    .B1(_198_),
    .B2(_342_),
    .C1(_352_),
    .Y(net59));
 sky130_fd_sc_hd__nand2_1 _795_ (.A(_233_),
    .B(_207_),
    .Y(_353_));
 sky130_fd_sc_hd__a32oi_1 _796_ (.A1(_070_),
    .A2(_099_),
    .A3(_232_),
    .B1(_310_),
    .B2(_348_),
    .Y(_354_));
 sky130_fd_sc_hd__o211ai_1 _797_ (.A1(_058_),
    .A2(_337_),
    .B1(_353_),
    .C1(_354_),
    .Y(net60));
 sky130_fd_sc_hd__nand3_1 _798_ (.A(_086_),
    .B(_071_),
    .C(_299_),
    .Y(_355_));
 sky130_fd_sc_hd__o21ai_0 _799_ (.A1(_071_),
    .A2(_298_),
    .B1(_355_),
    .Y(net61));
 sky130_fd_sc_hd__nand2_1 _800_ (.A(_103_),
    .B(_348_),
    .Y(_356_));
 sky130_fd_sc_hd__o22a_1 _801_ (.A1(_079_),
    .A2(_337_),
    .B1(_192_),
    .B2(_241_),
    .X(_357_));
 sky130_fd_sc_hd__o211ai_1 _802_ (.A1(_254_),
    .A2(_342_),
    .B1(_356_),
    .C1(_357_),
    .Y(net62));
 sky130_fd_sc_hd__nor2_1 _803_ (.A(_081_),
    .B(_337_),
    .Y(_358_));
 sky130_fd_sc_hd__a31oi_1 _804_ (.A1(net25),
    .A2(_170_),
    .A3(_348_),
    .B1(_358_),
    .Y(_359_));
 sky130_fd_sc_hd__o21ai_0 _805_ (.A1(_275_),
    .A2(_281_),
    .B1(_233_),
    .Y(_360_));
 sky130_fd_sc_hd__o211ai_1 _806_ (.A1(_270_),
    .A2(_342_),
    .B1(_359_),
    .C1(_360_),
    .Y(net63));
 sky130_fd_sc_hd__o22ai_1 _807_ (.A1(_296_),
    .A2(_301_),
    .B1(_303_),
    .B2(_071_),
    .Y(net64));
 sky130_fd_sc_hd__nand2_1 _808_ (.A(_068_),
    .B(_306_),
    .Y(_361_));
 sky130_fd_sc_hd__o21ai_0 _809_ (.A1(_071_),
    .A2(_305_),
    .B1(_361_),
    .Y(net65));
 sky130_fd_sc_hd__o22ai_1 _810_ (.A1(_071_),
    .A2(_312_),
    .B1(_314_),
    .B2(_296_),
    .Y(net66));
 sky130_fd_sc_hd__o22ai_1 _811_ (.A1(_071_),
    .A2(_316_),
    .B1(_317_),
    .B2(_296_),
    .Y(net67));
 sky130_fd_sc_hd__nand2_1 _812_ (.A(_046_),
    .B(_322_),
    .Y(_362_));
 sky130_fd_sc_hd__nand2_1 _813_ (.A(_068_),
    .B(_324_),
    .Y(_363_));
 sky130_fd_sc_hd__o21ai_0 _814_ (.A1(_321_),
    .A2(_362_),
    .B1(_363_),
    .Y(net68));
 sky130_fd_sc_hd__nor3_1 _815_ (.A(_035_),
    .B(_039_),
    .C(_046_),
    .Y(_364_));
 sky130_fd_sc_hd__nor2_1 _816_ (.A(_070_),
    .B(_328_),
    .Y(_365_));
 sky130_fd_sc_hd__mux2_1 _817_ (.A0(_027_),
    .A1(_056_),
    .S(_069_),
    .X(_366_));
 sky130_fd_sc_hd__o32ai_1 _818_ (.A1(_087_),
    .A2(_364_),
    .A3(_365_),
    .B1(_366_),
    .B2(_133_),
    .Y(net69));
 sky130_fd_sc_hd__nand2_1 _819_ (.A(_099_),
    .B(_341_),
    .Y(_367_));
 sky130_fd_sc_hd__o221ai_1 _820_ (.A1(_057_),
    .A2(_337_),
    .B1(_339_),
    .B2(_382_),
    .C1(_151_),
    .Y(_368_));
 sky130_fd_sc_hd__a32o_1 _821_ (.A1(_046_),
    .A2(_367_),
    .A3(_368_),
    .B1(_068_),
    .B2(_335_),
    .X(net70));
 sky130_fd_sc_hd__ha_1 _822_ (.A(_392_),
    .B(_393_),
    .COUT(_394_),
    .SUM(_395_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_69 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(data_in[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(data_in[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(data_in[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(data_in[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(data_in[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(data_in[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(data_in[15]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(data_in[16]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(data_in[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(data_in[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(data_in[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input12 (.A(data_in[1]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(data_in[20]),
    .X(net13));
 sky130_fd_sc_hd__dlymetal6s2s_1 input14 (.A(data_in[21]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(data_in[22]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(data_in[23]),
    .X(net16));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(data_in[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(data_in[25]),
    .X(net18));
 sky130_fd_sc_hd__dlymetal6s2s_1 input19 (.A(data_in[26]),
    .X(net19));
 sky130_fd_sc_hd__dlymetal6s2s_1 input20 (.A(data_in[27]),
    .X(net20));
 sky130_fd_sc_hd__dlymetal6s2s_1 input21 (.A(data_in[28]),
    .X(net21));
 sky130_fd_sc_hd__dlymetal6s2s_1 input22 (.A(data_in[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_2 input23 (.A(data_in[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_2 input24 (.A(data_in[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_2 input25 (.A(data_in[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_2 input26 (.A(data_in[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(data_in[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(data_in[5]),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 input29 (.A(data_in[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(data_in[7]),
    .X(net30));
 sky130_fd_sc_hd__dlymetal6s2s_1 input31 (.A(data_in[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(data_in[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_2 input33 (.A(direction),
    .X(net33));
 sky130_fd_sc_hd__buf_2 input34 (.A(rotate_amount[0]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(rotate_amount[1]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 input36 (.A(rotate_amount[2]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_4 input37 (.A(rotate_amount[3]),
    .X(net37));
 sky130_fd_sc_hd__buf_2 input38 (.A(rotate_amount[4]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 output39 (.A(net39),
    .X(data_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output40 (.A(net40),
    .X(data_out[10]));
 sky130_fd_sc_hd__clkbuf_1 output41 (.A(net41),
    .X(data_out[11]));
 sky130_fd_sc_hd__clkbuf_1 output42 (.A(net42),
    .X(data_out[12]));
 sky130_fd_sc_hd__clkbuf_1 output43 (.A(net43),
    .X(data_out[13]));
 sky130_fd_sc_hd__clkbuf_1 output44 (.A(net44),
    .X(data_out[14]));
 sky130_fd_sc_hd__clkbuf_1 output45 (.A(net45),
    .X(data_out[15]));
 sky130_fd_sc_hd__clkbuf_1 output46 (.A(net46),
    .X(data_out[16]));
 sky130_fd_sc_hd__clkbuf_1 output47 (.A(net47),
    .X(data_out[17]));
 sky130_fd_sc_hd__clkbuf_1 output48 (.A(net48),
    .X(data_out[18]));
 sky130_fd_sc_hd__clkbuf_1 output49 (.A(net49),
    .X(data_out[19]));
 sky130_fd_sc_hd__clkbuf_1 output50 (.A(net50),
    .X(data_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output51 (.A(net51),
    .X(data_out[20]));
 sky130_fd_sc_hd__clkbuf_1 output52 (.A(net52),
    .X(data_out[21]));
 sky130_fd_sc_hd__clkbuf_1 output53 (.A(net53),
    .X(data_out[22]));
 sky130_fd_sc_hd__clkbuf_1 output54 (.A(net54),
    .X(data_out[23]));
 sky130_fd_sc_hd__clkbuf_1 output55 (.A(net55),
    .X(data_out[24]));
 sky130_fd_sc_hd__clkbuf_1 output56 (.A(net56),
    .X(data_out[25]));
 sky130_fd_sc_hd__clkbuf_1 output57 (.A(net57),
    .X(data_out[26]));
 sky130_fd_sc_hd__clkbuf_1 output58 (.A(net58),
    .X(data_out[27]));
 sky130_fd_sc_hd__clkbuf_1 output59 (.A(net59),
    .X(data_out[28]));
 sky130_fd_sc_hd__clkbuf_1 output60 (.A(net60),
    .X(data_out[29]));
 sky130_fd_sc_hd__clkbuf_1 output61 (.A(net61),
    .X(data_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output62 (.A(net62),
    .X(data_out[30]));
 sky130_fd_sc_hd__clkbuf_1 output63 (.A(net63),
    .X(data_out[31]));
 sky130_fd_sc_hd__clkbuf_1 output64 (.A(net64),
    .X(data_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output65 (.A(net65),
    .X(data_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output66 (.A(net66),
    .X(data_out[5]));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net67),
    .X(data_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net68),
    .X(data_out[7]));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(net69),
    .X(data_out[8]));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net70),
    .X(data_out[9]));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_5 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_87 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_94 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_157 ();
endmodule
