
* cell clock_divider
* pin PWELL
* pin NWELL
* pin duty_cycle[7]
* pin duty_cycle[6]
* pin duty_cycle[5]
* pin clk_out
* pin clk_in
* pin duty_cycle[1]
* pin duty_cycle[3]
* pin duty_cycle[2]
* pin div_ratio[5]
* pin duty_cycle[4]
* pin div_ratio[4]
* pin duty_cycle[0]
* pin div_ratio[3]
* pin div_ratio[1]
* pin div_ratio[2]
* pin div_ratio[6]
* pin div_ratio[7]
* pin div_ratio[0]
* pin rst_n
.SUBCKT clock_divider 1 2 3 4 5 6 912 978 979 980 981 982 983 984 985 986 990
+ 991 993 994 995
* net 1 PWELL
* net 2 NWELL
* net 3 duty_cycle[7]
* net 4 duty_cycle[6]
* net 5 duty_cycle[5]
* net 6 clk_out
* net 912 clk_in
* net 978 duty_cycle[1]
* net 979 duty_cycle[3]
* net 980 duty_cycle[2]
* net 981 div_ratio[5]
* net 982 duty_cycle[4]
* net 983 div_ratio[4]
* net 984 duty_cycle[0]
* net 985 div_ratio[3]
* net 986 div_ratio[1]
* net 990 div_ratio[2]
* net 991 div_ratio[6]
* net 993 div_ratio[7]
* net 994 div_ratio[0]
* net 995 rst_n
* cell instance $1 m0 *1 238.07,463.4
X$1 987 2 848 1 BUF_X4
* cell instance $3 m0 *1 239.4,463.4
X$3 995 1 2 987 CLKBUF_X1
* cell instance $35 m0 *1 215.65,463.4
X$35 985 1 2 961 BUF_X1
* cell instance $39 m0 *1 217.93,463.4
X$39 990 1 2 963 BUF_X1
* cell instance $42 m0 *1 220.21,463.4
X$42 991 2 879 1 BUF_X4
* cell instance $43 m0 *1 221.54,463.4
X$43 993 1 2 497 BUF_X2
* cell instance $52 m0 *1 238.07,410.2
X$52 103 146 104 1 125 2 AOI21_X2
* cell instance $53 m0 *1 239.4,410.2
X$53 123 143 102 2 1 124 AND3_X1
* cell instance $96 m0 *1 220.4,410.2
X$96 1 118 106 62 94 44 2 AOI22_X4
* cell instance $100 r0 *1 220.59,410.2
X$100 118 106 1 222 2 NAND2_X4
* cell instance $103 r0 *1 224.2,410.2
X$103 85 119 140 1 2 121 NAND3_X2
* cell instance $104 r0 *1 225.53,410.2
X$104 140 119 85 2 1 148 AND3_X1
* cell instance $106 m0 *1 232.37,410.2
X$106 86 87 73 2 1 151 AND3_X1
* cell instance $107 m0 *1 231.61,410.2
X$107 73 87 86 1 2 105 NAND3_X1
* cell instance $111 m0 *1 235.79,410.2
X$111 123 121 102 2 1 149 AND3_X1
* cell instance $116 r0 *1 233.7,410.2
X$116 120 143 145 2 1 144 AND3_X1
* cell instance $118 r0 *1 236.17,410.2
X$118 121 123 105 1 122 2 AOI21_X2
* cell instance $119 r0 *1 237.5,410.2
X$119 143 120 1 2 103 NAND2_X1
* cell instance $121 r0 *1 238.83,410.2
X$121 102 121 123 1 2 146 NAND3_X1
* cell instance $454 m0 *1 210.52,463.4
X$454 986 1 2 752 BUF_X2
* cell instance $18268 m0 *1 203.49,407.4
X$18268 67 89 1 2 51 NOR2_X1
* cell instance $18269 m0 *1 203.11,407.4
X$18269 67 1 2 76 INV_X1
* cell instance $18270 m0 *1 204.06,407.4
X$18270 1 51 68 82 76 69 70 49 2 AOI222_X2
* cell instance $18272 m0 *1 206.91,407.4
X$18272 1 77 2 90 BUF_X8
* cell instance $18273 m0 *1 209.38,407.4
X$18273 67 83 53 1 2 80 MUX2_X1
* cell instance $18274 m0 *1 210.71,407.4
X$18274 67 70 77 1 53 2 AOI21_X1
* cell instance $18276 m0 *1 214.51,407.4
X$18276 99 14 2 1 79 AND2_X1
* cell instance $18277 m0 *1 215.27,407.4
X$18277 78 1 2 24 BUF_X2
* cell instance $18282 r0 *1 203.49,407.4
X$18282 133 81 1 2 69 NAND2_X1
* cell instance $18283 r0 *1 204.06,407.4
X$18283 77 1 2 92 BUF_X1
* cell instance $18284 r0 *1 204.63,407.4
X$18284 68 1 2 91 BUF_X2
* cell instance $18285 r0 *1 205.39,407.4
X$18285 1 17 91 109 70 77 2 AOI22_X4
* cell instance $18286 r0 *1 208.62,407.4
X$18286 1 92 36 95 97 93 2 AOI22_X4
* cell instance $18287 r0 *1 211.85,407.4
X$18287 81 18 11 2 1 93 OAI21_X2
* cell instance $18290 r0 *1 213.75,407.4
X$18290 40 38 108 1 2 NOR2_X4
* cell instance $18293 r0 *1 217.36,407.4
X$18293 84 52 79 71 2 1 117 AND4_X1
* cell instance $18295 m0 *1 220.21,407.4
X$18295 80 2 55 1 BUF_X4
* cell instance $18296 m0 *1 221.54,407.4
X$18296 44 94 71 65 2 1 58 AND4_X2
* cell instance $18299 r0 *1 221.92,407.4
X$18299 1 71 65 44 94 85 2 NAND4_X4
* cell instance $18300 m0 *1 224.39,407.4
X$18300 65 71 72 1 2 57 NAND3_X2
* cell instance $18301 m0 *1 223.25,407.4
X$18301 72 71 65 2 1 47 AND3_X2
* cell instance $18303 r0 *1 225.34,407.4
X$18303 1 47 45 120 74 85 2 AOI22_X4
* cell instance $18304 m0 *1 228.19,407.4
X$18304 56 1 2 88 BUF_X1
* cell instance $18305 m0 *1 226.1,407.4
X$18305 74 85 29 47 45 75 2 1 AOI221_X2
* cell instance $18306 m0 *1 228.76,407.4
X$18306 57 62 30 58 46 63 1 2 OAI221_X2
* cell instance $18307 m0 *1 230.85,407.4
X$18307 59 31 29 61 86 102 1 2 OAI221_X2
* cell instance $18312 r0 *1 228.95,407.4
X$18312 88 46 57 62 87 1 2 OAI211_X2
* cell instance $18313 r0 *1 230.66,407.4
X$18313 86 58 1 2 188 OR2_X2
* cell instance $18462 m0 *1 205.01,404.6
X$18462 1 38 10 35 40 34 2 NOR4_X4
* cell instance $18463 m0 *1 208.43,404.6
X$18463 41 1 2 35 BUF_X1
* cell instance $18464 m0 *1 209,404.6
X$18464 1 36 9 17 11 2 AOI21_X4
* cell instance $18465 m0 *1 211.47,404.6
X$18465 37 42 8 2 1 44 OAI21_X4
* cell instance $18466 m0 *1 213.94,404.6
X$18466 26 24 18 2 25 1 NOR3_X2
* cell instance $18467 m0 *1 215.27,404.6
X$18467 20 22 79 1 2 21 NAND3_X2
* cell instance $18468 m0 *1 216.6,404.6
X$18468 26 18 1 2 54 NOR2_X1
* cell instance $18469 m0 *1 217.17,404.6
X$18469 23 1 2 15 BUF_X1
* cell instance $18471 m0 *1 218.5,404.6
X$18471 19 52 36 2 1 33 AND3_X1
* cell instance $18472 m0 *1 219.45,404.6
X$18472 36 24 19 1 2 66 NAND3_X2
* cell instance $18474 m0 *1 220.97,404.6
X$18474 12 14 1 2 27 NOR2_X1
* cell instance $18475 m0 *1 221.54,404.6
X$18475 14 12 2 1 28 AND2_X1
* cell instance $18476 m0 *1 222.3,404.6
X$18476 13 33 32 2 1 30 OAI21_X2
* cell instance $18481 m0 *1 229.14,404.6
X$18481 56 29 58 30 31 1 2 OAI211_X2
* cell instance $18537 r0 *1 202.54,404.6
X$18537 50 1 2 14 BUF_X2
* cell instance $18540 r0 *1 204.25,404.6
X$18540 52 50 1 38 2 NAND2_X4
* cell instance $18541 r0 *1 205.96,404.6
X$18541 1 38 10 41 49 2 NOR3_X4
* cell instance $18542 r0 *1 208.62,404.6
X$18542 1 65 9 39 64 2 AOI21_X4
* cell instance $18543 r0 *1 211.09,404.6
X$18543 40 18 1 2 39 NAND2_X1
* cell instance $18545 r0 *1 212.04,404.6
X$18545 40 89 1 2 42 NOR2_X1
* cell instance $18546 r0 *1 212.61,404.6
X$18546 41 1 2 23 BUF_X2
* cell instance $18547 r0 *1 213.37,404.6
X$18547 38 41 12 1 43 2 AOI21_X1
* cell instance $18548 r0 *1 214.13,404.6
X$18548 10 43 36 1 48 2 AOI21_X1
* cell instance $18549 r0 *1 214.89,404.6
X$18549 1 29 25 24 21 2 AOI21_X4
* cell instance $18550 r0 *1 217.36,404.6
X$18550 54 21 24 2 1 46 MUX2_X2
* cell instance $18552 r0 *1 220.59,404.6
X$18552 1 74 27 66 28 2 AOI21_X4
* cell instance $18556 r0 *1 225.53,404.6
X$18556 45 47 1 2 59 NAND2_X1
* cell instance $18557 r0 *1 226.1,404.6
X$18557 45 29 47 55 1 2 73 NAND4_X1
* cell instance $18561 r0 *1 227.05,404.6
X$18561 55 2 56 1 BUF_X4
* cell instance $18562 r0 *1 228.38,404.6
X$18562 57 62 58 30 56 61 1 2 OAI221_X2
* cell instance $18563 r0 *1 230.47,404.6
X$18563 29 59 1 2 60 XNOR2_X2
* cell instance $19685 m0 *1 189.05,421.4
X$19685 216 1 2 201 INV_X2
* cell instance $19688 m0 *1 191.9,421.4
X$19688 301 248 300 1 2 246 NAND3_X1
* cell instance $19690 m0 *1 192.85,421.4
X$19690 217 249 302 248 301 218 2 1 AOI221_X2
* cell instance $19691 m0 *1 194.94,421.4
X$19691 300 1 2 268 INV_X1
* cell instance $19731 r0 *1 193.42,421.4
X$19731 1 267 302 248 301 2 AOI21_X4
* cell instance $19733 m0 *1 195.7,421.4
X$19733 268 291 267 1 269 2 AOI21_X1
* cell instance $19736 r0 *1 196.65,421.4
X$19736 268 500 325 267 2 1 260 AND4_X1
* cell instance $19737 m0 *1 197.79,421.4
X$19737 270 271 296 2 1 217 OAI21_X4
* cell instance $19746 r0 *1 202.16,421.4
X$19746 303 306 304 2 1 326 AND3_X1
* cell instance $19748 m0 *1 202.92,421.4
X$19748 326 2 17 1 BUF_X4
* cell instance $19749 m0 *1 205.77,421.4
X$19749 305 2 134 1 BUF_X4
* cell instance $19752 m0 *1 208.81,421.4
X$19752 250 219 272 115 177 328 1 2 OAI221_X2
* cell instance $19753 m0 *1 210.9,421.4
X$19753 34 1 2 272 BUF_X1
* cell instance $19756 m0 *1 215.27,421.4
X$19756 307 1 2 273 BUF_X1
* cell instance $19760 r0 *1 204.25,421.4
X$19760 303 306 304 11 2 1 376 AND4_X1
* cell instance $19763 r0 *1 205.96,421.4
X$19763 305 2 178 1 BUF_X4
* cell instance $19766 r0 *1 210.71,421.4
X$19766 81 250 219 2 1 341 OAI21_X2
* cell instance $19769 r0 *1 212.99,421.4
X$19769 328 134 2 332 1 XOR2_X2
* cell instance $19770 r0 *1 214.7,421.4
X$19770 1 307 353 332 314 274 2 OAI22_X4
* cell instance $19771 m0 *1 216.41,421.4
X$19771 95 134 1 2 308 NAND2_X1
* cell instance $19775 m0 *1 218.69,421.4
X$19775 307 308 1 2 278 OR2_X2
* cell instance $19779 r0 *1 218.31,421.4
X$19779 308 307 1 2 339 NOR2_X2
* cell instance $19782 m0 *1 220.97,421.4
X$19782 275 266 1 2 279 NOR2_X2
* cell instance $19785 m0 *1 222.11,421.4
X$19785 195 275 266 2 1 310 OAI21_X2
* cell instance $19788 r0 *1 221.92,421.4
X$19788 311 1 2 356 BUF_X1
* cell instance $19789 r0 *1 222.49,421.4
X$19789 276 1 2 335 BUF_X1
* cell instance $19790 r0 *1 223.06,421.4
X$19790 277 311 222 2 1 355 OAI21_X4
* cell instance $19791 m0 *1 226.48,421.4
X$19791 314 75 278 315 338 1 2 OAI211_X2
* cell instance $19792 m0 *1 223.82,421.4
X$19792 1 335 222 311 313 2 NOR3_X4
* cell instance $19793 m0 *1 228.19,421.4
X$19793 314 278 337 2 1 226 OAI21_X4
* cell instance $19798 r0 *1 226.86,421.4
X$19798 336 1 2 315 BUF_X1
* cell instance $19799 r0 *1 227.43,421.4
X$19799 1 449 354 338 317 316 2 OAI22_X4
* cell instance $19800 r0 *1 230.66,421.4
X$19800 1 316 63 330 334 2 NOR3_X4
* cell instance $19802 m0 *1 231.04,421.4
X$19802 225 252 226 297 313 279 1 2 333 OAI33_X1
* cell instance $19803 m0 *1 232.56,421.4
X$19803 164 86 280 1 331 2 AOI21_X1
* cell instance $19804 m0 *1 233.32,421.4
X$19804 226 1 2 295 BUF_X1
* cell instance $19808 r0 *1 233.32,421.4
X$19808 333 1 2 329 BUF_X2
* cell instance $19810 r0 *1 234.46,421.4
X$19810 331 230 327 1 324 2 AOI21_X2
* cell instance $19814 r0 *1 238.45,421.4
X$19814 231 166 344 2 320 1 OAI21_X1
* cell instance $19817 r0 *1 239.78,421.4
X$19817 231 166 211 2 406 1 OAI21_X1
* cell instance $19824 r0 *1 243.96,421.4
X$19824 317 230 1 2 345 NOR2_X1
* cell instance $19826 r0 *1 244.72,421.4
X$19826 318 286 345 1 2 319 NAND3_X1
* cell instance $19829 m0 *1 246.43,421.4
X$19829 255 283 1 2 323 OR2_X1
* cell instance $19832 m0 *1 247.95,421.4
X$19832 352 321 1 2 284 NOR2_X1
* cell instance $19871 r0 *1 246.62,421.4
X$19871 320 324 1 2 351 XOR2_X1
* cell instance $19873 r0 *1 247.95,421.4
X$19873 320 324 2 1 350 XNOR2_X1
* cell instance $19875 r0 *1 249.28,421.4
X$19875 253 283 1 2 397 XNOR2_X2
* cell instance $19876 r0 *1 251.18,421.4
X$19876 319 323 322 1 2 349 NAND3_X1
* cell instance $20029 m0 *1 184.11,449.4
X$20029 828 812 829 2 1 729 HA_X1
* cell instance $20030 m0 *1 183.35,449.4
X$20030 678 778 2 1 828 AND2_X1
* cell instance $20033 m0 *1 190.57,449.4
X$20033 486 732 2 1 815 AND2_X1
* cell instance $20034 m0 *1 191.33,449.4
X$20034 831 815 814 2 1 830 HA_X1
* cell instance $20038 r0 *1 185.25,449.4
X$20038 1 856 781 803 829 813 2 FA_X1
* cell instance $20042 r0 *1 190.76,449.4
X$20042 678 780 2 1 831 AND2_X1
* cell instance $20043 r0 *1 191.52,449.4
X$20043 1 908 832 833 814 872 2 FA_X1
* cell instance $20046 m0 *1 196.65,449.4
X$20046 833 1 2 816 INV_X1
* cell instance $20052 r0 *1 198.74,449.4
X$20052 1 871 818 836 835 876 2 FA_X1
* cell instance $20053 r0 *1 201.78,449.4
X$20053 836 1 2 839 INV_X2
* cell instance $20057 r0 *1 209.57,449.4
X$20057 844 1 2 843 INV_X1
* cell instance $20059 m0 *1 211.28,449.4
X$20059 849 752 2 1 846 AND2_X1
* cell instance $20061 m0 *1 212.04,449.4
X$20061 1 847 845 850 846 819 2 FA_X1
* cell instance $20062 m0 *1 215.08,449.4
X$20062 753 849 1 2 851 NAND2_X1
* cell instance $20068 r0 *1 212.99,449.4
X$20068 776 732 2 1 819 AND2_X1
* cell instance $20071 r0 *1 220.21,449.4
X$20071 903 566 2 866 1 XOR2_X2
* cell instance $20074 r0 *1 223.63,449.4
X$20074 632 866 820 2 1 859 HA_X1
* cell instance $20080 r0 *1 227.24,449.4
X$20080 854 865 2 1 821 XNOR2_X1
* cell instance $20081 m0 *1 227.62,449.4
X$20081 852 1 2 854 INV_X1
* cell instance $20089 r0 *1 230.47,449.4
X$20089 632 823 756 825 1 2 860 NAND4_X1
* cell instance $20092 m0 *1 232.18,449.4
X$20092 824 842 2 1 838 XNOR2_X1
* cell instance $20099 r0 *1 232.75,449.4
X$20099 888 823 756 825 1 2 842 NAND4_X1
* cell instance $20102 m0 *1 241.87,449.4
X$20102 825 718 797 2 1 791 HA_X1
* cell instance $20105 m0 *1 244.53,449.4
X$20105 862 794 798 2 1 827 HA_X1
* cell instance $20147 r0 *1 243.77,449.4
X$20147 826 792 827 1 863 2 AOI21_X2
* cell instance $20270 r0 *1 179.17,443.8
X$20270 484 778 2 1 796 AND2_X1
* cell instance $20272 m0 *1 185.06,443.8
X$20272 1 704 727 705 731 729 2 FA_X1
* cell instance $20277 r0 *1 186.58,443.8
X$20277 484 780 2 1 704 AND2_X1
* cell instance $20280 m0 *1 188.48,443.8
X$20280 485 732 2 1 731 AND2_X1
* cell instance $20283 r0 *1 189.43,443.8
X$20283 1 764 763 765 766 782 2 FA_X1
* cell instance $20284 m0 *1 189.81,443.8
X$20284 732 484 1 2 764 NAND2_X1
* cell instance $20286 m0 *1 190.38,443.8
X$20286 1 832 706 735 765 733 2 FA_X1
* cell instance $20289 m0 *1 195.7,443.8
X$20289 707 1 2 708 INV_X1
* cell instance $20293 m0 *1 201.4,443.8
X$20293 485 753 2 1 769 AND2_X1
* cell instance $20299 r0 *1 196.27,443.8
X$20299 747 485 1 2 766 NAND2_X1
* cell instance $20301 r0 *1 197.03,443.8
X$20301 484 747 2 1 783 AND2_X1
* cell instance $20305 r0 *1 200.26,443.8
X$20305 1 771 749 784 769 751 2 FA_X1
* cell instance $20306 r0 *1 203.3,443.8
X$20306 484 752 2 1 771 AND2_X1
* cell instance $20309 r0 *1 205.96,443.8
X$20309 678 752 2 1 811 AND2_X1
* cell instance $20311 m0 *1 207.29,443.8
X$20311 678 753 2 1 738 AND2_X1
* cell instance $20316 m0 *1 210.9,443.8
X$20316 780 710 2 1 739 AND2_X1
* cell instance $20318 m0 *1 211.66,443.8
X$20318 738 739 775 2 1 664 HA_X1
* cell instance $20319 m0 *1 213.56,443.8
X$20319 775 1 2 740 INV_X1
* cell instance $20320 m0 *1 213.94,443.8
X$20320 1 755 711 712 850 740 2 FA_X1
* cell instance $20322 m0 *1 220.02,443.8
X$20322 710 732 1 2 668 NAND2_X1
* cell instance $20324 m0 *1 220.78,443.8
X$20324 710 752 2 1 744 AND2_X1
* cell instance $20325 m0 *1 221.54,443.8
X$20325 776 753 2 1 743 AND2_X1
* cell instance $20327 m0 *1 222.49,443.8
X$20327 747 710 2 1 713 AND2_X1
* cell instance $20328 m0 *1 223.25,443.8
X$20328 743 744 624 2 1 714 HA_X1
* cell instance $20337 r0 *1 220.78,443.8
X$20337 776 752 2 1 777 AND2_X1
* cell instance $20338 r0 *1 221.54,443.8
X$20338 787 777 670 2 1 681 HA_X1
* cell instance $20343 r0 *1 234.84,443.8
X$20343 823 607 757 2 1 773 HA_X1
* cell instance $20344 r0 *1 236.74,443.8
X$20344 1 774 773 757 768 2 AOI21_X4
* cell instance $20346 m0 *1 236.93,443.8
X$20346 685 1 2 772 INV_X1
* cell instance $20347 m0 *1 237.5,443.8
X$20347 716 1 2 770 INV_X1
* cell instance $20350 m0 *1 238.83,443.8
X$20350 834 717 1 642 2 OR2_X4
* cell instance $20352 r0 *1 239.21,443.8
X$20352 770 772 767 2 1 768 OAI21_X4
* cell instance $20357 m0 *1 241.68,443.8
X$20357 1 759 642 758 717 737 762 800 2 OAI222_X2
* cell instance $20359 r0 *1 241.68,443.8
X$20359 699 801 1 2 758 NOR2_X1
* cell instance $20361 m0 *1 249.47,443.8
X$20361 620 1 2 722 BUF_X1
* cell instance $20362 m0 *1 247.76,443.8
X$20362 513 619 689 719 720 1 2 OAI211_X2
* cell instance $20363 m0 *1 250.04,443.8
X$20363 723 730 688 513 1 2 759 AOI22_X2
* cell instance $20365 m0 *1 252.51,443.8
X$20365 690 726 724 624 1 2 761 NOR4_X1
* cell instance $20403 r0 *1 248.33,443.8
X$20403 761 720 760 1 762 2 AOI21_X1
* cell instance $20405 r0 *1 249.47,443.8
X$20405 513 726 1 2 730 NOR2_X1
* cell instance $20551 m0 *1 178.22,446.6
X$20551 1 796 795 799 802 779 2 FA_X1
* cell instance $20556 m0 *1 183.73,446.6
X$20556 485 780 2 1 802 AND2_X1
* cell instance $20559 m0 *1 185.44,446.6
X$20559 781 1 2 745 INV_X1
* cell instance $20565 r0 *1 183.92,446.6
X$20565 486 780 2 1 812 AND2_X1
* cell instance $20569 m0 *1 190.76,446.6
X$20569 803 1 2 733 INV_X1
* cell instance $20571 m0 *1 195.7,446.6
X$20571 1 783 746 837 804 817 2 FA_X1
* cell instance $20573 r0 *1 191.14,446.6
X$20573 830 1 2 782 INV_X1
* cell instance $20576 r0 *1 196.08,446.6
X$20576 1 818 707 748 816 837 2 FA_X1
* cell instance $20579 m0 *1 199.12,446.6
X$20579 485 752 2 1 804 AND2_X1
* cell instance $20580 m0 *1 201.4,446.6
X$20580 1 807 750 808 839 784 2 FA_X1
* cell instance $20585 r0 *1 204.25,446.6
X$20585 486 753 2 1 841 AND2_X1
* cell instance $20586 m0 *1 207.86,446.6
X$20586 1 845 754 709 843 809 2 FA_X1
* cell instance $20587 m0 *1 204.82,446.6
X$20587 1 811 806 809 810 841 2 FA_X1
* cell instance $20592 r0 *1 205.39,446.6
X$20592 778 710 2 1 810 AND2_X1
* cell instance $20596 r0 *1 213.18,446.6
X$20596 785 747 2 1 847 AND2_X1
* cell instance $20598 m0 *1 218.88,446.6
X$20598 747 776 1 2 805 NAND2_X1
* cell instance $20599 m0 *1 215.84,446.6
X$20599 1 786 755 741 851 805 2 FA_X1
* cell instance $20604 r0 *1 217.55,446.6
X$20604 752 785 1 2 786 NAND2_X1
* cell instance $20608 r0 *1 220.78,446.6
X$20608 785 753 2 1 787 AND2_X1
* cell instance $20611 m0 *1 225.91,446.6
X$20611 1 788 852 638 853 848 2 DFFR_X1
* cell instance $20617 m0 *1 242.06,446.6
X$20617 1 789 800 848 997 7 2 DFFR_X2
* cell instance $20619 m0 *1 246.43,446.6
X$20619 720 726 2 1 794 AND2_X2
* cell instance $20661 r0 *1 227.62,446.6
X$20661 821 822 1 2 853 NOR2_X1
* cell instance $20665 r0 *1 229.52,446.6
X$20665 1 788 840 848 824 632 2 DFFR_X2
* cell instance $20666 r0 *1 233.7,446.6
X$20666 838 822 1 2 840 NOR2_X1
* cell instance $20669 r0 *1 241.87,446.6
X$20669 798 792 797 757 1 2 801 NAND4_X1
* cell instance $20670 r0 *1 242.82,446.6
X$20670 1 767 791 790 797 2 AOI21_X4
* cell instance $20671 r0 *1 245.29,446.6
X$20671 793 687 792 2 1 826 HA_X1
* cell instance $20796 r0 *1 178.6,441
X$20796 485 778 2 1 692 AND2_X1
* cell instance $20797 m0 *1 178.98,441
X$20797 633 646 693 2 1 575 HA_X1
* cell instance $20802 r0 *1 179.36,441
X$20802 1 855 523 647 799 693 2 FA_X1
* cell instance $20803 r0 *1 182.4,441
X$20803 497 678 2 1 646 AND2_X1
* cell instance $20806 r0 *1 183.73,441
X$20806 1 745 626 696 728 703 2 FA_X1
* cell instance $20808 m0 *1 185.06,441
X$20808 727 1 2 648 INV_X1
* cell instance $20813 m0 *1 187.34,441
X$20813 696 1 2 649 INV_X1
* cell instance $20814 m0 *1 190.76,441
X$20814 697 1 2 593 INV_X1
* cell instance $20819 r0 *1 187.34,441
X$20819 705 1 2 728 INV_X1
* cell instance $20823 r0 *1 189.81,441
X$20823 706 1 2 614 INV_X1
* cell instance $20826 r0 *1 192.47,441
X$20826 1 708 697 653 734 735 2 FA_X1
* cell instance $20827 r0 *1 195.51,441
X$20827 746 1 2 734 INV_X1
* cell instance $20829 r0 *1 196.65,441
X$20829 1 698 679 634 748 736 2 FA_X1
* cell instance $20830 r0 *1 199.69,441
X$20830 749 1 2 698 INV_X1
* cell instance $20832 m0 *1 199.88,441
X$20832 634 1 2 598 INV_X2
* cell instance $20833 m0 *1 203.49,441
X$20833 484 753 2 1 635 AND2_X1
* cell instance $20834 m0 *1 204.25,441
X$20834 635 806 661 2 1 658 HA_X1
* cell instance $20835 m0 *1 206.15,441
X$20835 1 754 659 660 857 661 2 FA_X1
* cell instance $20841 r0 *1 200.64,441
X$20841 750 1 2 736 INV_X1
* cell instance $20844 r0 *1 204.25,441
X$20844 808 1 2 680 INV_X2
* cell instance $20848 m0 *1 214.13,441
X$20848 711 1 2 636 INV_X1
* cell instance $20852 m0 *1 217.36,441
X$20852 712 1 2 637 INV_X1
* cell instance $20856 m0 *1 218.69,441
X$20856 667 1 2 615 INV_X1
* cell instance $20857 m0 *1 219.07,441
X$20857 1 702 667 669 741 668 2 FA_X1
* cell instance $20861 r0 *1 222.3,441
X$20861 753 710 1 2 641 NAND2_X1
* cell instance $20862 m0 *1 222.68,441
X$20862 670 713 671 2 1 604 HA_X1
* cell instance $20864 m0 *1 224.58,441
X$20864 714 671 682 2 1 605 HA_X1
* cell instance $20868 m0 *1 228.95,441
X$20868 638 389 675 2 1 701 HA_X1
* cell instance $20871 r0 *1 223.06,441
X$20871 681 1 2 702 INV_X1
* cell instance $20876 r0 *1 228.95,441
X$20876 899 701 1 2 742 NOR2_X1
* cell instance $20877 r0 *1 229.52,441
X$20877 639 774 683 2 1 700 OAI21_X4
* cell instance $20878 m0 *1 233.7,441
X$20878 617 674 685 675 1 2 699 NAND4_X1
* cell instance $20879 m0 *1 231.23,441
X$20879 1 684 640 674 700 2 AOI21_X4
* cell instance $20880 m0 *1 234.65,441
X$20880 675 1 2 715 INV_X1
* cell instance $20885 r0 *1 231.99,441
X$20885 742 715 684 2 1 717 OAI21_X4
* cell instance $20888 r0 *1 236.17,441
X$20888 756 510 685 2 1 716 HA_X1
* cell instance $20891 m0 *1 242.44,441
X$20891 641 642 676 1 2 677 OR3_X4
* cell instance $20892 m0 *1 244.72,441
X$20892 618 1 2 687 BUF_X1
* cell instance $20894 m0 *1 245.48,441
X$20894 1 694 677 631 665 2 AOI21_X4
* cell instance $20896 m0 *1 248.71,441
X$20896 619 1 2 663 BUF_X1
* cell instance $20897 m0 *1 249.28,441
X$20897 533 691 655 643 663 688 1 2 OAI221_X2
* cell instance $20898 m0 *1 251.37,441
X$20898 1 689 651 631 665 2 AOI21_X4
* cell instance $20899 m0 *1 253.84,441
X$20899 624 652 725 2 1 644 HA_X1
* cell instance $20900 m0 *1 255.74,441
X$20900 644 645 1 2 690 XOR2_X1
* cell instance $20937 r0 *1 244.91,441
X$20937 694 686 695 2 1 737 OAI21_X2
* cell instance $20938 r0 *1 246.24,441
X$20938 721 565 726 1 2 695 NOR3_X1
* cell instance $20940 r0 *1 247.19,441
X$20940 561 621 620 641 2 1 719 AND4_X1
* cell instance $20941 r0 *1 248.33,441
X$20941 620 621 1 2 721 NAND2_X1
* cell instance $20942 r0 *1 248.9,441
X$20942 721 533 1 2 760 NOR2_X1
* cell instance $20943 r0 *1 249.47,441
X$20943 619 561 621 722 2 1 723 AND4_X1
* cell instance $20944 r0 *1 250.61,441
X$20944 689 1 2 691 BUF_X1
* cell instance $20945 r0 *1 251.18,441
X$20945 533 1 2 726 INV_X1
* cell instance $20949 r0 *1 252.89,441
X$20949 725 1 2 724 INV_X1
* cell instance $21055 m0 *1 189.05,424.2
X$21055 202 147 216 2 340 1 OAI21_X1
* cell instance $21057 m0 *1 190,424.2
X$21057 159 357 201 2 375 1 NOR3_X2
* cell instance $21058 m0 *1 191.33,424.2
X$21058 357 201 1 2 407 NOR2_X1
* cell instance $21062 m0 *1 202.54,424.2
X$21062 306 303 304 1 89 2 NAND3_X4
* cell instance $21066 m0 *1 207.48,424.2
X$21066 1 376 377 312 443 71 2 NOR4_X4
* cell instance $21069 m0 *1 214.13,424.2
X$21069 134 328 1 2 378 XNOR2_X2
* cell instance $21070 m0 *1 216.03,424.2
X$21070 183 199 341 1 2 353 OR3_X1
* cell instance $21071 m0 *1 216.98,424.2
X$21071 341 199 183 2 379 1 NOR3_X2
* cell instance $21112 r0 *1 187.72,424.2
X$21112 436 1 2 216 CLKBUF_X2
* cell instance $21113 r0 *1 188.48,424.2
X$21113 403 1 2 383 INV_X1
* cell instance $21114 r0 *1 188.86,424.2
X$21114 302 147 300 1 2 381 NAND3_X1
* cell instance $21115 r0 *1 189.62,424.2
X$21115 357 383 340 2 1 405 AND3_X1
* cell instance $21116 r0 *1 190.57,424.2
X$21116 357 1 2 385 INV_X1
* cell instance $21117 r0 *1 190.95,424.2
X$21117 384 407 405 403 385 306 2 1 AOI221_X2
* cell instance $21121 r0 *1 200.83,424.2
X$21121 375 386 358 2 1 303 OAI21_X2
* cell instance $21123 r0 *1 202.35,424.2
X$21123 358 386 1 2 387 NOR2_X1
* cell instance $21126 r0 *1 203.49,424.2
X$21126 387 410 11 306 2 1 377 OAI22_X2
* cell instance $21127 r0 *1 205.2,424.2
X$21127 360 361 375 1 2 410 NAND3_X1
* cell instance $21128 r0 *1 205.96,424.2
X$21128 388 359 2 1 81 AND2_X2
* cell instance $21130 r0 *1 207.1,424.2
X$21130 359 388 1 2 135 NAND2_X1
* cell instance $21132 r0 *1 207.86,424.2
X$21132 360 361 1 11 2 NAND2_X4
* cell instance $21138 r0 *1 215.46,424.2
X$21138 341 307 1 2 394 NOR2_X2
* cell instance $21140 r0 *1 217.17,424.2
X$21140 274 1 2 389 INV_X2
* cell instance $21142 r0 *1 217.93,424.2
X$21142 1 362 379 366 378 389 2 AOI22_X4
* cell instance $21143 m0 *1 220.4,424.2
X$21143 1 183 199 312 390 2 NOR3_X4
* cell instance $21145 m0 *1 223.06,424.2
X$21145 356 222 1 2 363 NOR2_X1
* cell instance $21146 m0 *1 223.63,424.2
X$21146 310 364 142 277 312 354 2 1 AOI221_X2
* cell instance $21153 r0 *1 222.49,424.2
X$21153 95 184 362 1 365 2 AOI21_X2
* cell instance $21154 r0 *1 223.82,424.2
X$21154 172 184 1 2 364 NAND2_X1
* cell instance $21155 r0 *1 224.39,424.2
X$21155 312 277 1 2 392 NAND2_X1
* cell instance $21156 r0 *1 224.96,424.2
X$21156 142 195 1 2 393 NAND2_X1
* cell instance $21159 r0 *1 226.1,424.2
X$21159 1 145 365 355 394 2 AOI21_X4
* cell instance $21160 m0 *1 228.57,424.2
X$21160 1 143 366 355 339 2 AOI21_X4
* cell instance $21162 m0 *1 231.04,424.2
X$21162 336 1 2 337 BUF_X2
* cell instance $21164 m0 *1 231.99,424.2
X$21164 279 313 367 1 2 NOR2_X4
* cell instance $21165 m0 *1 233.7,424.2
X$21165 226 1 2 330 BUF_X1
* cell instance $21168 m0 *1 235.22,424.2
X$21168 1 342 329 343 211 2 NOR3_X4
* cell instance $21169 m0 *1 237.88,424.2
X$21169 317 343 368 342 1 2 344 NOR4_X1
* cell instance $21174 m0 *1 241.49,424.2
X$21174 283 253 2 369 1 XOR2_X2
* cell instance $21175 m0 *1 243.2,424.2
X$21175 1 255 213 346 347 370 2 NOR4_X4
* cell instance $21176 m0 *1 246.62,424.2
X$21176 347 346 232 317 1 2 352 NOR4_X1
* cell instance $21177 m0 *1 247.57,424.2
X$21177 145 284 351 1 2 348 MUX2_X1
* cell instance $21178 m0 *1 248.9,424.2
X$21178 401 351 234 1 2 371 OR3_X2
* cell instance $21179 m0 *1 250.04,424.2
X$21179 323 253 2 372 1 XOR2_X2
* cell instance $21180 m0 *1 251.75,424.2
X$21180 349 253 2 373 1 XOR2_X2
* cell instance $21218 r0 *1 228.57,424.2
X$21218 63 366 339 355 424 2 1 AOI211_X2
* cell instance $21219 r0 *1 230.28,424.2
X$21219 355 394 2 1 409 AND2_X1
* cell instance $21220 r0 *1 231.04,424.2
X$21220 409 365 1 2 230 OR2_X2
* cell instance $21221 r0 *1 231.99,424.2
X$21221 252 1 2 316 BUF_X1
* cell instance $21225 r0 *1 233.89,424.2
X$21225 367 195 342 1 2 NOR2_X4
* cell instance $21229 r0 *1 237.69,424.2
X$21229 329 1 2 368 BUF_X1
* cell instance $21230 r0 *1 238.26,424.2
X$21230 329 2 395 1 BUF_X4
* cell instance $21232 r0 *1 239.97,424.2
X$21232 168 406 2 1 446 AND2_X1
* cell instance $21234 r0 *1 241.49,424.2
X$21234 404 369 370 1 396 2 AOI21_X2
* cell instance $21235 r0 *1 242.82,424.2
X$21235 374 1 2 404 BUF_X1
* cell instance $21237 r0 *1 243.77,424.2
X$21237 370 369 1 2 322 NAND2_X2
* cell instance $21238 r0 *1 244.72,424.2
X$21238 345 1 2 255 INV_X2
* cell instance $21239 r0 *1 245.29,424.2
X$21239 1 398 255 346 213 402 2 OR4_X4
* cell instance $21240 r0 *1 247.76,424.2
X$21240 346 402 1 2 401 OR2_X2
* cell instance $21242 r0 *1 248.9,424.2
X$21242 232 401 397 398 350 400 1 2 OAI221_X2
* cell instance $21382 r0 *1 182.97,427
X$21382 487 1 2 435 INV_X1
* cell instance $21385 m0 *1 183.54,427
X$21385 463 535 434 2 1 433 HA_X1
* cell instance $21386 m0 *1 185.44,427
X$21386 433 1 2 202 BUF_X2
* cell instance $21387 m0 *1 186.2,427
X$21387 434 1 2 147 CLKBUF_X3
* cell instance $21390 m0 *1 188.1,427
X$21390 202 147 380 1 412 2 AOI21_X1
* cell instance $21392 r0 *1 186.39,427
X$21392 465 435 436 2 1 403 HA_X1
* cell instance $21393 r0 *1 188.29,427
X$21393 380 300 302 1 243 2 AOI21_X2
* cell instance $21394 m0 *1 190.19,427
X$21394 412 381 1 2 384 NAND2_X1
* cell instance $21395 m0 *1 189.24,427
X$21395 412 381 383 357 1 2 382 NAND4_X1
* cell instance $21399 m0 *1 191.33,427
X$21399 384 403 385 1 2 441 NOR3_X1
* cell instance $21403 r0 *1 192.09,427
X$21403 1 437 301 204 438 2 AOI21_X4
* cell instance $21404 m0 *1 192.66,427
X$21404 243 413 437 2 1 408 OAI21_X2
* cell instance $21408 r0 *1 194.56,427
X$21408 1 248 416 300 204 414 2 NAND4_X4
* cell instance $21409 m0 *1 197.6,427
X$21409 414 1 2 440 INV_X1
* cell instance $21410 m0 *1 195.13,427
X$21410 1 130 408 440 417 2 AOI21_X4
* cell instance $21412 m0 *1 198.74,427
X$21412 415 416 1 2 325 NAND2_X1
* cell instance $21413 m0 *1 199.31,427
X$21413 386 358 382 1 2 304 OR3_X2
* cell instance $21414 m0 *1 200.45,427
X$21414 416 417 2 305 1 XOR2_X2
* cell instance $21417 r0 *1 197.98,427
X$21417 1 270 438 416 415 2 AOI21_X4
* cell instance $21420 m0 *1 204.25,427
X$21420 387 441 361 360 2 1 443 AND4_X1
* cell instance $21423 m0 *1 206.15,427
X$21423 1 360 361 359 388 177 2 AND4_X4
* cell instance $21426 m0 *1 214.89,427
X$21426 172 133 1 2 419 NAND2_X1
* cell instance $21427 m0 *1 215.46,427
X$21427 419 447 109 2 1 307 MUX2_X2
* cell instance $21428 m0 *1 217.17,427
X$21428 172 11 1 2 447 NAND2_X1
* cell instance $21430 r0 *1 205.01,427
X$21430 442 271 418 1 2 388 OR3_X2
* cell instance $21431 r0 *1 206.15,427
X$21431 442 418 271 2 1 359 OAI21_X2
* cell instance $21432 r0 *1 207.48,427
X$21432 467 455 452 2 1 361 OAI21_X4
* cell instance $21434 r0 *1 210.33,427
X$21434 361 360 2 1 444 AND2_X1
* cell instance $21437 r0 *1 211.66,427
X$21437 444 1 2 133 CLKBUF_X3
* cell instance $21441 r0 *1 216.79,427
X$21441 312 11 1 2 420 NOR2_X1
* cell instance $21442 r0 *1 217.36,427
X$21442 312 133 1 2 421 NOR2_X1
* cell instance $21445 m0 *1 218.12,427
X$21445 109 133 1 2 276 XNOR2_X2
* cell instance $21446 m0 *1 222.49,427
X$21446 276 390 1 2 391 OR2_X1
* cell instance $21447 m0 *1 220.4,427
X$21447 184 172 309 390 276 411 1 2 OAI221_X2
* cell instance $21448 m0 *1 223.25,427
X$21448 391 363 309 392 449 2 1 AOI211_X2
* cell instance $21449 m0 *1 224.96,427
X$21449 423 390 393 363 1 2 450 NOR4_X1
* cell instance $21452 m0 *1 232.75,427
X$21452 367 334 450 2 327 1 OAI21_X1
* cell instance $21458 r0 *1 222.87,427
X$21458 390 276 1 2 422 NOR2_X1
* cell instance $21459 r0 *1 223.44,427
X$21459 171 422 310 423 448 1 2 OAI211_X2
* cell instance $21462 r0 *1 226.86,427
X$21462 1 448 411 168 424 207 2 AOI22_X4
* cell instance $21464 r0 *1 230.85,427
X$21464 207 424 457 281 60 507 2 1 AOI221_X2
* cell instance $21466 r0 *1 233.32,427
X$21466 1 231 334 60 281 2 AOI21_X4
* cell instance $21469 m0 *1 236.17,427
X$21469 342 343 395 1 2 425 OR3_X4
* cell instance $21471 r0 *1 236.74,427
X$21471 445 457 1 2 343 NAND2_X2
* cell instance $21474 r0 *1 238.26,427
X$21474 342 395 1 2 458 OR2_X1
* cell instance $21475 m0 *1 239.97,427
X$21475 395 342 1 2 426 NOR2_X2
* cell instance $21476 m0 *1 238.64,427
X$21476 425 2 210 1 BUF_X4
* cell instance $21485 r0 *1 241.68,427
X$21485 426 289 445 1 346 2 NAND3_X4
* cell instance $21487 m0 *1 243.96,427
X$21487 427 346 1 2 318 NOR2_X1
* cell instance $21489 m0 *1 246.81,427
X$21489 402 1 2 347 BUF_X1
* cell instance $21491 m0 *1 248.9,427
X$21491 397 439 321 1 2 NOR2_X4
* cell instance $21492 m0 *1 250.61,427
X$21492 398 2 439 1 BUF_X4
* cell instance $21493 m0 *1 251.94,427
X$21493 398 397 431 2 399 1 OAI21_X1
* cell instance $21495 m0 *1 252.89,427
X$21495 371 285 2 1 432 AND2_X1
* cell instance $21534 r0 *1 244.72,427
X$21534 402 1 2 427 BUF_X1
* cell instance $21536 r0 *1 246.81,427
X$21536 402 2 428 1 BUF_X4
* cell instance $21539 r0 *1 248.71,427
X$21539 399 429 285 371 430 2 1 AOI211_X2
* cell instance $21540 r0 *1 250.42,427
X$21540 1 483 321 285 371 2 AOI21_X4
* cell instance $21541 r0 *1 252.89,427
X$21541 285 371 1 2 460 NAND2_X1
* cell instance $21680 m0 *1 177.46,432.6
X$21680 494 1 2 515 INV_X1
* cell instance $21686 r0 *1 177.65,432.6
X$21686 1 523 535 538 795 534 2 FA_X1
* cell instance $21688 m0 *1 180.5,432.6
X$21688 495 1 2 496 INV_X1
* cell instance $21689 m0 *1 182.4,432.6
X$21689 484 497 2 1 518 AND2_X1
* cell instance $21697 m0 *1 185.82,432.6
X$21697 485 497 2 1 498 AND2_X1
* cell instance $21699 r0 *1 186.2,432.6
X$21699 538 539 537 2 1 380 HA_X1
* cell instance $21700 m0 *1 187.15,432.6
X$21700 537 1 2 300 CLKBUF_X3
* cell instance $21702 m0 *1 188.1,432.6
X$21702 499 2 248 1 BUF_X4
* cell instance $21708 r0 *1 190.19,432.6
X$21708 578 2 204 1 BUF_X4
* cell instance $21710 r0 *1 191.71,432.6
X$21710 580 1 2 301 CLKBUF_X3
* cell instance $21712 m0 *1 193.04,432.6
X$21712 301 1 2 524 INV_X1
* cell instance $21714 m0 *1 193.42,432.6
X$21714 248 1 2 540 INV_X1
* cell instance $21717 r0 *1 193.04,432.6
X$21717 540 525 524 1 544 2 AOI21_X1
* cell instance $21719 r0 *1 194.18,432.6
X$21719 438 416 204 2 525 1 OAI21_X1
* cell instance $21720 r0 *1 194.94,432.6
X$21720 1 542 541 131 525 501 543 544 2 AOI222_X2
* cell instance $21721 m0 *1 195.13,432.6
X$21721 301 248 1 2 501 NOR2_X1
* cell instance $21723 m0 *1 195.7,432.6
X$21723 500 451 501 2 1 542 AND3_X1
* cell instance $21724 m0 *1 196.65,432.6
X$21724 438 301 1 2 545 NOR2_X1
* cell instance $21725 m0 *1 197.22,432.6
X$21725 451 545 453 452 543 1 2 OAI211_X2
* cell instance $21726 m0 *1 198.93,432.6
X$21726 453 452 1 2 541 OR2_X2
* cell instance $21729 m0 *1 200.45,432.6
X$21729 1 451 415 503 502 2 AOI21_X4
* cell instance $21732 m0 *1 203.68,432.6
X$21732 1 454 503 470 453 504 2 OAI211_X4
* cell instance $21733 m0 *1 206.91,432.6
X$21733 520 2 502 1 BUF_X4
* cell instance $21737 m0 *1 216.03,432.6
X$21737 526 548 549 504 1 2 452 AOI211_X4
* cell instance $21738 m0 *1 218.12,432.6
X$21738 506 527 548 2 1 549 HA_X1
* cell instance $21747 r0 *1 206.34,432.6
X$21747 582 2 454 1 BUF_X4
* cell instance $21751 r0 *1 212.61,432.6
X$21751 546 1 2 470 CLKBUF_X3
* cell instance $21753 r0 *1 214.32,432.6
X$21753 547 2 504 1 BUF_X4
* cell instance $21756 r0 *1 216.79,432.6
X$21756 1 527 505 550 526 506 2 FA_X1
* cell instance $21759 r0 *1 220.78,432.6
X$21759 550 2 195 1 BUF_X4
* cell instance $21763 r0 *1 223.44,432.6
X$21763 588 553 554 2 1 526 HA_X1
* cell instance $21765 r0 *1 225.53,432.6
X$21765 605 590 555 2 1 553 HA_X1
* cell instance $21768 r0 *1 228,432.6
X$21768 554 1 2 457 CLKBUF_X3
* cell instance $21770 r0 *1 230.47,432.6
X$21770 556 1 2 587 BUF_X1
* cell instance $21771 r0 *1 231.04,432.6
X$21771 555 1 2 289 CLKBUF_X3
* cell instance $21772 m0 *1 231.99,432.6
X$21772 528 1 2 556 BUF_X1
* cell instance $21774 m0 *1 232.56,432.6
X$21774 259 456 195 367 457 557 1 2 OAI221_X2
* cell instance $21775 m0 *1 234.65,432.6
X$21775 492 557 508 165 522 1 2 OAI211_X2
* cell instance $21776 m0 *1 236.36,432.6
X$21776 425 1 2 508 BUF_X2
* cell instance $21778 m0 *1 237.31,432.6
X$21778 532 231 1 2 510 NOR2_X2
* cell instance $21780 m0 *1 238.45,432.6
X$21780 458 396 510 1 573 2 AOI21_X2
* cell instance $21781 m0 *1 239.78,432.6
X$21781 425 510 490 2 564 1 OAI21_X1
* cell instance $21784 r0 *1 232.37,432.6
X$21784 559 1 2 560 BUF_X1
* cell instance $21785 r0 *1 232.94,432.6
X$21785 558 1 2 559 BUF_X1
* cell instance $21786 r0 *1 233.51,432.6
X$21786 1 507 529 530 402 165 2 OAI22_X4
* cell instance $21787 r0 *1 236.74,432.6
X$21787 425 2 531 1 BUF_X4
* cell instance $21789 r0 *1 238.26,432.6
X$21789 457 473 231 2 1 563 OAI21_X2
* cell instance $21790 r0 *1 239.59,432.6
X$21790 426 231 473 1 576 2 AOI21_X2
* cell instance $21791 r0 *1 240.92,432.6
X$21791 168 564 2 1 676 XNOR2_X1
* cell instance $21795 m0 *1 241.49,432.6
X$21795 490 511 562 2 1 565 OAI21_X2
* cell instance $21797 m0 *1 243.01,432.6
X$21797 474 286 1 2 718 NOR2_X1
* cell instance $21799 m0 *1 244.34,432.6
X$21799 512 402 458 1 2 562 NOR3_X1
* cell instance $21800 m0 *1 245.1,432.6
X$21800 286 289 1 2 512 NAND2_X1
* cell instance $21805 m0 *1 246.81,432.6
X$21805 429 459 1 2 629 NOR2_X1
* cell instance $21808 m0 *1 249.09,432.6
X$21808 348 488 483 1 2 551 NAND3_X1
* cell instance $21809 m0 *1 248.52,432.6
X$21809 512 322 1 2 552 NAND2_X1
* cell instance $21811 r0 *1 249.66,432.6
X$21811 430 552 514 372 570 2 1 AOI211_X2
* cell instance $21812 m0 *1 250.42,432.6
X$21812 551 348 480 2 1 513 OAI21_X2
* cell instance $21814 m0 *1 251.75,432.6
X$21814 514 483 1 2 478 NAND2_X1
* cell instance $21817 r0 *1 251.75,432.6
X$21817 482 1 2 514 BUF_X2
* cell instance $21818 r0 *1 252.51,432.6
X$21818 1 622 483 482 372 2 AOI21_X4
* cell instance $21820 m0 *1 252.7,432.6
X$21820 372 482 429 460 1 2 623 AOI211_X4
* cell instance $21958 m0 *1 178.41,435.4
X$21958 566 484 2 1 571 AND2_X1
* cell instance $21959 m0 *1 179.17,435.4
X$21959 574 536 534 2 1 495 HA_X1
* cell instance $22010 r0 *1 177.27,435.4
X$22010 1 571 494 574 692 575 2 FA_X1
* cell instance $22012 m0 *1 182.97,435.4
X$22012 485 566 2 1 469 AND2_X1
* cell instance $22013 m0 *1 182.21,435.4
X$22013 497 486 2 1 536 AND2_X1
* cell instance $22017 m0 *1 187.34,435.4
X$22017 591 611 499 2 1 302 HA_X1
* cell instance $22024 r0 *1 190,435.4
X$22024 594 593 578 2 1 580 HA_X1
* cell instance $22028 m0 *1 193.42,435.4
X$22028 627 2 416 1 BUF_X4
* cell instance $22032 m0 *1 200.26,435.4
X$22032 567 2 503 1 BUF_X4
* cell instance $22039 r0 *1 194.75,435.4
X$22039 597 1 2 438 CLKBUF_X3
* cell instance $22043 r0 *1 199.88,435.4
X$22043 598 628 567 2 1 415 HA_X1
* cell instance $22048 r0 *1 206.15,435.4
X$22048 583 599 582 2 1 520 HA_X1
* cell instance $22050 r0 *1 211.09,435.4
X$22050 601 600 584 2 1 583 HA_X1
* cell instance $22052 m0 *1 212.61,435.4
X$22052 585 584 546 2 1 547 HA_X1
* cell instance $22060 r0 *1 221.35,435.4
X$22060 589 612 588 2 1 506 HA_X1
* cell instance $22061 r0 *1 223.25,435.4
X$22061 604 603 590 2 1 589 HA_X1
* cell instance $22062 r0 *1 225.15,435.4
X$22062 109 1 2 672 INV_X1
* cell instance $22068 m0 *1 231.8,435.4
X$22068 587 1 2 568 BUF_X1
* cell instance $22070 m0 *1 232.37,435.4
X$22070 586 1 2 528 BUF_X1
* cell instance $22071 m0 *1 232.94,435.4
X$22071 568 529 1 2 577 NOR2_X1
* cell instance $22073 m0 *1 234.46,435.4
X$22073 560 1 2 586 BUF_X1
* cell instance $22074 m0 *1 233.89,435.4
X$22074 581 1 2 558 BUF_X1
* cell instance $22075 m0 *1 235.03,435.4
X$22075 507 1 2 581 BUF_X1
* cell instance $22080 m0 *1 237.31,435.4
X$22080 165 569 1 2 532 NOR2_X1
* cell instance $22081 m0 *1 235.98,435.4
X$22081 531 2 530 1 BUF_X4
* cell instance $22082 m0 *1 237.88,435.4
X$22082 1 573 509 561 576 563 2 AOI22_X4
* cell instance $22087 m0 *1 249.66,435.4
X$22087 431 1 2 475 INV_X1
* cell instance $22125 r0 *1 235.98,435.4
X$22125 531 1 2 579 BUF_X1
* cell instance $22128 r0 *1 237.12,435.4
X$22128 579 1 2 569 BUF_X1
* cell instance $22129 r0 *1 237.69,435.4
X$22129 577 532 1 2 572 NOR2_X2
* cell instance $22133 r0 *1 245.86,435.4
X$22133 570 572 1 2 609 NAND2_X1
* cell instance $22224 m0 *1 182.4,429.8
X$22224 468 1 2 463 INV_X1
* cell instance $22260 r0 *1 170.24,429.8
X$22260 4 1 2 484 BUF_X2
* cell instance $22263 r0 *1 174.8,429.8
X$22263 5 1 2 486 BUF_X2
* cell instance $22264 r0 *1 175.56,429.8
X$22264 3 1 2 485 BUF_X2
* cell instance $22268 r0 *1 178.79,429.8
X$22268 1 496 487 468 515 516 2 FA_X1
* cell instance $22269 r0 *1 181.83,429.8
X$22269 517 1 2 516 INV_X1
* cell instance $22272 r0 *1 182.78,429.8
X$22272 469 518 517 2 1 464 HA_X1
* cell instance $22274 m0 *1 188.1,429.8
X$22274 466 1 2 357 CLKBUF_X2
* cell instance $22275 m0 *1 186.2,429.8
X$22275 464 498 465 2 1 466 HA_X1
* cell instance $22279 m0 *1 193.61,429.8
X$22279 248 300 1 2 413 NAND2_X2
* cell instance $22283 m0 *1 195.13,429.8
X$22283 1 451 414 437 358 413 2 OAI22_X4
* cell instance $22286 m0 *1 198.55,429.8
X$22286 453 452 414 2 386 1 NOR3_X2
* cell instance $22287 m0 *1 199.88,429.8
X$22287 451 452 453 2 1 417 OAI21_X2
* cell instance $22290 m0 *1 204.44,429.8
X$22290 503 1 2 442 INV_X1
* cell instance $22295 r0 *1 195.7,429.8
X$22295 438 1 2 500 INV_X1
* cell instance $22299 r0 *1 200.83,429.8
X$22299 1 503 416 502 296 454 2 OAI211_X4
* cell instance $22302 r0 *1 205.77,429.8
X$22302 520 454 1 2 418 NOR2_X1
* cell instance $22304 r0 *1 206.53,429.8
X$22304 504 520 505 470 521 2 1 AOI211_X2
* cell instance $22306 m0 *1 207.48,429.8
X$22306 454 1 2 467 INV_X1
* cell instance $22307 m0 *1 208.05,429.8
X$22307 455 452 467 1 2 360 OR3_X4
* cell instance $22310 r0 *1 208.24,429.8
X$22310 521 2 271 1 BUF_X4
* cell instance $22311 r0 *1 209.57,429.8
X$22311 504 470 1 2 455 NOR2_X2
* cell instance $22313 r0 *1 210.9,429.8
X$22313 470 505 1 2 312 XNOR2_X2
* cell instance $22315 r0 *1 212.99,429.8
X$22315 505 470 2 172 1 XOR2_X2
* cell instance $22317 m0 *1 216.79,429.8
X$22317 420 421 109 2 1 362 MUX2_X2
* cell instance $22323 m0 *1 224.01,429.8
X$22323 172 184 1 2 423 NOR2_X2
* cell instance $22324 m0 *1 224.96,429.8
X$22324 1 313 390 423 445 2 NOR3_X4
* cell instance $22325 m0 *1 227.62,429.8
X$22325 313 184 1 2 606 NOR2_X1
* cell instance $22334 r0 *1 231.23,429.8
X$22334 60 457 1 2 493 NAND2_X1
* cell instance $22335 r0 *1 231.8,429.8
X$22335 1 493 259 280 529 471 2 OAI22_X4
* cell instance $22336 m0 *1 233.7,429.8
X$22336 60 1 2 456 INV_X1
* cell instance $22337 m0 *1 232.37,429.8
X$22337 280 259 456 2 1 282 OAI21_X2
* cell instance $22338 m0 *1 234.08,429.8
X$22338 334 367 195 2 492 1 OAI21_X1
* cell instance $22342 r0 *1 235.03,429.8
X$22342 334 367 1 2 607 NOR2_X1
* cell instance $22344 r0 *1 235.98,429.8
X$22344 457 1 2 471 INV_X1
* cell instance $22346 r0 *1 236.74,429.8
X$22346 522 445 2 511 1 XOR2_X2
* cell instance $22347 r0 *1 238.45,429.8
X$22347 471 396 282 2 1 509 OAI21_X2
* cell instance $22349 m0 *1 239.97,429.8
X$22349 425 1 2 472 BUF_X1
* cell instance $22352 r0 *1 239.97,429.8
X$22352 168 472 282 1 2 491 NOR3_X1
* cell instance $22357 m0 *1 241.49,429.8
X$22357 374 1 2 473 BUF_X1
* cell instance $22360 r0 *1 240.92,429.8
X$22360 511 374 491 446 519 476 1 2 OAI221_X2
* cell instance $22362 m0 *1 243.39,429.8
X$22362 459 1 2 474 BUF_X1
* cell instance $22366 m0 *1 245.67,429.8
X$22366 286 289 1 2 429 XNOR2_X2
* cell instance $22369 m0 *1 248.52,429.8
X$22369 1 476 429 321 400 482 2 NOR4_X4
* cell instance $22371 r0 *1 243.2,429.8
X$22371 459 286 318 1 490 2 AOI21_X2
* cell instance $22373 r0 *1 244.91,429.8
X$22373 1 475 458 428 519 2 NOR3_X4
* cell instance $22374 r0 *1 247.57,429.8
X$22374 459 429 476 1 2 477 OR3_X1
* cell instance $22376 r0 *1 248.9,429.8
X$22376 321 1 2 459 BUF_X2
* cell instance $22377 r0 *1 249.66,429.8
X$22377 476 429 489 1 2 488 NOR3_X1
* cell instance $22378 r0 *1 250.42,429.8
X$22378 459 1 2 489 BUF_X1
* cell instance $22379 r0 *1 250.99,429.8
X$22379 322 475 1 2 481 NAND2_X1
* cell instance $22380 r0 *1 251.56,429.8
X$22380 478 482 373 2 1 533 OAI21_X2
* cell instance $22381 m0 *1 252.51,429.8
X$22381 460 322 1 2 479 NAND2_X1
* cell instance $22384 m0 *1 253.27,429.8
X$22384 429 431 1 2 462 NAND2_X1
* cell instance $22385 m0 *1 253.84,429.8
X$22385 429 481 462 432 2 1 461 OAI22_X2
* cell instance $22424 r0 *1 253.08,429.8
X$22424 477 479 373 1 480 2 AOI21_X1
* cell instance $22750 m0 *1 178.6,452.2
X$22750 486 778 2 1 864 AND2_X1
* cell instance $22751 m0 *1 179.36,452.2
X$22751 883 864 884 2 1 779 HA_X1
* cell instance $22752 m0 *1 181.26,452.2
X$22752 1 886 855 703 884 867 2 FA_X1
* cell instance $22753 m0 *1 184.3,452.2
X$22753 497 849 2 1 867 AND2_X1
* cell instance $22755 m0 *1 185.82,452.2
X$22755 874 870 813 2 1 886 HA_X1
* cell instance $22757 m0 *1 188.48,452.2
X$22757 497 785 2 1 870 AND2_X1
* cell instance $22761 m0 *1 198.55,452.2
X$22761 486 747 2 1 921 AND2_X1
* cell instance $22813 r0 *1 184.3,452.2
X$22813 873 678 2 1 883 AND2_X1
* cell instance $22815 r0 *1 185.82,452.2
X$22815 873 849 2 1 874 AND2_X1
* cell instance $22819 r0 *1 191.9,452.2
X$22819 497 776 2 1 918 AND2_X1
* cell instance $22822 r0 *1 194.56,452.2
X$22822 920 1 2 835 INV_X1
* cell instance $22826 r0 *1 197.41,452.2
X$22826 1 875 817 876 891 921 2 FA_X1
* cell instance $22828 r0 *1 201.97,452.2
X$22828 497 710 2 1 891 AND2_X1
* cell instance $22829 m0 *1 202.16,452.2
X$22829 486 752 2 1 892 AND2_X1
* cell instance $22832 m0 *1 203.11,452.2
X$22832 1 895 807 896 877 894 2 FA_X1
* cell instance $22834 m0 *1 206.91,452.2
X$22834 896 1 2 857 INV_X1
* cell instance $22835 m0 *1 207.29,452.2
X$22835 849 747 2 1 898 AND2_X1
* cell instance $22836 m0 *1 208.05,452.2
X$22836 780 776 2 1 897 AND2_X1
* cell instance $22837 m0 *1 208.81,452.2
X$22837 785 732 2 1 878 AND2_X1
* cell instance $22842 r0 *1 202.73,452.2
X$22842 1 922 751 877 892 923 2 FA_X1
* cell instance $22843 r0 *1 205.77,452.2
X$22843 873 710 2 1 923 AND2_X1
* cell instance $22845 r0 *1 207.29,452.2
X$22845 1 878 895 844 897 898 2 FA_X1
* cell instance $22848 r0 *1 214.13,452.2
X$22848 1 566 2 879 BUF_X8
* cell instance $22851 m0 *1 218.5,452.2
X$22851 497 858 2 1 869 XNOR2_X1
* cell instance $22853 m0 *1 219.64,452.2
X$22853 616 869 904 2 1 902 HA_X1
* cell instance $22854 m0 *1 221.54,452.2
X$22854 902 854 901 879 497 903 1 2 868 OAI33_X1
* cell instance $22855 m0 *1 222.87,452.2
X$22855 904 1 2 880 INV_X1
* cell instance $22856 m0 *1 223.25,452.2
X$22856 880 906 905 1 901 2 AOI21_X1
* cell instance $22859 r0 *1 218.5,452.2
X$22859 900 778 566 1 2 858 NOR3_X1
* cell instance $22861 r0 *1 222.3,452.2
X$22861 903 497 879 1 2 899 NOR3_X1
* cell instance $22864 r0 *1 224.01,452.2
X$22864 929 930 820 2 906 1 OAI21_X1
* cell instance $22867 m0 *1 225.15,452.2
X$22867 859 1 2 905 INV_X1
* cell instance $22870 m0 *1 228,452.2
X$22870 889 822 1 2 881 NOR2_X1
* cell instance $22877 r0 *1 227.24,452.2
X$22877 1 788 881 848 890 616 2 DFFR_X2
* cell instance $22878 m0 *1 229.14,452.2
X$22878 913 1 2 788 CLKBUF_X3
* cell instance $22881 m0 *1 231.04,452.2
X$22881 888 616 1 2 893 NAND2_X1
* cell instance $22882 m0 *1 230.47,452.2
X$22882 893 860 1 2 865 NOR2_X1
* cell instance $22884 m0 *1 231.8,452.2
X$22884 860 861 1 2 927 NOR2_X1
* cell instance $22888 r0 *1 231.61,452.2
X$22888 890 927 1 2 889 XOR2_X1
* cell instance $22890 r0 *1 233.51,452.2
X$22890 887 822 1 2 911 NOR2_X1
* cell instance $22891 r0 *1 234.08,452.2
X$22891 925 924 2 1 887 XNOR2_X1
* cell instance $22892 r0 *1 235.22,452.2
X$22892 885 756 825 1 2 924 NAND3_X1
* cell instance $22893 m0 *1 235.98,452.2
X$22893 862 793 834 1 2 861 NAND3_X2
* cell instance $22901 r0 *1 236.17,452.2
X$22901 868 1 2 822 INV_X2
* cell instance $22903 r0 *1 236.93,452.2
X$22903 861 1 2 885 INV_X1
* cell instance $22905 r0 *1 237.69,452.2
X$22905 882 822 1 2 914 NOR2_X1
* cell instance $22906 r0 *1 238.26,452.2
X$22906 915 861 2 1 882 XNOR2_X1
* cell instance $22909 m0 *1 243.2,452.2
X$22909 863 1 2 790 INV_X2
* cell instance $23035 m0 *1 186.96,455
X$23035 778 849 2 1 916 AND2_X1
* cell instance $23036 m0 *1 187.72,455
X$23036 1 907 856 917 918 916 2 FA_X1
* cell instance $23039 m0 *1 191.71,455
X$23039 917 1 2 872 INV_X1
* cell instance $23040 m0 *1 192.09,455
X$23040 778 785 2 1 909 AND2_X1
* cell instance $23041 m0 *1 192.85,455
X$23041 776 873 2 1 919 AND2_X1
* cell instance $23094 r0 *1 189.05,455
X$23094 873 785 2 1 907 AND2_X1
* cell instance $23097 r0 *1 191.71,455
X$23097 1 919 908 920 909 931 2 FA_X1
* cell instance $23099 m0 *1 198.74,455
X$23099 678 732 2 1 875 AND2_X1
* cell instance $23103 m0 *1 204.06,455
X$23103 678 747 2 1 922 AND2_X1
* cell instance $23108 m0 *1 218.69,455
X$23108 926 900 2 1 928 XNOR2_X1
* cell instance $23112 m0 *1 223.82,455
X$23112 823 928 910 2 1 930 HA_X1
* cell instance $23116 m0 *1 232.75,455
X$23116 1 788 911 848 925 823 2 DFFR_X2
* cell instance $23117 m0 *1 236.93,455
X$23117 1 789 914 848 915 825 2 DFFR_X2
* cell instance $23164 r0 *1 218.69,455
X$23164 778 1 2 926 INV_X1
* cell instance $23169 r0 *1 224.2,455
X$23169 910 1 2 943 INV_X1
* cell instance $23177 r0 *1 234.27,455
X$23177 912 1 2 913 CLKBUF_X3
* cell instance $23181 r0 *1 239.4,455
X$23181 913 1 2 789 CLKBUF_X3
* cell instance $23182 r0 *1 240.35,455
X$23182 789 1 2 996 CLKBUF_X1
* cell instance $23321 m0 *1 192.66,457.8
X$23321 849 780 2 1 931 AND2_X1
* cell instance $23330 r0 *1 201.4,457.8
X$23330 778 776 2 1 949 AND2_X1
* cell instance $23331 r0 *1 202.16,457.8
X$23331 1 950 871 932 949 944 2 FA_X1
* cell instance $23332 m0 *1 204.63,457.8
X$23332 932 1 2 894 INV_X1
* cell instance $23338 r0 *1 205.2,457.8
X$23338 785 780 2 1 950 AND2_X1
* cell instance $23340 r0 *1 209,457.8
X$23340 1 873 2 879 BUF_X8
* cell instance $23343 r0 *1 214.89,457.8
X$23343 753 752 747 1 2 952 NOR3_X1
* cell instance $23346 r0 *1 216.79,457.8
X$23346 963 2 747 1 BUF_X4
* cell instance $23348 m0 *1 218.5,457.8
X$23348 962 942 926 1 2 903 NAND3_X2
* cell instance $23352 m0 *1 224.39,457.8
X$23352 943 939 941 1 929 2 AOI21_X1
* cell instance $23357 r0 *1 218.69,457.8
X$23357 732 952 2 1 955 XNOR2_X1
* cell instance $23360 r0 *1 220.78,457.8
X$23360 747 942 2 1 960 XNOR2_X1
* cell instance $23361 r0 *1 221.92,457.8
X$23361 957 1 2 966 INV_X1
* cell instance $23362 r0 *1 222.3,457.8
X$23362 862 958 957 2 1 933 HA_X1
* cell instance $23363 r0 *1 224.2,457.8
X$23363 967 933 974 2 959 1 OAI21_X1
* cell instance $23365 r0 *1 225.72,457.8
X$23365 945 1 2 946 INV_X1
* cell instance $23366 r0 *1 226.1,457.8
X$23366 956 959 946 1 940 2 AOI21_X1
* cell instance $23372 r0 *1 227.43,457.8
X$23372 940 954 934 2 941 1 OAI21_X1
* cell instance $23373 m0 *1 228,457.8
X$23373 938 1 2 939 INV_X1
* cell instance $23376 m0 *1 228.57,457.8
X$23376 756 964 934 2 1 938 HA_X1
* cell instance $23380 r0 *1 228.19,457.8
X$23380 953 1 2 956 INV_X1
* cell instance $23382 r0 *1 228.76,457.8
X$23382 825 955 953 2 1 954 HA_X1
* cell instance $23387 r0 *1 233.51,457.8
X$23387 951 822 1 2 972 NOR2_X1
* cell instance $23388 r0 *1 234.08,457.8
X$23388 935 948 2 1 951 XNOR2_X1
* cell instance $23389 r0 *1 235.22,457.8
X$23389 888 825 1 2 948 NAND2_X1
* cell instance $23392 r0 *1 237.69,457.8
X$23392 947 793 2 1 888 AND2_X1
* cell instance $23394 m0 *1 238.64,457.8
X$23394 937 868 2 1 936 AND2_X1
* cell instance $23400 m0 *1 241.49,457.8
X$23400 1 789 936 848 998 862 2 DFFR_X2
* cell instance $23441 r0 *1 238.64,457.8
X$23441 834 862 937 2 1 947 HA_X1
* cell instance $23565 m0 *1 196.84,460.6
X$23565 980 2 785 1 BUF_X4
* cell instance $23566 m0 *1 198.17,460.6
X$23566 981 2 778 1 BUF_X4
* cell instance $23569 m0 *1 203.3,460.6
X$23569 849 732 2 1 944 AND2_X1
* cell instance $23573 m0 *1 214.7,460.6
X$23573 961 2 732 1 BUF_X4
* cell instance $23574 m0 *1 216.03,460.6
X$23574 963 961 780 2 962 1 NOR3_X2
* cell instance $23576 m0 *1 217.55,460.6
X$23576 780 989 2 1 964 XNOR2_X1
* cell instance $23578 m0 *1 218.88,460.6
X$23578 962 975 965 1 2 900 NAND3_X1
* cell instance $23579 m0 *1 219.64,460.6
X$23579 975 965 958 2 1 942 HA_X1
* cell instance $23581 m0 *1 222.3,460.6
X$23581 753 1 2 975 INV_X1
* cell instance $23635 r0 *1 197.03,460.6
X$23635 982 1 2 678 BUF_X2
* cell instance $23642 r0 *1 217.36,460.6
X$23642 942 1 2 988 INV_X1
* cell instance $23643 r0 *1 217.74,460.6
X$23643 988 963 732 1 2 989 NOR3_X1
* cell instance $23644 r0 *1 218.5,460.6
X$23644 752 1 2 965 INV_X1
* cell instance $23647 r0 *1 220.59,460.6
X$23647 994 1 2 753 BUF_X2
* cell instance $23650 m0 *1 223.25,460.6
X$23650 966 971 973 1 967 2 AOI21_X1
* cell instance $23653 r0 *1 223.63,460.6
X$23653 992 975 976 2 1 973 HA_X1
* cell instance $23654 m0 *1 224.77,460.6
X$23654 793 960 974 2 1 945 HA_X1
* cell instance $23655 m0 *1 224.39,460.6
X$23655 976 1 2 971 INV_X1
* cell instance $23658 m0 *1 231.23,460.6
X$23658 1 788 972 848 935 756 2 DFFR_X2
* cell instance $23666 r0 *1 235.03,460.6
X$23666 1 789 977 848 992 834 2 DFFR_X2
* cell instance $23667 m0 *1 235.98,460.6
X$23667 822 834 1 2 977 NOR2_X1
* cell instance $23673 m0 *1 239.4,460.6
X$23673 968 822 1 2 970 NOR2_X1
* cell instance $23675 m0 *1 239.97,460.6
X$23675 947 969 1 2 968 XOR2_X1
* cell instance $23677 m0 *1 241.3,460.6
X$23677 1 789 970 848 969 793 2 DFFR_X2
* cell instance $23840 r0 *1 178.6,438.2
X$23840 566 486 2 1 633 AND2_X1
* cell instance $23845 r0 *1 183.73,438.2
X$23845 1 626 613 650 648 647 2 FA_X1
* cell instance $23846 m0 *1 184.3,438.2
X$23846 613 1 2 539 INV_X1
* cell instance $23849 m0 *1 187.72,438.2
X$23849 592 1 2 611 INV_X1
* cell instance $23853 m0 *1 190.57,438.2
X$23853 595 1 2 594 INV_X1
* cell instance $23856 m0 *1 193.23,438.2
X$23856 596 654 627 2 1 597 HA_X1
* cell instance $23863 r0 *1 187.34,438.2
X$23863 650 1 2 591 INV_X1
* cell instance $23865 r0 *1 187.91,438.2
X$23865 1 614 592 595 763 649 2 FA_X1
* cell instance $23868 r0 *1 194.18,438.2
X$23868 653 1 2 596 INV_X1
* cell instance $23871 r0 *1 196.27,438.2
X$23871 679 1 2 654 INV_X1
* cell instance $23874 r0 *1 202.92,438.2
X$23874 1 659 628 657 680 658 2 FA_X1
* cell instance $23875 r0 *1 205.96,438.2
X$23875 657 1 2 599 INV_X2
* cell instance $23879 m0 *1 210.71,438.2
X$23879 660 1 2 600 INV_X1
* cell instance $23882 m0 *1 215.08,438.2
X$23882 630 602 527 2 1 585 HA_X1
* cell instance $23891 r0 *1 211.47,438.2
X$23891 709 1 2 662 INV_X1
* cell instance $23892 r0 *1 211.85,438.2
X$23892 1 636 601 666 662 664 2 FA_X1
* cell instance $23894 r0 *1 215.08,438.2
X$23894 666 1 2 602 INV_X1
* cell instance $23898 r0 *1 217.55,438.2
X$23898 615 637 612 2 1 630 HA_X1
* cell instance $23900 r0 *1 222.49,438.2
X$23900 669 1 2 603 INV_X1
* cell instance $23904 r0 *1 224.96,438.2
X$23904 682 1 2 431 BUF_X2
* cell instance $23907 r0 *1 227.43,438.2
X$23907 632 606 617 2 1 673 HA_X1
* cell instance $23909 r0 *1 229.71,438.2
X$23909 673 1 2 639 INV_X1
* cell instance $23910 r0 *1 230.09,438.2
X$23910 616 672 674 2 1 640 HA_X1
* cell instance $23911 r0 *1 231.99,438.2
X$23911 617 1 2 683 INV_X1
* cell instance $23922 r0 *1 243.58,438.2
X$23922 565 676 609 608 619 2 1 AOI211_X2
* cell instance $23923 m0 *1 246.05,438.2
X$23923 572 570 1 2 608 OR2_X2
* cell instance $23924 m0 *1 243.96,438.2
X$23924 610 618 426 1 2 631 OR3_X4
* cell instance $23925 m0 *1 247,438.2
X$23925 629 572 431 1 2 610 NAND3_X1
* cell instance $23926 m0 *1 247.76,438.2
X$23926 624 629 2 1 621 AND2_X1
* cell instance $23929 r0 *1 245.29,438.2
X$23929 625 565 608 609 1 2 686 AOI22_X1
* cell instance $23932 r0 *1 247.38,438.2
X$23932 561 618 610 2 1 665 OAI21_X2
* cell instance $23933 r0 *1 248.71,438.2
X$23933 620 621 561 533 1 2 625 NAND4_X1
* cell instance $23935 r0 *1 250.04,438.2
X$23935 431 618 561 621 2 1 643 AND4_X1
* cell instance $23937 m0 *1 250.42,438.2
X$23937 621 561 475 1 2 656 NAND3_X1
* cell instance $23940 r0 *1 251.37,438.2
X$23940 656 622 1 2 655 NOR2_X1
* cell instance $23941 r0 *1 251.94,438.2
X$23941 622 1 2 618 BUF_X2
* cell instance $23942 r0 *1 252.7,438.2
X$23942 622 431 1 2 652 XNOR2_X2
* cell instance $23944 m0 *1 253.08,438.2
X$23944 652 1 2 620 BUF_X1
* cell instance $23980 r0 *1 254.6,438.2
X$23980 644 461 623 2 1 651 OAI21_X4
* cell instance $23981 r0 *1 257.07,438.2
X$23981 461 623 1 2 645 NOR2_X1
* cell instance $24083 m0 *1 187.53,418.6
X$24083 242 257 244 2 1 173 MUX2_X2
* cell instance $24084 m0 *1 189.24,418.6
X$24084 216 200 243 246 2 1 258 AND4_X1
* cell instance $24085 m0 *1 190.38,418.6
X$24085 201 147 245 2 1 247 AND3_X1
* cell instance $24087 m0 *1 191.52,418.6
X$24087 258 247 217 2 1 175 MUX2_X2
* cell instance $24091 m0 *1 195.7,418.6
X$24091 268 218 1 2 157 XNOR2_X2
* cell instance $24132 r0 *1 187.91,418.6
X$24132 159 216 1 2 242 NOR2_X1
* cell instance $24135 r0 *1 189.05,418.6
X$24135 243 246 2 1 244 AND2_X1
* cell instance $24136 r0 *1 189.81,418.6
X$24136 245 202 201 1 2 257 NOR3_X1
* cell instance $24137 r0 *1 190.57,418.6
X$24137 300 204 248 2 1 245 AND3_X1
* cell instance $24140 r0 *1 193.42,418.6
X$24140 204 248 2 1 249 AND2_X1
* cell instance $24141 r0 *1 194.18,418.6
X$24141 249 300 1 2 293 NOR2_X1
* cell instance $24142 r0 *1 194.75,418.6
X$24142 248 204 1 2 291 NAND2_X1
* cell instance $24143 r0 *1 195.32,418.6
X$24143 1 260 292 160 267 293 294 269 2 AOI222_X2
* cell instance $24144 r0 *1 197.98,418.6
X$24144 270 267 271 296 294 1 2 OAI211_X2
* cell instance $24145 m0 *1 198.17,418.6
X$24145 204 217 1 2 67 XNOR2_X2
* cell instance $24150 m0 *1 207.1,418.6
X$24150 1 129 34 177 67 219 250 240 2 OAI222_X2
* cell instance $24151 m0 *1 209.76,418.6
X$24151 67 241 2 1 265 XNOR2_X1
* cell instance $24152 m0 *1 210.9,418.6
X$24152 83 1 2 241 BUF_X1
* cell instance $24155 r0 *1 199.69,418.6
X$24155 271 296 1 2 292 OR2_X2
* cell instance $24160 r0 *1 205.77,418.6
X$24160 89 2 115 1 BUF_X4
* cell instance $24163 r0 *1 208.05,418.6
X$24163 250 219 34 115 298 83 1 2 OAI221_X2
* cell instance $24164 r0 *1 210.14,418.6
X$24164 134 177 2 1 298 AND2_X1
* cell instance $24165 r0 *1 210.9,418.6
X$24165 250 219 1 2 274 NOR2_X2
* cell instance $24168 m0 *1 214.89,418.6
X$24168 95 94 44 134 1 2 299 NAND4_X1
* cell instance $24169 m0 *1 217.36,418.6
X$24169 221 251 1 2 275 NOR2_X2
* cell instance $24170 m0 *1 218.31,418.6
X$24170 251 221 1 2 264 OR2_X1
* cell instance $24172 r0 *1 214.89,418.6
X$24172 299 273 265 274 2 1 119 OAI22_X2
* cell instance $24174 m0 *1 219.45,418.6
X$24174 44 94 117 2 1 266 AND3_X2
* cell instance $24175 m0 *1 220.59,418.6
X$24175 126 48 266 276 222 182 1 2 262 OAI33_X1
* cell instance $24176 m0 *1 221.92,418.6
X$24176 117 94 44 1 2 223 NAND3_X1
* cell instance $24177 m0 *1 222.68,418.6
X$24177 94 44 1 2 277 NAND2_X2
* cell instance $24183 r0 *1 221.92,418.6
X$24183 297 264 223 1 309 2 AOI21_X2
* cell instance $24184 r0 *1 223.25,418.6
X$24184 182 1 2 311 BUF_X1
* cell instance $24188 r0 *1 225.15,418.6
X$24188 195 312 95 2 1 185 AND3_X2
* cell instance $24191 m0 *1 228.57,418.6
X$24191 263 224 187 2 1 252 MUX2_X2
* cell instance $24192 m0 *1 227.81,418.6
X$24192 262 1 2 86 CLKBUF_X2
* cell instance $24193 m0 *1 230.28,418.6
X$24193 261 1 2 336 BUF_X2
* cell instance $24194 m0 *1 231.04,418.6
X$24194 252 226 188 1 2 239 OR3_X2
* cell instance $24195 m0 *1 232.18,418.6
X$24195 164 226 61 188 2 281 1 OR4_X2
* cell instance $24196 m0 *1 233.51,418.6
X$24196 238 227 1 2 236 NAND2_X2
* cell instance $24201 r0 *1 228.38,418.6
X$24201 195 1 2 297 INV_X1
* cell instance $24202 r0 *1 228.76,418.6
X$24202 75 207 143 1 280 2 NAND3_X4
* cell instance $24203 r0 *1 231.23,418.6
X$24203 1 164 295 61 188 259 2 NOR4_X4
* cell instance $24204 r0 *1 234.65,418.6
X$24204 226 1 2 190 BUF_X1
* cell instance $24205 r0 *1 235.22,418.6
X$24205 226 1 2 256 BUF_X1
* cell instance $24209 r0 *1 237.12,418.6
X$24209 228 209 210 165 289 290 1 2 OAI221_X2
* cell instance $24210 r0 *1 239.21,418.6
X$24210 1 374 290 236 288 2 AOI21_X4
* cell instance $24212 m0 *1 239.4,418.6
X$24212 230 282 210 213 2 254 1 NOR4_X2
* cell instance $24213 m0 *1 241.3,418.6
X$24213 1 145 229 231 211 288 2 NAND4_X4
* cell instance $24215 m0 *1 244.91,418.6
X$24215 255 212 254 209 233 232 1 2 OAI221_X2
* cell instance $24254 r0 *1 241.68,418.6
X$24254 1 286 235 236 288 2 AOI21_X4
* cell instance $24255 r0 *1 244.15,418.6
X$24255 283 255 256 2 287 1 NOR3_X2
* cell instance $24258 r0 *1 246.43,418.6
X$24258 229 287 1 2 285 XNOR2_X2
* cell instance $24400 r0 *1 188.67,415.8
X$24400 202 1 2 200 INV_X1
* cell instance $24401 m0 *1 188.86,415.8
X$24401 200 216 1 2 174 NOR2_X2
* cell instance $24406 r0 *1 189.05,415.8
X$24406 1 201 147 202 176 2 NOR3_X4
* cell instance $24408 m0 *1 192.66,415.8
X$24408 1 173 175 176 174 203 2 NOR4_X4
* cell instance $24414 m0 *1 201.59,415.8
X$24414 131 1 2 50 BUF_X2
* cell instance $24416 m0 *1 202.54,415.8
X$24416 177 179 178 1 2 98 AND3_X4
* cell instance $24417 m0 *1 204.63,415.8
X$24417 179 178 177 1 40 2 NAND3_X4
* cell instance $24418 m0 *1 207.1,415.8
X$24418 72 112 240 2 1 182 OAI21_X4
* cell instance $24421 m0 *1 210.52,415.8
X$24421 98 17 1 2 215 NAND2_X1
* cell instance $24422 m0 *1 211.09,415.8
X$24422 134 81 179 2 1 99 AND3_X2
* cell instance $24424 m0 *1 212.42,415.8
X$24424 98 180 114 1 2 205 NAND3_X1
* cell instance $24425 m0 *1 213.18,415.8
X$24425 114 1 2 198 BUF_X2
* cell instance $24426 m0 *1 213.94,415.8
X$24426 1 183 181 215 197 2 AOI21_X4
* cell instance $24432 r0 *1 194.18,415.8
X$24432 203 2 41 1 BUF_X4
* cell instance $24436 r0 *1 197.98,415.8
X$24436 204 270 1 2 179 XNOR2_X2
* cell instance $24440 r0 *1 203.49,415.8
X$24440 81 178 179 1 9 2 NAND3_X4
* cell instance $24442 r0 *1 207.48,415.8
X$24442 100 114 180 1 250 2 NAND3_X4
* cell instance $24444 r0 *1 211.47,415.8
X$24444 99 89 1 2 219 NAND2_X2
* cell instance $24446 r0 *1 212.8,415.8
X$24446 115 205 100 1 251 2 AOI21_X2
* cell instance $24447 r0 *1 214.13,415.8
X$24447 115 99 133 114 220 1 2 OAI211_X2
* cell instance $24448 r0 *1 215.84,415.8
X$24448 220 181 108 100 2 1 221 OAI22_X2
* cell instance $24449 r0 *1 217.55,415.8
X$24449 11 109 2 1 206 XNOR2_X1
* cell instance $24452 m0 *1 220.59,415.8
X$24452 199 183 184 1 2 NOR2_X4
* cell instance $24457 r0 *1 224.2,415.8
X$24457 206 2 142 1 BUF_X4
* cell instance $24460 m0 *1 225.72,415.8
X$24460 195 172 95 2 1 141 AND3_X2
* cell instance $24461 r0 *1 226.29,415.8
X$24461 185 55 206 1 2 263 NAND3_X1
* cell instance $24463 m0 *1 228.19,415.8
X$24463 196 186 193 2 1 207 MUX2_X2
* cell instance $24464 m0 *1 227.24,415.8
X$24464 142 55 185 2 1 196 AND3_X1
* cell instance $24465 m0 *1 229.9,415.8
X$24465 187 1 2 193 BUF_X1
* cell instance $24467 m0 *1 230.66,415.8
X$24467 120 46 195 1 2 225 NAND3_X1
* cell instance $24468 m0 *1 231.42,415.8
X$24468 187 1 2 192 BUF_X1
* cell instance $24469 m0 *1 231.99,415.8
X$24469 120 1 2 208 INV_X1
* cell instance $24471 m0 *1 232.56,415.8
X$24471 61 190 1 2 189 NOR2_X2
* cell instance $24472 m0 *1 233.51,415.8
X$24472 214 189 1 2 238 NAND2_X1
* cell instance $24473 m0 *1 234.08,415.8
X$24473 190 164 188 2 1 191 OAI21_X2
* cell instance $24479 r0 *1 228.19,415.8
X$24479 141 55 142 1 2 224 NAND3_X1
* cell instance $24481 r0 *1 229.71,415.8
X$24481 187 1 2 261 BUF_X2
* cell instance $24483 r0 *1 230.66,415.8
X$24483 1 208 239 209 214 189 2 AOI22_X4
* cell instance $24484 r0 *1 233.89,415.8
X$24484 239 208 1 2 227 NAND2_X1
* cell instance $24487 r0 *1 236.36,415.8
X$24487 228 209 165 210 2 1 235 OAI22_X2
* cell instance $24488 r0 *1 238.07,415.8
X$24488 168 237 191 2 1 228 AND3_X1
* cell instance $24489 r0 *1 239.02,415.8
X$24489 191 237 1 253 2 NAND2_X4
* cell instance $24490 r0 *1 240.73,415.8
X$24490 211 231 125 2 1 283 OAI21_X4
* cell instance $24531 r0 *1 243.2,415.8
X$24531 125 211 1 2 212 NAND2_X1
* cell instance $24533 r0 *1 244.15,415.8
X$24533 209 254 228 230 212 2 1 234 OAI221_X1
* cell instance $24534 r0 *1 245.29,415.8
X$24534 209 228 1 2 233 OR2_X1
* cell instance $24640 m0 *1 192.09,413
X$24640 147 1 2 159 INV_X1
* cell instance $24683 r0 *1 193.61,413
X$24683 1 111 174 176 175 173 2 OR4_X4
* cell instance $24685 m0 *1 195.13,413
X$24685 159 130 1 2 10 XNOR2_X2
* cell instance $24691 r0 *1 199.69,413
X$24691 160 2 52 1 BUF_X4
* cell instance $24692 r0 *1 201.02,413
X$24692 160 1 2 78 BUF_X1
* cell instance $24693 m0 *1 201.4,413
X$24693 131 2 132 1 BUF_X4
* cell instance $24695 m0 *1 202.73,413
X$24695 133 132 1 2 161 NAND2_X1
* cell instance $24697 m0 *1 203.49,413
X$24697 161 17 157 9 1 2 113 AOI211_X4
* cell instance $24698 m0 *1 205.58,413
X$24698 134 81 132 2 1 170 AND3_X1
* cell instance $24699 m0 *1 206.53,413
X$24699 154 133 115 1 2 152 NAND3_X2
* cell instance $24701 m0 *1 208.05,413
X$24701 134 135 132 2 1 154 AND3_X1
* cell instance $24705 m0 *1 213.75,413
X$24705 41 40 181 2 1 94 OAI21_X4
* cell instance $24706 m0 *1 216.22,413
X$24706 1 137 172 100 127 155 2 NAND4_X4
* cell instance $24707 m0 *1 219.64,413
X$24707 155 156 1 2 138 NOR2_X2
* cell instance $24710 m0 *1 223.82,413
X$24710 139 138 142 1 2 140 NAND3_X1
* cell instance $24713 m0 *1 229.14,413
X$24713 141 142 1 2 163 NAND2_X1
* cell instance $24714 m0 *1 229.71,413
X$24714 142 141 2 1 169 AND2_X1
* cell instance $24717 m0 *1 233.7,413
X$24717 164 151 148 2 104 1 OAI21_X1
* cell instance $24718 m0 *1 234.46,413
X$24718 1 168 144 122 165 149 2 OAI211_X4
* cell instance $24719 m0 *1 237.69,413
X$24719 145 143 120 1 2 167 NAND3_X1
* cell instance $24720 m0 *1 238.45,413
X$24720 167 104 146 1 166 2 AOI21_X1
* cell instance $24721 m0 *1 239.21,413
X$24721 121 124 1 2 229 XNOR2_X2
* cell instance $24724 m0 *1 242.82,413
X$24724 148 124 1 2 213 XNOR2_X2
* cell instance $24762 r0 *1 201.59,413
X$24762 67 177 115 1 2 150 NAND3_X1
* cell instance $24763 r0 *1 202.35,413
X$24763 52 132 2 96 1 AND2_X4
* cell instance $24764 r0 *1 204.06,413
X$24764 96 2 180 1 BUF_X4
* cell instance $24766 r0 *1 205.77,413
X$24766 170 17 11 2 1 153 OAI21_X2
* cell instance $24767 r0 *1 207.1,413
X$24767 1 132 177 134 179 26 2 NAND4_X4
* cell instance $24769 r0 *1 211.28,413
X$24769 134 81 179 52 2 1 136 AND4_X1
* cell instance $24770 r0 *1 212.42,413
X$24770 114 99 89 1 2 197 NAND3_X2
* cell instance $24771 r0 *1 213.75,413
X$24771 180 100 1 2 181 NAND2_X2
* cell instance $24772 r0 *1 214.7,413
X$24772 180 1 2 158 BUF_X2
* cell instance $24774 r0 *1 215.84,413
X$24774 1 199 198 108 100 2 AOI21_X4
* cell instance $24776 r0 *1 219.07,413
X$24776 1 155 156 199 45 183 2 OAI22_X4
* cell instance $24777 r0 *1 222.3,413
X$24777 139 138 1 2 171 NAND2_X1
* cell instance $24778 r0 *1 222.87,413
X$24778 1 187 184 138 139 2 AOI21_X4
* cell instance $24781 r0 *1 227.05,413
X$24781 142 55 141 2 1 186 AND3_X1
* cell instance $24782 r0 *1 228,413
X$24782 142 185 2 1 194 AND2_X1
* cell instance $24783 r0 *1 228.76,413
X$24783 185 142 1 2 162 NAND2_X1
* cell instance $24784 r0 *1 229.33,413
X$24784 162 163 187 2 1 164 MUX2_X2
* cell instance $24785 r0 *1 231.04,413
X$24785 194 169 192 2 1 123 MUX2_X2
* cell instance $24786 r0 *1 232.75,413
X$24786 151 164 1 2 214 NOR2_X2
* cell instance $24791 r0 *1 238.07,413
X$24791 102 143 123 1 2 237 NAND3_X2
* cell instance $24935 r0 *1 194.37,410.2
X$24935 147 130 1 2 107 XNOR2_X2
* cell instance $24938 r0 *1 200.83,410.2
X$24938 111 2 114 1 BUF_X4
* cell instance $24939 m0 *1 204.25,410.2
X$24939 107 2 100 1 BUF_X4
* cell instance $24940 m0 *1 200.83,410.2
X$24940 1 111 98 96 107 68 2 NAND4_X4
* cell instance $24941 m0 *1 205.58,410.2
X$24941 76 69 18 2 112 1 NOR3_X2
* cell instance $24942 m0 *1 206.91,410.2
X$24942 9 17 1 2 70 NOR2_X2
* cell instance $24943 m0 *1 207.86,410.2
X$24943 49 1 2 90 BUF_X2
* cell instance $24945 r0 *1 202.16,410.2
X$24945 128 2 139 1 BUF_X4
* cell instance $24946 r0 *1 203.49,410.2
X$24946 1 150 82 128 152 153 19 113 2 AOI222_X2
* cell instance $24947 r0 *1 206.15,410.2
X$24947 1 152 153 72 113 19 2 AOI22_X4
* cell instance $24948 m0 *1 210.33,410.2
X$24948 76 18 1 2 129 NAND2_X1
* cell instance $24949 m0 *1 209,410.2
X$24949 133 135 115 1 2 97 NAND3_X2
* cell instance $24956 r0 *1 211.47,410.2
X$24956 100 114 115 136 1 116 2 NAND4_X2
* cell instance $24957 r0 *1 213.18,410.2
X$24957 114 99 115 158 1 137 2 NAND4_X2
* cell instance $24958 m0 *1 214.51,410.2
X$24958 12 38 100 1 2 126 NOR3_X1
* cell instance $24959 m0 *1 213.56,410.2
X$24959 98 115 1 2 12 NAND2_X2
* cell instance $24960 m0 *1 215.27,410.2
X$24960 10 110 18 2 101 1 OAI21_X1
* cell instance $24963 r0 *1 215.08,410.2
X$24963 157 18 26 2 1 127 OAI21_X2
* cell instance $24964 m0 *1 216.6,410.2
X$24964 100 114 1 2 84 NAND2_X1
* cell instance $24966 m0 *1 217.17,410.2
X$24966 101 116 108 1 2 106 NAND3_X2
* cell instance $24969 r0 *1 216.41,410.2
X$24969 41 1 2 110 BUF_X1
* cell instance $24970 r0 *1 216.98,410.2
X$24970 108 116 101 2 1 156 AND3_X1
* cell instance $24971 r0 *1 217.93,410.2
X$24971 100 127 137 172 2 1 118 AND4_X2
* cell instance $25223 m0 *1 213.56,401.8
X$25223 15 1 2 16 BUF_X1
* cell instance $25283 r0 *1 206.91,401.8
X$25283 49 1 2 64 BUF_X1
* cell instance $25286 r0 *1 208.43,401.8
X$25286 17 2 18 1 BUF_X4
* cell instance $25287 r0 *1 209.76,401.8
X$25287 23 9 17 2 8 1 NOR3_X2
* cell instance $25289 r0 *1 211.47,401.8
X$25289 38 10 1 2 37 NOR2_X1
* cell instance $25292 r0 *1 212.61,401.8
X$25292 10 15 19 1 2 NOR2_X4
* cell instance $25293 r0 *1 214.32,401.8
X$25293 18 11 10 16 2 1 20 OAI22_X2
* cell instance $25295 r0 *1 216.22,401.8
X$25295 11 18 1 2 22 NAND2_X1
* cell instance $25300 r0 *1 221.16,401.8
X$25300 14 12 1 2 13 OR2_X1
* cell instance $25301 r0 *1 221.92,401.8
X$25301 12 14 1 2 32 NAND2_X1
* cell instance $28793 r0 *1 458.66,264.6
X$28793 7 1 2 6 BUF_X1
* cell instance $32405 m0 *1 193.61,463.4
X$32405 1 776 2 978 BUF_X8
* cell instance $32406 m0 *1 196.08,463.4
X$32406 979 2 849 1 BUF_X4
* cell instance $32409 m0 *1 200.64,463.4
X$32409 1 780 2 983 BUF_X8
* cell instance $32412 m0 *1 209.38,463.4
X$32412 984 1 2 710 BUF_X2
.ENDS clock_divider

* cell AND3_X2
* pin A1
* pin A2
* pin A3
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND3_X2 1 2 3 5 6 7
* net 1 A1
* net 2 A2
* net 3 A3
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 5 1 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 4 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 4 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $6 r0 *1 0.17,0.2975 NMOS_VTL
M$6 9 1 4 6 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $7 r0 *1 0.36,0.2975 NMOS_VTL
M$7 8 2 9 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.55,0.2975 NMOS_VTL
M$8 6 3 8 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.74,0.2975 NMOS_VTL
M$9 7 4 6 6 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS AND3_X2

* cell NAND4_X2
* pin A3
* pin A2
* pin A1
* pin A4
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT NAND4_X2 1 2 3 4 5 6 7
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 A4
* net 5 PWELL,VSS
* net 6 ZN
* net 7 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 6 4 7 7 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.11025P PS=2.24U PD=2.24U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 7 1 6 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 6 2 7 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 7 3 6 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $9 r0 *1 0.21,0.2975 NMOS_VTL
M$9 13 4 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $10 r0 *1 0.4,0.2975 NMOS_VTL
M$10 12 1 13 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.59,0.2975 NMOS_VTL
M$11 11 2 12 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 0.78,0.2975 NMOS_VTL
M$12 6 3 11 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.97,0.2975 NMOS_VTL
M$13 8 3 6 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 1.16,0.2975 NMOS_VTL
M$14 10 2 8 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 1.35,0.2975 NMOS_VTL
M$15 9 1 10 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 1.54,0.2975 NMOS_VTL
M$16 5 4 9 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND4_X2

* cell AND4_X4
* pin PWELL,VSS
* pin A4
* pin A3
* pin A2
* pin A1
* pin ZN
* pin NWELL,VDD
.SUBCKT AND4_X4 1 2 3 4 6 7 14
* net 1 PWELL,VSS
* net 2 A4
* net 3 A3
* net 4 A2
* net 6 A1
* net 7 ZN
* net 14 NWELL,VDD
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 5 2 14 14 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 14 3 5 14 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $3 r0 *1 0.565,0.995 PMOS_VTL
M$3 5 4 14 14 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $4 r0 *1 0.755,0.995 PMOS_VTL
M$4 14 6 5 14 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $9 r0 *1 1.705,0.995 PMOS_VTL
M$9 7 5 14 14 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $13 r0 *1 0.185,0.2975 NMOS_VTL
M$13 8 2 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $14 r0 *1 0.375,0.2975 NMOS_VTL
M$14 9 3 8 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 0.565,0.2975 NMOS_VTL
M$15 10 4 9 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 0.755,0.2975 NMOS_VTL
M$16 5 6 10 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $17 r0 *1 0.945,0.2975 NMOS_VTL
M$17 12 6 5 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $18 r0 *1 1.135,0.2975 NMOS_VTL
M$18 11 4 12 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 1.325,0.2975 NMOS_VTL
M$19 13 3 11 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $20 r0 *1 1.515,0.2975 NMOS_VTL
M$20 1 2 13 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $21 r0 *1 1.705,0.2975 NMOS_VTL
M$21 7 5 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS AND4_X4

* cell AND4_X2
* pin A1
* pin A2
* pin A3
* pin A4
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND4_X2 1 2 3 4 6 7 8
* net 1 A1
* net 2 A2
* net 3 A3
* net 4 A4
* net 6 NWELL,VDD
* net 7 PWELL,VSS
* net 8 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 5 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 6 2 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 5 3 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 6 4 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 8 5 6 6 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $7 r0 *1 0.17,0.2975 NMOS_VTL
M$7 11 1 5 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $8 r0 *1 0.36,0.2975 NMOS_VTL
M$8 10 2 11 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.55,0.2975 NMOS_VTL
M$9 9 3 10 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.74,0.2975 NMOS_VTL
M$10 7 4 9 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.93,0.2975 NMOS_VTL
M$11 8 5 7 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS AND4_X2

* cell CLKBUF_X2
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT CLKBUF_X2 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.17,0.1875 NMOS_VTL
M$4 3 1 2 3 NMOS_VTL L=0.05U W=0.195U AS=0.020475P AD=0.01365P PS=0.6U PD=0.335U
* device instance $5 r0 *1 0.36,0.1875 NMOS_VTL
M$5 5 2 3 3 NMOS_VTL L=0.05U W=0.39U AS=0.0273P AD=0.034125P PS=0.67U PD=0.935U
.ENDS CLKBUF_X2

* cell DFFR_X1
* pin PWELL,VSS
* pin CK
* pin QN
* pin Q
* pin D
* pin RN
* pin NWELL,VDD
.SUBCKT DFFR_X1 1 3 8 9 16 18 19
* net 1 PWELL,VSS
* net 3 CK
* net 8 QN
* net 9 Q
* net 16 D
* net 18 RN
* net 19 NWELL,VDD
* device instance $1 r0 *1 3.41,0.995 PMOS_VTL
M$1 19 6 8 19 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 3.6,0.995 PMOS_VTL
M$2 9 7 19 19 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 2.455,1.04 PMOS_VTL
M$3 21 4 6 19 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.0063P PS=0.455U
+ PD=0.23U
* device instance $4 r0 *1 2.645,1.04 PMOS_VTL
M$4 19 7 21 19 PMOS_VTL L=0.05U W=0.09U AS=0.0063P AD=0.014175P PS=0.23U
+ PD=0.455U
* device instance $5 r0 *1 1.815,1.0125 PMOS_VTL
M$5 19 5 17 19 PMOS_VTL L=0.05U W=0.315U AS=0.03465P AD=0.033075P PS=0.85U
+ PD=0.525U
* device instance $6 r0 *1 2.075,1.0125 PMOS_VTL
M$6 23 5 19 19 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.525U
+ PD=0.455U
* device instance $7 r0 *1 2.265,1.0125 PMOS_VTL
M$7 6 2 23 19 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.014175P PS=0.455U
+ PD=0.455U
* device instance $8 r0 *1 2.835,1.1525 PMOS_VTL
M$8 7 18 19 19 PMOS_VTL L=0.05U W=0.315U AS=0.014175P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $9 r0 *1 3.025,1.1525 PMOS_VTL
M$9 19 6 7 19 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.033075P PS=0.455U
+ PD=0.84U
* device instance $10 r0 *1 1.08,1.065 PMOS_VTL
M$10 20 2 5 19 PMOS_VTL L=0.05U W=0.09U AS=0.01785P AD=0.0063P PS=0.56U PD=0.23U
* device instance $11 r0 *1 1.27,1.065 PMOS_VTL
M$11 19 17 20 19 PMOS_VTL L=0.05U W=0.09U AS=0.0063P AD=0.0063P PS=0.23U
+ PD=0.23U
* device instance $12 r0 *1 1.46,1.065 PMOS_VTL
M$12 20 18 19 19 PMOS_VTL L=0.05U W=0.09U AS=0.0063P AD=0.01035P PS=0.23U
+ PD=0.41U
* device instance $13 r0 *1 0.7,1.05 PMOS_VTL
M$13 22 16 19 19 PMOS_VTL L=0.05U W=0.42U AS=0.0441P AD=0.0294P PS=1.05U
+ PD=0.56U
* device instance $14 r0 *1 0.89,1.05 PMOS_VTL
M$14 5 4 22 19 PMOS_VTL L=0.05U W=0.42U AS=0.0294P AD=0.01785P PS=0.56U PD=0.56U
* device instance $15 r0 *1 0.17,1.1525 PMOS_VTL
M$15 19 3 2 19 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $16 r0 *1 0.36,1.1525 PMOS_VTL
M$16 4 2 19 19 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.033075P PS=0.455U
+ PD=0.84U
* device instance $17 r0 *1 3.41,0.2975 NMOS_VTL
M$17 1 6 8 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $18 r0 *1 3.6,0.2975 NMOS_VTL
M$18 9 7 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
* device instance $19 r0 *1 1.08,0.35 NMOS_VTL
M$19 12 4 5 1 NMOS_VTL L=0.05U W=0.09U AS=0.012775P AD=0.0063P PS=0.415U
+ PD=0.23U
* device instance $20 r0 *1 1.27,0.35 NMOS_VTL
M$20 11 17 12 1 NMOS_VTL L=0.05U W=0.09U AS=0.0063P AD=0.0063P PS=0.23U PD=0.23U
* device instance $21 r0 *1 1.46,0.35 NMOS_VTL
M$21 1 18 11 1 NMOS_VTL L=0.05U W=0.09U AS=0.0063P AD=0.00945P PS=0.23U PD=0.39U
* device instance $22 r0 *1 0.7,0.3525 NMOS_VTL
M$22 10 16 1 1 NMOS_VTL L=0.05U W=0.275U AS=0.028875P AD=0.01925P PS=0.76U
+ PD=0.415U
* device instance $23 r0 *1 0.89,0.3525 NMOS_VTL
M$23 5 2 10 1 NMOS_VTL L=0.05U W=0.275U AS=0.01925P AD=0.012775P PS=0.415U
+ PD=0.415U
* device instance $24 r0 *1 2.455,0.26 NMOS_VTL
M$24 15 2 6 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.0063P PS=0.35U PD=0.23U
* device instance $25 r0 *1 2.645,0.26 NMOS_VTL
M$25 1 7 15 1 NMOS_VTL L=0.05U W=0.09U AS=0.0063P AD=0.0105P PS=0.23U PD=0.35U
* device instance $26 r0 *1 1.815,0.32 NMOS_VTL
M$26 1 5 17 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.02205P PS=0.63U PD=0.42U
* device instance $27 r0 *1 2.075,0.32 NMOS_VTL
M$27 14 5 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.42U PD=0.35U
* device instance $28 r0 *1 2.265,0.32 NMOS_VTL
M$28 6 4 14 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0105P PS=0.35U PD=0.35U
* device instance $29 r0 *1 2.835,0.32 NMOS_VTL
M$29 13 18 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0105P AD=0.0147P PS=0.35U PD=0.35U
* device instance $30 r0 *1 3.025,0.32 NMOS_VTL
M$30 7 6 13 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.02205P PS=0.35U PD=0.63U
* device instance $31 r0 *1 0.17,0.245 NMOS_VTL
M$31 1 3 2 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $32 r0 *1 0.36,0.245 NMOS_VTL
M$32 4 2 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.02205P PS=0.35U PD=0.63U
.ENDS DFFR_X1

* cell BUF_X8
* pin PWELL,VSS
* pin Z
* pin NWELL,VDD
* pin A
.SUBCKT BUF_X8 1 3 4 5
* net 1 PWELL,VSS
* net 3 Z
* net 4 NWELL,VDD
* net 5 A
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 2 5 4 4 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 3 2 4 4 PMOS_VTL L=0.05U W=5.04U AS=0.3528P AD=0.37485P PS=6.16U PD=6.86U
* device instance $13 r0 *1 0.17,0.2975 NMOS_VTL
M$13 2 5 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $17 r0 *1 0.93,0.2975 NMOS_VTL
M$17 3 2 1 1 NMOS_VTL L=0.05U W=3.32U AS=0.2324P AD=0.246925P PS=4.44U PD=4.925U
.ENDS BUF_X8

* cell OAI33_X1
* pin B3
* pin B2
* pin B1
* pin A1
* pin A2
* pin A3
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OAI33_X1 1 2 3 4 5 6 7 8 10
* net 1 B3
* net 2 B2
* net 3 B1
* net 4 A1
* net 5 A2
* net 6 A3
* net 7 PWELL,VSS
* net 8 NWELL,VDD
* net 10 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 14 1 8 8 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 13 2 14 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.565,0.995 PMOS_VTL
M$3 10 3 13 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.755,0.995 PMOS_VTL
M$4 12 4 10 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.945,0.995 PMOS_VTL
M$5 11 5 12 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.135,0.995 PMOS_VTL
M$6 8 6 11 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.185,0.2975 NMOS_VTL
M$7 9 1 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $8 r0 *1 0.375,0.2975 NMOS_VTL
M$8 7 2 9 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.565,0.2975 NMOS_VTL
M$9 9 3 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.755,0.2975 NMOS_VTL
M$10 10 4 9 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.945,0.2975 NMOS_VTL
M$11 9 5 10 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 1.135,0.2975 NMOS_VTL
M$12 10 6 9 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI33_X1

* cell FA_X1
* pin PWELL,VSS
* pin B
* pin CO
* pin S
* pin CI
* pin A
* pin NWELL,VDD
.SUBCKT FA_X1 1 2 3 8 11 12 14
* net 1 PWELL,VSS
* net 2 B
* net 3 CO
* net 8 S
* net 11 CI
* net 12 A
* net 14 NWELL,VDD
* device instance $1 r0 *1 0.385,1.0275 PMOS_VTL
M$1 17 2 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $2 r0 *1 0.575,1.0275 PMOS_VTL
M$2 4 12 17 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.765,1.0275 PMOS_VTL
M$3 15 11 4 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02265P PS=0.455U
+ PD=0.535U
* device instance $4 r0 *1 0.96,1.1025 PMOS_VTL
M$4 14 12 15 14 PMOS_VTL L=0.05U W=0.315U AS=0.02265P AD=0.02205P PS=0.535U
+ PD=0.455U
* device instance $5 r0 *1 1.15,1.1025 PMOS_VTL
M$5 15 2 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.033075P PS=0.455U
+ PD=0.84U
* device instance $6 r0 *1 0.195,0.995 PMOS_VTL
M$6 14 4 3 14 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.033075P PS=1.47U
+ PD=0.77U
* device instance $7 r0 *1 1.49,1.1525 PMOS_VTL
M$7 16 2 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $8 r0 *1 1.68,1.1525 PMOS_VTL
M$8 14 11 16 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $9 r0 *1 1.87,1.1525 PMOS_VTL
M$9 16 12 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $10 r0 *1 2.06,1.1525 PMOS_VTL
M$10 7 4 16 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.023625P PS=0.455U
+ PD=0.465U
* device instance $11 r0 *1 2.26,1.1525 PMOS_VTL
M$11 18 11 7 14 PMOS_VTL L=0.05U W=0.315U AS=0.023625P AD=0.02205P PS=0.465U
+ PD=0.455U
* device instance $12 r0 *1 2.45,1.1525 PMOS_VTL
M$12 19 2 18 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $13 r0 *1 2.64,1.1525 PMOS_VTL
M$13 19 12 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $14 r0 *1 2.83,0.995 PMOS_VTL
M$14 8 7 14 14 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U
+ PD=1.47U
* device instance $15 r0 *1 1.49,0.195 NMOS_VTL
M$15 6 2 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $16 r0 *1 1.68,0.195 NMOS_VTL
M$16 1 11 6 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $17 r0 *1 1.87,0.195 NMOS_VTL
M$17 6 12 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $18 r0 *1 2.06,0.195 NMOS_VTL
M$18 7 4 6 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.01575P PS=0.35U PD=0.36U
* device instance $19 r0 *1 2.26,0.195 NMOS_VTL
M$19 9 11 7 1 NMOS_VTL L=0.05U W=0.21U AS=0.01575P AD=0.0147P PS=0.36U PD=0.35U
* device instance $20 r0 *1 2.45,0.195 NMOS_VTL
M$20 10 2 9 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $21 r0 *1 2.64,0.195 NMOS_VTL
M$21 1 12 10 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
* device instance $22 r0 *1 2.83,0.2975 NMOS_VTL
M$22 8 7 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
* device instance $23 r0 *1 0.385,0.32 NMOS_VTL
M$23 13 2 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.021875P AD=0.0147P PS=0.555U
+ PD=0.35U
* device instance $24 r0 *1 0.575,0.32 NMOS_VTL
M$24 4 12 13 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $25 r0 *1 0.765,0.32 NMOS_VTL
M$25 5 11 4 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.015225P PS=0.35U
+ PD=0.355U
* device instance $26 r0 *1 0.96,0.32 NMOS_VTL
M$26 1 12 5 1 NMOS_VTL L=0.05U W=0.21U AS=0.015225P AD=0.0147P PS=0.355U
+ PD=0.35U
* device instance $27 r0 *1 1.15,0.32 NMOS_VTL
M$27 5 2 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.02205P PS=0.35U PD=0.63U
* device instance $28 r0 *1 0.195,0.2975 NMOS_VTL
M$28 1 4 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.021875P PS=1.04U
+ PD=0.555U
.ENDS FA_X1

* cell AND3_X4
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT AND3_X4 1 2 3 5 6 7
* net 1 A3
* net 2 A2
* net 3 A1
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 6 6 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 6 2 4 6 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 4 3 6 6 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $7 r0 *1 1.31,0.995 PMOS_VTL
M$7 7 4 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $11 r0 *1 0.17,0.2975 NMOS_VTL
M$11 11 1 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $12 r0 *1 0.36,0.2975 NMOS_VTL
M$12 10 2 11 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.55,0.2975 NMOS_VTL
M$13 4 3 10 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 0.74,0.2975 NMOS_VTL
M$14 8 3 4 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 0.93,0.2975 NMOS_VTL
M$15 9 2 8 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 1.12,0.2975 NMOS_VTL
M$16 5 1 9 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $17 r0 *1 1.31,0.2975 NMOS_VTL
M$17 7 4 5 5 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS AND3_X4

* cell AND2_X4
* pin A2
* pin A1
* pin NWELL,VDD
* pin ZN
* pin PWELL,VSS
.SUBCKT AND2_X4 1 2 4 5 6
* net 1 A2
* net 2 A1
* net 4 NWELL,VDD
* net 5 ZN
* net 6 PWELL,VSS
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 3 1 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 4 2 3 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 5 3 4 4 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $9 r0 *1 0.17,0.2975 NMOS_VTL
M$9 8 1 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $10 r0 *1 0.36,0.2975 NMOS_VTL
M$10 3 2 8 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.55,0.2975 NMOS_VTL
M$11 7 2 3 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 0.74,0.2975 NMOS_VTL
M$12 6 1 7 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.93,0.2975 NMOS_VTL
M$13 5 3 6 6 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS AND2_X4

* cell AOI222_X2
* pin PWELL,VSS
* pin C2
* pin C1
* pin ZN
* pin B2
* pin B1
* pin A1
* pin A2
* pin NWELL,VDD
.SUBCKT AOI222_X2 1 2 3 4 5 6 8 9 16
* net 1 PWELL,VSS
* net 2 C2
* net 3 C1
* net 4 ZN
* net 5 B2
* net 6 B1
* net 8 A1
* net 9 A2
* net 16 NWELL,VDD
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 16 2 15 16 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 15 3 16 16 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 17 5 15 16 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 15 6 17 16 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $9 r0 *1 1.875,0.995 PMOS_VTL
M$9 4 8 17 16 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $11 r0 *1 2.255,0.995 PMOS_VTL
M$11 4 9 17 16 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $13 r0 *1 1.875,0.2975 NMOS_VTL
M$13 4 8 7 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $14 r0 *1 2.065,0.2975 NMOS_VTL
M$14 11 8 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 2.255,0.2975 NMOS_VTL
M$15 1 9 11 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 2.445,0.2975 NMOS_VTL
M$16 7 9 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
* device instance $17 r0 *1 0.17,0.2975 NMOS_VTL
M$17 10 2 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $18 r0 *1 0.36,0.2975 NMOS_VTL
M$18 4 3 10 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 0.55,0.2975 NMOS_VTL
M$19 12 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $20 r0 *1 0.74,0.2975 NMOS_VTL
M$20 1 2 12 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $21 r0 *1 0.93,0.2975 NMOS_VTL
M$21 13 5 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $22 r0 *1 1.12,0.2975 NMOS_VTL
M$22 4 6 13 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $23 r0 *1 1.31,0.2975 NMOS_VTL
M$23 14 6 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $24 r0 *1 1.5,0.2975 NMOS_VTL
M$24 1 5 14 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI222_X2

* cell NOR3_X2
* pin A3
* pin A2
* pin A1
* pin NWELL,VDD
* pin ZN
* pin PWELL,VSS
.SUBCKT NOR3_X2 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 NWELL,VDD
* net 5 ZN
* net 6 PWELL,VSS
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 10 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 9 2 10 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 5 3 9 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 8 3 5 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 7 2 8 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 4 1 7 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.21,0.2975 NMOS_VTL
M$7 5 1 6 6 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.072625P PS=1.595U
+ PD=1.595U
* device instance $8 r0 *1 0.4,0.2975 NMOS_VTL
M$8 6 2 5 6 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $9 r0 *1 0.59,0.2975 NMOS_VTL
M$9 5 3 6 6 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
.ENDS NOR3_X2

* cell OAI221_X1
* pin B2
* pin B1
* pin A
* pin C2
* pin C1
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT OAI221_X1 1 2 3 4 5 7 8 9
* net 1 B2
* net 2 B1
* net 3 A
* net 4 C2
* net 5 C1
* net 7 NWELL,VDD
* net 8 PWELL,VSS
* net 9 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 12 1 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 9 2 12 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 7 3 9 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 11 4 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 9 5 11 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.17,0.2975 NMOS_VTL
M$6 8 1 6 8 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $7 r0 *1 0.36,0.2975 NMOS_VTL
M$7 6 2 8 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.55,0.2975 NMOS_VTL
M$8 10 3 6 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.74,0.2975 NMOS_VTL
M$9 9 4 10 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.93,0.2975 NMOS_VTL
M$10 10 5 9 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI221_X1

* cell NOR4_X2
* pin A3
* pin A2
* pin A1
* pin A4
* pin NWELL,VDD
* pin ZN
* pin PWELL,VSS
.SUBCKT NOR4_X2 1 2 3 4 5 6 7
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 A4
* net 5 NWELL,VDD
* net 6 ZN
* net 7 PWELL,VSS
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 12 4 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 11 1 12 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 10 2 11 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 6 3 10 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 9 3 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 13 2 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.35,0.995 PMOS_VTL
M$7 8 1 13 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.54,0.995 PMOS_VTL
M$8 5 4 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 0.21,0.2975 NMOS_VTL
M$9 6 4 7 7 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.072625P PS=1.595U
+ PD=1.595U
* device instance $10 r0 *1 0.4,0.2975 NMOS_VTL
M$10 7 1 6 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $11 r0 *1 0.59,0.2975 NMOS_VTL
M$11 6 2 7 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $12 r0 *1 0.78,0.2975 NMOS_VTL
M$12 7 3 6 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
.ENDS NOR4_X2

* cell OAI211_X4
* pin PWELL,VSS
* pin A
* pin B
* pin C2
* pin ZN
* pin C1
* pin NWELL,VDD
.SUBCKT OAI211_X4 1 3 4 5 6 7 12
* net 1 PWELL,VSS
* net 3 A
* net 4 B
* net 5 C2
* net 6 ZN
* net 7 C1
* net 12 NWELL,VDD
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 6 3 12 12 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 12 4 6 12 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.1764P PS=3.08U PD=3.08U
* device instance $9 r0 *1 1.69,0.995 PMOS_VTL
M$9 13 5 12 12 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $10 r0 *1 1.88,0.995 PMOS_VTL
M$10 6 7 13 12 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $11 r0 *1 2.07,0.995 PMOS_VTL
M$11 15 7 6 12 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $12 r0 *1 2.26,0.995 PMOS_VTL
M$12 12 5 15 12 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $13 r0 *1 2.45,0.995 PMOS_VTL
M$13 14 5 12 12 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $14 r0 *1 2.64,0.995 PMOS_VTL
M$14 6 7 14 12 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $15 r0 *1 2.83,0.995 PMOS_VTL
M$15 16 7 6 12 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $16 r0 *1 3.02,0.995 PMOS_VTL
M$16 12 5 16 12 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U
+ PD=1.47U
* device instance $17 r0 *1 0.17,0.2975 NMOS_VTL
M$17 8 3 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $18 r0 *1 0.36,0.2975 NMOS_VTL
M$18 1 4 8 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 0.55,0.2975 NMOS_VTL
M$19 10 4 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $20 r0 *1 0.74,0.2975 NMOS_VTL
M$20 2 3 10 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $21 r0 *1 0.93,0.2975 NMOS_VTL
M$21 9 3 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $22 r0 *1 1.12,0.2975 NMOS_VTL
M$22 1 4 9 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $23 r0 *1 1.31,0.2975 NMOS_VTL
M$23 11 4 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $24 r0 *1 1.5,0.2975 NMOS_VTL
M$24 2 3 11 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $25 r0 *1 1.69,0.2975 NMOS_VTL
M$25 6 5 2 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
* device instance $26 r0 *1 1.88,0.2975 NMOS_VTL
M$26 2 7 6 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.1162P PS=2.22U PD=2.22U
.ENDS OAI211_X4

* cell NAND4_X4
* pin PWELL,VSS
* pin A3
* pin A4
* pin A1
* pin A2
* pin ZN
* pin NWELL,VDD
.SUBCKT NAND4_X4 1 2 3 7 8 9 10
* net 1 PWELL,VSS
* net 2 A3
* net 3 A4
* net 7 A1
* net 8 A2
* net 9 ZN
* net 10 NWELL,VDD
* device instance $1 r0 *1 0.215,0.995 PMOS_VTL
M$1 10 7 9 10 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.975,0.995 PMOS_VTL
M$5 10 8 9 10 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.22365P PS=3.08U PD=3.23U
* device instance $9 r0 *1 1.885,0.995 PMOS_VTL
M$9 10 2 9 10 PMOS_VTL L=0.05U W=2.52U AS=0.22365P AD=0.1764P PS=3.23U PD=3.08U
* device instance $13 r0 *1 2.645,0.995 PMOS_VTL
M$13 10 3 9 10 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $17 r0 *1 1.885,0.2975 NMOS_VTL
M$17 5 2 6 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $21 r0 *1 2.645,0.2975 NMOS_VTL
M$21 1 3 6 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
* device instance $25 r0 *1 0.215,0.2975 NMOS_VTL
M$25 9 7 4 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $29 r0 *1 0.975,0.2975 NMOS_VTL
M$29 5 8 4 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS NAND4_X4

* cell NAND2_X4
* pin A2
* pin A1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT NAND2_X4 1 2 4 5 6
* net 1 A2
* net 2 A1
* net 4 PWELL,VSS
* net 5 ZN
* net 6 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 5 1 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 5 2 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $9 r0 *1 0.21,0.2975 NMOS_VTL
M$9 4 1 3 4 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $13 r0 *1 0.97,0.2975 NMOS_VTL
M$13 5 2 3 4 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS NAND2_X4

* cell NAND2_X2
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND2_X2 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.195,0.995 PMOS_VTL
M$1 5 1 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.11025P PS=2.24U PD=2.24U
* device instance $2 r0 *1 0.385,0.995 PMOS_VTL
M$2 4 2 5 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $5 r0 *1 0.195,0.2975 NMOS_VTL
M$5 7 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.385,0.2975 NMOS_VTL
M$6 5 2 7 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.575,0.2975 NMOS_VTL
M$7 6 2 5 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.765,0.2975 NMOS_VTL
M$8 3 1 6 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND2_X2

* cell NAND3_X4
* pin A2
* pin A1
* pin A3
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT NAND3_X4 1 2 3 4 5 6
* net 1 A2
* net 2 A1
* net 3 A3
* net 4 PWELL,VSS
* net 5 ZN
* net 6 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 5 3 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.19845P PS=3.78U PD=3.78U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 6 1 5 6 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.1764P PS=3.08U PD=3.08U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 5 2 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.1764P PS=3.08U PD=3.08U
* device instance $13 r0 *1 0.21,0.2975 NMOS_VTL
M$13 13 3 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $14 r0 *1 0.4,0.2975 NMOS_VTL
M$14 12 1 13 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 0.59,0.2975 NMOS_VTL
M$15 5 2 12 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 0.78,0.2975 NMOS_VTL
M$16 10 2 5 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $17 r0 *1 0.97,0.2975 NMOS_VTL
M$17 8 1 10 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $18 r0 *1 1.16,0.2975 NMOS_VTL
M$18 4 3 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 1.35,0.2975 NMOS_VTL
M$19 9 3 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $20 r0 *1 1.54,0.2975 NMOS_VTL
M$20 7 1 9 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $21 r0 *1 1.73,0.2975 NMOS_VTL
M$21 5 2 7 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $22 r0 *1 1.92,0.2975 NMOS_VTL
M$22 14 2 5 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $23 r0 *1 2.11,0.2975 NMOS_VTL
M$23 11 1 14 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $24 r0 *1 2.3,0.2975 NMOS_VTL
M$24 4 3 11 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND3_X4

* cell OR3_X1
* pin A1
* pin A2
* pin A3
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR3_X1 1 2 3 5 6 7
* net 1 A1
* net 2 A2
* net 3 A3
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 9 1 4 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 8 2 9 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 8 3 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 4 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.195 NMOS_VTL
M$5 5 1 4 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $6 r0 *1 0.36,0.195 NMOS_VTL
M$6 4 2 5 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $7 r0 *1 0.55,0.195 NMOS_VTL
M$7 5 3 4 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $8 r0 *1 0.74,0.2975 NMOS_VTL
M$8 7 4 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OR3_X1

* cell MUX2_X1
* pin A
* pin S
* pin B
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT MUX2_X1 1 2 3 5 6 8
* net 1 A
* net 2 S
* net 3 B
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 8 Z
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 6 2 4 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 9 1 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 7 2 9 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $4 r0 *1 0.74,1.1525 PMOS_VTL
M$4 10 4 7 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $5 r0 *1 0.93,1.1525 PMOS_VTL
M$5 10 3 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 8 7 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.17,0.195 NMOS_VTL
M$7 5 2 4 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $8 r0 *1 0.36,0.195 NMOS_VTL
M$8 12 1 5 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $9 r0 *1 0.55,0.195 NMOS_VTL
M$9 7 4 12 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $10 r0 *1 0.74,0.195 NMOS_VTL
M$10 11 2 7 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $11 r0 *1 0.93,0.195 NMOS_VTL
M$11 5 3 11 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
* device instance $12 r0 *1 1.12,0.2975 NMOS_VTL
M$12 8 7 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS MUX2_X1

* cell OAI22_X2
* pin B2
* pin B1
* pin A2
* pin A1
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT OAI22_X2 1 2 3 4 6 7 8
* net 1 B2
* net 2 B1
* net 3 A2
* net 4 A1
* net 6 NWELL,VDD
* net 7 PWELL,VSS
* net 8 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 10 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 8 2 10 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 9 2 8 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 6 1 9 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 12 3 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 8 4 12 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.31,0.995 PMOS_VTL
M$7 11 4 8 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.5,0.995 PMOS_VTL
M$8 6 3 11 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 0.17,0.2975 NMOS_VTL
M$9 7 1 5 7 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $10 r0 *1 0.36,0.2975 NMOS_VTL
M$10 5 2 7 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $13 r0 *1 0.93,0.2975 NMOS_VTL
M$13 8 3 5 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $14 r0 *1 1.12,0.2975 NMOS_VTL
M$14 5 4 8 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
.ENDS OAI22_X2

* cell XOR2_X2
* pin B
* pin A
* pin NWELL,VDD
* pin Z
* pin PWELL,VSS
.SUBCKT XOR2_X2 1 2 4 5 7
* net 1 B
* net 2 A
* net 4 NWELL,VDD
* net 5 Z
* net 7 PWELL,VSS
* device instance $1 r0 *1 0.2,0.995 PMOS_VTL
M$1 8 2 3 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.39,0.995 PMOS_VTL
M$2 4 1 8 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.58,0.995 PMOS_VTL
M$3 6 3 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.77,0.995 PMOS_VTL
M$4 5 2 6 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $5 r0 *1 0.96,0.995 PMOS_VTL
M$5 6 1 5 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $9 r0 *1 0.2,0.2975 NMOS_VTL
M$9 3 2 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $10 r0 *1 0.39,0.2975 NMOS_VTL
M$10 7 1 3 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.58,0.2975 NMOS_VTL
M$11 5 3 7 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $12 r0 *1 0.77,0.2975 NMOS_VTL
M$12 10 2 5 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.96,0.2975 NMOS_VTL
M$13 7 1 10 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 1.15,0.2975 NMOS_VTL
M$14 9 1 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 1.34,0.2975 NMOS_VTL
M$15 5 2 9 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
.ENDS XOR2_X2

* cell OR3_X2
* pin A1
* pin A2
* pin A3
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR3_X2 1 2 3 5 6 7
* net 1 A1
* net 2 A2
* net 3 A3
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 9 1 4 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 8 2 9 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 8 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 4 6 6 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $6 r0 *1 0.17,0.2975 NMOS_VTL
M$6 5 1 4 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $7 r0 *1 0.36,0.2975 NMOS_VTL
M$7 4 2 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.55,0.2975 NMOS_VTL
M$8 5 3 4 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.74,0.2975 NMOS_VTL
M$9 7 4 5 5 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS OR3_X2

* cell AOI211_X4
* pin C1
* pin C2
* pin B
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT AOI211_X4 1 2 3 4 8 9 10
* net 1 C1
* net 2 C2
* net 3 B
* net 4 A
* net 8 PWELL,VSS
* net 9 NWELL,VDD
* net 10 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 6 1 7 9 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 7 2 6 9 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 11 3 7 9 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 9 4 11 9 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 5 6 9 9 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $7 r0 *1 1.31,0.995 PMOS_VTL
M$7 10 5 9 9 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $11 r0 *1 0.17,0.2975 NMOS_VTL
M$11 12 1 6 8 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $12 r0 *1 0.36,0.2975 NMOS_VTL
M$12 8 2 12 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.55,0.2975 NMOS_VTL
M$13 6 3 8 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 0.74,0.2975 NMOS_VTL
M$14 8 4 6 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 0.93,0.2975 NMOS_VTL
M$15 5 6 8 8 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $17 r0 *1 1.31,0.2975 NMOS_VTL
M$17 10 5 8 8 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U
+ PD=2.705U
.ENDS AOI211_X4

* cell OR2_X1
* pin A1
* pin A2
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR2_X1 1 2 3 5 6
* net 1 A1
* net 2 A2
* net 3 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 7 1 4 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 7 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 4 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.195 NMOS_VTL
M$4 4 1 3 3 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $5 r0 *1 0.36,0.195 NMOS_VTL
M$5 3 2 4 3 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 4 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OR2_X1

* cell OR4_X4
* pin PWELL,VSS
* pin ZN
* pin A4
* pin A3
* pin A2
* pin A1
* pin NWELL,VDD
.SUBCKT OR4_X4 1 3 4 5 6 7 8
* net 1 PWELL,VSS
* net 3 ZN
* net 4 A4
* net 5 A3
* net 6 A2
* net 7 A1
* net 8 NWELL,VDD
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 10 4 8 8 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 9 5 10 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 11 6 9 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 2 7 11 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 13 7 2 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 14 6 13 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.31,0.995 PMOS_VTL
M$7 12 5 14 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.5,0.995 PMOS_VTL
M$8 8 4 12 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $9 r0 *1 1.69,0.995 PMOS_VTL
M$9 3 2 8 8 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $13 r0 *1 0.17,0.2975 NMOS_VTL
M$13 2 4 1 1 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $14 r0 *1 0.36,0.2975 NMOS_VTL
M$14 1 5 2 1 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $15 r0 *1 0.55,0.2975 NMOS_VTL
M$15 2 6 1 1 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $16 r0 *1 0.74,0.2975 NMOS_VTL
M$16 1 7 2 1 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $21 r0 *1 1.69,0.2975 NMOS_VTL
M$21 3 2 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS OR4_X4

* cell BUF_X2
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT BUF_X2 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 4 1 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.21,0.2975 NMOS_VTL
M$4 3 1 2 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.4,0.2975 NMOS_VTL
M$5 5 2 3 3 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS BUF_X2

* cell XNOR2_X2
* pin A
* pin B
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT XNOR2_X2 2 3 4 5 7
* net 2 A
* net 3 B
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 1.135,0.995 PMOS_VTL
M$1 7 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 1.325,0.995 PMOS_VTL
M$2 9 2 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 1.515,0.995 PMOS_VTL
M$3 5 3 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 1.705,0.995 PMOS_VTL
M$4 8 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.18,0.995 PMOS_VTL
M$5 7 1 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $7 r0 *1 0.56,0.995 PMOS_VTL
M$7 1 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 0.75,0.995 PMOS_VTL
M$8 5 2 1 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 1.135,0.2975 NMOS_VTL
M$9 6 2 7 4 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $11 r0 *1 1.515,0.2975 NMOS_VTL
M$11 6 3 7 4 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $13 r0 *1 0.18,0.2975 NMOS_VTL
M$13 6 1 4 4 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $15 r0 *1 0.56,0.2975 NMOS_VTL
M$15 10 3 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 0.75,0.2975 NMOS_VTL
M$16 1 2 10 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS XNOR2_X2

* cell AOI22_X2
* pin B2
* pin B1
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT AOI22_X2 1 2 3 4 5 7 8
* net 1 B2
* net 2 B1
* net 3 A2
* net 4 A1
* net 5 PWELL,VSS
* net 7 NWELL,VDD
* net 8 ZN
* device instance $1 r0 *1 0.175,0.995 PMOS_VTL
M$1 7 1 6 7 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $2 r0 *1 0.365,0.995 PMOS_VTL
M$2 6 2 7 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $5 r0 *1 0.935,0.995 PMOS_VTL
M$5 8 3 6 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $6 r0 *1 1.125,0.995 PMOS_VTL
M$6 6 4 8 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $9 r0 *1 0.175,0.2975 NMOS_VTL
M$9 12 1 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $10 r0 *1 0.365,0.2975 NMOS_VTL
M$10 8 2 12 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.555,0.2975 NMOS_VTL
M$11 10 2 8 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 0.745,0.2975 NMOS_VTL
M$12 5 1 10 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.935,0.2975 NMOS_VTL
M$13 11 3 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 1.125,0.2975 NMOS_VTL
M$14 8 4 11 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 1.315,0.2975 NMOS_VTL
M$15 9 4 8 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 1.505,0.2975 NMOS_VTL
M$16 5 3 9 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI22_X2

* cell NOR4_X1
* pin A4
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NOR4_X1 1 2 3 4 5 6 7
* net 1 A4
* net 2 A3
* net 3 A2
* net 4 A1
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 10 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 9 2 10 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 8 3 9 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 4 8 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 7 1 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.36,0.2975 NMOS_VTL
M$6 5 2 7 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.55,0.2975 NMOS_VTL
M$7 7 3 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.74,0.2975 NMOS_VTL
M$8 5 4 7 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NOR4_X1

* cell OAI211_X2
* pin A
* pin B
* pin C2
* pin C1
* pin ZN
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT OAI211_X2 1 2 3 4 6 7 8
* net 1 A
* net 2 B
* net 3 C2
* net 4 C1
* net 6 ZN
* net 7 PWELL,VSS
* net 8 NWELL,VDD
* device instance $1 r0 *1 0.205,0.995 PMOS_VTL
M$1 6 1 8 8 PMOS_VTL L=0.05U W=1.26U AS=0.111825P AD=0.0882P PS=2.245U PD=1.54U
* device instance $2 r0 *1 0.395,0.995 PMOS_VTL
M$2 8 2 6 8 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.089775P PS=1.54U PD=1.545U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 10 3 8 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 6 4 10 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.35,0.995 PMOS_VTL
M$7 9 4 6 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.54,0.995 PMOS_VTL
M$8 8 3 9 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 0.205,0.2975 NMOS_VTL
M$9 12 1 5 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $10 r0 *1 0.395,0.2975 NMOS_VTL
M$10 7 2 12 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.585,0.2975 NMOS_VTL
M$11 11 2 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.0300875P PS=0.555U
+ PD=0.56U
* device instance $12 r0 *1 0.78,0.2975 NMOS_VTL
M$12 5 1 11 7 NMOS_VTL L=0.05U W=0.415U AS=0.0300875P AD=0.02905P PS=0.56U
+ PD=0.555U
* device instance $13 r0 *1 0.97,0.2975 NMOS_VTL
M$13 6 3 5 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $14 r0 *1 1.16,0.2975 NMOS_VTL
M$14 5 4 6 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
.ENDS OAI211_X2

* cell AOI22_X1
* pin B2
* pin B1
* pin A1
* pin A2
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT AOI22_X1 1 2 3 4 5 7 8
* net 1 B2
* net 2 B1
* net 3 A1
* net 4 A2
* net 5 PWELL,VSS
* net 7 NWELL,VDD
* net 8 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 7 1 6 7 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 6 2 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.565,0.995 PMOS_VTL
M$3 8 3 6 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.755,0.995 PMOS_VTL
M$4 6 4 8 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.185,0.2975 NMOS_VTL
M$5 10 1 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.375,0.2975 NMOS_VTL
M$6 8 2 10 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.565,0.2975 NMOS_VTL
M$7 9 3 8 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.755,0.2975 NMOS_VTL
M$8 5 4 9 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI22_X1

* cell OR2_X4
* pin A2
* pin A1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT OR2_X4 1 2 3 5 6
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 5 ZN
* net 6 NWELL,VDD
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 8 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 4 2 8 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 7 2 4 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 6 1 7 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 5 4 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $9 r0 *1 0.17,0.2975 NMOS_VTL
M$9 4 1 3 3 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $10 r0 *1 0.36,0.2975 NMOS_VTL
M$10 3 2 4 3 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $13 r0 *1 0.93,0.2975 NMOS_VTL
M$13 5 4 3 3 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS OR2_X4

* cell OAI222_X2
* pin PWELL,VSS
* pin C1
* pin C2
* pin B1
* pin B2
* pin A1
* pin A2
* pin ZN
* pin NWELL,VDD
.SUBCKT OAI222_X2 1 4 5 6 7 8 9 10 11
* net 1 PWELL,VSS
* net 4 C1
* net 5 C2
* net 6 B1
* net 7 B2
* net 8 A1
* net 9 A2
* net 10 ZN
* net 11 NWELL,VDD
* device instance $1 r0 *1 0.215,0.995 PMOS_VTL
M$1 12 4 10 11 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.405,0.995 PMOS_VTL
M$2 11 5 12 11 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.595,0.995 PMOS_VTL
M$3 13 5 11 11 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.785,0.995 PMOS_VTL
M$4 10 4 13 11 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.975,0.995 PMOS_VTL
M$5 14 6 10 11 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.165,0.995 PMOS_VTL
M$6 11 7 14 11 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.355,0.995 PMOS_VTL
M$7 15 7 11 11 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.545,0.995 PMOS_VTL
M$8 10 6 15 11 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0945P PS=0.77U PD=0.93U
* device instance $9 r0 *1 1.895,0.995 PMOS_VTL
M$9 16 8 10 11 PMOS_VTL L=0.05U W=0.63U AS=0.0945P AD=0.0441P PS=0.93U PD=0.77U
* device instance $10 r0 *1 2.085,0.995 PMOS_VTL
M$10 11 9 16 11 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $11 r0 *1 2.275,0.995 PMOS_VTL
M$11 17 9 11 11 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $12 r0 *1 2.465,0.995 PMOS_VTL
M$12 10 8 17 11 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0693P PS=0.77U PD=1.48U
* device instance $13 r0 *1 1.895,0.2975 NMOS_VTL
M$13 10 8 3 1 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.072625P PS=1.595U
+ PD=1.595U
* device instance $14 r0 *1 2.085,0.2975 NMOS_VTL
M$14 3 9 10 1 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $17 r0 *1 0.215,0.2975 NMOS_VTL
M$17 1 4 2 1 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $18 r0 *1 0.405,0.2975 NMOS_VTL
M$18 2 5 1 1 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $21 r0 *1 0.975,0.2975 NMOS_VTL
M$21 3 6 2 1 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $22 r0 *1 1.165,0.2975 NMOS_VTL
M$22 2 7 3 1 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
.ENDS OAI222_X2

* cell OR3_X4
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR3_X4 1 2 3 5 6 7
* net 1 A3
* net 2 A2
* net 3 A1
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.205,0.995 PMOS_VTL
M$1 11 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.395,0.995 PMOS_VTL
M$2 10 2 11 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.585,0.995 PMOS_VTL
M$3 4 3 10 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.775,0.995 PMOS_VTL
M$4 9 3 4 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.965,0.995 PMOS_VTL
M$5 8 2 9 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.155,0.995 PMOS_VTL
M$6 6 1 8 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.345,0.995 PMOS_VTL
M$7 7 4 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.177975P AD=0.200025P PS=3.085U
+ PD=3.785U
* device instance $11 r0 *1 0.205,0.2975 NMOS_VTL
M$11 4 1 5 5 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $12 r0 *1 0.395,0.2975 NMOS_VTL
M$12 5 2 4 5 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $13 r0 *1 0.585,0.2975 NMOS_VTL
M$13 4 3 5 5 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $17 r0 *1 1.345,0.2975 NMOS_VTL
M$17 7 4 5 5 NMOS_VTL L=0.05U W=1.66U AS=0.1172375P AD=0.1317625P PS=2.225U
+ PD=2.71U
.ENDS OR3_X4

* cell OR2_X2
* pin A1
* pin A2
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR2_X2 1 2 3 5 6
* net 1 A1
* net 2 A2
* net 3 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 1 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 4 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 4 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.36,0.2975 NMOS_VTL
M$6 3 2 4 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.55,0.2975 NMOS_VTL
M$7 6 4 3 3 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS OR2_X2

* cell NOR3_X1
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NOR3_X1 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 8 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 7 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.2975 NMOS_VTL
M$4 6 1 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.36,0.2975 NMOS_VTL
M$5 4 2 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 3 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NOR3_X1

* cell AOI211_X2
* pin B
* pin A
* pin C2
* pin C1
* pin ZN
* pin NWELL,VDD
* pin PWELL,VSS
.SUBCKT AOI211_X2 1 2 3 4 6 7 8
* net 1 B
* net 2 A
* net 3 C2
* net 4 C1
* net 6 ZN
* net 7 NWELL,VDD
* net 8 PWELL,VSS
* device instance $1 r0 *1 0.175,0.995 PMOS_VTL
M$1 10 1 5 7 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.365,0.995 PMOS_VTL
M$2 7 2 10 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.555,0.995 PMOS_VTL
M$3 9 2 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.745,0.995 PMOS_VTL
M$4 5 1 9 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.055125P PS=0.77U PD=0.805U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 6 3 5 7 PMOS_VTL L=0.05U W=1.26U AS=0.099225P AD=0.11025P PS=1.575U PD=2.24U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 5 4 6 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $9 r0 *1 0.175,0.2975 NMOS_VTL
M$9 6 1 8 8 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0653625P PS=1.595U
+ PD=1.145U
* device instance $10 r0 *1 0.365,0.2975 NMOS_VTL
M$10 8 2 6 8 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $13 r0 *1 0.97,0.2975 NMOS_VTL
M$13 11 3 8 8 NMOS_VTL L=0.05U W=0.415U AS=0.0363125P AD=0.02905P PS=0.59U
+ PD=0.555U
* device instance $14 r0 *1 1.16,0.2975 NMOS_VTL
M$14 6 4 11 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 1.35,0.2975 NMOS_VTL
M$15 12 4 6 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 1.54,0.2975 NMOS_VTL
M$16 8 3 12 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI211_X2

* cell CLKBUF_X1
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT CLKBUF_X1 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.19,1.1525 PMOS_VTL
M$1 2 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.033075P PS=0.77U
+ PD=0.84U
* device instance $2 r0 *1 0.38,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.19,0.2075 NMOS_VTL
M$3 3 1 2 3 NMOS_VTL L=0.05U W=0.095U AS=0.009975P AD=0.01015P PS=0.4U PD=0.335U
* device instance $4 r0 *1 0.38,0.2575 NMOS_VTL
M$4 5 2 3 3 NMOS_VTL L=0.05U W=0.195U AS=0.01015P AD=0.020475P PS=0.335U PD=0.6U
.ENDS CLKBUF_X1

* cell NAND3_X2
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND3_X2 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 6 1 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.11025P PS=2.24U PD=2.24U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 5 2 6 5 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 6 3 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $7 r0 *1 0.21,0.2975 NMOS_VTL
M$7 10 1 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $8 r0 *1 0.4,0.2975 NMOS_VTL
M$8 9 2 10 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.59,0.2975 NMOS_VTL
M$9 6 3 9 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.78,0.2975 NMOS_VTL
M$10 8 3 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.97,0.2975 NMOS_VTL
M$11 7 2 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 1.16,0.2975 NMOS_VTL
M$12 4 1 7 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND3_X2

* cell AOI21_X2
* pin A
* pin B2
* pin B1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT AOI21_X2 1 2 3 4 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 4 PWELL,VSS
* net 6 ZN
* net 7 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 7 1 5 7 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 6 2 5 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 5 3 6 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $7 r0 *1 0.21,0.2975 NMOS_VTL
M$7 6 1 4 4 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $9 r0 *1 0.59,0.2975 NMOS_VTL
M$9 9 2 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.78,0.2975 NMOS_VTL
M$10 6 3 9 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.97,0.2975 NMOS_VTL
M$11 8 3 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 1.16,0.2975 NMOS_VTL
M$12 4 2 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI21_X2

* cell CLKBUF_X3
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT CLKBUF_X3 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=1.89U AS=0.1323P AD=0.15435P PS=2.31U PD=3.01U
* device instance $5 r0 *1 0.17,0.1875 NMOS_VTL
M$5 3 1 2 3 NMOS_VTL L=0.05U W=0.195U AS=0.020475P AD=0.01365P PS=0.6U PD=0.335U
* device instance $6 r0 *1 0.36,0.1875 NMOS_VTL
M$6 5 2 3 3 NMOS_VTL L=0.05U W=0.585U AS=0.04095P AD=0.047775P PS=1.005U
+ PD=1.27U
.ENDS CLKBUF_X3

* cell INV_X2
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT INV_X2 1 2 3 4
* net 1 A
* net 2 PWELL,VSS
* net 3 NWELL,VDD
* net 4 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 4 1 3 3 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.11025P PS=2.24U PD=2.24U
* device instance $3 r0 *1 0.185,0.2975 NMOS_VTL
M$3 4 1 2 2 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.072625P PS=1.595U
+ PD=1.595U
.ENDS INV_X2

* cell NAND2_X1
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND2_X1 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 5 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 4 2 5 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.185,0.2975 NMOS_VTL
M$3 6 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $4 r0 *1 0.375,0.2975 NMOS_VTL
M$4 5 2 6 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND2_X1

* cell AND2_X1
* pin A1
* pin A2
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND2_X1 1 2 4 5 6
* net 1 A1
* net 2 A2
* net 4 NWELL,VDD
* net 5 PWELL,VSS
* net 6 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 3 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 3 2 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.195 NMOS_VTL
M$4 7 1 3 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $5 r0 *1 0.36,0.195 NMOS_VTL
M$5 5 2 7 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 3 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AND2_X1

* cell HA_X1
* pin A
* pin B
* pin S
* pin NWELL,VDD
* pin PWELL,VSS
* pin CO
.SUBCKT HA_X1 1 2 4 5 6 9
* net 1 A
* net 2 B
* net 4 S
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 9 CO
* device instance $1 r0 *1 0.785,1.0275 PMOS_VTL
M$1 10 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.0338625P AD=0.02205P PS=0.775U
+ PD=0.455U
* device instance $2 r0 *1 0.975,1.0275 PMOS_VTL
M$2 7 1 10 5 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.033075P PS=0.455U
+ PD=0.84U
* device instance $3 r0 *1 0.21,0.995 PMOS_VTL
M$3 4 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $4 r0 *1 0.4,0.995 PMOS_VTL
M$4 3 1 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.59,0.995 PMOS_VTL
M$5 5 7 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0338625P PS=0.77U PD=0.775U
* device instance $6 r0 *1 1.345,1.0275 PMOS_VTL
M$6 8 1 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $7 r0 *1 1.535,1.0275 PMOS_VTL
M$7 8 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $8 r0 *1 1.725,0.995 PMOS_VTL
M$8 9 8 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 0.785,0.195 NMOS_VTL
M$9 7 2 6 6 NMOS_VTL L=0.05U W=0.21U AS=0.0224P AD=0.0147P PS=0.56U PD=0.35U
* device instance $10 r0 *1 0.975,0.195 NMOS_VTL
M$10 6 1 7 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.02205P PS=0.35U PD=0.63U
* device instance $11 r0 *1 0.21,0.2975 NMOS_VTL
M$11 11 2 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $12 r0 *1 0.4,0.2975 NMOS_VTL
M$12 4 1 11 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.59,0.2975 NMOS_VTL
M$13 6 7 4 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.0224P PS=0.555U PD=0.56U
* device instance $14 r0 *1 1.345,0.195 NMOS_VTL
M$14 12 1 8 6 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $15 r0 *1 1.535,0.195 NMOS_VTL
M$15 6 2 12 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
* device instance $16 r0 *1 1.725,0.2975 NMOS_VTL
M$16 9 8 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS HA_X1

* cell AND4_X1
* pin A1
* pin A2
* pin A3
* pin A4
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND4_X1 1 2 3 4 6 7 8
* net 1 A1
* net 2 A2
* net 3 A3
* net 4 A4
* net 6 NWELL,VDD
* net 7 PWELL,VSS
* net 8 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 5 1 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 6 2 5 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 5 3 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $4 r0 *1 0.74,1.1525 PMOS_VTL
M$4 5 4 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 8 5 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.17,0.195 NMOS_VTL
M$6 10 1 5 7 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $7 r0 *1 0.36,0.195 NMOS_VTL
M$7 11 2 10 7 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $8 r0 *1 0.55,0.195 NMOS_VTL
M$8 9 3 11 7 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $9 r0 *1 0.74,0.195 NMOS_VTL
M$9 7 4 9 7 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $10 r0 *1 0.93,0.2975 NMOS_VTL
M$10 8 5 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AND4_X1

* cell AND2_X2
* pin A1
* pin A2
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND2_X2 1 2 4 5 6
* net 1 A1
* net 2 A2
* net 4 NWELL,VDD
* net 5 PWELL,VSS
* net 6 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 3 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 4 2 3 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 7 1 3 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.36,0.2975 NMOS_VTL
M$6 5 2 7 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.55,0.2975 NMOS_VTL
M$7 6 3 5 5 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS AND2_X2

* cell NAND3_X1
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND3_X1 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 6 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.2975 NMOS_VTL
M$4 8 1 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.36,0.2975 NMOS_VTL
M$5 7 2 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 3 7 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND3_X1

* cell NOR2_X1
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NOR2_X1 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 6 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 5 2 6 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.185,0.2975 NMOS_VTL
M$3 5 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $4 r0 *1 0.375,0.2975 NMOS_VTL
M$4 3 2 5 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NOR2_X1

* cell INV_X1
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT INV_X1 1 2 3 4
* net 1 A
* net 2 PWELL,VSS
* net 3 NWELL,VDD
* net 4 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 3 3 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.06615P PS=1.47U PD=1.47U
* device instance $2 r0 *1 0.17,0.2975 NMOS_VTL
M$2 4 1 2 2 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.043575P PS=1.04U
+ PD=1.04U
.ENDS INV_X1

* cell BUF_X4
* pin A
* pin NWELL,VDD
* pin Z
* pin PWELL,VSS
.SUBCKT BUF_X4 1 3 4 5
* net 1 A
* net 3 NWELL,VDD
* net 4 Z
* net 5 PWELL,VSS
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 2 1 3 3 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 4 2 3 3 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $7 r0 *1 0.17,0.2975 NMOS_VTL
M$7 2 1 5 5 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $9 r0 *1 0.55,0.2975 NMOS_VTL
M$9 4 2 5 5 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS BUF_X4

* cell BUF_X1
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT BUF_X1 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 2 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.033075P PS=0.77U
+ PD=0.84U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.17,0.195 NMOS_VTL
M$3 3 1 2 3 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.021875P PS=0.63U PD=0.555U
* device instance $4 r0 *1 0.36,0.2975 NMOS_VTL
M$4 5 2 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS BUF_X1

* cell DFFR_X2
* pin PWELL,VSS
* pin CK
* pin D
* pin RN
* pin QN
* pin Q
* pin NWELL,VDD
.SUBCKT DFFR_X2 1 3 5 9 11 12 19
* net 1 PWELL,VSS
* net 3 CK
* net 5 D
* net 9 RN
* net 11 QN
* net 12 Q
* net 19 NWELL,VDD
* device instance $1 r0 *1 2.51,1.025 PMOS_VTL
M$1 23 4 8 19 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.0063P PS=0.455U
+ PD=0.23U
* device instance $2 r0 *1 2.7,1.025 PMOS_VTL
M$2 23 10 19 19 PMOS_VTL L=0.05U W=0.09U AS=0.0252P AD=0.0063P PS=0.77U PD=0.23U
* device instance $3 r0 *1 1.875,1.0125 PMOS_VTL
M$3 19 6 7 19 PMOS_VTL L=0.05U W=0.315U AS=0.04725P AD=0.0322875P PS=0.93U
+ PD=0.52U
* device instance $4 r0 *1 2.13,1.0125 PMOS_VTL
M$4 22 6 19 19 PMOS_VTL L=0.05U W=0.315U AS=0.0322875P AD=0.02205P PS=0.52U
+ PD=0.455U
* device instance $5 r0 *1 2.32,1.0125 PMOS_VTL
M$5 8 2 22 19 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.014175P PS=0.455U
+ PD=0.455U
* device instance $6 r0 *1 2.89,0.995 PMOS_VTL
M$6 10 9 19 19 PMOS_VTL L=0.05U W=0.63U AS=0.0252P AD=0.048825P PS=0.77U
+ PD=0.785U
* device instance $7 r0 *1 3.095,0.995 PMOS_VTL
M$7 19 8 10 19 PMOS_VTL L=0.05U W=0.63U AS=0.048825P AD=0.06615P PS=0.785U
+ PD=0.84U
* device instance $8 r0 *1 3.355,0.995 PMOS_VTL
M$8 11 8 19 19 PMOS_VTL L=0.05U W=1.26U AS=0.1323P AD=0.11025P PS=1.68U PD=1.61U
* device instance $10 r0 *1 3.805,0.995 PMOS_VTL
M$10 12 10 19 19 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U
+ PD=2.24U
* device instance $12 r0 *1 1.1,1.065 PMOS_VTL
M$12 20 2 6 19 PMOS_VTL L=0.05U W=0.09U AS=0.01785P AD=0.0063P PS=0.56U PD=0.23U
* device instance $13 r0 *1 1.29,1.065 PMOS_VTL
M$13 19 7 20 19 PMOS_VTL L=0.05U W=0.09U AS=0.0063P AD=0.0063P PS=0.23U PD=0.23U
* device instance $14 r0 *1 1.48,1.065 PMOS_VTL
M$14 20 9 19 19 PMOS_VTL L=0.05U W=0.09U AS=0.0063P AD=0.01035P PS=0.23U
+ PD=0.41U
* device instance $15 r0 *1 0.72,1.05 PMOS_VTL
M$15 21 5 19 19 PMOS_VTL L=0.05U W=0.42U AS=0.0441P AD=0.0294P PS=1.05U PD=0.56U
* device instance $16 r0 *1 0.91,1.05 PMOS_VTL
M$16 6 4 21 19 PMOS_VTL L=0.05U W=0.42U AS=0.0294P AD=0.01785P PS=0.56U PD=0.56U
* device instance $17 r0 *1 0.19,1.0325 PMOS_VTL
M$17 19 3 2 19 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $18 r0 *1 0.38,1.0325 PMOS_VTL
M$18 4 2 19 19 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.033075P PS=0.455U
+ PD=0.84U
* device instance $19 r0 *1 3.425,0.2975 NMOS_VTL
M$19 11 8 1 1 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U
+ PD=1.11U
* device instance $21 r0 *1 3.805,0.2975 NMOS_VTL
M$21 12 10 1 1 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U
+ PD=1.595U
* device instance $23 r0 *1 2.445,0.26 NMOS_VTL
M$23 18 2 8 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.0063P PS=0.35U PD=0.23U
* device instance $24 r0 *1 2.635,0.26 NMOS_VTL
M$24 18 10 1 1 NMOS_VTL L=0.05U W=0.09U AS=0.017675P AD=0.0063P PS=0.555U
+ PD=0.23U
* device instance $25 r0 *1 1.875,0.32 NMOS_VTL
M$25 1 6 7 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $26 r0 *1 2.065,0.32 NMOS_VTL
M$26 16 6 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $27 r0 *1 2.255,0.32 NMOS_VTL
M$27 8 4 16 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0105P PS=0.35U PD=0.35U
* device instance $28 r0 *1 2.825,0.2975 NMOS_VTL
M$28 17 9 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.017675P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $29 r0 *1 3.015,0.2975 NMOS_VTL
M$29 10 8 17 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
* device instance $30 r0 *1 0.19,0.245 NMOS_VTL
M$30 1 3 2 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $31 r0 *1 0.38,0.245 NMOS_VTL
M$31 4 2 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.02205P PS=0.35U PD=0.63U
* device instance $32 r0 *1 1.1,0.35 NMOS_VTL
M$32 15 4 6 1 NMOS_VTL L=0.05U W=0.09U AS=0.012775P AD=0.0063P PS=0.415U
+ PD=0.23U
* device instance $33 r0 *1 1.29,0.35 NMOS_VTL
M$33 14 7 15 1 NMOS_VTL L=0.05U W=0.09U AS=0.0063P AD=0.0063P PS=0.23U PD=0.23U
* device instance $34 r0 *1 1.48,0.35 NMOS_VTL
M$34 1 9 14 1 NMOS_VTL L=0.05U W=0.09U AS=0.0063P AD=0.00945P PS=0.23U PD=0.39U
* device instance $35 r0 *1 0.72,0.3525 NMOS_VTL
M$35 13 5 1 1 NMOS_VTL L=0.05U W=0.275U AS=0.028875P AD=0.01925P PS=0.76U
+ PD=0.415U
* device instance $36 r0 *1 0.91,0.3525 NMOS_VTL
M$36 6 2 13 1 NMOS_VTL L=0.05U W=0.275U AS=0.01925P AD=0.012775P PS=0.415U
+ PD=0.415U
.ENDS DFFR_X2

* cell XOR2_X1
* pin A
* pin B
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT XOR2_X1 1 3 4 5 6
* net 1 A
* net 3 B
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 Z
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 8 1 2 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 8 3 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.0338625P AD=0.02205P PS=0.775U
+ PD=0.455U
* device instance $3 r0 *1 0.555,0.995 PMOS_VTL
M$3 7 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0338625P AD=0.0441P PS=0.775U PD=0.77U
* device instance $4 r0 *1 0.745,0.995 PMOS_VTL
M$4 6 1 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.935,0.995 PMOS_VTL
M$5 7 3 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.17,0.195 NMOS_VTL
M$6 2 1 4 4 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $7 r0 *1 0.36,0.195 NMOS_VTL
M$7 4 3 2 4 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0224P PS=0.35U PD=0.56U
* device instance $8 r0 *1 0.555,0.2975 NMOS_VTL
M$8 6 2 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.0224P AD=0.02905P PS=0.56U PD=0.555U
* device instance $9 r0 *1 0.745,0.2975 NMOS_VTL
M$9 9 1 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.935,0.2975 NMOS_VTL
M$10 4 3 9 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS XOR2_X1

* cell OR4_X2
* pin A1
* pin A2
* pin A3
* pin A4
* pin NWELL,VDD
* pin ZN
* pin PWELL,VSS
.SUBCKT OR4_X2 1 2 3 4 6 7 8
* net 1 A1
* net 2 A2
* net 3 A3
* net 4 A4
* net 6 NWELL,VDD
* net 7 ZN
* net 8 PWELL,VSS
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 11 1 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 10 2 11 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 9 3 10 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 6 4 9 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 7 5 6 6 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $7 r0 *1 0.17,0.2975 NMOS_VTL
M$7 5 1 8 8 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $8 r0 *1 0.36,0.2975 NMOS_VTL
M$8 8 2 5 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.55,0.2975 NMOS_VTL
M$9 5 3 8 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.74,0.2975 NMOS_VTL
M$10 8 4 5 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.93,0.2975 NMOS_VTL
M$11 7 5 8 8 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS OR4_X2

* cell OAI221_X2
* pin C2
* pin C1
* pin B1
* pin B2
* pin A
* pin ZN
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT OAI221_X2 1 2 3 4 5 7 9 10
* net 1 C2
* net 2 C1
* net 3 B1
* net 4 B2
* net 5 A
* net 7 ZN
* net 9 PWELL,VSS
* net 10 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 12 1 10 10 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 7 2 12 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 11 2 7 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 10 1 11 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 7 5 10 10 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 14 3 7 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.35,0.995 PMOS_VTL
M$7 10 4 14 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.54,0.995 PMOS_VTL
M$8 13 4 10 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $9 r0 *1 1.73,0.995 PMOS_VTL
M$9 7 3 13 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $11 r0 *1 0.21,0.2975 NMOS_VTL
M$11 7 1 6 9 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $12 r0 *1 0.4,0.2975 NMOS_VTL
M$12 6 2 7 9 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $15 r0 *1 0.97,0.2975 NMOS_VTL
M$15 8 5 6 9 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $16 r0 *1 1.16,0.2975 NMOS_VTL
M$16 9 3 8 9 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $17 r0 *1 1.35,0.2975 NMOS_VTL
M$17 8 4 9 9 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
.ENDS OAI221_X2

* cell XNOR2_X1
* pin A
* pin B
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT XNOR2_X1 1 2 4 5 7
* net 1 A
* net 2 B
* net 4 NWELL,VDD
* net 5 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.18,1.1525 PMOS_VTL
M$1 3 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.37,1.1525 PMOS_VTL
M$2 3 2 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.0338625P AD=0.02205P PS=0.775U
+ PD=0.455U
* device instance $3 r0 *1 0.565,0.995 PMOS_VTL
M$3 7 3 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.0338625P AD=0.0441P PS=0.775U PD=0.77U
* device instance $4 r0 *1 0.755,0.995 PMOS_VTL
M$4 8 1 7 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.945,0.995 PMOS_VTL
M$5 4 2 8 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.18,0.195 NMOS_VTL
M$6 9 1 3 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $7 r0 *1 0.37,0.195 NMOS_VTL
M$7 5 2 9 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0224P PS=0.35U PD=0.56U
* device instance $8 r0 *1 0.565,0.2975 NMOS_VTL
M$8 6 3 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.0224P AD=0.02905P PS=0.56U PD=0.555U
* device instance $9 r0 *1 0.755,0.2975 NMOS_VTL
M$9 7 1 6 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.945,0.2975 NMOS_VTL
M$10 6 2 7 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS XNOR2_X1

* cell NOR2_X4
* pin A2
* pin A1
* pin ZN
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT NOR2_X4 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 ZN
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 9 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 3 2 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 8 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 5 1 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 7 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 3 2 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.35,0.995 PMOS_VTL
M$7 6 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.54,0.995 PMOS_VTL
M$8 5 1 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 0.21,0.2975 NMOS_VTL
M$9 3 1 4 4 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.130725P PS=2.705U
+ PD=2.705U
* device instance $10 r0 *1 0.4,0.2975 NMOS_VTL
M$10 4 2 3 4 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.1162P PS=2.22U PD=2.22U
.ENDS NOR2_X4

* cell AOI22_X4
* pin PWELL,VSS
* pin B2
* pin B1
* pin ZN
* pin A2
* pin A1
* pin NWELL,VDD
.SUBCKT AOI22_X4 1 2 3 4 5 6 16
* net 1 PWELL,VSS
* net 2 B2
* net 3 B1
* net 4 ZN
* net 5 A2
* net 6 A1
* net 16 NWELL,VDD
* device instance $1 r0 *1 0.175,0.995 PMOS_VTL
M$1 16 2 15 16 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $2 r0 *1 0.365,0.995 PMOS_VTL
M$2 15 3 16 16 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.1764P PS=3.08U PD=3.08U
* device instance $9 r0 *1 1.695,0.995 PMOS_VTL
M$9 4 5 15 16 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $10 r0 *1 1.885,0.995 PMOS_VTL
M$10 15 6 4 16 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.1764P PS=3.08U PD=3.08U
* device instance $17 r0 *1 0.175,0.2975 NMOS_VTL
M$17 7 2 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $18 r0 *1 0.365,0.2975 NMOS_VTL
M$18 4 3 7 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 0.555,0.2975 NMOS_VTL
M$19 10 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $20 r0 *1 0.745,0.2975 NMOS_VTL
M$20 1 2 10 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $21 r0 *1 0.935,0.2975 NMOS_VTL
M$21 8 2 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $22 r0 *1 1.125,0.2975 NMOS_VTL
M$22 4 3 8 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $23 r0 *1 1.315,0.2975 NMOS_VTL
M$23 12 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $24 r0 *1 1.505,0.2975 NMOS_VTL
M$24 1 2 12 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $25 r0 *1 1.695,0.2975 NMOS_VTL
M$25 13 5 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $26 r0 *1 1.885,0.2975 NMOS_VTL
M$26 4 6 13 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $27 r0 *1 2.075,0.2975 NMOS_VTL
M$27 11 6 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $28 r0 *1 2.265,0.2975 NMOS_VTL
M$28 1 5 11 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $29 r0 *1 2.455,0.2975 NMOS_VTL
M$29 14 5 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $30 r0 *1 2.645,0.2975 NMOS_VTL
M$30 4 6 14 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $31 r0 *1 2.835,0.2975 NMOS_VTL
M$31 9 6 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $32 r0 *1 3.025,0.2975 NMOS_VTL
M$32 1 5 9 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI22_X4

* cell NOR4_X4
* pin PWELL,VSS
* pin A1
* pin A2
* pin A3
* pin A4
* pin ZN
* pin NWELL,VDD
.SUBCKT NOR4_X4 1 2 3 4 5 6 10
* net 1 PWELL,VSS
* net 2 A1
* net 3 A2
* net 4 A3
* net 5 A4
* net 6 ZN
* net 10 NWELL,VDD
* device instance $1 r0 *1 1.92,0.995 PMOS_VTL
M$1 8 4 9 10 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 2.68,0.995 PMOS_VTL
M$5 10 5 9 10 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $9 r0 *1 0.17,0.995 PMOS_VTL
M$9 6 2 7 10 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $13 r0 *1 0.93,0.995 PMOS_VTL
M$13 8 3 7 10 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $17 r0 *1 0.17,0.2975 NMOS_VTL
M$17 6 2 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $21 r0 *1 0.93,0.2975 NMOS_VTL
M$21 6 3 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
* device instance $25 r0 *1 1.92,0.2975 NMOS_VTL
M$25 1 4 6 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $29 r0 *1 2.68,0.2975 NMOS_VTL
M$29 1 5 6 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS NOR4_X4

* cell NOR2_X2
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NOR2_X2 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 7 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 5 2 7 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 6 2 5 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 4 1 6 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.21,0.2975 NMOS_VTL
M$5 5 1 3 3 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.072625P PS=1.595U
+ PD=1.595U
* device instance $6 r0 *1 0.4,0.2975 NMOS_VTL
M$6 3 2 5 3 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
.ENDS NOR2_X2

* cell NOR3_X4
* pin PWELL,VSS
* pin A1
* pin A2
* pin A3
* pin ZN
* pin NWELL,VDD
.SUBCKT NOR3_X4 1 2 3 4 5 8
* net 1 PWELL,VSS
* net 2 A1
* net 3 A2
* net 4 A3
* net 5 ZN
* net 8 NWELL,VDD
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 5 2 7 8 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 6 3 7 8 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $9 r0 *1 1.875,0.995 PMOS_VTL
M$9 6 4 8 8 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.19845P PS=3.78U PD=3.78U
* device instance $13 r0 *1 1.875,0.2975 NMOS_VTL
M$13 5 4 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.130725P PS=2.705U
+ PD=2.705U
* device instance $17 r0 *1 0.17,0.2975 NMOS_VTL
M$17 5 2 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $21 r0 *1 0.93,0.2975 NMOS_VTL
M$21 5 3 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS NOR3_X4

* cell MUX2_X2
* pin A
* pin B
* pin S
* pin NWELL,VDD
* pin PWELL,VSS
* pin Z
.SUBCKT MUX2_X2 1 2 3 6 7 8
* net 1 A
* net 2 B
* net 3 S
* net 6 NWELL,VDD
* net 7 PWELL,VSS
* net 8 Z
* device instance $1 r0 *1 1.16,0.995 PMOS_VTL
M$1 8 4 6 6 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.077175P PS=2.24U PD=1.54U
* device instance $3 r0 *1 1.54,1.1525 PMOS_VTL
M$3 9 3 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.033075P PS=0.77U
+ PD=0.84U
* device instance $4 r0 *1 0.215,0.995 PMOS_VTL
M$4 6 1 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $5 r0 *1 0.405,0.995 PMOS_VTL
M$5 5 9 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 0.595,0.995 PMOS_VTL
M$6 4 2 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.045675P PS=0.77U PD=0.775U
* device instance $7 r0 *1 0.79,0.995 PMOS_VTL
M$7 5 3 4 6 PMOS_VTL L=0.05U W=0.63U AS=0.045675P AD=0.0693P PS=0.775U PD=1.48U
* device instance $8 r0 *1 1.54,0.195 NMOS_VTL
M$8 9 3 7 7 NMOS_VTL L=0.05U W=0.21U AS=0.021875P AD=0.02205P PS=0.555U PD=0.63U
* device instance $9 r0 *1 1.16,0.2975 NMOS_VTL
M$9 8 4 7 7 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.050925P PS=1.595U
+ PD=1.11U
* device instance $11 r0 *1 0.215,0.2975 NMOS_VTL
M$11 11 1 4 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $12 r0 *1 0.405,0.2975 NMOS_VTL
M$12 7 9 11 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.595,0.2975 NMOS_VTL
M$13 10 2 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.0300875P PS=0.555U
+ PD=0.56U
* device instance $14 r0 *1 0.79,0.2975 NMOS_VTL
M$14 4 3 10 7 NMOS_VTL L=0.05U W=0.415U AS=0.0300875P AD=0.043575P PS=0.56U
+ PD=1.04U
.ENDS MUX2_X2

* cell OAI21_X4
* pin A
* pin B2
* pin B1
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT OAI21_X4 1 2 3 5 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 1 5 5 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 11 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 7 3 11 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.31,0.995 PMOS_VTL
M$7 10 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.5,0.995 PMOS_VTL
M$8 5 2 10 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $9 r0 *1 1.69,0.995 PMOS_VTL
M$9 9 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $10 r0 *1 1.88,0.995 PMOS_VTL
M$10 7 3 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $11 r0 *1 2.07,0.995 PMOS_VTL
M$11 8 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $12 r0 *1 2.26,0.995 PMOS_VTL
M$12 5 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $13 r0 *1 0.17,0.2975 NMOS_VTL
M$13 6 1 4 6 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $17 r0 *1 0.93,0.2975 NMOS_VTL
M$17 7 2 4 6 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
* device instance $18 r0 *1 1.12,0.2975 NMOS_VTL
M$18 4 3 7 6 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.1162P PS=2.22U PD=2.22U
.ENDS OAI21_X4

* cell NAND4_X1
* pin A4
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND4_X1 1 2 3 4 5 6 7
* net 1 A4
* net 2 A3
* net 3 A2
* net 4 A1
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 6 2 7 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 7 3 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 6 4 7 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 10 1 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.36,0.2975 NMOS_VTL
M$6 9 2 10 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.55,0.2975 NMOS_VTL
M$7 8 3 9 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.74,0.2975 NMOS_VTL
M$8 7 4 8 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND4_X1

* cell AOI221_X2
* pin B1
* pin B2
* pin A
* pin C2
* pin C1
* pin ZN
* pin NWELL,VDD
* pin PWELL,VSS
.SUBCKT AOI221_X2 1 2 3 4 5 6 8 9
* net 1 B1
* net 2 B2
* net 3 A
* net 4 C2
* net 5 C1
* net 6 ZN
* net 8 NWELL,VDD
* net 9 PWELL,VSS
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 3 10 8 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.09135P PS=2.24U PD=1.55U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 8 1 7 8 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 7 2 8 8 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $7 r0 *1 1.32,0.995 PMOS_VTL
M$7 6 4 10 8 PMOS_VTL L=0.05U W=1.26U AS=0.09135P AD=0.11025P PS=1.55U PD=2.24U
* device instance $8 r0 *1 1.51,0.995 PMOS_VTL
M$8 10 5 6 8 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $11 r0 *1 0.17,0.2975 NMOS_VTL
M$11 6 3 9 9 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.060175P PS=1.595U
+ PD=1.12U
* device instance $12 r0 *1 0.36,0.2975 NMOS_VTL
M$12 14 1 6 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.55,0.2975 NMOS_VTL
M$13 9 2 14 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 0.74,0.2975 NMOS_VTL
M$14 13 2 9 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 0.93,0.2975 NMOS_VTL
M$15 6 1 13 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $17 r0 *1 1.32,0.2975 NMOS_VTL
M$17 12 4 9 9 NMOS_VTL L=0.05U W=0.415U AS=0.031125P AD=0.02905P PS=0.565U
+ PD=0.555U
* device instance $18 r0 *1 1.51,0.2975 NMOS_VTL
M$18 6 5 12 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 1.7,0.2975 NMOS_VTL
M$19 11 5 6 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $20 r0 *1 1.89,0.2975 NMOS_VTL
M$20 9 4 11 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI221_X2

* cell AOI21_X1
* pin A
* pin B2
* pin B1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT AOI21_X1 1 2 3 4 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 4 PWELL,VSS
* net 6 ZN
* net 7 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 6 2 5 7 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 5 3 6 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 7 1 5 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.21,0.2975 NMOS_VTL
M$4 8 2 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.4,0.2975 NMOS_VTL
M$5 6 3 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.59,0.2975 NMOS_VTL
M$6 4 1 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI21_X1

* cell AND3_X1
* pin A1
* pin A2
* pin A3
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND3_X1 1 2 3 5 6 7
* net 1 A1
* net 2 A2
* net 3 A3
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 5 1 4 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 4 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 4 3 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 4 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.195 NMOS_VTL
M$5 8 1 4 6 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $6 r0 *1 0.36,0.195 NMOS_VTL
M$6 9 2 8 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $7 r0 *1 0.55,0.195 NMOS_VTL
M$7 6 3 9 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $8 r0 *1 0.74,0.2975 NMOS_VTL
M$8 7 4 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AND3_X1

* cell OAI21_X1
* pin B2
* pin B1
* pin A
* pin NWELL,VDD
* pin ZN
* pin PWELL,VSS
.SUBCKT OAI21_X1 1 2 3 5 6 7
* net 1 B2
* net 2 B1
* net 3 A
* net 5 NWELL,VDD
* net 6 ZN
* net 7 PWELL,VSS
* device instance $1 r0 *1 0.195,0.995 PMOS_VTL
M$1 8 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.385,0.995 PMOS_VTL
M$2 6 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.575,0.995 PMOS_VTL
M$3 5 3 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.195,0.2975 NMOS_VTL
M$4 6 1 4 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.385,0.2975 NMOS_VTL
M$5 4 2 6 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.575,0.2975 NMOS_VTL
M$6 7 3 4 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI21_X1

* cell OAI21_X2
* pin A
* pin B2
* pin B1
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT OAI21_X2 1 2 3 5 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 1 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 8 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 3 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 9 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 5 2 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.17,0.2975 NMOS_VTL
M$7 6 1 4 6 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $9 r0 *1 0.55,0.2975 NMOS_VTL
M$9 7 2 4 6 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $10 r0 *1 0.74,0.2975 NMOS_VTL
M$10 4 3 7 6 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
.ENDS OAI21_X2

* cell OAI22_X4
* pin PWELL,VSS
* pin B2
* pin B1
* pin A2
* pin ZN
* pin A1
* pin NWELL,VDD
.SUBCKT OAI22_X4 1 3 4 5 6 7 8
* net 1 PWELL,VSS
* net 3 B2
* net 4 B1
* net 5 A2
* net 6 ZN
* net 7 A1
* net 8 NWELL,VDD
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 9 3 8 8 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 6 4 9 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 11 4 6 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 8 3 11 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 10 3 8 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 6 4 10 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.31,0.995 PMOS_VTL
M$7 12 4 6 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.5,0.995 PMOS_VTL
M$8 8 3 12 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $9 r0 *1 1.69,0.995 PMOS_VTL
M$9 13 5 8 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $10 r0 *1 1.88,0.995 PMOS_VTL
M$10 6 7 13 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $11 r0 *1 2.07,0.995 PMOS_VTL
M$11 14 7 6 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $12 r0 *1 2.26,0.995 PMOS_VTL
M$12 8 5 14 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $13 r0 *1 2.45,0.995 PMOS_VTL
M$13 15 5 8 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $14 r0 *1 2.64,0.995 PMOS_VTL
M$14 6 7 15 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $15 r0 *1 2.83,0.995 PMOS_VTL
M$15 16 7 6 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $16 r0 *1 3.02,0.995 PMOS_VTL
M$16 8 5 16 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $17 r0 *1 0.17,0.2975 NMOS_VTL
M$17 1 3 2 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $18 r0 *1 0.36,0.2975 NMOS_VTL
M$18 2 4 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.1162P PS=2.22U PD=2.22U
* device instance $25 r0 *1 1.69,0.2975 NMOS_VTL
M$25 6 5 2 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
* device instance $26 r0 *1 1.88,0.2975 NMOS_VTL
M$26 2 7 6 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.1162P PS=2.22U PD=2.22U
.ENDS OAI22_X4

* cell AOI21_X4
* pin PWELL,VSS
* pin ZN
* pin A
* pin B2
* pin B1
* pin NWELL,VDD
.SUBCKT AOI21_X4 1 2 3 4 5 11
* net 1 PWELL,VSS
* net 2 ZN
* net 3 A
* net 4 B2
* net 5 B1
* net 11 NWELL,VDD
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 11 3 10 11 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.945,0.995 PMOS_VTL
M$5 2 4 10 11 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $6 r0 *1 1.135,0.995 PMOS_VTL
M$6 10 5 2 11 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.1764P PS=3.08U PD=3.08U
* device instance $13 r0 *1 0.185,0.2975 NMOS_VTL
M$13 2 3 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $17 r0 *1 0.945,0.2975 NMOS_VTL
M$17 8 4 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $18 r0 *1 1.135,0.2975 NMOS_VTL
M$18 2 5 8 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 1.325,0.2975 NMOS_VTL
M$19 9 5 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $20 r0 *1 1.515,0.2975 NMOS_VTL
M$20 1 4 9 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $21 r0 *1 1.705,0.2975 NMOS_VTL
M$21 6 4 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $22 r0 *1 1.895,0.2975 NMOS_VTL
M$22 2 5 6 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $23 r0 *1 2.085,0.2975 NMOS_VTL
M$23 7 5 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $24 r0 *1 2.275,0.2975 NMOS_VTL
M$24 1 4 7 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI21_X4
