
* cell configurable_param_fifo
* pin wr_data[5]
* pin rd_data[5]
* pin rd_data[6]
* pin wr_data[1]
* pin wr_data[6]
* pin wr_en
* pin PWELL
* pin NWELL
* pin wr_data[4]
* pin wr_data[2]
* pin clk
* pin rst_n
* pin full
* pin rd_data[4]
* pin rd_data[7]
* pin rd_data[1]
* pin rd_data[2]
* pin almost_full
* pin empty
* pin almost_empty
* pin rd_en
* pin wr_data[7]
* pin wr_data[3]
* pin wr_data[0]
* pin rd_data[3]
* pin rd_data[0]
.SUBCKT configurable_param_fifo 1 2 3 4 5 6 7 8 48 81 149 305 312 321 322 407
+ 431 455 475 496 497 613 617 618 621 622
* net 1 wr_data[5]
* net 2 rd_data[5]
* net 3 rd_data[6]
* net 4 wr_data[1]
* net 5 wr_data[6]
* net 6 wr_en
* net 7 PWELL
* net 8 NWELL
* net 48 wr_data[4]
* net 81 wr_data[2]
* net 149 clk
* net 305 rst_n
* net 312 full
* net 321 rd_data[4]
* net 322 rd_data[7]
* net 407 rd_data[1]
* net 431 rd_data[2]
* net 455 almost_full
* net 475 empty
* net 496 almost_empty
* net 497 rd_en
* net 613 wr_data[7]
* net 617 wr_data[3]
* net 618 wr_data[0]
* net 621 rd_data[3]
* net 622 rd_data[0]
* cell instance $3 m0 *1 249.66,211.4
X$3 1 7 8 15 BUF_X2
* cell instance $8 m0 *1 251.94,4.2
X$8 104 7 8 2 BUF_X1
* cell instance $14 r0 *1 257.07,1.4
X$14 103 7 8 3 BUF_X1
* cell instance $20 m0 *1 255.93,208.6
X$20 4 7 8 16 BUF_X2
* cell instance $28 m0 *1 260.3,208.6
X$28 5 7 8 11 BUF_X2
* cell instance $34 m0 *1 272.27,4.2
X$34 6 8 207 7 BUF_X4
* cell instance $39 m0 *1 271.7,245
X$39 275 268 329 7 8 345 NAND3_X1
* cell instance $44 m0 *1 277.78,245
X$44 344 270 379 8 7 346 HA_X1
* cell instance $45 m0 *1 279.68,245
X$45 346 7 8 359 INV_X1
* cell instance $80 m0 *1 260.11,245
X$80 7 328 361 331 344 8 DFF_X2
* cell instance $82 m0 *1 263.72,245
X$82 344 8 162 7 BUF_X4
* cell instance $85 r0 *1 259.92,245
X$85 123 7 8 358 INV_X2
* cell instance $88 r0 *1 261.06,245
X$88 50 128 362 7 8 375 MUX2_X1
* cell instance $89 r0 *1 262.39,245
X$89 344 369 362 8 7 427 HA_X1
* cell instance $93 r0 *1 269.61,245
X$93 360 358 7 8 376 NOR2_X1
* cell instance $95 r0 *1 270.94,245
X$95 277 296 345 7 8 391 OR3_X1
* cell instance $96 r0 *1 271.89,245
X$96 345 296 277 8 377 7 OAI21_X1
* cell instance $99 r0 *1 276.45,245
X$99 502 292 262 8 378 7 OAI21_X1
* cell instance $101 r0 *1 277.97,245
X$101 380 7 8 384 INV_X1
* cell instance $103 r0 *1 278.54,245
X$103 7 268 381 383 359 386 8 FA_X1
* cell instance $160 m0 *1 272.08,247.8
X$160 358 391 377 7 393 8 AOI21_X1
* cell instance $161 m0 *1 268.47,247.8
X$161 7 376 361 772 329 8 DFF_X2
* cell instance $164 m0 *1 276.64,247.8
X$164 386 268 388 8 7 380 HA_X1
* cell instance $166 m0 *1 279.3,247.8
X$166 388 7 8 385 INV_X1
* cell instance $206 m0 *1 249.09,247.8
X$206 308 172 370 7 8 394 MUX2_X1
* cell instance $207 m0 *1 247.76,247.8
X$207 369 8 122 7 BUF_X4
* cell instance $208 m0 *1 250.42,247.8
X$208 370 162 373 7 8 365 MUX2_X1
* cell instance $209 m0 *1 251.75,247.8
X$209 372 389 395 7 396 8 AOI21_X1
* cell instance $212 r0 *1 247.95,247.8
X$212 7 690 370 394 327 8 DFF_X1
* cell instance $216 r0 *1 252.51,247.8
X$216 146 374 262 8 372 7 OAI21_X1
* cell instance $218 m0 *1 252.89,247.8
X$218 308 165 373 7 8 364 MUX2_X1
* cell instance $224 r0 *1 255.36,247.8
X$224 7 694 374 396 361 8 DFF_X1
* cell instance $226 m0 *1 262.2,247.8
X$226 7 397 361 386 369 8 DFF_X2
* cell instance $227 m0 *1 261.44,247.8
X$227 262 375 8 7 397 AND2_X1
* cell instance $233 r0 *1 272.27,247.8
X$233 401 7 8 390 BUF_X1
* cell instance $237 r0 *1 277.02,247.8
X$237 379 388 390 404 8 7 317 AND4_X2
* cell instance $239 r0 *1 278.54,247.8
X$239 434 382 378 8 413 7 OAI21_X1
* cell instance $240 r0 *1 279.3,247.8
X$240 379 7 8 405 INV_X1
* cell instance $241 r0 *1 279.68,247.8
X$241 346 385 384 8 411 7 OAI21_X1
* cell instance $243 r0 *1 280.82,247.8
X$243 383 405 406 7 409 8 AOI21_X1
* cell instance $295 m0 *1 254.41,228.2
X$295 7 687 204 211 51 8 DFF_X1
* cell instance $297 m0 *1 257.64,228.2
X$297 7 658 187 210 51 8 DFF_X1
* cell instance $336 m0 *1 231.23,228.2
X$336 34 182 160 7 8 199 MUX2_X1
* cell instance $338 m0 *1 232.56,228.2
X$338 183 7 8 765 INV_X1
* cell instance $341 m0 *1 236.17,228.2
X$341 7 666 184 190 183 8 DFF_X1
* cell instance $347 m0 *1 244.53,228.2
X$347 184 122 185 7 8 219 MUX2_X1
* cell instance $350 r0 *1 231.04,228.2
X$350 7 721 160 199 183 8 DFF_X1
* cell instance $351 r0 *1 234.27,228.2
X$351 147 7 8 183 CLKBUF_X3
* cell instance $355 r0 *1 243.2,228.2
X$355 35 121 185 7 8 220 MUX2_X1
* cell instance $357 m0 *1 247.19,228.2
X$357 200 188 202 221 7 8 189 AOI22_X1
* cell instance $359 m0 *1 248.14,228.2
X$359 200 214 202 219 7 8 131 AOI22_X1
* cell instance $363 r0 *1 248.33,228.2
X$363 201 7 8 762 INV_X2
* cell instance $364 r0 *1 248.9,228.2
X$364 7 698 203 217 201 8 DFF_X1
* cell instance $366 m0 *1 250.23,228.2
X$366 35 172 203 7 8 217 MUX2_X1
* cell instance $368 m0 *1 252.51,228.2
X$368 35 165 204 7 8 211 MUX2_X1
* cell instance $370 r0 *1 252.13,228.2
X$370 203 162 204 7 8 214 MUX2_X1
* cell instance $375 r0 *1 264.29,228.2
X$375 147 7 8 205 CLKBUF_X3
* cell instance $376 r0 *1 265.24,228.2
X$376 205 7 8 767 INV_X4
* cell instance $438 m0 *1 251.37,217
X$438 35 67 41 7 8 39 MUX2_X1
* cell instance $440 m0 *1 252.7,217
X$440 41 68 40 7 8 53 MUX2_X1
* cell instance $444 m0 *1 256.5,217
X$444 34 38 69 7 8 52 MUX2_X1
* cell instance $445 m0 *1 257.83,217
X$445 7 667 69 52 51 8 DFF_X1
* cell instance $484 m0 *1 232.18,217
X$484 7 655 64 63 32 8 DFF_X1
* cell instance $491 r0 *1 232.18,217
X$491 34 61 64 7 8 63 MUX2_X1
* cell instance $492 r0 *1 233.51,217
X$492 64 59 20 7 8 87 MUX2_X1
* cell instance $497 m0 *1 244.91,217
X$497 10 50 80 7 8 79 MUX2_X1
* cell instance $498 m0 *1 241.68,217
X$498 7 663 80 37 27 8 DFF_X1
* cell instance $506 r0 *1 246.81,217
X$506 65 53 66 54 7 8 107 AOI22_X1
* cell instance $507 r0 *1 247.76,217
X$507 65 76 66 79 7 8 88 AOI22_X1
* cell instance $510 r0 *1 249.85,217
X$510 65 73 66 44 7 8 89 AOI22_X1
* cell instance $513 r0 *1 257.26,217
X$513 34 67 90 7 8 94 MUX2_X1
* cell instance $514 r0 *1 258.59,217
X$514 90 68 69 7 8 76 MUX2_X1
* cell instance $515 r0 *1 259.92,217
X$515 71 68 70 7 8 73 MUX2_X1
* cell instance $517 r0 *1 261.44,217
X$517 25 67 71 7 8 72 MUX2_X1
* cell instance $519 r0 *1 263.15,217
X$519 7 722 71 72 51 8 DFF_X1
* cell instance $1165 m0 *1 1.9,245
X$1165 347 7 8 322 BUF_X1
* cell instance $1201 m0 *1 206.15,245
X$1201 7 674 336 348 315 8 DFF_X1
* cell instance $1244 m0 *1 209.95,245
X$1244 336 151 367 7 8 337 MUX2_X1
* cell instance $1247 m0 *1 211.47,245
X$1247 337 142 349 7 8 352 MUX2_X1
* cell instance $1252 m0 *1 213.94,245
X$1252 285 7 8 308 BUF_X2
* cell instance $1255 m0 *1 217.17,245
X$1255 7 656 338 351 315 8 DFF_X1
* cell instance $1258 r0 *1 215.46,245
X$1258 308 182 355 7 8 363 MUX2_X1
* cell instance $1259 r0 *1 216.79,245
X$1259 7 701 355 363 315 8 DFF_X1
* cell instance $1260 r0 *1 220.02,245
X$1260 355 159 338 7 8 366 MUX2_X1
* cell instance $1262 m0 *1 224.01,245
X$1262 7 680 339 333 309 8 DFF_X1
* cell instance $1264 m0 *1 227.24,245
X$1264 323 96 97 7 8 340 NOR3_X1
* cell instance $1265 m0 *1 228,245
X$1265 340 115 7 8 341 NOR2_X1
* cell instance $1269 m0 *1 232.56,245
X$1269 59 8 56 7 BUF_X4
* cell instance $1272 m0 *1 235.6,245
X$1272 392 102 8 7 347 AND2_X2
* cell instance $1277 r0 *1 225.34,245
X$1277 59 8 151 7 BUF_X4
* cell instance $1278 r0 *1 226.67,245
X$1278 352 158 366 157 341 389 7 8 OAI221_X2
* cell instance $1283 r0 *1 237.5,245
X$1283 7 749 357 356 309 8 DFF_X1
* cell instance $1285 m0 *1 237.69,245
X$1285 285 139 357 7 8 356 MUX2_X1
* cell instance $1293 r0 *1 241.87,245
X$1293 7 699 342 354 327 8 DFF_X1
* cell instance $1294 m0 *1 242.63,245
X$1294 308 121 342 7 8 354 MUX2_X1
* cell instance $1296 m0 *1 243.96,245
X$1296 357 122 342 7 8 353 MUX2_X1
* cell instance $1304 r0 *1 247.95,245
X$1304 369 7 8 142 INV_X4
* cell instance $1306 r0 *1 249.28,245
X$1306 200 365 202 353 7 8 371 AOI22_X1
* cell instance $1307 r0 *1 250.23,245
X$1307 128 343 371 8 7 395 AND3_X1
* cell instance $1309 m0 *1 250.23,245
X$1309 65 350 66 335 7 8 343 AOI22_X1
* cell instance $1315 r0 *1 251.75,245
X$1315 7 697 373 364 327 8 DFF_X1
* cell instance $1334 m0 *1 241.11,491.4
X$1334 577 7 8 622 BUF_X1
* cell instance $1364 m0 *1 273.79,239.4
X$1364 267 8 258 7 BUF_X4
* cell instance $1366 m0 *1 276.07,239.4
X$1366 298 296 268 7 8 299 MUX2_X1
* cell instance $1367 m0 *1 277.4,239.4
X$1367 262 299 8 7 251 AND2_X1
* cell instance $1369 m0 *1 278.35,239.4
X$1369 270 268 769 8 7 297 HA_X1
* cell instance $1370 m0 *1 280.25,239.4
X$1370 297 8 261 7 BUF_X4
* cell instance $1406 r0 *1 273.79,239.4
X$1406 7 300 205 270 275 8 DFF_X2
* cell instance $8104 r0 *1 196.08,231
X$8104 48 7 8 222 CLKBUF_X2
* cell instance $8111 r0 *1 209.95,231
X$8111 7 720 195 196 180 8 DFF_X1
* cell instance $8127 m0 *1 242.44,231
X$8127 7 648 185 220 201 8 DFF_X1
* cell instance $8131 m0 *1 249.47,231
X$8131 147 7 8 201 CLKBUF_X3
* cell instance $8137 r0 *1 260.3,231
X$8137 7 759 206 208 205 8 DFF_X1
* cell instance $13143 r0 *1 214.7,264.6
X$13143 7 691 586 574 469 8 DFF_X1
* cell instance $13146 r0 *1 218.88,264.6
X$13146 586 159 587 7 8 492 MUX2_X1
* cell instance $13149 r0 *1 220.97,264.6
X$13149 412 182 575 7 8 583 MUX2_X1
* cell instance $13150 r0 *1 222.3,264.6
X$13150 7 736 575 583 469 8 DFF_X1
* cell instance $13151 r0 *1 225.53,264.6
X$13151 575 159 591 7 8 510 MUX2_X1
* cell instance $13156 r0 *1 231.8,264.6
X$13156 594 159 576 7 8 584 MUX2_X1
* cell instance $13160 r0 *1 236.93,264.6
X$13160 490 139 578 7 8 585 MUX2_X1
* cell instance $13163 r0 *1 238.45,264.6
X$13163 7 709 578 585 511 8 DFF_X1
* cell instance $13164 m0 *1 239.21,264.6
X$13164 554 102 8 7 577 AND2_X2
* cell instance $13171 m0 *1 243.01,264.6
X$13171 570 102 8 7 579 AND2_X2
* cell instance $13176 r0 *1 244.53,264.6
X$13176 7 700 556 557 538 8 DFF_X1
* cell instance $13178 m0 *1 244.91,264.6
X$13178 421 121 556 7 8 557 MUX2_X1
* cell instance $13181 m0 *1 247.19,264.6
X$13181 122 8 50 7 BUF_X4
* cell instance $13182 r0 *1 247.76,264.6
X$13182 578 50 556 7 8 582 MUX2_X1
* cell instance $13184 r0 *1 249.09,264.6
X$13184 588 200 202 582 7 8 581 AOI22_X1
* cell instance $13188 r0 *1 252.51,264.6
X$13188 421 165 580 7 8 589 MUX2_X1
* cell instance $13189 r0 *1 253.84,264.6
X$13189 601 162 580 7 8 588 MUX2_X1
* cell instance $16321 r0 *1 243.58,488.6
X$16321 579 7 8 621 BUF_X1
* cell instance $18595 m0 *1 211.09,261.8
X$18595 7 628 531 546 469 8 DFF_X1
* cell instance $18598 m0 *1 221.92,261.8
X$18598 7 653 533 565 469 8 DFF_X1
* cell instance $18602 m0 *1 227.62,261.8
X$18602 7 649 444 527 511 8 DFF_X1
* cell instance $18651 r0 *1 235.41,261.8
X$18651 7 706 554 553 511 8 DFF_X1
* cell instance $18652 m0 *1 235.98,261.8
X$18652 567 534 568 7 553 8 AOI21_X1
* cell instance $18657 r0 *1 238.64,261.8
X$18657 146 554 262 8 567 7 OAI21_X1
* cell instance $18663 m0 *1 242.25,261.8
X$18663 555 524 573 7 569 8 AOI21_X1
* cell instance $18664 m0 *1 243.01,261.8
X$18664 146 570 262 8 555 7 OAI21_X1
* cell instance $18667 r0 *1 240.92,261.8
X$18667 7 718 570 569 538 8 DFF_X1
* cell instance $18669 m0 *1 247.38,261.8
X$18669 128 571 558 8 7 573 AND3_X1
* cell instance $18672 m0 *1 249.09,261.8
X$18672 146 537 581 8 7 568 AND3_X1
* cell instance $18677 m0 *1 252.13,261.8
X$18677 421 38 572 7 8 559 MUX2_X1
* cell instance $18679 m0 *1 253.46,261.8
X$18679 7 626 540 539 538 8 DFF_X1
* cell instance $18683 r0 *1 252.13,261.8
X$18683 7 714 572 559 538 8 DFF_X1
* cell instance $18688 m0 *1 259.35,261.8
X$18688 7 637 560 561 516 8 DFF_X1
* cell instance $18689 m0 *1 264.1,261.8
X$18689 542 38 7 8 564 XOR2_X1
* cell instance $18690 m0 *1 265.24,261.8
X$18690 564 358 7 8 563 NOR2_X1
* cell instance $18691 m0 *1 265.81,261.8
X$18691 7 563 516 771 542 8 DFF_X2
* cell instance $18729 r0 *1 259.35,261.8
X$18729 412 38 566 7 8 562 MUX2_X1
* cell instance $18730 r0 *1 260.68,261.8
X$18730 7 710 566 562 516 8 DFF_X1
* cell instance $18889 r0 *1 213.18,267.4
X$18889 472 7 8 400 CLKBUF_X3
* cell instance $18892 m0 *1 214.51,267.4
X$18892 421 182 586 7 8 574 MUX2_X1
* cell instance $18894 m0 *1 219.07,267.4
X$18894 490 133 587 7 8 597 MUX2_X1
* cell instance $18900 r0 *1 217.74,267.4
X$18900 7 723 587 597 469 8 DFF_X1
* cell instance $18905 r0 *1 223.82,267.4
X$18905 7 729 591 599 511 8 DFF_X1
* cell instance $18906 m0 *1 224.77,267.4
X$18906 532 133 591 7 8 599 MUX2_X1
* cell instance $18910 m0 *1 227.81,267.4
X$18910 490 7 8 421 BUF_X2
* cell instance $18916 m0 *1 228.95,267.4
X$18916 400 182 594 7 8 600 MUX2_X1
* cell instance $18917 r0 *1 229.33,267.4
X$18917 7 717 594 600 511 8 DFF_X1
* cell instance $18918 m0 *1 231.99,267.4
X$18918 7 629 576 593 511 8 DFF_X1
* cell instance $18919 m0 *1 230.66,267.4
X$18919 472 133 576 7 8 593 MUX2_X1
* cell instance $18933 m0 *1 247.19,267.4
X$18933 200 590 202 592 7 8 449 AOI22_X1
* cell instance $18935 m0 *1 248.14,267.4
X$18935 200 598 202 603 7 8 558 AOI22_X1
* cell instance $18940 r0 *1 249.47,267.4
X$18940 612 162 605 7 8 590 MUX2_X1
* cell instance $18942 m0 *1 251.18,267.4
X$18942 7 625 580 589 538 8 DFF_X1
* cell instance $18988 r0 *1 250.99,267.4
X$18988 7 711 601 602 538 8 DFF_X1
* cell instance $18989 r0 *1 254.22,267.4
X$18989 421 172 601 7 8 602 MUX2_X1
* cell instance $18993 r0 *1 258.02,267.4
X$18993 606 162 595 7 8 598 MUX2_X1
* cell instance $18997 r0 *1 261.82,267.4
X$18997 7 708 595 596 516 8 DFF_X1
* cell instance $19167 r0 *1 217.17,273
X$19167 613 7 8 472 BUF_X2
* cell instance $19168 m0 *1 217.74,273
X$19168 618 7 8 490 BUF_X2
* cell instance $19180 r0 *1 226.1,273
X$19180 617 7 8 532 BUF_X2
* cell instance $19195 m0 *1 242.44,273
X$19195 7 627 611 619 538 8 DFF_X1
* cell instance $19392 m0 *1 222.11,270.2
X$19392 532 7 8 412 BUF_X2
* cell instance $19400 m0 *1 233.89,270.2
X$19400 532 139 609 7 8 616 MUX2_X1
* cell instance $19404 r0 *1 235.03,270.2
X$19404 7 712 609 616 511 8 DFF_X1
* cell instance $19406 r0 *1 238.45,270.2
X$19406 7 713 610 620 511 8 DFF_X1
* cell instance $19407 m0 *1 238.83,270.2
X$19407 472 139 610 7 8 620 MUX2_X1
* cell instance $19413 m0 *1 242.06,270.2
X$19413 400 121 608 7 8 604 MUX2_X1
* cell instance $19414 m0 *1 243.39,270.2
X$19414 610 122 608 7 8 592 MUX2_X1
* cell instance $19415 m0 *1 244.72,270.2
X$19415 609 122 611 7 8 603 MUX2_X1
* cell instance $19418 m0 *1 249.28,270.2
X$19418 400 172 612 7 8 615 MUX2_X1
* cell instance $19420 m0 *1 250.8,270.2
X$19420 400 165 605 7 8 614 MUX2_X1
* cell instance $19424 r0 *1 241.68,270.2
X$19424 7 705 608 604 538 8 DFF_X1
* cell instance $19425 r0 *1 244.91,270.2
X$19425 412 121 611 7 8 619 MUX2_X1
* cell instance $19427 r0 *1 246.62,270.2
X$19427 7 716 612 615 538 8 DFF_X1
* cell instance $19428 r0 *1 249.85,270.2
X$19428 7 715 605 614 538 8 DFF_X1
* cell instance $19430 m0 *1 258.4,270.2
X$19430 7 665 606 607 516 8 DFF_X1
* cell instance $19431 m0 *1 257.07,270.2
X$19431 412 172 606 7 8 607 MUX2_X1
* cell instance $19432 m0 *1 261.63,270.2
X$19432 412 165 595 7 8 596 MUX2_X1
* cell instance $19624 m0 *1 208.43,259
X$19624 7 633 507 529 469 8 DFF_X1
* cell instance $19625 m0 *1 211.85,259
X$19625 490 33 530 7 8 544 MUX2_X1
* cell instance $19627 r0 *1 208.43,259
X$19627 400 82 507 7 8 529 MUX2_X1
* cell instance $19630 r0 *1 210.71,259
X$19630 7 727 530 544 469 8 DFF_X1
* cell instance $19632 m0 *1 213.56,259
X$19632 531 56 530 7 8 521 MUX2_X1
* cell instance $19635 r0 *1 213.94,259
X$19635 421 82 531 7 8 546 MUX2_X1
* cell instance $19637 r0 *1 218.31,259
X$19637 7 693 547 545 469 8 DFF_X1
* cell instance $19638 m0 *1 219.26,259
X$19638 532 33 547 7 8 545 MUX2_X1
* cell instance $19640 m0 *1 220.59,259
X$19640 533 56 547 7 8 508 MUX2_X1
* cell instance $19644 m0 *1 225.91,259
X$19644 490 13 509 7 8 549 MUX2_X1
* cell instance $19647 r0 *1 221.54,259
X$19647 412 82 533 7 8 565 MUX2_X1
* cell instance $19651 r0 *1 225.53,259
X$19651 7 735 509 549 511 8 DFF_X1
* cell instance $19652 m0 *1 228.57,259
X$19652 532 13 444 7 8 527 MUX2_X1
* cell instance $19658 m0 *1 235.41,259
X$19658 7 642 513 535 511 8 DFF_X1
* cell instance $19659 m0 *1 234.08,259
X$19659 490 9 513 7 8 535 MUX2_X1
* cell instance $19668 m0 *1 245.67,259
X$19668 513 122 536 7 8 552 MUX2_X1
* cell instance $19669 m0 *1 242.44,259
X$19669 7 638 536 514 327 8 DFF_X1
* cell instance $19673 m0 *1 259.35,259
X$19673 162 8 68 7 BUF_X4
* cell instance $19676 m0 *1 267.52,259
X$19676 517 520 7 8 548 XOR2_X1
* cell instance $19677 m0 *1 268.66,259
X$19677 548 358 7 8 541 NOR2_X1
* cell instance $19681 r0 *1 247.19,259
X$19681 65 550 66 522 7 8 571 AOI22_X1
* cell instance $19684 r0 *1 249.09,259
X$19684 552 66 65 551 7 8 537 AOI22_X1
* cell instance $19687 r0 *1 250.61,259
X$19687 147 7 8 538 CLKBUF_X3
* cell instance $19688 r0 *1 251.56,259
X$19688 538 7 8 CLKBUF_X1
* cell instance $19690 r0 *1 252.51,259
X$19690 540 68 572 7 8 551 MUX2_X1
* cell instance $19691 r0 *1 253.84,259
X$19691 421 67 540 7 8 539 MUX2_X1
* cell instance $19696 r0 *1 258.02,259
X$19696 560 68 566 7 8 550 MUX2_X1
* cell instance $19697 r0 *1 259.35,259
X$19697 412 67 560 7 8 561 MUX2_X1
* cell instance $19701 r0 *1 268.66,259
X$19701 7 541 516 774 517 8 DFF_X2
* cell instance $19703 m0 *1 270.56,259
X$19703 517 542 8 318 7 XOR2_X2
* cell instance $19707 m0 *1 273.6,259
X$19707 543 7 8 102 CLKBUF_X3
* cell instance $19711 m0 *1 276.83,259
X$19711 456 7 8 476 INV_X4
* cell instance $19712 m0 *1 277.78,259
X$19712 7 646 543 519 516 8 DFF_X1
* cell instance $19900 m0 *1 206.72,256.2
X$19900 7 632 489 498 469 8 DFF_X1
* cell instance $19901 m0 *1 205.39,256.2
X$19901 472 33 489 7 8 498 MUX2_X1
* cell instance $19905 m0 *1 212.04,256.2
X$19905 7 623 468 467 469 8 DFF_X1
* cell instance $19909 m0 *1 216.98,256.2
X$19909 501 96 521 7 8 503 MUX2_X1
* cell instance $19912 m0 *1 221.54,256.2
X$19912 491 142 508 7 8 523 MUX2_X1
* cell instance $19916 m0 *1 225.34,256.2
X$19916 503 158 157 492 504 534 7 8 OAI221_X2
* cell instance $19918 m0 *1 227.62,256.2
X$19918 493 115 7 8 504 NOR2_X1
* cell instance $19920 m0 *1 228.95,256.2
X$19920 471 115 7 8 526 NOR2_X1
* cell instance $19928 r0 *1 225.91,256.2
X$19928 523 158 510 157 526 524 7 8 OAI221_X2
* cell instance $19931 m0 *1 232.37,256.2
X$19931 147 7 8 511 CLKBUF_X3
* cell instance $19932 m0 *1 230.66,256.2
X$19932 96 158 7 157 8 NAND2_X4
* cell instance $19939 m0 *1 242.25,256.2
X$19939 421 24 536 7 8 514 MUX2_X1
* cell instance $19943 m0 *1 248.33,256.2
X$19943 7 158 56 451 202 8 NOR3_X4
* cell instance $19944 m0 *1 250.99,256.2
X$19944 7 68 56 451 66 8 NOR3_X4
* cell instance $19948 m0 *1 262.01,256.2
X$19948 494 7 8 128 CLKBUF_X3
* cell instance $19952 r0 *1 233.32,256.2
X$19952 532 9 512 7 8 528 MUX2_X1
* cell instance $19953 r0 *1 234.65,256.2
X$19953 7 740 512 528 511 8 DFF_X1
* cell instance $19955 r0 *1 239.4,256.2
X$19955 412 24 515 7 8 525 MUX2_X1
* cell instance $19956 r0 *1 240.73,256.2
X$19956 7 758 515 525 327 8 DFF_X1
* cell instance $19957 r0 *1 243.96,256.2
X$19957 512 50 515 7 8 522 MUX2_X1
* cell instance $19962 r0 *1 249.66,256.2
X$19962 147 7 8 327 CLKBUF_X3
* cell instance $19963 r0 *1 250.61,256.2
X$19963 327 7 8 764 INV_X2
* cell instance $19966 m0 *1 263.53,256.2
X$19966 494 427 115 159 7 8 520 NAND4_X1
* cell instance $19968 m0 *1 264.48,256.2
X$19968 505 358 7 8 484 NOR2_X1
* cell instance $19973 r0 *1 265.05,256.2
X$19973 147 7 8 516 CLKBUF_X3
* cell instance $19974 r0 *1 266,256.2
X$19974 516 7 8 763 INV_X2
* cell instance $19975 m0 *1 266.38,256.2
X$19975 147 7 8 361 CLKBUF_X3
* cell instance $19977 m0 *1 267.33,256.2
X$19977 361 7 8 CLKBUF_X1
* cell instance $19983 r0 *1 270.37,256.2
X$19983 542 517 7 8 452 XNOR2_X2
* cell instance $19985 m0 *1 273.03,256.2
X$19985 518 317 452 7 494 8 AOI21_X2
* cell instance $19993 m0 *1 277.21,256.2
X$19993 433 502 7 8 495 OR2_X1
* cell instance $19994 m0 *1 277.97,256.2
X$19994 476 358 7 8 500 NOR2_X1
* cell instance $19999 r0 *1 278.16,256.2
X$19999 476 518 358 7 8 519 NOR3_X1
* cell instance $20002 m0 *1 285.19,256.2
X$20002 499 7 8 518 INV_X1
* cell instance $20080 m0 *1 484.69,256.2
X$20080 497 7 8 499 CLKBUF_X3
* cell instance $20179 m0 *1 203.3,253.4
X$20179 7 635 420 432 315 8 DFF_X1
* cell instance $20186 r0 *1 209.38,253.4
X$20186 507 151 489 7 8 466 MUX2_X1
* cell instance $20187 r0 *1 210.71,253.4
X$20187 479 142 466 7 8 480 MUX2_X1
* cell instance $20189 m0 *1 212.42,253.4
X$20189 7 624 422 435 315 8 DFF_X1
* cell instance $20192 m0 *1 216.41,253.4
X$20192 147 7 8 315 CLKBUF_X3
* cell instance $20196 r0 *1 212.42,253.4
X$20196 490 141 468 7 8 467 MUX2_X1
* cell instance $20198 r0 *1 214.13,253.4
X$20198 468 151 422 7 8 501 MUX2_X1
* cell instance $20201 r0 *1 216.6,253.4
X$20201 147 7 8 469 CLKBUF_X3
* cell instance $20202 r0 *1 217.55,253.4
X$20202 7 733 470 458 469 8 DFF_X1
* cell instance $20204 m0 *1 220.02,253.4
X$20204 532 141 470 7 8 458 MUX2_X1
* cell instance $20206 r0 *1 220.78,253.4
X$20206 470 151 423 7 8 491 MUX2_X1
* cell instance $20210 r0 *1 226.1,253.4
X$20210 438 151 509 7 8 485 MUX2_X1
* cell instance $20212 r0 *1 227.62,253.4
X$20212 485 96 97 7 8 493 NOR3_X1
* cell instance $20213 m0 *1 228,253.4
X$20213 414 59 444 7 8 445 MUX2_X1
* cell instance $20216 m0 *1 229.52,253.4
X$20216 7 645 446 487 309 8 DFF_X1
* cell instance $20217 m0 *1 232.75,253.4
X$20217 415 59 446 7 8 463 MUX2_X1
* cell instance $20218 m0 *1 234.08,253.4
X$20218 463 96 97 7 8 447 NOR3_X1
* cell instance $20220 m0 *1 237.88,253.4
X$20220 7 640 448 440 309 8 DFF_X1
* cell instance $20224 m0 *1 243.58,253.4
X$20224 448 50 442 7 8 465 MUX2_X1
* cell instance $20226 m0 *1 246.43,253.4
X$20226 65 461 66 465 7 8 464 AOI22_X1
* cell instance $20227 m0 *1 247.38,253.4
X$20227 128 464 449 8 7 443 AND3_X1
* cell instance $20228 m0 *1 248.33,253.4
X$20228 7 142 426 451 65 8 NOR3_X4
* cell instance $20230 m0 *1 251.18,253.4
X$20230 400 67 450 7 8 462 MUX2_X1
* cell instance $20233 r0 *1 228.76,253.4
X$20233 445 96 97 7 8 471 NOR3_X1
* cell instance $20235 r0 *1 229.9,253.4
X$20235 472 13 446 7 8 487 MUX2_X1
* cell instance $20237 r0 *1 231.42,253.4
X$20237 309 7 8 766 INV_X1
* cell instance $20238 r0 *1 231.8,253.4
X$20238 147 7 8 309 CLKBUF_X3
* cell instance $20239 r0 *1 232.75,253.4
X$20239 157 584 488 480 158 8 7 424 OAI221_X1
* cell instance $20240 r0 *1 233.89,253.4
X$20240 447 115 7 8 488 NOR2_X1
* cell instance $20245 r0 *1 248.33,253.4
X$20245 7 122 426 451 200 8 NOR3_X4
* cell instance $20246 r0 *1 250.99,253.4
X$20246 7 731 450 462 327 8 DFF_X1
* cell instance $20247 m0 *1 253.08,253.4
X$20247 450 68 473 7 8 461 MUX2_X1
* cell instance $20251 r0 *1 254.22,253.4
X$20251 400 38 473 7 8 486 MUX2_X1
* cell instance $20254 r0 *1 256.12,253.4
X$20254 7 732 473 486 361 8 DFF_X1
* cell instance $20255 m0 *1 256.5,253.4
X$20255 115 7 8 451 INV_X4
* cell instance $20257 m0 *1 257.45,253.4
X$20257 59 7 8 426 INV_X2
* cell instance $20260 m0 *1 261.82,253.4
X$20260 426 460 8 7 441 XNOR2_X1
* cell instance $20261 m0 *1 262.96,253.4
X$20261 128 427 7 8 460 NAND2_X1
* cell instance $20265 m0 *1 272.84,253.4
X$20265 459 7 8 404 BUF_X2
* cell instance $20269 r0 *1 261.63,253.4
X$20269 494 159 50 97 7 8 506 NAND4_X1
* cell instance $20270 r0 *1 262.58,253.4
X$20270 451 506 8 7 505 XNOR2_X1
* cell instance $20272 r0 *1 264.1,253.4
X$20272 483 8 115 7 BUF_X4
* cell instance $20273 r0 *1 265.43,253.4
X$20273 7 482 483 484 361 8 DFF_X1
* cell instance $20276 r0 *1 271.89,253.4
X$20276 482 428 459 8 7 481 HA_X1
* cell instance $20278 m0 *1 274.74,253.4
X$20278 317 452 7 8 456 NAND2_X1
* cell instance $20279 m0 *1 273.98,253.4
X$20279 481 403 404 7 457 8 AOI21_X1
* cell instance $20282 m0 *1 277.02,253.4
X$20282 404 429 8 7 478 XNOR2_X1
* cell instance $20286 r0 *1 274.93,253.4
X$20286 457 453 7 8 474 NAND2_X1
* cell instance $20288 r0 *1 275.69,253.4
X$20288 318 474 8 7 502 XNOR2_X1
* cell instance $20291 r0 *1 277.78,253.4
X$20291 478 495 500 8 477 7 OAI21_X1
* cell instance $20292 r0 *1 278.54,253.4
X$20292 7 477 361 775 454 8 DFF_X2
* cell instance $20293 m0 *1 279.49,253.4
X$20293 454 410 430 8 433 7 OAI21_X1
* cell instance $20375 r0 *1 484.88,253.4
X$20375 454 7 8 496 BUF_X1
* cell instance $20379 r0 *1 486.78,253.4
X$20379 476 7 8 475 BUF_X1
* cell instance $20380 m0 *1 487.16,253.4
X$20380 406 7 8 455 BUF_X1
* cell instance $20456 m0 *1 207.48,247.8
X$20456 7 630 367 387 315 8 DFF_X1
* cell instance $20457 m0 *1 210.71,247.8
X$20457 367 179 308 7 8 387 MUX2_X1
* cell instance $20522 r0 *1 230.85,247.8
X$20522 7 746 415 399 309 8 DFF_X1
* cell instance $20524 r0 *1 234.27,247.8
X$20524 7 741 392 425 309 8 DFF_X1
* cell instance $20526 m0 *1 235.22,247.8
X$20526 146 392 123 8 368 7 OAI21_X1
* cell instance $20625 m0 *1 204.82,250.6
X$20625 7 631 398 408 315 8 DFF_X1
* cell instance $20627 m0 *1 208.05,250.6
X$20627 398 179 400 7 8 408 MUX2_X1
* cell instance $20632 m0 *1 224.77,250.6
X$20632 421 61 438 7 8 437 MUX2_X1
* cell instance $20634 m0 *1 226.29,250.6
X$20634 412 61 414 7 8 439 MUX2_X1
* cell instance $20637 m0 *1 231.42,250.6
X$20637 400 61 415 7 8 399 MUX2_X1
* cell instance $20643 r0 *1 204.82,250.6
X$20643 472 141 420 7 8 432 MUX2_X1
* cell instance $20645 r0 *1 206.91,250.6
X$20645 420 151 398 7 8 479 MUX2_X1
* cell instance $20648 r0 *1 214.51,250.6
X$20648 422 179 421 7 8 435 MUX2_X1
* cell instance $20651 r0 *1 217.55,250.6
X$20651 7 695 423 436 315 8 DFF_X1
* cell instance $20652 r0 *1 220.78,250.6
X$20652 423 179 412 7 8 436 MUX2_X1
* cell instance $20654 r0 *1 222.3,250.6
X$20654 7 730 438 437 315 8 DFF_X1
* cell instance $20656 r0 *1 225.72,250.6
X$20656 7 696 414 439 309 8 DFF_X1
* cell instance $20661 r0 *1 235.03,250.6
X$20661 368 424 443 7 425 8 AOI21_X1
* cell instance $20665 r0 *1 238.26,250.6
X$20665 472 9 448 7 8 440 MUX2_X1
* cell instance $20667 r0 *1 241.11,250.6
X$20667 7 752 442 417 327 8 DFF_X1
* cell instance $20668 m0 *1 241.87,250.6
X$20668 400 24 442 7 8 417 MUX2_X1
* cell instance $20674 m0 *1 258.59,250.6
X$20674 418 8 59 7 BUF_X4
* cell instance $20678 m0 *1 262.39,250.6
X$20678 7 416 418 419 361 8 DFF_X1
* cell instance $20681 m0 *1 266.57,250.6
X$20681 374 102 8 7 402 AND2_X2
* cell instance $20688 r0 *1 262.58,250.6
X$20688 441 358 7 8 419 NOR2_X1
* cell instance $20690 r0 *1 269.23,250.6
X$20690 7 704 428 393 361 8 DFF_X1
* cell instance $20691 m0 *1 271.89,250.6
X$20691 416 329 401 8 7 403 HA_X1
* cell instance $20696 r0 *1 272.46,250.6
X$20696 428 8 277 7 BUF_X4
* cell instance $20699 r0 *1 274.93,250.6
X$20699 404 390 381 7 8 453 NAND3_X1
* cell instance $20702 r0 *1 276.26,250.6
X$20702 404 429 7 8 434 XOR2_X1
* cell instance $20704 m0 *1 276.64,250.6
X$20704 403 411 390 7 429 8 AOI21_X2
* cell instance $20705 m0 *1 277.97,250.6
X$20705 7 413 361 773 406 8 DFF_X2
* cell instance $20706 m0 *1 281.58,250.6
X$20706 383 405 7 8 410 NAND2_X1
* cell instance $20742 r0 *1 277.4,250.6
X$20742 381 390 8 7 430 XNOR2_X1
* cell instance $20744 r0 *1 278.73,250.6
X$20744 358 430 409 7 8 382 OR3_X1
* cell instance $20796 m0 *1 484.31,250.6
X$20796 271 7 8 407 BUF_X1
* cell instance $20801 r0 *1 484.31,250.6
X$20801 402 7 8 431 BUF_X1
* cell instance $20923 m0 *1 205.58,219.8
X$20923 7 641 92 93 22 8 DFF_X1
* cell instance $20925 m0 *1 208.81,219.8
X$20925 35 82 92 7 8 93 MUX2_X1
* cell instance $20931 m0 *1 227.05,219.8
X$20931 7 668 62 85 32 8 DFF_X1
* cell instance $20945 r0 *1 208.43,219.8
X$20945 92 56 75 7 8 116 MUX2_X1
* cell instance $20955 r0 *1 243.2,219.8
X$20955 7 702 124 111 27 8 DFF_X1
* cell instance $20958 r0 *1 248.33,219.8
X$20958 7 703 105 100 27 8 DFF_X1
* cell instance $20962 m0 *1 257.64,219.8
X$20962 7 670 90 94 51 8 DFF_X1
* cell instance $20963 m0 *1 261.44,219.8
X$20963 25 38 70 7 8 91 MUX2_X1
* cell instance $20966 m0 *1 262.96,219.8
X$20966 7 664 70 91 51 8 DFF_X1
* cell instance $21309 m0 *1 206.72,233.8
X$21309 222 141 232 7 8 233 MUX2_X1
* cell instance $21311 m0 *1 208.81,233.8
X$21311 232 151 195 7 8 194 MUX2_X1
* cell instance $21312 m0 *1 210.14,233.8
X$21312 195 179 223 7 8 196 MUX2_X1
* cell instance $21315 m0 *1 212.42,233.8
X$21315 222 7 8 223 BUF_X2
* cell instance $21364 r0 *1 204.63,233.8
X$21364 222 33 240 7 8 272 MUX2_X1
* cell instance $21365 r0 *1 205.96,233.8
X$21365 7 707 232 233 180 8 DFF_X1
* cell instance $21367 r0 *1 209.57,233.8
X$21367 194 142 253 7 8 235 MUX2_X1
* cell instance $21370 r0 *1 215.46,233.8
X$21370 223 182 224 7 8 197 MUX2_X1
* cell instance $21371 m0 *1 216.03,233.8
X$21371 7 660 224 197 180 8 DFF_X1
* cell instance $21376 m0 *1 227.62,233.8
X$21376 222 13 198 7 8 226 MUX2_X1
* cell instance $21381 r0 *1 217.93,233.8
X$21381 222 133 225 7 8 242 MUX2_X1
* cell instance $21383 r0 *1 220.02,233.8
X$21383 224 159 225 7 8 255 MUX2_X1
* cell instance $21387 r0 *1 224.96,233.8
X$21387 235 158 255 157 256 244 7 8 OAI221_X2
* cell instance $21389 r0 *1 227.05,233.8
X$21389 7 738 198 226 183 8 DFF_X1
* cell instance $21392 m0 *1 232.37,233.8
X$21392 56 8 159 7 BUF_X4
* cell instance $21393 m0 *1 234.46,233.8
X$21393 7 634 227 239 183 8 DFF_X1
* cell instance $21397 r0 *1 234.08,233.8
X$21397 222 139 227 7 8 239 MUX2_X1
* cell instance $21398 r0 *1 235.41,233.8
X$21398 222 9 257 7 8 280 MUX2_X1
* cell instance $21404 m0 *1 251.94,233.8
X$21404 128 8 146 7 BUF_X4
* cell instance $21405 m0 *1 253.27,233.8
X$21405 223 67 229 7 8 236 MUX2_X1
* cell instance $21408 m0 *1 261.44,233.8
X$21408 223 165 206 7 8 208 MUX2_X1
* cell instance $21409 m0 *1 262.77,233.8
X$21409 231 162 206 7 8 230 MUX2_X1
* cell instance $21451 r0 *1 244.15,233.8
X$21451 223 121 238 7 8 248 MUX2_X1
* cell instance $21454 r0 *1 246.43,233.8
X$21454 227 122 238 7 8 237 MUX2_X1
* cell instance $21455 r0 *1 247.76,233.8
X$21455 200 230 202 237 7 8 249 AOI22_X1
* cell instance $21456 r0 *1 248.71,233.8
X$21456 254 176 186 7 228 8 AOI21_X1
* cell instance $21460 r0 *1 251.94,233.8
X$21460 7 760 229 236 201 8 DFF_X1
* cell instance $21464 r0 *1 259.16,233.8
X$21464 223 172 231 7 8 234 MUX2_X1
* cell instance $21465 r0 *1 260.49,233.8
X$21465 7 739 231 234 205 8 DFF_X1
* cell instance $21569 m0 *1 203.49,236.6
X$21569 7 654 240 272 180 8 DFF_X1
* cell instance $21573 m0 *1 209.19,236.6
X$21573 241 56 240 7 8 253 MUX2_X1
* cell instance $21574 m0 *1 210.52,236.6
X$21574 223 82 241 7 8 273 MUX2_X1
* cell instance $21576 m0 *1 217.93,236.6
X$21576 7 661 225 242 180 8 DFF_X1
* cell instance $21580 m0 *1 223.63,236.6
X$21580 7 662 260 243 180 8 DFF_X1
* cell instance $21622 r0 *1 209.76,236.6
X$21622 7 689 241 273 180 8 DFF_X1
* cell instance $21625 r0 *1 217.55,236.6
X$21625 142 8 96 7 BUF_X4
* cell instance $21630 r0 *1 224.39,236.6
X$21630 223 61 260 7 8 243 MUX2_X1
* cell instance $21632 m0 *1 227.43,236.6
X$21632 260 59 198 7 8 279 MUX2_X1
* cell instance $21634 m0 *1 228.76,236.6
X$21634 279 96 97 7 8 278 NOR3_X1
* cell instance $21635 m0 *1 229.52,236.6
X$21635 278 115 7 8 256 NOR2_X1
* cell instance $21641 r0 *1 231.99,236.6
X$21641 288 261 7 61 8 NAND2_X4
* cell instance $21644 m0 *1 235.79,236.6
X$21644 7 652 257 280 183 8 DFF_X1
* cell instance $21645 m0 *1 239.78,236.6
X$21645 223 24 246 7 8 263 MUX2_X1
* cell instance $21648 m0 *1 241.49,236.6
X$21648 257 50 246 7 8 247 MUX2_X1
* cell instance $21654 r0 *1 238.07,236.6
X$21654 123 7 8 262 CLKBUF_X3
* cell instance $21658 r0 *1 240.35,236.6
X$21658 7 756 246 263 183 8 DFF_X1
* cell instance $21660 m0 *1 244.15,236.6
X$21660 7 657 238 248 201 8 DFF_X1
* cell instance $21662 m0 *1 247.38,236.6
X$21662 128 283 249 8 7 245 AND3_X1
* cell instance $21663 m0 *1 248.33,236.6
X$21663 65 282 66 247 7 8 283 AOI22_X1
* cell instance $21670 r0 *1 248.71,236.6
X$21670 7 737 264 228 201 8 DFF_X1
* cell instance $21671 r0 *1 251.94,236.6
X$21671 146 264 262 8 254 7 OAI21_X1
* cell instance $21673 m0 *1 254.41,236.6
X$21673 229 68 250 7 8 282 MUX2_X1
* cell instance $21675 m0 *1 255.74,236.6
X$21675 223 38 250 7 8 281 MUX2_X1
* cell instance $21676 m0 *1 257.07,236.6
X$21676 7 672 250 281 205 8 DFF_X1
* cell instance $21683 r0 *1 260.68,236.6
X$21683 265 261 7 67 8 NAND2_X4
* cell instance $21685 r0 *1 262.77,236.6
X$21685 265 252 7 38 8 NAND2_X4
* cell instance $21689 m0 *1 271.51,236.6
X$21689 275 268 768 8 7 276 HA_X1
* cell instance $21690 m0 *1 273.41,236.6
X$21690 276 8 252 7 BUF_X4
* cell instance $21692 m0 *1 276.26,236.6
X$21692 7 251 205 269 268 8 DFF_X2
* cell instance $21729 r0 *1 272.65,236.6
X$21729 275 269 770 8 7 267 HA_X1
* cell instance $21730 r0 *1 274.55,236.6
X$21730 274 8 289 7 BUF_X4
* cell instance $21734 r0 *1 277.21,236.6
X$21734 270 269 298 8 7 274 HA_X1
* cell instance $21899 m0 *1 207.86,217
X$21899 7 643 75 55 22 8 DFF_X1
* cell instance $21902 m0 *1 211.28,217
X$21902 7 644 57 74 22 8 DFF_X1
* cell instance $21904 m0 *1 216.03,217
X$21904 11 7 8 25 BUF_X2
* cell instance $21907 m0 *1 217.74,217
X$21907 7 671 58 77 22 8 DFF_X1
* cell instance $21910 r0 *1 207.86,217
X$21910 15 33 75 7 8 55 MUX2_X1
* cell instance $21914 r0 *1 211.85,217
X$21914 25 82 57 7 8 74 MUX2_X1
* cell instance $21915 r0 *1 213.18,217
X$21915 57 56 49 7 8 150 MUX2_X1
* cell instance $21919 r0 *1 218.5,217
X$21919 34 82 58 7 8 77 MUX2_X1
* cell instance $21920 r0 *1 219.83,217
X$21920 58 56 46 7 8 83 MUX2_X1
* cell instance $21922 m0 *1 223.06,217
X$21922 7 683 60 78 22 8 DFF_X1
* cell instance $21928 r0 *1 224.2,217
X$21928 35 61 60 7 8 78 MUX2_X1
* cell instance $21929 r0 *1 225.53,217
X$21929 60 59 31 7 8 84 MUX2_X1
* cell instance $21930 r0 *1 226.86,217
X$21930 25 61 62 7 8 85 MUX2_X1
* cell instance $21936 r0 *1 228.76,217
X$21936 62 59 14 7 8 86 MUX2_X1
* cell instance $21975 m0 *1 206.53,225.4
X$21975 15 141 156 7 8 169 MUX2_X1
* cell instance $22018 r0 *1 203.49,225.4
X$22018 7 745 156 169 180 8 DFF_X1
* cell instance $22020 r0 *1 207.1,225.4
X$22020 156 151 193 7 8 170 MUX2_X1
* cell instance $22022 r0 *1 209.19,225.4
X$22022 170 142 116 7 8 173 MUX2_X1
* cell instance $22024 m0 *1 212.23,225.4
X$22024 117 151 212 7 8 143 MUX2_X1
* cell instance $22026 m0 *1 213.56,225.4
X$22026 143 142 150 7 8 134 MUX2_X1
* cell instance $22030 m0 *1 218.88,225.4
X$22030 95 151 181 7 8 152 MUX2_X1
* cell instance $22034 r0 *1 217.17,225.4
X$22034 147 7 8 180 CLKBUF_X3
* cell instance $22037 r0 *1 218.69,225.4
X$22037 147 7 8 22 CLKBUF_X3
* cell instance $22039 m0 *1 220.78,225.4
X$22039 152 142 83 7 8 155 MUX2_X1
* cell instance $22044 m0 *1 226.1,225.4
X$22044 7 678 144 154 32 8 DFF_X1
* cell instance $22045 m0 *1 224.77,225.4
X$22045 191 159 132 7 8 153 MUX2_X1
* cell instance $22046 m0 *1 229.33,225.4
X$22046 15 133 144 7 8 154 MUX2_X1
* cell instance $22051 r0 *1 226.67,225.4
X$22051 173 158 174 157 113 109 7 8 OAI221_X2
* cell instance $22052 r0 *1 228.76,225.4
X$22052 218 159 144 7 8 174 MUX2_X1
* cell instance $22055 r0 *1 231.99,225.4
X$22055 155 158 177 157 145 176 7 8 OAI221_X2
* cell instance $22056 m0 *1 233.51,225.4
X$22056 119 115 7 8 145 NOR2_X1
* cell instance $22057 m0 *1 232.56,225.4
X$22057 147 7 8 32 CLKBUF_X3
* cell instance $22065 m0 *1 249.66,225.4
X$22065 147 7 8 27 CLKBUF_X3
* cell instance $22066 m0 *1 250.61,225.4
X$22066 27 7 8 CLKBUF_X1
* cell instance $22070 r0 *1 234.08,225.4
X$22070 160 159 138 7 8 177 MUX2_X1
* cell instance $22075 r0 *1 238.26,225.4
X$22075 15 139 184 7 8 190 MUX2_X1
* cell instance $22077 r0 *1 240.35,225.4
X$22077 7 724 161 178 32 8 DFF_X1
* cell instance $22078 r0 *1 243.58,225.4
X$22078 34 121 161 7 8 178 MUX2_X1
* cell instance $22079 r0 *1 244.91,225.4
X$22079 120 122 161 7 8 221 MUX2_X1
* cell instance $22082 r0 *1 247.95,225.4
X$22082 146 88 189 8 7 186 AND3_X1
* cell instance $22084 r0 *1 249.28,225.4
X$22084 200 171 202 130 7 8 175 AOI22_X1
* cell instance $22088 m0 *1 253.84,225.4
X$22088 7 677 163 148 27 8 DFF_X1
* cell instance $22091 m0 *1 259.54,225.4
X$22091 51 7 8 761 INV_X2
* cell instance $22092 m0 *1 260.11,225.4
X$22092 147 7 8 51 CLKBUF_X3
* cell instance $22093 m0 *1 261.06,225.4
X$22093 7 650 164 168 51 8 DFF_X1
* cell instance $22139 r0 *1 254.6,225.4
X$22139 34 172 163 7 8 148 MUX2_X1
* cell instance $22140 r0 *1 255.93,225.4
X$22140 163 162 187 7 8 188 MUX2_X1
* cell instance $22141 r0 *1 257.26,225.4
X$22141 34 165 187 7 8 210 MUX2_X1
* cell instance $22145 r0 *1 259.92,225.4
X$22145 164 162 166 7 8 171 MUX2_X1
* cell instance $22146 r0 *1 261.25,225.4
X$22146 25 172 164 7 8 168 MUX2_X1
* cell instance $22147 r0 *1 262.58,225.4
X$22147 25 165 166 7 8 167 MUX2_X1
* cell instance $22150 r0 *1 265.05,225.4
X$22150 7 734 166 167 205 8 DFF_X1
* cell instance $22294 m0 *1 204.82,228.2
X$22294 7 639 193 209 180 8 DFF_X1
* cell instance $22296 m0 *1 208.05,228.2
X$22296 193 179 35 7 8 209 MUX2_X1
* cell instance $22300 m0 *1 211.85,228.2
X$22300 212 179 25 7 8 213 MUX2_X1
* cell instance $22302 m0 *1 216.22,228.2
X$22302 7 659 181 215 180 8 DFF_X1
* cell instance $22303 m0 *1 219.45,228.2
X$22303 181 179 34 7 8 215 MUX2_X1
* cell instance $22304 m0 *1 220.78,228.2
X$22304 25 182 191 7 8 216 MUX2_X1
* cell instance $22305 m0 *1 222.11,228.2
X$22305 7 675 191 216 183 8 DFF_X1
* cell instance $22306 m0 *1 225.34,228.2
X$22306 7 679 218 192 183 8 DFF_X1
* cell instance $22307 m0 *1 228.57,228.2
X$22307 35 182 218 7 8 192 MUX2_X1
* cell instance $22314 r0 *1 210.71,228.2
X$22314 7 743 212 213 180 8 DFF_X1
* cell instance $22413 r0 *1 210.52,222.6
X$22413 7 744 117 129 22 8 DFF_X1
* cell instance $22414 m0 *1 211.66,222.6
X$22414 11 141 117 7 8 129 MUX2_X1
* cell instance $22420 m0 *1 216.41,222.6
X$22420 7 669 95 108 22 8 DFF_X1
* cell instance $22422 m0 *1 221.35,222.6
X$22422 7 676 132 110 22 8 DFF_X1
* cell instance $22426 m0 *1 227.05,222.6
X$22426 84 96 97 7 8 114 NOR3_X1
* cell instance $22427 m0 *1 227.81,222.6
X$22427 114 115 7 8 113 NOR2_X1
* cell instance $22432 r0 *1 217.74,222.6
X$22432 16 141 95 7 8 108 MUX2_X1
* cell instance $22436 r0 *1 222.68,222.6
X$22436 11 133 132 7 8 110 MUX2_X1
* cell instance $22440 r0 *1 226.1,222.6
X$22440 134 158 153 157 135 118 7 8 OAI221_X2
* cell instance $22442 r0 *1 228.57,222.6
X$22442 136 115 7 8 135 NOR2_X1
* cell instance $22444 m0 *1 229.71,222.6
X$22444 86 96 97 7 8 136 NOR3_X1
* cell instance $22450 r0 *1 230.47,222.6
X$22450 16 133 138 7 8 137 MUX2_X1
* cell instance $22451 r0 *1 231.8,222.6
X$22451 7 726 138 137 32 8 DFF_X1
* cell instance $22453 m0 *1 233.89,222.6
X$22453 87 96 97 7 8 119 NOR3_X1
* cell instance $22459 r0 *1 237.88,222.6
X$22459 16 139 120 7 8 140 MUX2_X1
* cell instance $22460 r0 *1 239.21,222.6
X$22460 7 725 120 140 32 8 DFF_X1
* cell instance $22463 m0 *1 241.87,222.6
X$22463 7 688 98 112 27 8 DFF_X1
* cell instance $22466 m0 *1 248.14,222.6
X$22466 99 109 106 7 100 8 AOI21_X1
* cell instance $22470 m0 *1 251.37,222.6
X$22470 105 102 8 7 104 AND2_X2
* cell instance $22474 r0 *1 242.44,222.6
X$22474 11 139 98 7 8 112 MUX2_X1
* cell instance $22476 r0 *1 243.96,222.6
X$22476 25 121 124 7 8 111 MUX2_X1
* cell instance $22477 r0 *1 245.29,222.6
X$22477 98 122 124 7 8 130 MUX2_X1
* cell instance $22480 r0 *1 247.76,222.6
X$22480 128 107 131 8 7 106 AND3_X1
* cell instance $22482 r0 *1 249.47,222.6
X$22482 146 105 123 8 99 7 OAI21_X1
* cell instance $22484 r0 *1 250.42,222.6
X$22484 128 89 175 8 7 125 AND3_X1
* cell instance $22485 r0 *1 251.37,222.6
X$22485 101 118 125 7 127 8 AOI21_X1
* cell instance $22487 r0 *1 252.32,222.6
X$22487 146 126 123 8 101 7 OAI21_X1
* cell instance $22488 r0 *1 253.08,222.6
X$22488 7 750 126 127 27 8 DFF_X1
* cell instance $22489 m0 *1 255.17,222.6
X$22489 68 8 97 7 BUF_X4
* cell instance $22491 m0 *1 256.5,222.6
X$22491 126 102 8 7 103 AND2_X2
* cell instance $23692 m0 *1 227.81,211.4
X$23692 11 13 14 7 8 19 MUX2_X1
* cell instance $23751 r0 *1 222.11,211.4
X$23751 7 728 31 30 22 8 DFF_X1
* cell instance $23752 r0 *1 225.34,211.4
X$23752 15 13 31 7 8 30 MUX2_X1
* cell instance $23757 r0 *1 227.43,211.4
X$23757 7 753 14 19 32 8 DFF_X1
* cell instance $23760 r0 *1 231.61,211.4
X$23760 7 692 20 21 32 8 DFF_X1
* cell instance $23761 m0 *1 231.99,211.4
X$23761 16 13 20 7 8 21 MUX2_X1
* cell instance $23767 m0 *1 241.3,211.4
X$23767 16 9 10 7 8 12 MUX2_X1
* cell instance $23773 r0 *1 236.93,211.4
X$23773 15 9 23 7 8 29 MUX2_X1
* cell instance $23777 m0 *1 244.53,211.4
X$23777 7 686 18 17 27 8 DFF_X1
* cell instance $23781 r0 *1 246.43,211.4
X$23781 7 719 28 26 27 8 DFF_X1
* cell instance $23989 r0 *1 239.21,208.6
X$23989 7 757 10 12 32 8 DFF_X1
* cell instance $24000 r0 *1 243.58,208.6
X$24000 11 9 18 7 8 17 MUX2_X1
* cell instance $24559 m0 *1 212.8,214.2
X$24559 15 7 8 35 CLKBUF_X3
* cell instance $24604 r0 *1 211.28,214.2
X$24604 7 748 49 42 22 8 DFF_X1
* cell instance $24606 r0 *1 214.7,214.2
X$24606 11 33 49 7 8 42 MUX2_X1
* cell instance $24609 r0 *1 217.74,214.2
X$24609 7 751 46 45 22 8 DFF_X1
* cell instance $24611 m0 *1 218.69,214.2
X$24611 16 33 46 7 8 45 MUX2_X1
* cell instance $24616 m0 *1 236.17,214.2
X$24616 7 636 23 29 32 8 DFF_X1
* cell instance $24617 m0 *1 239.4,214.2
X$24617 35 24 36 7 8 47 MUX2_X1
* cell instance $24622 r0 *1 224.58,214.2
X$24622 16 7 8 34 BUF_X2
* cell instance $24626 r0 *1 237.88,214.2
X$24626 7 747 36 47 32 8 DFF_X1
* cell instance $24627 r0 *1 241.11,214.2
X$24627 23 50 36 7 8 54 MUX2_X1
* cell instance $24631 m0 *1 245.86,214.2
X$24631 25 24 28 7 8 26 MUX2_X1
* cell instance $24636 r0 *1 243.58,214.2
X$24636 34 24 80 7 8 37 MUX2_X1
* cell instance $24639 m0 *1 249.66,214.2
X$24639 7 682 40 43 27 8 DFF_X1
* cell instance $24640 m0 *1 248.33,214.2
X$24640 18 50 28 7 8 44 MUX2_X1
* cell instance $24687 r0 *1 250.61,214.2
X$24687 35 38 40 7 8 43 MUX2_X1
* cell instance $24688 r0 *1 251.94,214.2
X$24688 7 742 41 39 27 8 DFF_X1
* cell instance $24798 m0 *1 201.4,239.4
X$24798 81 7 8 285 CLKBUF_X2
* cell instance $24858 m0 *1 219.45,239.4
X$24858 259 258 7 33 8 NAND2_X4
* cell instance $24860 m0 *1 221.16,239.4
X$24860 252 259 8 7 284 AND2_X1
* cell instance $24861 m0 *1 221.92,239.4
X$24861 288 258 7 82 8 NAND2_X4
* cell instance $24865 r0 *1 219.64,239.4
X$24865 288 252 7 141 8 NAND2_X4
* cell instance $24866 r0 *1 221.35,239.4
X$24866 7 179 8 284 BUF_X8
* cell instance $24871 r0 *1 226.67,239.4
X$24871 285 13 287 7 8 286 MUX2_X1
* cell instance $24875 m0 *1 229.52,239.4
X$24875 288 289 7 182 8 NAND2_X4
* cell instance $24876 m0 *1 227.81,239.4
X$24876 259 289 7 133 8 NAND2_X4
* cell instance $24877 m0 *1 231.23,239.4
X$24877 259 261 7 13 8 NAND2_X4
* cell instance $24879 m0 *1 234.46,239.4
X$24879 303 244 245 7 301 8 AOI21_X1
* cell instance $24881 m0 *1 235.41,239.4
X$24881 146 290 262 8 303 7 OAI21_X1
* cell instance $24889 r0 *1 232.37,239.4
X$24889 7 755 290 301 183 8 DFF_X1
* cell instance $24890 r0 *1 235.6,239.4
X$24890 290 102 8 7 302 AND2_X2
* cell instance $24893 r0 *1 240.35,239.4
X$24893 291 258 7 139 8 NAND2_X4
* cell instance $24896 m0 *1 241.49,239.4
X$24896 291 289 7 9 8 NAND2_X4
* cell instance $24899 m0 *1 244.91,239.4
X$24899 291 261 7 24 8 NAND2_X4
* cell instance $24903 m0 *1 256.5,239.4
X$24903 264 102 8 7 271 AND2_X2
* cell instance $24905 m0 *1 260.49,239.4
X$24905 265 289 7 172 8 NAND2_X4
* cell instance $24906 m0 *1 262.2,239.4
X$24906 265 258 7 165 8 NAND2_X4
* cell instance $24912 r0 *1 243.77,239.4
X$24912 291 252 7 121 8 NAND2_X4
* cell instance $24915 r0 *1 249.28,239.4
X$24915 162 7 8 158 INV_X4
* cell instance $24920 m0 *1 266.57,239.4
X$24920 7 277 292 304 288 8 NOR3_X4
* cell instance $24921 m0 *1 269.23,239.4
X$24921 7 277 292 266 259 8 NOR3_X4
* cell instance $24926 r0 *1 267.9,239.4
X$24926 7 293 292 304 291 8 NOR3_X4
* cell instance $24927 r0 *1 270.56,239.4
X$24927 295 252 207 7 8 294 NAND3_X1
* cell instance $24930 r0 *1 271.89,239.4
X$24930 295 7 8 292 INV_X4
* cell instance $24931 r0 *1 272.84,239.4
X$24931 295 207 7 8 296 NAND2_X1
* cell instance $24934 m0 *1 5.51,242.2
X$24934 302 7 8 321 BUF_X1
* cell instance $24967 m0 *1 203.68,242.2
X$24967 7 647 306 314 315 8 DFF_X1
* cell instance $24968 m0 *1 206.91,242.2
X$24968 285 33 306 7 8 314 MUX2_X1
* cell instance $24970 m0 *1 209.76,242.2
X$24970 7 673 307 316 315 8 DFF_X1
* cell instance $24971 m0 *1 212.99,242.2
X$24971 308 82 307 7 8 316 MUX2_X1
* cell instance $24977 m0 *1 225.91,242.2
X$24977 7 681 287 286 309 8 DFF_X1
* cell instance $25037 r0 *1 207.1,242.2
X$25037 285 141 336 7 8 348 MUX2_X1
* cell instance $25041 r0 *1 210.52,242.2
X$25041 307 56 306 7 8 349 MUX2_X1
* cell instance $25044 r0 *1 218.12,242.2
X$25044 285 133 338 7 8 351 MUX2_X1
* cell instance $25049 r0 *1 224.96,242.2
X$25049 308 61 339 7 8 333 MUX2_X1
* cell instance $25050 r0 *1 226.29,242.2
X$25050 339 59 287 7 8 323 MUX2_X1
* cell instance $25058 r0 *1 231.99,242.2
X$25058 305 7 8 123 BUF_X2
* cell instance $25062 r0 *1 237.69,242.2
X$25062 285 9 310 7 8 324 MUX2_X1
* cell instance $25064 m0 *1 237.88,242.2
X$25064 7 651 310 324 309 8 DFF_X1
* cell instance $25067 m0 *1 242.25,242.2
X$25067 149 7 8 147 CLKBUF_X3
* cell instance $25069 m0 *1 244.72,242.2
X$25069 7 685 326 325 201 8 DFF_X1
* cell instance $25075 r0 *1 244.53,242.2
X$25075 308 24 326 7 8 325 MUX2_X1
* cell instance $25076 r0 *1 245.86,242.2
X$25076 310 50 326 7 8 335 MUX2_X1
* cell instance $25078 m0 *1 251.56,242.2
X$25078 308 38 320 7 8 319 MUX2_X1
* cell instance $25079 m0 *1 248.33,242.2
X$25079 7 684 320 319 201 8 DFF_X1
* cell instance $25080 m0 *1 252.89,242.2
X$25080 308 67 311 7 8 334 MUX2_X1
* cell instance $25088 r0 *1 251.94,242.2
X$25088 311 68 320 7 8 350 MUX2_X1
* cell instance $25089 r0 *1 253.27,242.2
X$25089 7 754 311 334 327 8 DFF_X1
* cell instance $25092 r0 *1 260.3,242.2
X$25092 262 332 8 7 328 AND2_X1
* cell instance $25093 r0 *1 261.06,242.2
X$25093 97 128 331 7 8 332 MUX2_X1
* cell instance $25098 m0 *1 269.04,242.2
X$25098 277 7 8 293 INV_X1
* cell instance $25099 r0 *1 269.04,242.2
X$25099 330 294 8 7 360 XNOR2_X1
* cell instance $25101 m0 *1 269.8,242.2
X$25101 330 207 7 8 304 NAND2_X2
* cell instance $25103 r0 *1 270.94,242.2
X$25103 329 7 8 330 INV_X1
* cell instance $25105 m0 *1 271.13,242.2
X$25105 317 318 266 293 7 8 265 AOI211_X4
* cell instance $25108 r0 *1 271.51,242.2
X$25108 329 207 7 8 266 NAND2_X1
* cell instance $25111 m0 *1 274.36,242.2
X$25111 317 318 7 8 295 NAND2_X2
* cell instance $25112 m0 *1 275.5,242.2
X$25112 262 313 8 7 300 AND2_X1
* cell instance $25113 m0 *1 276.26,242.2
X$25113 270 296 275 7 8 313 MUX2_X1
* cell instance $25202 m0 *1 484.5,242.2
X$25202 292 7 8 312 BUF_X1
.ENDS configurable_param_fifo

* cell NAND2_X2
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND2_X2 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.195,0.995 PMOS_VTL
M$1 5 1 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.11025P PS=2.24U PD=2.24U
* device instance $2 r0 *1 0.385,0.995 PMOS_VTL
M$2 4 2 5 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $5 r0 *1 0.195,0.2975 NMOS_VTL
M$5 7 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.385,0.2975 NMOS_VTL
M$6 5 2 7 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.575,0.2975 NMOS_VTL
M$7 6 2 5 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.765,0.2975 NMOS_VTL
M$8 3 1 6 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND2_X2

* cell AOI211_X4
* pin C1
* pin C2
* pin B
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT AOI211_X4 1 2 3 4 8 9 10
* net 1 C1
* net 2 C2
* net 3 B
* net 4 A
* net 8 PWELL,VSS
* net 9 NWELL,VDD
* net 10 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 6 1 7 9 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 7 2 6 9 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 11 3 7 9 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 9 4 11 9 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 5 6 9 9 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $7 r0 *1 1.31,0.995 PMOS_VTL
M$7 10 5 9 9 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $11 r0 *1 0.17,0.2975 NMOS_VTL
M$11 12 1 6 8 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $12 r0 *1 0.36,0.2975 NMOS_VTL
M$12 8 2 12 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.55,0.2975 NMOS_VTL
M$13 6 3 8 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 0.74,0.2975 NMOS_VTL
M$14 8 4 6 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 0.93,0.2975 NMOS_VTL
M$15 5 6 8 8 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $17 r0 *1 1.31,0.2975 NMOS_VTL
M$17 10 5 8 8 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U
+ PD=2.705U
.ENDS AOI211_X4

* cell CLKBUF_X2
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT CLKBUF_X2 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.17,0.1875 NMOS_VTL
M$4 3 1 2 3 NMOS_VTL L=0.05U W=0.195U AS=0.020475P AD=0.01365P PS=0.6U PD=0.335U
* device instance $5 r0 *1 0.36,0.1875 NMOS_VTL
M$5 5 2 3 3 NMOS_VTL L=0.05U W=0.39U AS=0.0273P AD=0.034125P PS=0.67U PD=0.935U
.ENDS CLKBUF_X2

* cell BUF_X8
* pin PWELL,VSS
* pin Z
* pin NWELL,VDD
* pin A
.SUBCKT BUF_X8 1 3 4 5
* net 1 PWELL,VSS
* net 3 Z
* net 4 NWELL,VDD
* net 5 A
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 2 5 4 4 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 3 2 4 4 PMOS_VTL L=0.05U W=5.04U AS=0.3528P AD=0.37485P PS=6.16U PD=6.86U
* device instance $13 r0 *1 0.17,0.2975 NMOS_VTL
M$13 2 5 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $17 r0 *1 0.93,0.2975 NMOS_VTL
M$17 3 2 1 1 NMOS_VTL L=0.05U W=3.32U AS=0.2324P AD=0.246925P PS=4.44U PD=4.925U
.ENDS BUF_X8

* cell OAI221_X1
* pin B2
* pin B1
* pin A
* pin C2
* pin C1
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT OAI221_X1 1 2 3 4 5 7 8 9
* net 1 B2
* net 2 B1
* net 3 A
* net 4 C2
* net 5 C1
* net 7 NWELL,VDD
* net 8 PWELL,VSS
* net 9 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 12 1 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 9 2 12 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 7 3 9 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 11 4 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 9 5 11 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.17,0.2975 NMOS_VTL
M$6 8 1 6 8 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $7 r0 *1 0.36,0.2975 NMOS_VTL
M$7 6 2 8 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.55,0.2975 NMOS_VTL
M$8 10 3 6 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.74,0.2975 NMOS_VTL
M$9 9 4 10 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.93,0.2975 NMOS_VTL
M$10 10 5 9 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI221_X1

* cell NOR3_X1
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NOR3_X1 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 8 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 7 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.2975 NMOS_VTL
M$4 6 1 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.36,0.2975 NMOS_VTL
M$5 4 2 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 3 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NOR3_X1

* cell NAND2_X1
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND2_X1 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 5 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 4 2 5 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.185,0.2975 NMOS_VTL
M$3 6 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $4 r0 *1 0.375,0.2975 NMOS_VTL
M$4 5 2 6 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND2_X1

* cell XNOR2_X2
* pin A
* pin B
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT XNOR2_X2 2 3 4 5 7
* net 2 A
* net 3 B
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 1.135,0.995 PMOS_VTL
M$1 7 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 1.325,0.995 PMOS_VTL
M$2 9 2 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 1.515,0.995 PMOS_VTL
M$3 5 3 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 1.705,0.995 PMOS_VTL
M$4 8 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.18,0.995 PMOS_VTL
M$5 7 1 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $7 r0 *1 0.56,0.995 PMOS_VTL
M$7 1 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 0.75,0.995 PMOS_VTL
M$8 5 2 1 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 1.135,0.2975 NMOS_VTL
M$9 6 2 7 4 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $11 r0 *1 1.515,0.2975 NMOS_VTL
M$11 6 3 7 4 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $13 r0 *1 0.18,0.2975 NMOS_VTL
M$13 6 1 4 4 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $15 r0 *1 0.56,0.2975 NMOS_VTL
M$15 10 3 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 0.75,0.2975 NMOS_VTL
M$16 1 2 10 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS XNOR2_X2

* cell AND2_X2
* pin A1
* pin A2
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND2_X2 1 2 4 5 6
* net 1 A1
* net 2 A2
* net 4 NWELL,VDD
* net 5 PWELL,VSS
* net 6 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 3 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 4 2 3 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 7 1 3 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.36,0.2975 NMOS_VTL
M$6 5 2 7 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.55,0.2975 NMOS_VTL
M$7 6 3 5 5 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS AND2_X2

* cell BUF_X2
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT BUF_X2 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 4 1 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.21,0.2975 NMOS_VTL
M$4 3 1 2 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.4,0.2975 NMOS_VTL
M$5 5 2 3 3 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS BUF_X2

* cell BUF_X1
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT BUF_X1 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 2 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.033075P PS=0.77U
+ PD=0.84U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.17,0.195 NMOS_VTL
M$3 3 1 2 3 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.021875P PS=0.63U PD=0.555U
* device instance $4 r0 *1 0.36,0.2975 NMOS_VTL
M$4 5 2 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS BUF_X1

* cell XOR2_X2
* pin B
* pin A
* pin NWELL,VDD
* pin Z
* pin PWELL,VSS
.SUBCKT XOR2_X2 1 2 4 5 7
* net 1 B
* net 2 A
* net 4 NWELL,VDD
* net 5 Z
* net 7 PWELL,VSS
* device instance $1 r0 *1 0.2,0.995 PMOS_VTL
M$1 8 2 3 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.39,0.995 PMOS_VTL
M$2 4 1 8 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.58,0.995 PMOS_VTL
M$3 6 3 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.77,0.995 PMOS_VTL
M$4 5 2 6 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $5 r0 *1 0.96,0.995 PMOS_VTL
M$5 6 1 5 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $9 r0 *1 0.2,0.2975 NMOS_VTL
M$9 3 2 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $10 r0 *1 0.39,0.2975 NMOS_VTL
M$10 7 1 3 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.58,0.2975 NMOS_VTL
M$11 5 3 7 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $12 r0 *1 0.77,0.2975 NMOS_VTL
M$12 10 2 5 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.96,0.2975 NMOS_VTL
M$13 7 1 10 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 1.15,0.2975 NMOS_VTL
M$14 9 1 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 1.34,0.2975 NMOS_VTL
M$15 5 2 9 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
.ENDS XOR2_X2

* cell NAND3_X1
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND3_X1 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 6 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.2975 NMOS_VTL
M$4 8 1 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.36,0.2975 NMOS_VTL
M$5 7 2 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 3 7 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND3_X1

* cell CLKBUF_X1
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT CLKBUF_X1 1 3 4
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.19,1.1525 PMOS_VTL
M$1 2 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.033075P PS=0.77U
+ PD=0.84U
* device instance $2 r0 *1 0.38,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.19,0.2075 NMOS_VTL
M$3 3 1 2 3 NMOS_VTL L=0.05U W=0.095U AS=0.009975P AD=0.01015P PS=0.4U PD=0.335U
* device instance $4 r0 *1 0.38,0.2575 NMOS_VTL
M$4 5 2 3 3 NMOS_VTL L=0.05U W=0.195U AS=0.01015P AD=0.020475P PS=0.335U PD=0.6U
.ENDS CLKBUF_X1

* cell CLKBUF_X3
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT CLKBUF_X3 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=1.89U AS=0.1323P AD=0.15435P PS=2.31U PD=3.01U
* device instance $5 r0 *1 0.17,0.1875 NMOS_VTL
M$5 3 1 2 3 NMOS_VTL L=0.05U W=0.195U AS=0.020475P AD=0.01365P PS=0.6U PD=0.335U
* device instance $6 r0 *1 0.36,0.1875 NMOS_VTL
M$6 5 2 3 3 NMOS_VTL L=0.05U W=0.585U AS=0.04095P AD=0.047775P PS=1.005U
+ PD=1.27U
.ENDS CLKBUF_X3

* cell NOR3_X4
* pin PWELL,VSS
* pin A1
* pin A2
* pin A3
* pin ZN
* pin NWELL,VDD
.SUBCKT NOR3_X4 1 2 3 4 5 8
* net 1 PWELL,VSS
* net 2 A1
* net 3 A2
* net 4 A3
* net 5 ZN
* net 8 NWELL,VDD
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 5 2 7 8 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 6 3 7 8 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $9 r0 *1 1.875,0.995 PMOS_VTL
M$9 6 4 8 8 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.19845P PS=3.78U PD=3.78U
* device instance $13 r0 *1 1.875,0.2975 NMOS_VTL
M$13 5 4 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.130725P PS=2.705U
+ PD=2.705U
* device instance $17 r0 *1 0.17,0.2975 NMOS_VTL
M$17 5 2 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $21 r0 *1 0.93,0.2975 NMOS_VTL
M$21 5 3 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS NOR3_X4

* cell NAND4_X1
* pin A4
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND4_X1 1 2 3 4 5 6 7
* net 1 A4
* net 2 A3
* net 3 A2
* net 4 A1
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 6 2 7 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 7 3 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 6 4 7 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 10 1 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.36,0.2975 NMOS_VTL
M$6 9 2 10 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.55,0.2975 NMOS_VTL
M$7 8 3 9 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.74,0.2975 NMOS_VTL
M$8 7 4 8 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND4_X1

* cell XOR2_X1
* pin A
* pin B
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT XOR2_X1 1 3 4 5 6
* net 1 A
* net 3 B
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 Z
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 8 1 2 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 8 3 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.0338625P AD=0.02205P PS=0.775U
+ PD=0.455U
* device instance $3 r0 *1 0.555,0.995 PMOS_VTL
M$3 7 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0338625P AD=0.0441P PS=0.775U PD=0.77U
* device instance $4 r0 *1 0.745,0.995 PMOS_VTL
M$4 6 1 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.935,0.995 PMOS_VTL
M$5 7 3 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.17,0.195 NMOS_VTL
M$6 2 1 4 4 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $7 r0 *1 0.36,0.195 NMOS_VTL
M$7 4 3 2 4 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0224P PS=0.35U PD=0.56U
* device instance $8 r0 *1 0.555,0.2975 NMOS_VTL
M$8 6 2 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.0224P AD=0.02905P PS=0.56U PD=0.555U
* device instance $9 r0 *1 0.745,0.2975 NMOS_VTL
M$9 9 1 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.935,0.2975 NMOS_VTL
M$10 4 3 9 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS XOR2_X1

* cell AOI21_X2
* pin A
* pin B2
* pin B1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT AOI21_X2 1 2 3 4 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 4 PWELL,VSS
* net 6 ZN
* net 7 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 7 1 5 7 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 6 2 5 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 5 3 6 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $7 r0 *1 0.21,0.2975 NMOS_VTL
M$7 6 1 4 4 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $9 r0 *1 0.59,0.2975 NMOS_VTL
M$9 9 2 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.78,0.2975 NMOS_VTL
M$10 6 3 9 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.97,0.2975 NMOS_VTL
M$11 8 3 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 1.16,0.2975 NMOS_VTL
M$12 4 2 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI21_X2

* cell OR2_X1
* pin A1
* pin A2
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR2_X1 1 2 3 5 6
* net 1 A1
* net 2 A2
* net 3 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 7 1 4 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 7 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 4 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.195 NMOS_VTL
M$4 4 1 3 3 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $5 r0 *1 0.36,0.195 NMOS_VTL
M$5 3 2 4 3 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 4 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OR2_X1

* cell XNOR2_X1
* pin A
* pin B
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT XNOR2_X1 1 2 4 5 7
* net 1 A
* net 2 B
* net 4 NWELL,VDD
* net 5 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.18,1.1525 PMOS_VTL
M$1 3 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.37,1.1525 PMOS_VTL
M$2 3 2 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.0338625P AD=0.02205P PS=0.775U
+ PD=0.455U
* device instance $3 r0 *1 0.565,0.995 PMOS_VTL
M$3 7 3 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.0338625P AD=0.0441P PS=0.775U PD=0.77U
* device instance $4 r0 *1 0.755,0.995 PMOS_VTL
M$4 8 1 7 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.945,0.995 PMOS_VTL
M$5 4 2 8 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.18,0.195 NMOS_VTL
M$6 9 1 3 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $7 r0 *1 0.37,0.195 NMOS_VTL
M$7 5 2 9 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0224P PS=0.35U PD=0.56U
* device instance $8 r0 *1 0.565,0.2975 NMOS_VTL
M$8 6 3 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.0224P AD=0.02905P PS=0.56U PD=0.555U
* device instance $9 r0 *1 0.755,0.2975 NMOS_VTL
M$9 7 1 6 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.945,0.2975 NMOS_VTL
M$10 6 2 7 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS XNOR2_X1

* cell AND4_X2
* pin A1
* pin A2
* pin A3
* pin A4
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND4_X2 1 2 3 4 6 7 8
* net 1 A1
* net 2 A2
* net 3 A3
* net 4 A4
* net 6 NWELL,VDD
* net 7 PWELL,VSS
* net 8 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 5 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 6 2 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 5 3 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 6 4 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 8 5 6 6 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $7 r0 *1 0.17,0.2975 NMOS_VTL
M$7 11 1 5 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $8 r0 *1 0.36,0.2975 NMOS_VTL
M$8 10 2 11 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.55,0.2975 NMOS_VTL
M$9 9 3 10 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.74,0.2975 NMOS_VTL
M$10 7 4 9 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.93,0.2975 NMOS_VTL
M$11 8 5 7 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS AND4_X2

* cell DFF_X1
* pin PWELL,VSS
* pin QN
* pin Q
* pin D
* pin CK
* pin NWELL,VDD
.SUBCKT DFF_X1 1 8 9 14 15 16
* net 1 PWELL,VSS
* net 8 QN
* net 9 Q
* net 14 D
* net 15 CK
* net 16 NWELL,VDD
* device instance $1 r0 *1 2.85,0.995 PMOS_VTL
M$1 16 6 8 16 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 3.04,0.995 PMOS_VTL
M$2 9 7 16 16 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.185,0.9425 PMOS_VTL
M$3 16 5 2 16 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.014175P PS=0.84U
+ PD=0.455U
* device instance $4 r0 *1 0.375,1.055 PMOS_VTL
M$4 17 3 16 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.0063P PS=0.455U
+ PD=0.23U
* device instance $5 r0 *1 0.565,1.055 PMOS_VTL
M$5 17 5 4 16 PMOS_VTL L=0.05U W=0.09U AS=0.018075P AD=0.0063P PS=0.565U
+ PD=0.23U
* device instance $6 r0 *1 0.76,0.975 PMOS_VTL
M$6 18 2 4 16 PMOS_VTL L=0.05U W=0.42U AS=0.018075P AD=0.0294P PS=0.565U
+ PD=0.56U
* device instance $7 r0 *1 0.95,0.975 PMOS_VTL
M$7 16 14 18 16 PMOS_VTL L=0.05U W=0.42U AS=0.0294P AD=0.025725P PS=0.56U
+ PD=0.56U
* device instance $8 r0 *1 1.14,1.0275 PMOS_VTL
M$8 3 4 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.025725P AD=0.0567P PS=0.56U
+ PD=0.99U
* device instance $9 r0 *1 1.555,1.0275 PMOS_VTL
M$9 16 15 5 16 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $10 r0 *1 1.745,1.0275 PMOS_VTL
M$10 19 4 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $11 r0 *1 1.935,1.0275 PMOS_VTL
M$11 6 5 19 16 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.014175P PS=0.455U
+ PD=0.455U
* device instance $12 r0 *1 2.125,1.14 PMOS_VTL
M$12 20 2 6 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.006525P PS=0.455U
+ PD=0.235U
* device instance $13 r0 *1 2.32,1.14 PMOS_VTL
M$13 20 7 16 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.006525P PS=0.455U
+ PD=0.235U
* device instance $14 r0 *1 2.51,1.0275 PMOS_VTL
M$14 7 6 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.014175P AD=0.033075P PS=0.455U
+ PD=0.84U
* device instance $15 r0 *1 2.85,0.2975 NMOS_VTL
M$15 1 6 8 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $16 r0 *1 3.04,0.2975 NMOS_VTL
M$16 9 7 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
* device instance $17 r0 *1 0.185,0.285 NMOS_VTL
M$17 1 5 2 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0105P PS=0.63U PD=0.35U
* device instance $18 r0 *1 0.375,0.345 NMOS_VTL
M$18 10 3 1 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.0063P PS=0.35U PD=0.23U
* device instance $19 r0 *1 0.565,0.345 NMOS_VTL
M$19 10 2 4 1 NMOS_VTL L=0.05U W=0.09U AS=0.013P AD=0.0063P PS=0.42U PD=0.23U
* device instance $20 r0 *1 1.14,0.285 NMOS_VTL
M$20 3 4 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.016975P AD=0.02205P PS=0.415U
+ PD=0.63U
* device instance $21 r0 *1 0.76,0.3175 NMOS_VTL
M$21 11 5 4 1 NMOS_VTL L=0.05U W=0.275U AS=0.013P AD=0.01925P PS=0.42U PD=0.415U
* device instance $22 r0 *1 0.95,0.3175 NMOS_VTL
M$22 1 14 11 1 NMOS_VTL L=0.05U W=0.275U AS=0.01925P AD=0.016975P PS=0.415U
+ PD=0.415U
* device instance $23 r0 *1 2.125,0.345 NMOS_VTL
M$23 12 5 6 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.006525P PS=0.35U
+ PD=0.235U
* device instance $24 r0 *1 2.32,0.345 NMOS_VTL
M$24 12 7 1 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.006525P PS=0.35U
+ PD=0.235U
* device instance $25 r0 *1 1.555,0.36 NMOS_VTL
M$25 1 15 5 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $26 r0 *1 1.745,0.36 NMOS_VTL
M$26 13 4 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $27 r0 *1 1.935,0.36 NMOS_VTL
M$27 6 2 13 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0105P PS=0.35U PD=0.35U
* device instance $28 r0 *1 2.51,0.36 NMOS_VTL
M$28 7 6 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0105P AD=0.02205P PS=0.35U PD=0.63U
.ENDS DFF_X1

* cell DFF_X2
* pin PWELL,VSS
* pin D
* pin CK
* pin QN
* pin Q
* pin NWELL,VDD
.SUBCKT DFF_X2 1 6 8 10 11 16
* net 1 PWELL,VSS
* net 6 D
* net 8 CK
* net 10 QN
* net 11 Q
* net 16 NWELL,VDD
* device instance $1 r0 *1 2.855,0.995 PMOS_VTL
M$1 10 9 16 16 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $3 r0 *1 3.235,0.995 PMOS_VTL
M$3 11 2 16 16 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $5 r0 *1 0.2,0.9275 PMOS_VTL
M$5 16 7 3 16 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.014175P PS=0.84U
+ PD=0.455U
* device instance $6 r0 *1 0.39,1.04 PMOS_VTL
M$6 17 4 16 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.0063P PS=0.455U
+ PD=0.23U
* device instance $7 r0 *1 0.58,1.04 PMOS_VTL
M$7 17 7 5 16 PMOS_VTL L=0.05U W=0.09U AS=0.01785P AD=0.0063P PS=0.56U PD=0.23U
* device instance $8 r0 *1 0.77,0.975 PMOS_VTL
M$8 18 3 5 16 PMOS_VTL L=0.05U W=0.42U AS=0.01785P AD=0.0294P PS=0.56U PD=0.56U
* device instance $9 r0 *1 0.96,0.975 PMOS_VTL
M$9 16 6 18 16 PMOS_VTL L=0.05U W=0.42U AS=0.0294P AD=0.025725P PS=0.56U
+ PD=0.56U
* device instance $10 r0 *1 1.15,1.0275 PMOS_VTL
M$10 4 5 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.025725P AD=0.0567P PS=0.56U
+ PD=0.99U
* device instance $11 r0 *1 2.135,0.915 PMOS_VTL
M$11 20 3 9 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.0063P PS=0.455U
+ PD=0.23U
* device instance $12 r0 *1 2.325,0.915 PMOS_VTL
M$12 20 2 16 16 PMOS_VTL L=0.05U W=0.09U AS=0.0252P AD=0.0063P PS=0.77U PD=0.23U
* device instance $13 r0 *1 1.565,1.0275 PMOS_VTL
M$13 16 8 7 16 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $14 r0 *1 1.755,1.0275 PMOS_VTL
M$14 19 5 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $15 r0 *1 1.945,1.0275 PMOS_VTL
M$15 9 7 19 16 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.014175P PS=0.455U
+ PD=0.455U
* device instance $16 r0 *1 2.515,0.995 PMOS_VTL
M$16 2 9 16 16 PMOS_VTL L=0.05U W=0.63U AS=0.0252P AD=0.06615P PS=0.77U PD=1.47U
* device instance $17 r0 *1 2.855,0.2975 NMOS_VTL
M$17 10 9 1 1 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U
+ PD=1.11U
* device instance $19 r0 *1 3.235,0.2975 NMOS_VTL
M$19 11 2 1 1 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U
+ PD=1.595U
* device instance $21 r0 *1 0.39,0.31 NMOS_VTL
M$21 12 4 1 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.0063P PS=0.35U PD=0.23U
* device instance $22 r0 *1 0.58,0.31 NMOS_VTL
M$22 12 3 5 1 NMOS_VTL L=0.05U W=0.09U AS=0.012775P AD=0.0063P PS=0.415U
+ PD=0.23U
* device instance $23 r0 *1 1.15,0.25 NMOS_VTL
M$23 4 5 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.016975P AD=0.02205P PS=0.415U
+ PD=0.63U
* device instance $24 r0 *1 0.77,0.2825 NMOS_VTL
M$24 13 7 5 1 NMOS_VTL L=0.05U W=0.275U AS=0.012775P AD=0.01925P PS=0.415U
+ PD=0.415U
* device instance $25 r0 *1 0.96,0.2825 NMOS_VTL
M$25 1 6 13 1 NMOS_VTL L=0.05U W=0.275U AS=0.01925P AD=0.016975P PS=0.415U
+ PD=0.415U
* device instance $26 r0 *1 0.2,0.37 NMOS_VTL
M$26 1 7 3 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0105P PS=0.63U PD=0.35U
* device instance $27 r0 *1 1.565,0.35 NMOS_VTL
M$27 1 8 7 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $28 r0 *1 1.755,0.35 NMOS_VTL
M$28 14 5 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $29 r0 *1 1.945,0.35 NMOS_VTL
M$29 9 3 14 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0105P PS=0.35U PD=0.35U
* device instance $30 r0 *1 2.135,0.41 NMOS_VTL
M$30 15 7 9 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.0063P PS=0.35U PD=0.23U
* device instance $31 r0 *1 2.325,0.41 NMOS_VTL
M$31 15 2 1 1 NMOS_VTL L=0.05U W=0.09U AS=0.017675P AD=0.0063P PS=0.555U
+ PD=0.23U
* device instance $32 r0 *1 2.515,0.2975 NMOS_VTL
M$32 2 9 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.017675P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS DFF_X2

* cell HA_X1
* pin A
* pin B
* pin S
* pin NWELL,VDD
* pin PWELL,VSS
* pin CO
.SUBCKT HA_X1 1 2 4 5 6 9
* net 1 A
* net 2 B
* net 4 S
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 9 CO
* device instance $1 r0 *1 0.785,1.0275 PMOS_VTL
M$1 10 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.0338625P AD=0.02205P PS=0.775U
+ PD=0.455U
* device instance $2 r0 *1 0.975,1.0275 PMOS_VTL
M$2 7 1 10 5 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.033075P PS=0.455U
+ PD=0.84U
* device instance $3 r0 *1 0.21,0.995 PMOS_VTL
M$3 4 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $4 r0 *1 0.4,0.995 PMOS_VTL
M$4 3 1 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.59,0.995 PMOS_VTL
M$5 5 7 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0338625P PS=0.77U PD=0.775U
* device instance $6 r0 *1 1.345,1.0275 PMOS_VTL
M$6 8 1 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $7 r0 *1 1.535,1.0275 PMOS_VTL
M$7 8 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $8 r0 *1 1.725,0.995 PMOS_VTL
M$8 9 8 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 0.785,0.195 NMOS_VTL
M$9 7 2 6 6 NMOS_VTL L=0.05U W=0.21U AS=0.0224P AD=0.0147P PS=0.56U PD=0.35U
* device instance $10 r0 *1 0.975,0.195 NMOS_VTL
M$10 6 1 7 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.02205P PS=0.35U PD=0.63U
* device instance $11 r0 *1 0.21,0.2975 NMOS_VTL
M$11 11 2 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $12 r0 *1 0.4,0.2975 NMOS_VTL
M$12 4 1 11 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.59,0.2975 NMOS_VTL
M$13 6 7 4 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.0224P PS=0.555U PD=0.56U
* device instance $14 r0 *1 1.345,0.195 NMOS_VTL
M$14 12 1 8 6 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $15 r0 *1 1.535,0.195 NMOS_VTL
M$15 6 2 12 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
* device instance $16 r0 *1 1.725,0.2975 NMOS_VTL
M$16 9 8 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS HA_X1

* cell FA_X1
* pin PWELL,VSS
* pin B
* pin CO
* pin S
* pin CI
* pin A
* pin NWELL,VDD
.SUBCKT FA_X1 1 2 3 8 11 12 14
* net 1 PWELL,VSS
* net 2 B
* net 3 CO
* net 8 S
* net 11 CI
* net 12 A
* net 14 NWELL,VDD
* device instance $1 r0 *1 0.385,1.0275 PMOS_VTL
M$1 17 2 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $2 r0 *1 0.575,1.0275 PMOS_VTL
M$2 4 12 17 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.765,1.0275 PMOS_VTL
M$3 15 11 4 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02265P PS=0.455U
+ PD=0.535U
* device instance $4 r0 *1 0.96,1.1025 PMOS_VTL
M$4 14 12 15 14 PMOS_VTL L=0.05U W=0.315U AS=0.02265P AD=0.02205P PS=0.535U
+ PD=0.455U
* device instance $5 r0 *1 1.15,1.1025 PMOS_VTL
M$5 15 2 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.033075P PS=0.455U
+ PD=0.84U
* device instance $6 r0 *1 0.195,0.995 PMOS_VTL
M$6 14 4 3 14 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.033075P PS=1.47U
+ PD=0.77U
* device instance $7 r0 *1 1.49,1.1525 PMOS_VTL
M$7 16 2 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $8 r0 *1 1.68,1.1525 PMOS_VTL
M$8 14 11 16 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $9 r0 *1 1.87,1.1525 PMOS_VTL
M$9 16 12 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $10 r0 *1 2.06,1.1525 PMOS_VTL
M$10 7 4 16 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.023625P PS=0.455U
+ PD=0.465U
* device instance $11 r0 *1 2.26,1.1525 PMOS_VTL
M$11 18 11 7 14 PMOS_VTL L=0.05U W=0.315U AS=0.023625P AD=0.02205P PS=0.465U
+ PD=0.455U
* device instance $12 r0 *1 2.45,1.1525 PMOS_VTL
M$12 19 2 18 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $13 r0 *1 2.64,1.1525 PMOS_VTL
M$13 19 12 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $14 r0 *1 2.83,0.995 PMOS_VTL
M$14 8 7 14 14 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U
+ PD=1.47U
* device instance $15 r0 *1 1.49,0.195 NMOS_VTL
M$15 6 2 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $16 r0 *1 1.68,0.195 NMOS_VTL
M$16 1 11 6 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $17 r0 *1 1.87,0.195 NMOS_VTL
M$17 6 12 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $18 r0 *1 2.06,0.195 NMOS_VTL
M$18 7 4 6 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.01575P PS=0.35U PD=0.36U
* device instance $19 r0 *1 2.26,0.195 NMOS_VTL
M$19 9 11 7 1 NMOS_VTL L=0.05U W=0.21U AS=0.01575P AD=0.0147P PS=0.36U PD=0.35U
* device instance $20 r0 *1 2.45,0.195 NMOS_VTL
M$20 10 2 9 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $21 r0 *1 2.64,0.195 NMOS_VTL
M$21 1 12 10 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
* device instance $22 r0 *1 2.83,0.2975 NMOS_VTL
M$22 8 7 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
* device instance $23 r0 *1 0.385,0.32 NMOS_VTL
M$23 13 2 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.021875P AD=0.0147P PS=0.555U
+ PD=0.35U
* device instance $24 r0 *1 0.575,0.32 NMOS_VTL
M$24 4 12 13 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $25 r0 *1 0.765,0.32 NMOS_VTL
M$25 5 11 4 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.015225P PS=0.35U
+ PD=0.355U
* device instance $26 r0 *1 0.96,0.32 NMOS_VTL
M$26 1 12 5 1 NMOS_VTL L=0.05U W=0.21U AS=0.015225P AD=0.0147P PS=0.355U
+ PD=0.35U
* device instance $27 r0 *1 1.15,0.32 NMOS_VTL
M$27 5 2 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.02205P PS=0.35U PD=0.63U
* device instance $28 r0 *1 0.195,0.2975 NMOS_VTL
M$28 1 4 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.021875P PS=1.04U
+ PD=0.555U
.ENDS FA_X1

* cell OAI221_X2
* pin C2
* pin C1
* pin B1
* pin B2
* pin A
* pin ZN
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT OAI221_X2 1 2 3 4 5 7 9 10
* net 1 C2
* net 2 C1
* net 3 B1
* net 4 B2
* net 5 A
* net 7 ZN
* net 9 PWELL,VSS
* net 10 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 12 1 10 10 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 7 2 12 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 11 2 7 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 10 1 11 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 7 5 10 10 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 14 3 7 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.35,0.995 PMOS_VTL
M$7 10 4 14 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.54,0.995 PMOS_VTL
M$8 13 4 10 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $9 r0 *1 1.73,0.995 PMOS_VTL
M$9 7 3 13 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $11 r0 *1 0.21,0.2975 NMOS_VTL
M$11 7 1 6 9 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $12 r0 *1 0.4,0.2975 NMOS_VTL
M$12 6 2 7 9 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $15 r0 *1 0.97,0.2975 NMOS_VTL
M$15 8 5 6 9 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $16 r0 *1 1.16,0.2975 NMOS_VTL
M$16 9 3 8 9 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $17 r0 *1 1.35,0.2975 NMOS_VTL
M$17 8 4 9 9 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
.ENDS OAI221_X2

* cell AND3_X1
* pin A1
* pin A2
* pin A3
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND3_X1 1 2 3 5 6 7
* net 1 A1
* net 2 A2
* net 3 A3
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 5 1 4 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 4 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 4 3 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 4 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.195 NMOS_VTL
M$5 8 1 4 6 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $6 r0 *1 0.36,0.195 NMOS_VTL
M$6 9 2 8 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $7 r0 *1 0.55,0.195 NMOS_VTL
M$7 6 3 9 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $8 r0 *1 0.74,0.2975 NMOS_VTL
M$8 7 4 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AND3_X1

* cell AOI22_X1
* pin B2
* pin B1
* pin A1
* pin A2
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT AOI22_X1 1 2 3 4 5 7 8
* net 1 B2
* net 2 B1
* net 3 A1
* net 4 A2
* net 5 PWELL,VSS
* net 7 NWELL,VDD
* net 8 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 7 1 6 7 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 6 2 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.565,0.995 PMOS_VTL
M$3 8 3 6 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.755,0.995 PMOS_VTL
M$4 6 4 8 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.185,0.2975 NMOS_VTL
M$5 10 1 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.375,0.2975 NMOS_VTL
M$6 8 2 10 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.565,0.2975 NMOS_VTL
M$7 9 3 8 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.755,0.2975 NMOS_VTL
M$8 5 4 9 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI22_X1

* cell OR3_X1
* pin A1
* pin A2
* pin A3
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR3_X1 1 2 3 5 6 7
* net 1 A1
* net 2 A2
* net 3 A3
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 9 1 4 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 8 2 9 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 8 3 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 4 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.195 NMOS_VTL
M$5 5 1 4 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $6 r0 *1 0.36,0.195 NMOS_VTL
M$6 4 2 5 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $7 r0 *1 0.55,0.195 NMOS_VTL
M$7 5 3 4 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $8 r0 *1 0.74,0.2975 NMOS_VTL
M$8 7 4 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OR3_X1

* cell AOI21_X1
* pin A
* pin B2
* pin B1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT AOI21_X1 1 2 3 4 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 4 PWELL,VSS
* net 6 ZN
* net 7 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 6 2 5 7 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 5 3 6 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 7 1 5 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.21,0.2975 NMOS_VTL
M$4 8 2 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.4,0.2975 NMOS_VTL
M$5 6 3 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.59,0.2975 NMOS_VTL
M$6 4 1 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI21_X1

* cell OAI21_X1
* pin B2
* pin B1
* pin A
* pin NWELL,VDD
* pin ZN
* pin PWELL,VSS
.SUBCKT OAI21_X1 1 2 3 5 6 7
* net 1 B2
* net 2 B1
* net 3 A
* net 5 NWELL,VDD
* net 6 ZN
* net 7 PWELL,VSS
* device instance $1 r0 *1 0.195,0.995 PMOS_VTL
M$1 8 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.385,0.995 PMOS_VTL
M$2 6 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.575,0.995 PMOS_VTL
M$3 5 3 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.195,0.2975 NMOS_VTL
M$4 6 1 4 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.385,0.2975 NMOS_VTL
M$5 4 2 6 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.575,0.2975 NMOS_VTL
M$6 7 3 4 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI21_X1

* cell NOR2_X1
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NOR2_X1 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 6 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 5 2 6 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.185,0.2975 NMOS_VTL
M$3 5 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $4 r0 *1 0.375,0.2975 NMOS_VTL
M$4 3 2 5 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NOR2_X1

* cell INV_X2
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT INV_X2 1 2 3 4
* net 1 A
* net 2 PWELL,VSS
* net 3 NWELL,VDD
* net 4 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 4 1 3 3 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.11025P PS=2.24U PD=2.24U
* device instance $3 r0 *1 0.185,0.2975 NMOS_VTL
M$3 4 1 2 2 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.072625P PS=1.595U
+ PD=1.595U
.ENDS INV_X2

* cell AND2_X1
* pin A1
* pin A2
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND2_X1 1 2 4 5 6
* net 1 A1
* net 2 A2
* net 4 NWELL,VDD
* net 5 PWELL,VSS
* net 6 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 3 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 3 2 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.195 NMOS_VTL
M$4 7 1 3 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $5 r0 *1 0.36,0.195 NMOS_VTL
M$5 5 2 7 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 3 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AND2_X1

* cell MUX2_X1
* pin A
* pin S
* pin B
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT MUX2_X1 1 2 3 5 6 8
* net 1 A
* net 2 S
* net 3 B
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 8 Z
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 6 2 4 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 9 1 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 7 2 9 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $4 r0 *1 0.74,1.1525 PMOS_VTL
M$4 10 4 7 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $5 r0 *1 0.93,1.1525 PMOS_VTL
M$5 10 3 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 8 7 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.17,0.195 NMOS_VTL
M$7 5 2 4 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $8 r0 *1 0.36,0.195 NMOS_VTL
M$8 12 1 5 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $9 r0 *1 0.55,0.195 NMOS_VTL
M$9 7 4 12 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $10 r0 *1 0.74,0.195 NMOS_VTL
M$10 11 2 7 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $11 r0 *1 0.93,0.195 NMOS_VTL
M$11 5 3 11 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
* device instance $12 r0 *1 1.12,0.2975 NMOS_VTL
M$12 8 7 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS MUX2_X1

* cell NAND2_X4
* pin A2
* pin A1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT NAND2_X4 1 2 4 5 6
* net 1 A2
* net 2 A1
* net 4 PWELL,VSS
* net 5 ZN
* net 6 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 5 1 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 5 2 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $9 r0 *1 0.21,0.2975 NMOS_VTL
M$9 4 1 3 4 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $13 r0 *1 0.97,0.2975 NMOS_VTL
M$13 5 2 3 4 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS NAND2_X4

* cell BUF_X4
* pin A
* pin NWELL,VDD
* pin Z
* pin PWELL,VSS
.SUBCKT BUF_X4 1 3 4 5
* net 1 A
* net 3 NWELL,VDD
* net 4 Z
* net 5 PWELL,VSS
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 2 1 3 3 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 4 2 3 3 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $7 r0 *1 0.17,0.2975 NMOS_VTL
M$7 2 1 5 5 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $9 r0 *1 0.55,0.2975 NMOS_VTL
M$9 4 2 5 5 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS BUF_X4

* cell INV_X1
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT INV_X1 1 2 3 4
* net 1 A
* net 2 PWELL,VSS
* net 3 NWELL,VDD
* net 4 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 3 3 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.06615P PS=1.47U PD=1.47U
* device instance $2 r0 *1 0.17,0.2975 NMOS_VTL
M$2 4 1 2 2 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.043575P PS=1.04U
+ PD=1.04U
.ENDS INV_X1

* cell INV_X4
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT INV_X4 1 2 3 4
* net 1 A
* net 2 PWELL,VSS
* net 3 NWELL,VDD
* net 4 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 3 3 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.19845P PS=3.78U PD=3.78U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 4 1 2 2 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.130725P PS=2.705U
+ PD=2.705U
.ENDS INV_X4
