module axi_lite_master (arready,
    arvalid,
    awready,
    awvalid,
    bready,
    bvalid,
    clk,
    read_done,
    read_req,
    rready,
    rst_n,
    rvalid,
    wready,
    write_done,
    write_req,
    wvalid,
    araddr,
    awaddr,
    bresp,
    rdata,
    read_addr,
    read_data,
    rresp,
    wdata,
    write_addr,
    write_data,
    write_strb,
    wstrb);
 input arready;
 output arvalid;
 input awready;
 output awvalid;
 output bready;
 input bvalid;
 input clk;
 output read_done;
 input read_req;
 output rready;
 input rst_n;
 input rvalid;
 input wready;
 output write_done;
 input write_req;
 output wvalid;
 output [31:0] araddr;
 output [31:0] awaddr;
 input [1:0] bresp;
 input [31:0] rdata;
 input [31:0] read_addr;
 output [31:0] read_data;
 input [1:0] rresp;
 output [31:0] wdata;
 input [31:0] write_addr;
 input [31:0] write_data;
 input [3:0] write_strb;
 output [3:0] wstrb;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire \state_r[0] ;
 wire \state_r[1] ;
 wire \state_r[2] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;

 sky130_fd_sc_hd__buf_2 _207_ (.A(\state_r[0] ),
    .X(_142_));
 sky130_fd_sc_hd__nor3_1 _208_ (.A(\state_r[2] ),
    .B(\state_r[1] ),
    .C(_142_),
    .Y(_143_));
 sky130_fd_sc_hd__and2_0 _209_ (.A(net69),
    .B(_143_),
    .X(_144_));
 sky130_fd_sc_hd__clkbuf_2 _210_ (.A(_144_),
    .X(_145_));
 sky130_fd_sc_hd__buf_4 _211_ (.A(_145_),
    .X(_146_));
 sky130_fd_sc_hd__mux2_1 _212_ (.A0(net141),
    .A1(net37),
    .S(_146_),
    .X(_000_));
 sky130_fd_sc_hd__mux2_1 _213_ (.A0(net142),
    .A1(net38),
    .S(_146_),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _214_ (.A0(net143),
    .A1(net39),
    .S(_146_),
    .X(_002_));
 sky130_fd_sc_hd__mux2_1 _215_ (.A0(net144),
    .A1(net40),
    .S(_146_),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _216_ (.A0(net145),
    .A1(net41),
    .S(_146_),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _217_ (.A0(net146),
    .A1(net42),
    .S(_146_),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _218_ (.A0(net147),
    .A1(net43),
    .S(_146_),
    .X(_006_));
 sky130_fd_sc_hd__mux2_1 _219_ (.A0(net148),
    .A1(net44),
    .S(_146_),
    .X(_007_));
 sky130_fd_sc_hd__mux2_1 _220_ (.A0(net149),
    .A1(net45),
    .S(_146_),
    .X(_008_));
 sky130_fd_sc_hd__mux2_1 _221_ (.A0(net150),
    .A1(net46),
    .S(_146_),
    .X(_009_));
 sky130_fd_sc_hd__buf_4 _222_ (.A(_145_),
    .X(_147_));
 sky130_fd_sc_hd__mux2_1 _223_ (.A0(net151),
    .A1(net47),
    .S(_147_),
    .X(_010_));
 sky130_fd_sc_hd__mux2_1 _224_ (.A0(net152),
    .A1(net48),
    .S(_147_),
    .X(_011_));
 sky130_fd_sc_hd__mux2_1 _225_ (.A0(net153),
    .A1(net49),
    .S(_147_),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _226_ (.A0(net154),
    .A1(net50),
    .S(_147_),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _227_ (.A0(net155),
    .A1(net51),
    .S(_147_),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _228_ (.A0(net156),
    .A1(net52),
    .S(_147_),
    .X(_015_));
 sky130_fd_sc_hd__mux2_1 _229_ (.A0(net157),
    .A1(net53),
    .S(_147_),
    .X(_016_));
 sky130_fd_sc_hd__mux2_1 _230_ (.A0(net158),
    .A1(net54),
    .S(_147_),
    .X(_017_));
 sky130_fd_sc_hd__mux2_1 _231_ (.A0(net159),
    .A1(net55),
    .S(_147_),
    .X(_018_));
 sky130_fd_sc_hd__mux2_1 _232_ (.A0(net160),
    .A1(net56),
    .S(_147_),
    .X(_019_));
 sky130_fd_sc_hd__buf_4 _233_ (.A(_145_),
    .X(_148_));
 sky130_fd_sc_hd__mux2_1 _234_ (.A0(net161),
    .A1(net57),
    .S(_148_),
    .X(_020_));
 sky130_fd_sc_hd__mux2_1 _235_ (.A0(net162),
    .A1(net58),
    .S(_148_),
    .X(_021_));
 sky130_fd_sc_hd__mux2_1 _236_ (.A0(net163),
    .A1(net59),
    .S(_148_),
    .X(_022_));
 sky130_fd_sc_hd__mux2_1 _237_ (.A0(net164),
    .A1(net60),
    .S(_148_),
    .X(_023_));
 sky130_fd_sc_hd__mux2_1 _238_ (.A0(net165),
    .A1(net61),
    .S(_148_),
    .X(_024_));
 sky130_fd_sc_hd__mux2_1 _239_ (.A0(net166),
    .A1(net62),
    .S(_148_),
    .X(_025_));
 sky130_fd_sc_hd__mux2_1 _240_ (.A0(net167),
    .A1(net63),
    .S(_148_),
    .X(_026_));
 sky130_fd_sc_hd__mux2_1 _241_ (.A0(net168),
    .A1(net64),
    .S(_148_),
    .X(_027_));
 sky130_fd_sc_hd__mux2_1 _242_ (.A0(net169),
    .A1(net65),
    .S(_148_),
    .X(_028_));
 sky130_fd_sc_hd__mux2_1 _243_ (.A0(net170),
    .A1(net66),
    .S(_148_),
    .X(_029_));
 sky130_fd_sc_hd__mux2_1 _244_ (.A0(net171),
    .A1(net67),
    .S(_145_),
    .X(_030_));
 sky130_fd_sc_hd__mux2_1 _245_ (.A0(net172),
    .A1(net68),
    .S(_145_),
    .X(_031_));
 sky130_fd_sc_hd__buf_2 _246_ (.A(\state_r[2] ),
    .X(_149_));
 sky130_fd_sc_hd__buf_2 _247_ (.A(_149_),
    .X(_150_));
 sky130_fd_sc_hd__buf_2 _248_ (.A(\state_r[1] ),
    .X(_151_));
 sky130_fd_sc_hd__buf_2 _249_ (.A(_142_),
    .X(_152_));
 sky130_fd_sc_hd__nor2_1 _250_ (.A(_151_),
    .B(_152_),
    .Y(_153_));
 sky130_fd_sc_hd__a21oi_1 _251_ (.A1(net69),
    .A2(_153_),
    .B1(net173),
    .Y(_154_));
 sky130_fd_sc_hd__inv_1 _252_ (.A(\state_r[1] ),
    .Y(_155_));
 sky130_fd_sc_hd__nand2b_1 _253_ (.A_N(_142_),
    .B(net2),
    .Y(_156_));
 sky130_fd_sc_hd__nand3_1 _254_ (.A(_155_),
    .B(net173),
    .C(_156_),
    .Y(_157_));
 sky130_fd_sc_hd__o21ai_0 _255_ (.A1(_150_),
    .A2(_154_),
    .B1(_157_),
    .Y(_032_));
 sky130_fd_sc_hd__and2_0 _256_ (.A(net136),
    .B(_143_),
    .X(_158_));
 sky130_fd_sc_hd__clkbuf_2 _257_ (.A(_158_),
    .X(_159_));
 sky130_fd_sc_hd__buf_6 _258_ (.A(_159_),
    .X(_160_));
 sky130_fd_sc_hd__buf_6 _259_ (.A(_160_),
    .X(_161_));
 sky130_fd_sc_hd__mux2_1 _260_ (.A0(net174),
    .A1(net72),
    .S(_161_),
    .X(_033_));
 sky130_fd_sc_hd__mux2_1 _261_ (.A0(net175),
    .A1(net73),
    .S(_161_),
    .X(_034_));
 sky130_fd_sc_hd__mux2_1 _262_ (.A0(net176),
    .A1(net74),
    .S(_161_),
    .X(_035_));
 sky130_fd_sc_hd__mux2_1 _263_ (.A0(net177),
    .A1(net75),
    .S(_161_),
    .X(_036_));
 sky130_fd_sc_hd__mux2_1 _264_ (.A0(net178),
    .A1(net76),
    .S(_161_),
    .X(_037_));
 sky130_fd_sc_hd__mux2_1 _265_ (.A0(net179),
    .A1(net77),
    .S(_161_),
    .X(_038_));
 sky130_fd_sc_hd__mux2_1 _266_ (.A0(net180),
    .A1(net78),
    .S(_161_),
    .X(_039_));
 sky130_fd_sc_hd__mux2_1 _267_ (.A0(net181),
    .A1(net79),
    .S(_161_),
    .X(_040_));
 sky130_fd_sc_hd__mux2_1 _268_ (.A0(net182),
    .A1(net80),
    .S(_161_),
    .X(_041_));
 sky130_fd_sc_hd__mux2_1 _269_ (.A0(net183),
    .A1(net81),
    .S(_161_),
    .X(_042_));
 sky130_fd_sc_hd__buf_6 _270_ (.A(_160_),
    .X(_162_));
 sky130_fd_sc_hd__mux2_1 _271_ (.A0(net184),
    .A1(net82),
    .S(_162_),
    .X(_043_));
 sky130_fd_sc_hd__mux2_1 _272_ (.A0(net185),
    .A1(net83),
    .S(_162_),
    .X(_044_));
 sky130_fd_sc_hd__mux2_1 _273_ (.A0(net186),
    .A1(net84),
    .S(_162_),
    .X(_045_));
 sky130_fd_sc_hd__mux2_1 _274_ (.A0(net187),
    .A1(net85),
    .S(_162_),
    .X(_046_));
 sky130_fd_sc_hd__mux2_1 _275_ (.A0(net188),
    .A1(net86),
    .S(_162_),
    .X(_047_));
 sky130_fd_sc_hd__mux2_1 _276_ (.A0(net189),
    .A1(net87),
    .S(_162_),
    .X(_048_));
 sky130_fd_sc_hd__mux2_1 _277_ (.A0(net190),
    .A1(net88),
    .S(_162_),
    .X(_049_));
 sky130_fd_sc_hd__mux2_1 _278_ (.A0(net191),
    .A1(net89),
    .S(_162_),
    .X(_050_));
 sky130_fd_sc_hd__mux2_1 _279_ (.A0(net192),
    .A1(net90),
    .S(_162_),
    .X(_051_));
 sky130_fd_sc_hd__mux2_1 _280_ (.A0(net193),
    .A1(net91),
    .S(_162_),
    .X(_052_));
 sky130_fd_sc_hd__buf_4 _281_ (.A(_159_),
    .X(_163_));
 sky130_fd_sc_hd__mux2_1 _282_ (.A0(net194),
    .A1(net92),
    .S(_163_),
    .X(_053_));
 sky130_fd_sc_hd__mux2_1 _283_ (.A0(net195),
    .A1(net93),
    .S(_163_),
    .X(_054_));
 sky130_fd_sc_hd__mux2_1 _284_ (.A0(net196),
    .A1(net94),
    .S(_163_),
    .X(_055_));
 sky130_fd_sc_hd__mux2_1 _285_ (.A0(net197),
    .A1(net95),
    .S(_163_),
    .X(_056_));
 sky130_fd_sc_hd__mux2_1 _286_ (.A0(net198),
    .A1(net96),
    .S(_163_),
    .X(_057_));
 sky130_fd_sc_hd__mux2_1 _287_ (.A0(net199),
    .A1(net97),
    .S(_163_),
    .X(_058_));
 sky130_fd_sc_hd__mux2_1 _288_ (.A0(net200),
    .A1(net98),
    .S(_163_),
    .X(_059_));
 sky130_fd_sc_hd__mux2_1 _289_ (.A0(net201),
    .A1(net99),
    .S(_163_),
    .X(_060_));
 sky130_fd_sc_hd__mux2_1 _290_ (.A0(net202),
    .A1(net100),
    .S(_163_),
    .X(_061_));
 sky130_fd_sc_hd__mux2_1 _291_ (.A0(net203),
    .A1(net101),
    .S(_163_),
    .X(_062_));
 sky130_fd_sc_hd__buf_4 _292_ (.A(_159_),
    .X(_164_));
 sky130_fd_sc_hd__mux2_1 _293_ (.A0(net204),
    .A1(net102),
    .S(_164_),
    .X(_063_));
 sky130_fd_sc_hd__mux2_1 _294_ (.A0(net205),
    .A1(net103),
    .S(_164_),
    .X(_064_));
 sky130_fd_sc_hd__nor2_1 _295_ (.A(_149_),
    .B(_152_),
    .Y(_165_));
 sky130_fd_sc_hd__a22oi_1 _296_ (.A1(_150_),
    .A2(net206),
    .B1(_165_),
    .B2(net136),
    .Y(_166_));
 sky130_fd_sc_hd__inv_1 _297_ (.A(net206),
    .Y(_167_));
 sky130_fd_sc_hd__a311o_1 _298_ (.A1(_155_),
    .A2(_142_),
    .A3(net3),
    .B1(_167_),
    .C1(_149_),
    .X(_168_));
 sky130_fd_sc_hd__o21ai_0 _299_ (.A1(_151_),
    .A2(_166_),
    .B1(_168_),
    .Y(_065_));
 sky130_fd_sc_hd__inv_1 _300_ (.A(net4),
    .Y(_169_));
 sky130_fd_sc_hd__a31oi_1 _301_ (.A1(_151_),
    .A2(net279),
    .A3(net71),
    .B1(net207),
    .Y(_170_));
 sky130_fd_sc_hd__nor2_1 _302_ (.A(_152_),
    .B(_170_),
    .Y(_171_));
 sky130_fd_sc_hd__a21oi_1 _303_ (.A1(net207),
    .A2(_169_),
    .B1(_171_),
    .Y(_172_));
 sky130_fd_sc_hd__o2bb2ai_1 _304_ (.A1_N(_155_),
    .A2_N(net207),
    .B1(_172_),
    .B2(_150_),
    .Y(_066_));
 sky130_fd_sc_hd__nand3_2 _305_ (.A(_142_),
    .B(net241),
    .C(net70),
    .Y(_173_));
 sky130_fd_sc_hd__nor3b_4 _306_ (.A(\state_r[1] ),
    .B(_173_),
    .C_N(\state_r[2] ),
    .Y(_174_));
 sky130_fd_sc_hd__buf_4 _307_ (.A(_174_),
    .X(_175_));
 sky130_fd_sc_hd__mux2_1 _308_ (.A0(net208),
    .A1(net5),
    .S(_175_),
    .X(_067_));
 sky130_fd_sc_hd__mux2_1 _309_ (.A0(net209),
    .A1(net6),
    .S(_175_),
    .X(_068_));
 sky130_fd_sc_hd__mux2_1 _310_ (.A0(net210),
    .A1(net7),
    .S(_175_),
    .X(_069_));
 sky130_fd_sc_hd__mux2_1 _311_ (.A0(net211),
    .A1(net8),
    .S(_175_),
    .X(_070_));
 sky130_fd_sc_hd__mux2_1 _312_ (.A0(net212),
    .A1(net9),
    .S(_175_),
    .X(_071_));
 sky130_fd_sc_hd__mux2_1 _313_ (.A0(net213),
    .A1(net10),
    .S(_175_),
    .X(_072_));
 sky130_fd_sc_hd__mux2_1 _314_ (.A0(net214),
    .A1(net11),
    .S(_175_),
    .X(_073_));
 sky130_fd_sc_hd__mux2_1 _315_ (.A0(net215),
    .A1(net12),
    .S(_175_),
    .X(_074_));
 sky130_fd_sc_hd__mux2_1 _316_ (.A0(net216),
    .A1(net13),
    .S(_175_),
    .X(_075_));
 sky130_fd_sc_hd__mux2_1 _317_ (.A0(net217),
    .A1(net14),
    .S(_175_),
    .X(_076_));
 sky130_fd_sc_hd__buf_4 _318_ (.A(_174_),
    .X(_176_));
 sky130_fd_sc_hd__mux2_1 _319_ (.A0(net218),
    .A1(net15),
    .S(_176_),
    .X(_077_));
 sky130_fd_sc_hd__mux2_1 _320_ (.A0(net219),
    .A1(net16),
    .S(_176_),
    .X(_078_));
 sky130_fd_sc_hd__mux2_1 _321_ (.A0(net220),
    .A1(net17),
    .S(_176_),
    .X(_079_));
 sky130_fd_sc_hd__mux2_1 _322_ (.A0(net221),
    .A1(net18),
    .S(_176_),
    .X(_080_));
 sky130_fd_sc_hd__mux2_1 _323_ (.A0(net222),
    .A1(net19),
    .S(_176_),
    .X(_081_));
 sky130_fd_sc_hd__mux2_1 _324_ (.A0(net223),
    .A1(net20),
    .S(_176_),
    .X(_082_));
 sky130_fd_sc_hd__mux2_1 _325_ (.A0(net224),
    .A1(net21),
    .S(_176_),
    .X(_083_));
 sky130_fd_sc_hd__mux2_1 _326_ (.A0(net225),
    .A1(net22),
    .S(_176_),
    .X(_084_));
 sky130_fd_sc_hd__mux2_1 _327_ (.A0(net226),
    .A1(net23),
    .S(_176_),
    .X(_085_));
 sky130_fd_sc_hd__mux2_1 _328_ (.A0(net227),
    .A1(net24),
    .S(_176_),
    .X(_086_));
 sky130_fd_sc_hd__buf_4 _329_ (.A(_174_),
    .X(_177_));
 sky130_fd_sc_hd__mux2_1 _330_ (.A0(net228),
    .A1(net25),
    .S(_177_),
    .X(_087_));
 sky130_fd_sc_hd__mux2_1 _331_ (.A0(net229),
    .A1(net26),
    .S(_177_),
    .X(_088_));
 sky130_fd_sc_hd__mux2_1 _332_ (.A0(net230),
    .A1(net27),
    .S(_177_),
    .X(_089_));
 sky130_fd_sc_hd__mux2_1 _333_ (.A0(net231),
    .A1(net28),
    .S(_177_),
    .X(_090_));
 sky130_fd_sc_hd__mux2_1 _334_ (.A0(net232),
    .A1(net29),
    .S(_177_),
    .X(_091_));
 sky130_fd_sc_hd__mux2_1 _335_ (.A0(net233),
    .A1(net30),
    .S(_177_),
    .X(_092_));
 sky130_fd_sc_hd__mux2_1 _336_ (.A0(net234),
    .A1(net31),
    .S(_177_),
    .X(_093_));
 sky130_fd_sc_hd__mux2_1 _337_ (.A0(net235),
    .A1(net32),
    .S(_177_),
    .X(_094_));
 sky130_fd_sc_hd__mux2_1 _338_ (.A0(net236),
    .A1(net33),
    .S(_177_),
    .X(_095_));
 sky130_fd_sc_hd__mux2_1 _339_ (.A0(net237),
    .A1(net34),
    .S(_177_),
    .X(_096_));
 sky130_fd_sc_hd__mux2_1 _340_ (.A0(net238),
    .A1(net35),
    .S(_174_),
    .X(_097_));
 sky130_fd_sc_hd__mux2_1 _341_ (.A0(net239),
    .A1(net36),
    .S(_174_),
    .X(_098_));
 sky130_fd_sc_hd__a41o_1 _342_ (.A1(_155_),
    .A2(_152_),
    .A3(net241),
    .A4(net70),
    .B1(net240),
    .X(_178_));
 sky130_fd_sc_hd__nand2_1 _343_ (.A(_150_),
    .B(_178_),
    .Y(_179_));
 sky130_fd_sc_hd__o21ai_0 _344_ (.A1(_151_),
    .A2(_152_),
    .B1(net240),
    .Y(_180_));
 sky130_fd_sc_hd__nand2_1 _345_ (.A(_179_),
    .B(_180_),
    .Y(_099_));
 sky130_fd_sc_hd__inv_1 _346_ (.A(net241),
    .Y(_181_));
 sky130_fd_sc_hd__a31oi_1 _347_ (.A1(_149_),
    .A2(net173),
    .A3(net2),
    .B1(net241),
    .Y(_182_));
 sky130_fd_sc_hd__o22a_1 _348_ (.A1(_181_),
    .A2(net70),
    .B1(_182_),
    .B2(_152_),
    .X(_183_));
 sky130_fd_sc_hd__o22ai_1 _349_ (.A1(_150_),
    .A2(_181_),
    .B1(_183_),
    .B2(_151_),
    .Y(_100_));
 sky130_fd_sc_hd__nor3_1 _350_ (.A(_149_),
    .B(_151_),
    .C(net136),
    .Y(_184_));
 sky130_fd_sc_hd__a211oi_1 _351_ (.A1(_149_),
    .A2(_151_),
    .B1(_152_),
    .C1(_184_),
    .Y(_185_));
 sky130_fd_sc_hd__a211oi_1 _352_ (.A1(net206),
    .A2(net3),
    .B1(_149_),
    .C1(\state_r[1] ),
    .Y(_186_));
 sky130_fd_sc_hd__nor2_1 _353_ (.A(net136),
    .B(net69),
    .Y(_187_));
 sky130_fd_sc_hd__a22oi_1 _354_ (.A1(_142_),
    .A2(_186_),
    .B1(_187_),
    .B2(_143_),
    .Y(_188_));
 sky130_fd_sc_hd__nand3b_1 _355_ (.A_N(_142_),
    .B(net279),
    .C(net71),
    .Y(_189_));
 sky130_fd_sc_hd__nand3_1 _356_ (.A(_142_),
    .B(net207),
    .C(net4),
    .Y(_190_));
 sky130_fd_sc_hd__nand4b_1 _357_ (.A_N(_149_),
    .B(\state_r[1] ),
    .C(_189_),
    .D(_190_),
    .Y(_191_));
 sky130_fd_sc_hd__inv_1 _358_ (.A(net173),
    .Y(_192_));
 sky130_fd_sc_hd__o2111ai_1 _359_ (.A1(_192_),
    .A2(_156_),
    .B1(_173_),
    .C1(_155_),
    .D1(_149_),
    .Y(_193_));
 sky130_fd_sc_hd__nand3_1 _360_ (.A(_188_),
    .B(_191_),
    .C(_193_),
    .Y(_194_));
 sky130_fd_sc_hd__mux2_1 _361_ (.A0(_185_),
    .A1(_152_),
    .S(_194_),
    .X(_101_));
 sky130_fd_sc_hd__xnor2_1 _362_ (.A(_151_),
    .B(_152_),
    .Y(_195_));
 sky130_fd_sc_hd__o31ai_1 _363_ (.A1(_150_),
    .A2(_194_),
    .A3(_195_),
    .B1(_191_),
    .Y(_102_));
 sky130_fd_sc_hd__inv_1 _364_ (.A(net136),
    .Y(_196_));
 sky130_fd_sc_hd__o21ai_0 _365_ (.A1(_150_),
    .A2(_196_),
    .B1(_153_),
    .Y(_197_));
 sky130_fd_sc_hd__o21ai_0 _366_ (.A1(_194_),
    .A2(_197_),
    .B1(_193_),
    .Y(_103_));
 sky130_fd_sc_hd__mux2_1 _367_ (.A0(net242),
    .A1(net104),
    .S(_164_),
    .X(_104_));
 sky130_fd_sc_hd__mux2_1 _368_ (.A0(net243),
    .A1(net105),
    .S(_164_),
    .X(_105_));
 sky130_fd_sc_hd__mux2_1 _369_ (.A0(net244),
    .A1(net106),
    .S(_164_),
    .X(_106_));
 sky130_fd_sc_hd__mux2_1 _370_ (.A0(net245),
    .A1(net107),
    .S(_164_),
    .X(_107_));
 sky130_fd_sc_hd__mux2_1 _371_ (.A0(net246),
    .A1(net108),
    .S(_164_),
    .X(_108_));
 sky130_fd_sc_hd__mux2_1 _372_ (.A0(net247),
    .A1(net109),
    .S(_164_),
    .X(_109_));
 sky130_fd_sc_hd__mux2_1 _373_ (.A0(net248),
    .A1(net110),
    .S(_164_),
    .X(_110_));
 sky130_fd_sc_hd__mux2_1 _374_ (.A0(net249),
    .A1(net111),
    .S(_164_),
    .X(_111_));
 sky130_fd_sc_hd__clkbuf_4 _375_ (.A(_159_),
    .X(_198_));
 sky130_fd_sc_hd__mux2_1 _376_ (.A0(net250),
    .A1(net112),
    .S(_198_),
    .X(_112_));
 sky130_fd_sc_hd__mux2_1 _377_ (.A0(net251),
    .A1(net113),
    .S(_198_),
    .X(_113_));
 sky130_fd_sc_hd__mux2_1 _378_ (.A0(net252),
    .A1(net114),
    .S(_198_),
    .X(_114_));
 sky130_fd_sc_hd__mux2_1 _379_ (.A0(net253),
    .A1(net115),
    .S(_198_),
    .X(_115_));
 sky130_fd_sc_hd__mux2_1 _380_ (.A0(net254),
    .A1(net116),
    .S(_198_),
    .X(_116_));
 sky130_fd_sc_hd__mux2_1 _381_ (.A0(net255),
    .A1(net117),
    .S(_198_),
    .X(_117_));
 sky130_fd_sc_hd__mux2_1 _382_ (.A0(net256),
    .A1(net118),
    .S(_198_),
    .X(_118_));
 sky130_fd_sc_hd__mux2_1 _383_ (.A0(net257),
    .A1(net119),
    .S(_198_),
    .X(_119_));
 sky130_fd_sc_hd__mux2_1 _384_ (.A0(net258),
    .A1(net120),
    .S(_198_),
    .X(_120_));
 sky130_fd_sc_hd__mux2_1 _385_ (.A0(net259),
    .A1(net121),
    .S(_198_),
    .X(_121_));
 sky130_fd_sc_hd__clkbuf_4 _386_ (.A(_159_),
    .X(_199_));
 sky130_fd_sc_hd__mux2_1 _387_ (.A0(net260),
    .A1(net122),
    .S(_199_),
    .X(_122_));
 sky130_fd_sc_hd__mux2_1 _388_ (.A0(net261),
    .A1(net123),
    .S(_199_),
    .X(_123_));
 sky130_fd_sc_hd__mux2_1 _389_ (.A0(net262),
    .A1(net124),
    .S(_199_),
    .X(_124_));
 sky130_fd_sc_hd__mux2_1 _390_ (.A0(net263),
    .A1(net125),
    .S(_199_),
    .X(_125_));
 sky130_fd_sc_hd__mux2_1 _391_ (.A0(net264),
    .A1(net126),
    .S(_199_),
    .X(_126_));
 sky130_fd_sc_hd__mux2_1 _392_ (.A0(net265),
    .A1(net127),
    .S(_199_),
    .X(_127_));
 sky130_fd_sc_hd__mux2_1 _393_ (.A0(net266),
    .A1(net128),
    .S(_199_),
    .X(_128_));
 sky130_fd_sc_hd__mux2_1 _394_ (.A0(net267),
    .A1(net129),
    .S(_199_),
    .X(_129_));
 sky130_fd_sc_hd__mux2_1 _395_ (.A0(net268),
    .A1(net130),
    .S(_199_),
    .X(_130_));
 sky130_fd_sc_hd__mux2_1 _396_ (.A0(net269),
    .A1(net131),
    .S(_199_),
    .X(_131_));
 sky130_fd_sc_hd__mux2_1 _397_ (.A0(net270),
    .A1(net132),
    .S(_160_),
    .X(_132_));
 sky130_fd_sc_hd__mux2_1 _398_ (.A0(net271),
    .A1(net133),
    .S(_160_),
    .X(_133_));
 sky130_fd_sc_hd__mux2_1 _399_ (.A0(net272),
    .A1(net134),
    .S(_160_),
    .X(_134_));
 sky130_fd_sc_hd__mux2_1 _400_ (.A0(net273),
    .A1(net135),
    .S(_160_),
    .X(_135_));
 sky130_fd_sc_hd__o21ai_0 _401_ (.A1(_150_),
    .A2(_152_),
    .B1(net274),
    .Y(_200_));
 sky130_fd_sc_hd__nor2_1 _402_ (.A(_150_),
    .B(_190_),
    .Y(_201_));
 sky130_fd_sc_hd__o21ai_0 _403_ (.A1(net274),
    .A2(_201_),
    .B1(_151_),
    .Y(_202_));
 sky130_fd_sc_hd__nand2_1 _404_ (.A(_200_),
    .B(_202_),
    .Y(_136_));
 sky130_fd_sc_hd__mux2_1 _405_ (.A0(net275),
    .A1(net137),
    .S(_160_),
    .X(_137_));
 sky130_fd_sc_hd__mux2_1 _406_ (.A0(net276),
    .A1(net138),
    .S(_160_),
    .X(_138_));
 sky130_fd_sc_hd__mux2_1 _407_ (.A0(net277),
    .A1(net139),
    .S(_160_),
    .X(_139_));
 sky130_fd_sc_hd__mux2_1 _408_ (.A0(net278),
    .A1(net140),
    .S(_160_),
    .X(_140_));
 sky130_fd_sc_hd__nor3b_1 _409_ (.A(_149_),
    .B(_186_),
    .C_N(_142_),
    .Y(_203_));
 sky130_fd_sc_hd__nor2_1 _410_ (.A(net279),
    .B(_203_),
    .Y(_204_));
 sky130_fd_sc_hd__nand2b_1 _411_ (.A_N(_142_),
    .B(net71),
    .Y(_205_));
 sky130_fd_sc_hd__nand3b_1 _412_ (.A_N(_150_),
    .B(net279),
    .C(_205_),
    .Y(_206_));
 sky130_fd_sc_hd__o21ai_0 _413_ (.A1(_151_),
    .A2(_204_),
    .B1(_206_),
    .Y(_141_));
 sky130_fd_sc_hd__dfrtp_1 \araddr[0]$_DFFE_PN0P_  (.D(_000_),
    .Q(net141),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[10]$_DFFE_PN0P_  (.D(_001_),
    .Q(net142),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[11]$_DFFE_PN0P_  (.D(_002_),
    .Q(net143),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[12]$_DFFE_PN0P_  (.D(_003_),
    .Q(net144),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[13]$_DFFE_PN0P_  (.D(_004_),
    .Q(net145),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[14]$_DFFE_PN0P_  (.D(_005_),
    .Q(net146),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[15]$_DFFE_PN0P_  (.D(_006_),
    .Q(net147),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[16]$_DFFE_PN0P_  (.D(_007_),
    .Q(net148),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[17]$_DFFE_PN0P_  (.D(_008_),
    .Q(net149),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[18]$_DFFE_PN0P_  (.D(_009_),
    .Q(net150),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[19]$_DFFE_PN0P_  (.D(_010_),
    .Q(net151),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[1]$_DFFE_PN0P_  (.D(_011_),
    .Q(net152),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[20]$_DFFE_PN0P_  (.D(_012_),
    .Q(net153),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[21]$_DFFE_PN0P_  (.D(_013_),
    .Q(net154),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[22]$_DFFE_PN0P_  (.D(_014_),
    .Q(net155),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[23]$_DFFE_PN0P_  (.D(_015_),
    .Q(net156),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[24]$_DFFE_PN0P_  (.D(_016_),
    .Q(net157),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[25]$_DFFE_PN0P_  (.D(_017_),
    .Q(net158),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[26]$_DFFE_PN0P_  (.D(_018_),
    .Q(net159),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[27]$_DFFE_PN0P_  (.D(_019_),
    .Q(net160),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[28]$_DFFE_PN0P_  (.D(_020_),
    .Q(net161),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[29]$_DFFE_PN0P_  (.D(_021_),
    .Q(net162),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[2]$_DFFE_PN0P_  (.D(_022_),
    .Q(net163),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[30]$_DFFE_PN0P_  (.D(_023_),
    .Q(net164),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[31]$_DFFE_PN0P_  (.D(_024_),
    .Q(net165),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[3]$_DFFE_PN0P_  (.D(_025_),
    .Q(net166),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[4]$_DFFE_PN0P_  (.D(_026_),
    .Q(net167),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[5]$_DFFE_PN0P_  (.D(_027_),
    .Q(net168),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[6]$_DFFE_PN0P_  (.D(_028_),
    .Q(net169),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[7]$_DFFE_PN0P_  (.D(_029_),
    .Q(net170),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[8]$_DFFE_PN0P_  (.D(_030_),
    .Q(net171),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \araddr[9]$_DFFE_PN0P_  (.D(_031_),
    .Q(net172),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \arvalid$_DFFE_PN0P_  (.D(_032_),
    .Q(net173),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[0]$_DFFE_PN0P_  (.D(_033_),
    .Q(net174),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[10]$_DFFE_PN0P_  (.D(_034_),
    .Q(net175),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[11]$_DFFE_PN0P_  (.D(_035_),
    .Q(net176),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[12]$_DFFE_PN0P_  (.D(_036_),
    .Q(net177),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[13]$_DFFE_PN0P_  (.D(_037_),
    .Q(net178),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[14]$_DFFE_PN0P_  (.D(_038_),
    .Q(net179),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[15]$_DFFE_PN0P_  (.D(_039_),
    .Q(net180),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[16]$_DFFE_PN0P_  (.D(_040_),
    .Q(net181),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[17]$_DFFE_PN0P_  (.D(_041_),
    .Q(net182),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[18]$_DFFE_PN0P_  (.D(_042_),
    .Q(net183),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[19]$_DFFE_PN0P_  (.D(_043_),
    .Q(net184),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[1]$_DFFE_PN0P_  (.D(_044_),
    .Q(net185),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[20]$_DFFE_PN0P_  (.D(_045_),
    .Q(net186),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[21]$_DFFE_PN0P_  (.D(_046_),
    .Q(net187),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[22]$_DFFE_PN0P_  (.D(_047_),
    .Q(net188),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[23]$_DFFE_PN0P_  (.D(_048_),
    .Q(net189),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[24]$_DFFE_PN0P_  (.D(_049_),
    .Q(net190),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[25]$_DFFE_PN0P_  (.D(_050_),
    .Q(net191),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[26]$_DFFE_PN0P_  (.D(_051_),
    .Q(net192),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[27]$_DFFE_PN0P_  (.D(_052_),
    .Q(net193),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[28]$_DFFE_PN0P_  (.D(_053_),
    .Q(net194),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[29]$_DFFE_PN0P_  (.D(_054_),
    .Q(net195),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[2]$_DFFE_PN0P_  (.D(_055_),
    .Q(net196),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[30]$_DFFE_PN0P_  (.D(_056_),
    .Q(net197),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[31]$_DFFE_PN0P_  (.D(_057_),
    .Q(net198),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[3]$_DFFE_PN0P_  (.D(_058_),
    .Q(net199),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[4]$_DFFE_PN0P_  (.D(_059_),
    .Q(net200),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[5]$_DFFE_PN0P_  (.D(_060_),
    .Q(net201),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[6]$_DFFE_PN0P_  (.D(_061_),
    .Q(net202),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[7]$_DFFE_PN0P_  (.D(_062_),
    .Q(net203),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[8]$_DFFE_PN0P_  (.D(_063_),
    .Q(net204),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awaddr[9]$_DFFE_PN0P_  (.D(_064_),
    .Q(net205),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \awvalid$_DFFE_PN0P_  (.D(_065_),
    .Q(net206),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \bready$_DFFE_PN0P_  (.D(_066_),
    .Q(net207),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[0]$_DFFE_PN0P_  (.D(_067_),
    .Q(net208),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[10]$_DFFE_PN0P_  (.D(_068_),
    .Q(net209),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[11]$_DFFE_PN0P_  (.D(_069_),
    .Q(net210),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[12]$_DFFE_PN0P_  (.D(_070_),
    .Q(net211),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[13]$_DFFE_PN0P_  (.D(_071_),
    .Q(net212),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[14]$_DFFE_PN0P_  (.D(_072_),
    .Q(net213),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[15]$_DFFE_PN0P_  (.D(_073_),
    .Q(net214),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[16]$_DFFE_PN0P_  (.D(_074_),
    .Q(net215),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[17]$_DFFE_PN0P_  (.D(_075_),
    .Q(net216),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[18]$_DFFE_PN0P_  (.D(_076_),
    .Q(net217),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[19]$_DFFE_PN0P_  (.D(_077_),
    .Q(net218),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[1]$_DFFE_PN0P_  (.D(_078_),
    .Q(net219),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[20]$_DFFE_PN0P_  (.D(_079_),
    .Q(net220),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[21]$_DFFE_PN0P_  (.D(_080_),
    .Q(net221),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[22]$_DFFE_PN0P_  (.D(_081_),
    .Q(net222),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[23]$_DFFE_PN0P_  (.D(_082_),
    .Q(net223),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[24]$_DFFE_PN0P_  (.D(_083_),
    .Q(net224),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[25]$_DFFE_PN0P_  (.D(_084_),
    .Q(net225),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[26]$_DFFE_PN0P_  (.D(_085_),
    .Q(net226),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[27]$_DFFE_PN0P_  (.D(_086_),
    .Q(net227),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[28]$_DFFE_PN0P_  (.D(_087_),
    .Q(net228),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[29]$_DFFE_PN0P_  (.D(_088_),
    .Q(net229),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[2]$_DFFE_PN0P_  (.D(_089_),
    .Q(net230),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[30]$_DFFE_PN0P_  (.D(_090_),
    .Q(net231),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[31]$_DFFE_PN0P_  (.D(_091_),
    .Q(net232),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[3]$_DFFE_PN0P_  (.D(_092_),
    .Q(net233),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[4]$_DFFE_PN0P_  (.D(_093_),
    .Q(net234),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[5]$_DFFE_PN0P_  (.D(_094_),
    .Q(net235),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[6]$_DFFE_PN0P_  (.D(_095_),
    .Q(net236),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[7]$_DFFE_PN0P_  (.D(_096_),
    .Q(net237),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[8]$_DFFE_PN0P_  (.D(_097_),
    .Q(net238),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[9]$_DFFE_PN0P_  (.D(_098_),
    .Q(net239),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_done_r$_DFFE_PN0P_  (.D(_099_),
    .Q(net240),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rready$_DFFE_PN0P_  (.D(_100_),
    .Q(net241),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \state_r[0]$_DFFE_PN0P_  (.D(_101_),
    .Q(\state_r[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \state_r[1]$_DFFE_PN0P_  (.D(_102_),
    .Q(\state_r[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \state_r[2]$_DFFE_PN0P_  (.D(_103_),
    .Q(\state_r[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[0]$_DFFE_PN0P_  (.D(_104_),
    .Q(net242),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[10]$_DFFE_PN0P_  (.D(_105_),
    .Q(net243),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[11]$_DFFE_PN0P_  (.D(_106_),
    .Q(net244),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[12]$_DFFE_PN0P_  (.D(_107_),
    .Q(net245),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[13]$_DFFE_PN0P_  (.D(_108_),
    .Q(net246),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[14]$_DFFE_PN0P_  (.D(_109_),
    .Q(net247),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[15]$_DFFE_PN0P_  (.D(_110_),
    .Q(net248),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[16]$_DFFE_PN0P_  (.D(_111_),
    .Q(net249),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[17]$_DFFE_PN0P_  (.D(_112_),
    .Q(net250),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[18]$_DFFE_PN0P_  (.D(_113_),
    .Q(net251),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[19]$_DFFE_PN0P_  (.D(_114_),
    .Q(net252),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[1]$_DFFE_PN0P_  (.D(_115_),
    .Q(net253),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[20]$_DFFE_PN0P_  (.D(_116_),
    .Q(net254),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[21]$_DFFE_PN0P_  (.D(_117_),
    .Q(net255),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[22]$_DFFE_PN0P_  (.D(_118_),
    .Q(net256),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[23]$_DFFE_PN0P_  (.D(_119_),
    .Q(net257),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[24]$_DFFE_PN0P_  (.D(_120_),
    .Q(net258),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[25]$_DFFE_PN0P_  (.D(_121_),
    .Q(net259),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[26]$_DFFE_PN0P_  (.D(_122_),
    .Q(net260),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[27]$_DFFE_PN0P_  (.D(_123_),
    .Q(net261),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[28]$_DFFE_PN0P_  (.D(_124_),
    .Q(net262),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[29]$_DFFE_PN0P_  (.D(_125_),
    .Q(net263),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[2]$_DFFE_PN0P_  (.D(_126_),
    .Q(net264),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[30]$_DFFE_PN0P_  (.D(_127_),
    .Q(net265),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[31]$_DFFE_PN0P_  (.D(_128_),
    .Q(net266),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[3]$_DFFE_PN0P_  (.D(_129_),
    .Q(net267),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[4]$_DFFE_PN0P_  (.D(_130_),
    .Q(net268),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[5]$_DFFE_PN0P_  (.D(_131_),
    .Q(net269),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[6]$_DFFE_PN0P_  (.D(_132_),
    .Q(net270),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[7]$_DFFE_PN0P_  (.D(_133_),
    .Q(net271),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[8]$_DFFE_PN0P_  (.D(_134_),
    .Q(net272),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wdata[9]$_DFFE_PN0P_  (.D(_135_),
    .Q(net273),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \write_done_r$_DFFE_PN0P_  (.D(_136_),
    .Q(net274),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wstrb[0]$_DFFE_PN0P_  (.D(_137_),
    .Q(net275),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wstrb[1]$_DFFE_PN0P_  (.D(_138_),
    .Q(net276),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wstrb[2]$_DFFE_PN0P_  (.D(_139_),
    .Q(net277),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wstrb[3]$_DFFE_PN0P_  (.D(_140_),
    .Q(net278),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wvalid$_DFFE_PN0P_  (.D(_141_),
    .Q(net279),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__buf_16 hold1 (.A(net280),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_132 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(arready),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(awready),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(bvalid),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(net315),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(net310),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(net336),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(net313),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(net331),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(net350),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(net380),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(net338),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(net366),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(net354),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(net292),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(net328),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(net343),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(net381),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(net295),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(net314),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(net282),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(net369),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(net323),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(net370),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(net388),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(net351),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(net359),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(net403),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(net360),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(net399),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(net404),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(net301),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(net385),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(net297),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(net290),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(net289),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(net337),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(net371),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(net361),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(net358),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(net333),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(net363),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(net412),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(net326),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(net382),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(net334),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(net393),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(net364),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(net325),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(net302),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(net340),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(net389),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(net299),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(net407),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(net368),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(net339),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(net402),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(net346),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(net375),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(net320),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(net397),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(net410),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(net394),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(net309),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(net352),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(net378),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(net392),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(net408),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(read_req),
    .X(net69));
 sky130_fd_sc_hd__dlymetal6s2s_1 input69 (.A(rvalid),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(wready),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(net305),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(net347),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(net317),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(net377),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(net391),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(net332),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(net357),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(net330),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(net285),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 input80 (.A(net311),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(net353),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(net362),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(net284),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(net308),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(net365),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(net349),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(net345),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(net329),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(net288),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input90 (.A(net306),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(net379),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 input92 (.A(net390),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(net312),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 input94 (.A(net341),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 input95 (.A(net409),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 input96 (.A(net319),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(net400),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 input98 (.A(net356),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 input99 (.A(net294),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(net304),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 input101 (.A(net303),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 input102 (.A(net286),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 input103 (.A(net367),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 input104 (.A(net291),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 input105 (.A(net374),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 input106 (.A(net321),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 input107 (.A(net316),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 input108 (.A(net335),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 input109 (.A(net287),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_1 input110 (.A(net372),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 input111 (.A(net307),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 input112 (.A(net384),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 input113 (.A(net344),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 input114 (.A(net298),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_1 input115 (.A(net348),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 input116 (.A(net376),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_1 input117 (.A(net296),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 input118 (.A(net300),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 input119 (.A(net373),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 input120 (.A(net327),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 input121 (.A(net342),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 input122 (.A(net281),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(net322),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 input124 (.A(net387),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 input125 (.A(net386),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 input126 (.A(net355),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 input127 (.A(net318),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 input128 (.A(net293),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 input129 (.A(net283),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 input130 (.A(net396),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 input131 (.A(net324),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 input132 (.A(net406),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 input133 (.A(net405),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 input134 (.A(net395),
    .X(net135));
 sky130_fd_sc_hd__dlymetal6s2s_1 input135 (.A(write_req),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 input136 (.A(net398),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 input137 (.A(net411),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 input138 (.A(net383),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_1 input139 (.A(net401),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 output140 (.A(net141),
    .X(araddr[0]));
 sky130_fd_sc_hd__clkbuf_1 output141 (.A(net142),
    .X(araddr[10]));
 sky130_fd_sc_hd__clkbuf_1 output142 (.A(net143),
    .X(araddr[11]));
 sky130_fd_sc_hd__clkbuf_1 output143 (.A(net144),
    .X(araddr[12]));
 sky130_fd_sc_hd__clkbuf_1 output144 (.A(net145),
    .X(araddr[13]));
 sky130_fd_sc_hd__clkbuf_1 output145 (.A(net146),
    .X(araddr[14]));
 sky130_fd_sc_hd__clkbuf_1 output146 (.A(net147),
    .X(araddr[15]));
 sky130_fd_sc_hd__clkbuf_1 output147 (.A(net148),
    .X(araddr[16]));
 sky130_fd_sc_hd__clkbuf_1 output148 (.A(net149),
    .X(araddr[17]));
 sky130_fd_sc_hd__clkbuf_1 output149 (.A(net150),
    .X(araddr[18]));
 sky130_fd_sc_hd__clkbuf_1 output150 (.A(net151),
    .X(araddr[19]));
 sky130_fd_sc_hd__clkbuf_1 output151 (.A(net152),
    .X(araddr[1]));
 sky130_fd_sc_hd__clkbuf_1 output152 (.A(net153),
    .X(araddr[20]));
 sky130_fd_sc_hd__clkbuf_1 output153 (.A(net154),
    .X(araddr[21]));
 sky130_fd_sc_hd__clkbuf_1 output154 (.A(net155),
    .X(araddr[22]));
 sky130_fd_sc_hd__clkbuf_1 output155 (.A(net156),
    .X(araddr[23]));
 sky130_fd_sc_hd__clkbuf_1 output156 (.A(net157),
    .X(araddr[24]));
 sky130_fd_sc_hd__clkbuf_1 output157 (.A(net158),
    .X(araddr[25]));
 sky130_fd_sc_hd__clkbuf_1 output158 (.A(net159),
    .X(araddr[26]));
 sky130_fd_sc_hd__clkbuf_1 output159 (.A(net160),
    .X(araddr[27]));
 sky130_fd_sc_hd__clkbuf_1 output160 (.A(net161),
    .X(araddr[28]));
 sky130_fd_sc_hd__clkbuf_1 output161 (.A(net162),
    .X(araddr[29]));
 sky130_fd_sc_hd__clkbuf_1 output162 (.A(net163),
    .X(araddr[2]));
 sky130_fd_sc_hd__clkbuf_1 output163 (.A(net164),
    .X(araddr[30]));
 sky130_fd_sc_hd__clkbuf_1 output164 (.A(net165),
    .X(araddr[31]));
 sky130_fd_sc_hd__clkbuf_1 output165 (.A(net166),
    .X(araddr[3]));
 sky130_fd_sc_hd__clkbuf_1 output166 (.A(net167),
    .X(araddr[4]));
 sky130_fd_sc_hd__clkbuf_1 output167 (.A(net168),
    .X(araddr[5]));
 sky130_fd_sc_hd__clkbuf_1 output168 (.A(net169),
    .X(araddr[6]));
 sky130_fd_sc_hd__clkbuf_1 output169 (.A(net170),
    .X(araddr[7]));
 sky130_fd_sc_hd__clkbuf_1 output170 (.A(net171),
    .X(araddr[8]));
 sky130_fd_sc_hd__clkbuf_1 output171 (.A(net172),
    .X(araddr[9]));
 sky130_fd_sc_hd__clkbuf_1 output172 (.A(net173),
    .X(arvalid));
 sky130_fd_sc_hd__clkbuf_1 output173 (.A(net174),
    .X(awaddr[0]));
 sky130_fd_sc_hd__clkbuf_1 output174 (.A(net175),
    .X(awaddr[10]));
 sky130_fd_sc_hd__clkbuf_1 output175 (.A(net176),
    .X(awaddr[11]));
 sky130_fd_sc_hd__clkbuf_1 output176 (.A(net177),
    .X(awaddr[12]));
 sky130_fd_sc_hd__clkbuf_1 output177 (.A(net178),
    .X(awaddr[13]));
 sky130_fd_sc_hd__clkbuf_1 output178 (.A(net179),
    .X(awaddr[14]));
 sky130_fd_sc_hd__clkbuf_1 output179 (.A(net180),
    .X(awaddr[15]));
 sky130_fd_sc_hd__clkbuf_1 output180 (.A(net181),
    .X(awaddr[16]));
 sky130_fd_sc_hd__clkbuf_1 output181 (.A(net182),
    .X(awaddr[17]));
 sky130_fd_sc_hd__clkbuf_1 output182 (.A(net183),
    .X(awaddr[18]));
 sky130_fd_sc_hd__clkbuf_1 output183 (.A(net184),
    .X(awaddr[19]));
 sky130_fd_sc_hd__clkbuf_1 output184 (.A(net185),
    .X(awaddr[1]));
 sky130_fd_sc_hd__clkbuf_1 output185 (.A(net186),
    .X(awaddr[20]));
 sky130_fd_sc_hd__clkbuf_1 output186 (.A(net187),
    .X(awaddr[21]));
 sky130_fd_sc_hd__clkbuf_1 output187 (.A(net188),
    .X(awaddr[22]));
 sky130_fd_sc_hd__clkbuf_1 output188 (.A(net189),
    .X(awaddr[23]));
 sky130_fd_sc_hd__clkbuf_1 output189 (.A(net190),
    .X(awaddr[24]));
 sky130_fd_sc_hd__clkbuf_1 output190 (.A(net191),
    .X(awaddr[25]));
 sky130_fd_sc_hd__clkbuf_1 output191 (.A(net192),
    .X(awaddr[26]));
 sky130_fd_sc_hd__clkbuf_1 output192 (.A(net193),
    .X(awaddr[27]));
 sky130_fd_sc_hd__clkbuf_1 output193 (.A(net194),
    .X(awaddr[28]));
 sky130_fd_sc_hd__clkbuf_1 output194 (.A(net195),
    .X(awaddr[29]));
 sky130_fd_sc_hd__clkbuf_1 output195 (.A(net196),
    .X(awaddr[2]));
 sky130_fd_sc_hd__clkbuf_1 output196 (.A(net197),
    .X(awaddr[30]));
 sky130_fd_sc_hd__clkbuf_1 output197 (.A(net198),
    .X(awaddr[31]));
 sky130_fd_sc_hd__clkbuf_1 output198 (.A(net199),
    .X(awaddr[3]));
 sky130_fd_sc_hd__clkbuf_1 output199 (.A(net200),
    .X(awaddr[4]));
 sky130_fd_sc_hd__clkbuf_1 output200 (.A(net201),
    .X(awaddr[5]));
 sky130_fd_sc_hd__clkbuf_1 output201 (.A(net202),
    .X(awaddr[6]));
 sky130_fd_sc_hd__clkbuf_1 output202 (.A(net203),
    .X(awaddr[7]));
 sky130_fd_sc_hd__clkbuf_1 output203 (.A(net204),
    .X(awaddr[8]));
 sky130_fd_sc_hd__clkbuf_1 output204 (.A(net205),
    .X(awaddr[9]));
 sky130_fd_sc_hd__clkbuf_1 output205 (.A(net206),
    .X(awvalid));
 sky130_fd_sc_hd__clkbuf_1 output206 (.A(net207),
    .X(bready));
 sky130_fd_sc_hd__clkbuf_1 output207 (.A(net208),
    .X(read_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output208 (.A(net209),
    .X(read_data[10]));
 sky130_fd_sc_hd__clkbuf_1 output209 (.A(net210),
    .X(read_data[11]));
 sky130_fd_sc_hd__clkbuf_1 output210 (.A(net211),
    .X(read_data[12]));
 sky130_fd_sc_hd__clkbuf_1 output211 (.A(net212),
    .X(read_data[13]));
 sky130_fd_sc_hd__clkbuf_1 output212 (.A(net213),
    .X(read_data[14]));
 sky130_fd_sc_hd__clkbuf_1 output213 (.A(net214),
    .X(read_data[15]));
 sky130_fd_sc_hd__clkbuf_1 output214 (.A(net215),
    .X(read_data[16]));
 sky130_fd_sc_hd__clkbuf_1 output215 (.A(net216),
    .X(read_data[17]));
 sky130_fd_sc_hd__clkbuf_1 output216 (.A(net217),
    .X(read_data[18]));
 sky130_fd_sc_hd__clkbuf_1 output217 (.A(net218),
    .X(read_data[19]));
 sky130_fd_sc_hd__clkbuf_1 output218 (.A(net219),
    .X(read_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output219 (.A(net220),
    .X(read_data[20]));
 sky130_fd_sc_hd__clkbuf_1 output220 (.A(net221),
    .X(read_data[21]));
 sky130_fd_sc_hd__clkbuf_1 output221 (.A(net222),
    .X(read_data[22]));
 sky130_fd_sc_hd__clkbuf_1 output222 (.A(net223),
    .X(read_data[23]));
 sky130_fd_sc_hd__clkbuf_1 output223 (.A(net224),
    .X(read_data[24]));
 sky130_fd_sc_hd__clkbuf_1 output224 (.A(net225),
    .X(read_data[25]));
 sky130_fd_sc_hd__clkbuf_1 output225 (.A(net226),
    .X(read_data[26]));
 sky130_fd_sc_hd__clkbuf_1 output226 (.A(net227),
    .X(read_data[27]));
 sky130_fd_sc_hd__clkbuf_1 output227 (.A(net228),
    .X(read_data[28]));
 sky130_fd_sc_hd__clkbuf_1 output228 (.A(net229),
    .X(read_data[29]));
 sky130_fd_sc_hd__clkbuf_1 output229 (.A(net230),
    .X(read_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output230 (.A(net231),
    .X(read_data[30]));
 sky130_fd_sc_hd__clkbuf_1 output231 (.A(net232),
    .X(read_data[31]));
 sky130_fd_sc_hd__clkbuf_1 output232 (.A(net233),
    .X(read_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output233 (.A(net234),
    .X(read_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output234 (.A(net235),
    .X(read_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output235 (.A(net236),
    .X(read_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output236 (.A(net237),
    .X(read_data[7]));
 sky130_fd_sc_hd__clkbuf_1 output237 (.A(net238),
    .X(read_data[8]));
 sky130_fd_sc_hd__clkbuf_1 output238 (.A(net239),
    .X(read_data[9]));
 sky130_fd_sc_hd__clkbuf_1 output239 (.A(net240),
    .X(read_done));
 sky130_fd_sc_hd__clkbuf_1 output240 (.A(net241),
    .X(rready));
 sky130_fd_sc_hd__clkbuf_1 output241 (.A(net242),
    .X(wdata[0]));
 sky130_fd_sc_hd__clkbuf_1 output242 (.A(net243),
    .X(wdata[10]));
 sky130_fd_sc_hd__clkbuf_1 output243 (.A(net244),
    .X(wdata[11]));
 sky130_fd_sc_hd__clkbuf_1 output244 (.A(net245),
    .X(wdata[12]));
 sky130_fd_sc_hd__clkbuf_1 output245 (.A(net246),
    .X(wdata[13]));
 sky130_fd_sc_hd__clkbuf_1 output246 (.A(net247),
    .X(wdata[14]));
 sky130_fd_sc_hd__clkbuf_1 output247 (.A(net248),
    .X(wdata[15]));
 sky130_fd_sc_hd__clkbuf_1 output248 (.A(net249),
    .X(wdata[16]));
 sky130_fd_sc_hd__clkbuf_1 output249 (.A(net250),
    .X(wdata[17]));
 sky130_fd_sc_hd__clkbuf_1 output250 (.A(net251),
    .X(wdata[18]));
 sky130_fd_sc_hd__clkbuf_1 output251 (.A(net252),
    .X(wdata[19]));
 sky130_fd_sc_hd__clkbuf_1 output252 (.A(net253),
    .X(wdata[1]));
 sky130_fd_sc_hd__clkbuf_1 output253 (.A(net254),
    .X(wdata[20]));
 sky130_fd_sc_hd__clkbuf_1 output254 (.A(net255),
    .X(wdata[21]));
 sky130_fd_sc_hd__clkbuf_1 output255 (.A(net256),
    .X(wdata[22]));
 sky130_fd_sc_hd__clkbuf_1 output256 (.A(net257),
    .X(wdata[23]));
 sky130_fd_sc_hd__clkbuf_1 output257 (.A(net258),
    .X(wdata[24]));
 sky130_fd_sc_hd__clkbuf_1 output258 (.A(net259),
    .X(wdata[25]));
 sky130_fd_sc_hd__clkbuf_1 output259 (.A(net260),
    .X(wdata[26]));
 sky130_fd_sc_hd__clkbuf_1 output260 (.A(net261),
    .X(wdata[27]));
 sky130_fd_sc_hd__clkbuf_1 output261 (.A(net262),
    .X(wdata[28]));
 sky130_fd_sc_hd__clkbuf_1 output262 (.A(net263),
    .X(wdata[29]));
 sky130_fd_sc_hd__clkbuf_1 output263 (.A(net264),
    .X(wdata[2]));
 sky130_fd_sc_hd__clkbuf_1 output264 (.A(net265),
    .X(wdata[30]));
 sky130_fd_sc_hd__clkbuf_1 output265 (.A(net266),
    .X(wdata[31]));
 sky130_fd_sc_hd__clkbuf_1 output266 (.A(net267),
    .X(wdata[3]));
 sky130_fd_sc_hd__clkbuf_1 output267 (.A(net268),
    .X(wdata[4]));
 sky130_fd_sc_hd__clkbuf_1 output268 (.A(net269),
    .X(wdata[5]));
 sky130_fd_sc_hd__clkbuf_1 output269 (.A(net270),
    .X(wdata[6]));
 sky130_fd_sc_hd__clkbuf_1 output270 (.A(net271),
    .X(wdata[7]));
 sky130_fd_sc_hd__clkbuf_1 output271 (.A(net272),
    .X(wdata[8]));
 sky130_fd_sc_hd__clkbuf_1 output272 (.A(net273),
    .X(wdata[9]));
 sky130_fd_sc_hd__clkbuf_1 output273 (.A(net274),
    .X(write_done));
 sky130_fd_sc_hd__clkbuf_1 output274 (.A(net275),
    .X(wstrb[0]));
 sky130_fd_sc_hd__clkbuf_1 output275 (.A(net276),
    .X(wstrb[1]));
 sky130_fd_sc_hd__clkbuf_1 output276 (.A(net277),
    .X(wstrb[2]));
 sky130_fd_sc_hd__clkbuf_1 output277 (.A(net278),
    .X(wstrb[3]));
 sky130_fd_sc_hd__clkbuf_1 output278 (.A(net279),
    .X(wvalid));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload0 (.A(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload1 (.A(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload2 (.A(clknet_4_2_0_clk));
 sky130_fd_sc_hd__inv_6 clkload3 (.A(clknet_4_3_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload4 (.A(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload5 (.A(clknet_4_6_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload6 (.A(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload7 (.A(clknet_4_8_0_clk));
 sky130_fd_sc_hd__inv_6 clkload8 (.A(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload9 (.A(clknet_4_11_0_clk));
 sky130_fd_sc_hd__inv_6 clkload10 (.A(clknet_4_12_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload11 (.A(clknet_4_13_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload12 (.A(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(write_data[27]),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(rdata[24]),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(write_data[4]),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(write_addr[20]),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(write_addr[17]),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(write_addr[9]),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(write_data[15]),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(write_addr[26]),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(rdata[9]),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(rdata[8]),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(write_data[10]),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(rdata[19]),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(write_data[3]),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(write_addr[6]),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(rdata[22]),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(write_data[22]),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(rdata[7]),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(write_data[1]),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(read_addr[24]),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(write_data[23]),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(rdata[5]),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(read_addr[21]),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(write_addr[8]),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(write_addr[7]),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(write_addr[0]),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(write_addr[27]),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(write_data[17]),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(write_addr[21]),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(read_addr[5]),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(rdata[10]),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(write_addr[18]),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(write_addr[2]),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(rdata[12]),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(rdata[23]),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(rdata[0]),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(write_data[13]),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(write_addr[11]),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(write_data[31]),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(write_addr[3]),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(read_addr[30]),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(write_data[12]),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(write_data[28]),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(rdata[26]),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(write_data[6]),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(read_addr[20]),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(read_addr[16]),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(write_data[25]),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(rdata[1]),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(write_addr[25]),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(write_addr[16]),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(rdata[13]),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(write_addr[14]),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(read_addr[13]),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(read_addr[18]),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(write_data[14]),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(rdata[11]),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(read_addr[0]),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(rdata[16]),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(read_addr[27]),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(read_addr[22]),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(write_addr[30]),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(write_data[26]),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(rdata[20]),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(write_data[19]),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(write_addr[24]),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(read_addr[29]),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(write_addr[10]),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(write_data[20]),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(write_addr[23]),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(rdata[14]),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(rdata[29]),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(read_addr[6]),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(write_addr[19]),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(rdata[18]),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(write_data[30]),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(write_addr[5]),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(write_addr[15]),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(read_addr[12]),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(rdata[2]),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(rdata[31]),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(read_addr[11]),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(write_addr[1]),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(read_addr[14]),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(read_addr[1]),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(write_addr[22]),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(rdata[17]),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(write_data[0]),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(read_addr[26]),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(rdata[25]),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(rdata[27]),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(read_addr[10]),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(write_data[16]),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(write_data[24]),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(write_data[11]),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(read_addr[2]),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(write_data[21]),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(write_addr[12]),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(read_addr[7]),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(write_addr[28]),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(rdata[15]),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(rdata[21]),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(read_addr[17]),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(write_strb[2]),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(write_data[18]),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(rdata[6]),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(write_data[2]),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(write_data[29]),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(rdata[28]),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(read_addr[23]),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(write_addr[29]),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(write_addr[13]),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(read_addr[8]),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(read_addr[19]),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(read_addr[4]),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(write_data[9]),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(write_data[5]),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(read_addr[31]),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(write_strb[0]),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(rdata[3]),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(write_addr[4]),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(write_strb[3]),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(read_addr[28]),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(rdata[30]),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(rdata[4]),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(write_data[8]),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(write_data[7]),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(read_addr[25]),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(read_addr[9]),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(write_addr[31]),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(read_addr[3]),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(write_strb[1]),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(read_addr[15]),
    .X(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(read_addr[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(read_addr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(rst_n));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(write_addr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(write_addr[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(write_addr[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(write_addr[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(write_addr[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(write_addr[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(write_addr[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(write_addr[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(write_addr[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(write_data[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(read_addr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(read_addr[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(write_addr[1]));
 sky130_fd_sc_hd__fill_1 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_217 ();
endmodule
