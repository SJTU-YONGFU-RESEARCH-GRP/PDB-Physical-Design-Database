module sine_cosine_generator (clk,
    enable,
    rst_n,
    valid_out,
    cosine_out,
    phase_in,
    sine_out);
 input clk;
 input enable;
 input rst_n;
 output valid_out;
 output [15:0] cosine_out;
 input [15:0] phase_in;
 output [15:0] sine_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net51;

 sky130_fd_sc_hd__clkbuf_2 _237_ (.A(net6),
    .X(_196_));
 sky130_fd_sc_hd__inv_1 _238_ (.A(_196_),
    .Y(_223_));
 sky130_fd_sc_hd__inv_1 _239_ (.A(net7),
    .Y(_224_));
 sky130_fd_sc_hd__clkbuf_4 _240_ (.A(net2),
    .X(_197_));
 sky130_fd_sc_hd__clkbuf_4 _241_ (.A(_197_),
    .X(_198_));
 sky130_fd_sc_hd__clkbuf_4 _242_ (.A(_198_),
    .X(_199_));
 sky130_fd_sc_hd__clkbuf_4 _243_ (.A(_225_),
    .X(_200_));
 sky130_fd_sc_hd__and2_0 _244_ (.A(net8),
    .B(_233_),
    .X(_201_));
 sky130_fd_sc_hd__buf_2 _245_ (.A(_201_),
    .X(_202_));
 sky130_fd_sc_hd__buf_4 _246_ (.A(phase_in[15]),
    .X(_203_));
 sky130_fd_sc_hd__inv_1 _247_ (.A(_203_),
    .Y(_204_));
 sky130_fd_sc_hd__o21a_1 _248_ (.A1(_200_),
    .A2(_202_),
    .B1(_204_),
    .X(_205_));
 sky130_fd_sc_hd__buf_2 _249_ (.A(_204_),
    .X(_206_));
 sky130_fd_sc_hd__buf_2 _250_ (.A(net8),
    .X(_207_));
 sky130_fd_sc_hd__clkbuf_4 _251_ (.A(_235_),
    .X(_208_));
 sky130_fd_sc_hd__nand2b_2 _252_ (.A_N(_207_),
    .B(_208_),
    .Y(_209_));
 sky130_fd_sc_hd__buf_2 _253_ (.A(_207_),
    .X(_210_));
 sky130_fd_sc_hd__clkbuf_4 _254_ (.A(_229_),
    .X(_211_));
 sky130_fd_sc_hd__a21oi_1 _255_ (.A1(_210_),
    .A2(_200_),
    .B1(_211_),
    .Y(_212_));
 sky130_fd_sc_hd__o21ai_0 _256_ (.A1(_206_),
    .A2(_209_),
    .B1(_212_),
    .Y(_213_));
 sky130_fd_sc_hd__nor4_1 _257_ (.A(net9),
    .B(net3),
    .C(net11),
    .D(net12),
    .Y(_214_));
 sky130_fd_sc_hd__nor4_1 _258_ (.A(net10),
    .B(net13),
    .C(net15),
    .D(net4),
    .Y(_215_));
 sky130_fd_sc_hd__nor4_2 _259_ (.A(net14),
    .B(net17),
    .C(net16),
    .D(net5),
    .Y(_216_));
 sky130_fd_sc_hd__and3_1 _260_ (.A(_214_),
    .B(_215_),
    .C(_216_),
    .X(_217_));
 sky130_fd_sc_hd__buf_2 _261_ (.A(_217_),
    .X(_218_));
 sky130_fd_sc_hd__o21ai_1 _262_ (.A1(_205_),
    .A2(_213_),
    .B1(_218_),
    .Y(_219_));
 sky130_fd_sc_hd__buf_2 _263_ (.A(_210_),
    .X(_220_));
 sky130_fd_sc_hd__nand2_1 _264_ (.A(_220_),
    .B(_196_),
    .Y(_221_));
 sky130_fd_sc_hd__o21ai_0 _265_ (.A1(_231_),
    .A2(_220_),
    .B1(_221_),
    .Y(_222_));
 sky130_fd_sc_hd__nand3_4 _266_ (.A(_214_),
    .B(_215_),
    .C(_216_),
    .Y(_022_));
 sky130_fd_sc_hd__nand4_2 _267_ (.A(net9),
    .B(net14),
    .C(net17),
    .D(net16),
    .Y(_023_));
 sky130_fd_sc_hd__nand3_1 _268_ (.A(net5),
    .B(net4),
    .C(_225_),
    .Y(_024_));
 sky130_fd_sc_hd__nand4_2 _269_ (.A(net11),
    .B(net10),
    .C(net13),
    .D(net12),
    .Y(_025_));
 sky130_fd_sc_hd__nand4b_2 _270_ (.A_N(net8),
    .B(net3),
    .C(net15),
    .D(_203_),
    .Y(_026_));
 sky130_fd_sc_hd__or4_1 _271_ (.A(_023_),
    .B(_024_),
    .C(_025_),
    .D(_026_),
    .X(_027_));
 sky130_fd_sc_hd__nand2b_1 _272_ (.A_N(net8),
    .B(_200_),
    .Y(_028_));
 sky130_fd_sc_hd__buf_2 _273_ (.A(_233_),
    .X(_029_));
 sky130_fd_sc_hd__nand2b_1 _274_ (.A_N(net8),
    .B(_203_),
    .Y(_030_));
 sky130_fd_sc_hd__a21oi_1 _275_ (.A1(_029_),
    .A2(_030_),
    .B1(_208_),
    .Y(_031_));
 sky130_fd_sc_hd__a22oi_1 _276_ (.A1(_022_),
    .A2(_027_),
    .B1(_028_),
    .B2(_031_),
    .Y(_032_));
 sky130_fd_sc_hd__a21oi_1 _277_ (.A1(_219_),
    .A2(_222_),
    .B1(_032_),
    .Y(_033_));
 sky130_fd_sc_hd__clkbuf_4 _278_ (.A(_197_),
    .X(_034_));
 sky130_fd_sc_hd__nor2_1 _279_ (.A(net18),
    .B(_034_),
    .Y(_035_));
 sky130_fd_sc_hd__a21oi_1 _280_ (.A1(_199_),
    .A2(_033_),
    .B1(_035_),
    .Y(_000_));
 sky130_fd_sc_hd__nor2_1 _281_ (.A(_211_),
    .B(_235_),
    .Y(_036_));
 sky130_fd_sc_hd__nor3_1 _282_ (.A(_204_),
    .B(_210_),
    .C(_036_),
    .Y(_037_));
 sky130_fd_sc_hd__o21ai_0 _283_ (.A1(_233_),
    .A2(_211_),
    .B1(_210_),
    .Y(_038_));
 sky130_fd_sc_hd__nor2_1 _284_ (.A(_203_),
    .B(_038_),
    .Y(_039_));
 sky130_fd_sc_hd__o21ai_1 _285_ (.A1(_037_),
    .A2(_039_),
    .B1(_218_),
    .Y(_040_));
 sky130_fd_sc_hd__a2111o_4 _286_ (.A1(_233_),
    .A2(_030_),
    .B1(_225_),
    .C1(_235_),
    .D1(_211_),
    .X(_041_));
 sky130_fd_sc_hd__nor4_4 _287_ (.A(_023_),
    .B(_024_),
    .C(_025_),
    .D(_026_),
    .Y(_042_));
 sky130_fd_sc_hd__a21oi_4 _288_ (.A1(_218_),
    .A2(_041_),
    .B1(_042_),
    .Y(_043_));
 sky130_fd_sc_hd__buf_2 _289_ (.A(_203_),
    .X(_044_));
 sky130_fd_sc_hd__buf_2 _290_ (.A(_207_),
    .X(_045_));
 sky130_fd_sc_hd__nand3_1 _291_ (.A(_044_),
    .B(_045_),
    .C(_208_),
    .Y(_046_));
 sky130_fd_sc_hd__nor2_1 _292_ (.A(_233_),
    .B(_200_),
    .Y(_047_));
 sky130_fd_sc_hd__or2_0 _293_ (.A(_203_),
    .B(_207_),
    .X(_048_));
 sky130_fd_sc_hd__or2_0 _294_ (.A(_047_),
    .B(_048_),
    .X(_049_));
 sky130_fd_sc_hd__a21oi_2 _295_ (.A1(_046_),
    .A2(_049_),
    .B1(_022_),
    .Y(_050_));
 sky130_fd_sc_hd__nor3b_1 _296_ (.A(_043_),
    .B(_050_),
    .C_N(_197_),
    .Y(_051_));
 sky130_fd_sc_hd__clkbuf_4 _297_ (.A(_203_),
    .X(_052_));
 sky130_fd_sc_hd__nand2_1 _298_ (.A(_045_),
    .B(_226_),
    .Y(_053_));
 sky130_fd_sc_hd__o21ai_0 _299_ (.A1(_045_),
    .A2(net7),
    .B1(_053_),
    .Y(_054_));
 sky130_fd_sc_hd__nand2_1 _300_ (.A(_207_),
    .B(_235_),
    .Y(_055_));
 sky130_fd_sc_hd__nand2b_1 _301_ (.A_N(_210_),
    .B(net7),
    .Y(_056_));
 sky130_fd_sc_hd__nand3_1 _302_ (.A(_052_),
    .B(_055_),
    .C(_056_),
    .Y(_057_));
 sky130_fd_sc_hd__o21ai_0 _303_ (.A1(_052_),
    .A2(_054_),
    .B1(_057_),
    .Y(_058_));
 sky130_fd_sc_hd__nor2_1 _304_ (.A(_197_),
    .B(net19),
    .Y(_059_));
 sky130_fd_sc_hd__a31oi_1 _305_ (.A1(_198_),
    .A2(_043_),
    .A3(_058_),
    .B1(_059_),
    .Y(_060_));
 sky130_fd_sc_hd__a21boi_0 _306_ (.A1(_040_),
    .A2(_051_),
    .B1_N(_060_),
    .Y(_001_));
 sky130_fd_sc_hd__buf_6 _307_ (.A(_043_),
    .X(_061_));
 sky130_fd_sc_hd__buf_2 _308_ (.A(_052_),
    .X(_062_));
 sky130_fd_sc_hd__xnor2_1 _309_ (.A(_220_),
    .B(_196_),
    .Y(_063_));
 sky130_fd_sc_hd__inv_1 _310_ (.A(_045_),
    .Y(_064_));
 sky130_fd_sc_hd__nand2_1 _311_ (.A(_064_),
    .B(_196_),
    .Y(_065_));
 sky130_fd_sc_hd__nand2_1 _312_ (.A(_045_),
    .B(_211_),
    .Y(_066_));
 sky130_fd_sc_hd__nand3_1 _313_ (.A(_062_),
    .B(_065_),
    .C(_066_),
    .Y(_067_));
 sky130_fd_sc_hd__o21ai_1 _314_ (.A1(_062_),
    .A2(_063_),
    .B1(_067_),
    .Y(_068_));
 sky130_fd_sc_hd__clkinvlp_4 _315_ (.A(_211_),
    .Y(_069_));
 sky130_fd_sc_hd__nor2_1 _316_ (.A(_210_),
    .B(_069_),
    .Y(_070_));
 sky130_fd_sc_hd__nand3_1 _317_ (.A(_052_),
    .B(_209_),
    .C(_066_),
    .Y(_071_));
 sky130_fd_sc_hd__clkbuf_4 _318_ (.A(_218_),
    .X(_072_));
 sky130_fd_sc_hd__o311a_1 _319_ (.A1(_044_),
    .A2(_202_),
    .A3(_070_),
    .B1(_071_),
    .C1(_072_),
    .X(_073_));
 sky130_fd_sc_hd__a21o_1 _320_ (.A1(_028_),
    .A2(_055_),
    .B1(_203_),
    .X(_074_));
 sky130_fd_sc_hd__nand4_2 _321_ (.A(_197_),
    .B(_218_),
    .C(_041_),
    .D(_074_),
    .Y(_075_));
 sky130_fd_sc_hd__o22ai_1 _322_ (.A1(_198_),
    .A2(net20),
    .B1(_073_),
    .B2(_075_),
    .Y(_076_));
 sky130_fd_sc_hd__a31oi_1 _323_ (.A1(_199_),
    .A2(_061_),
    .A3(_068_),
    .B1(_076_),
    .Y(_002_));
 sky130_fd_sc_hd__o211ai_1 _324_ (.A1(_029_),
    .A2(_211_),
    .B1(_044_),
    .C1(_045_),
    .Y(_077_));
 sky130_fd_sc_hd__o31a_1 _325_ (.A1(_044_),
    .A2(_210_),
    .A3(_036_),
    .B1(_077_),
    .X(_078_));
 sky130_fd_sc_hd__nand2b_1 _326_ (.A_N(_078_),
    .B(_072_),
    .Y(_079_));
 sky130_fd_sc_hd__buf_2 _327_ (.A(_197_),
    .X(_080_));
 sky130_fd_sc_hd__a21o_1 _328_ (.A1(_218_),
    .A2(_041_),
    .B1(_042_),
    .X(_081_));
 sky130_fd_sc_hd__clkbuf_4 _329_ (.A(_206_),
    .X(_082_));
 sky130_fd_sc_hd__nand2b_1 _330_ (.A_N(_227_),
    .B(_207_),
    .Y(_083_));
 sky130_fd_sc_hd__o211ai_1 _331_ (.A1(_082_),
    .A2(_083_),
    .B1(_048_),
    .C1(_198_),
    .Y(_084_));
 sky130_fd_sc_hd__o22ai_1 _332_ (.A1(_080_),
    .A2(net21),
    .B1(_081_),
    .B2(_084_),
    .Y(_085_));
 sky130_fd_sc_hd__a21oi_1 _333_ (.A1(_051_),
    .A2(_079_),
    .B1(_085_),
    .Y(_003_));
 sky130_fd_sc_hd__inv_1 _334_ (.A(net22),
    .Y(_086_));
 sky130_fd_sc_hd__nand3_1 _335_ (.A(_206_),
    .B(_209_),
    .C(_066_),
    .Y(_087_));
 sky130_fd_sc_hd__o311a_1 _336_ (.A1(_206_),
    .A2(_202_),
    .A3(_070_),
    .B1(_087_),
    .C1(_072_),
    .X(_088_));
 sky130_fd_sc_hd__nor3_1 _337_ (.A(_043_),
    .B(_050_),
    .C(_088_),
    .Y(_089_));
 sky130_fd_sc_hd__nand2_1 _338_ (.A(_064_),
    .B(_211_),
    .Y(_090_));
 sky130_fd_sc_hd__o211a_1 _339_ (.A1(_231_),
    .A2(_220_),
    .B1(_066_),
    .C1(_206_),
    .X(_091_));
 sky130_fd_sc_hd__a31oi_1 _340_ (.A1(_062_),
    .A2(_221_),
    .A3(_090_),
    .B1(_091_),
    .Y(_092_));
 sky130_fd_sc_hd__o21ai_0 _341_ (.A1(_081_),
    .A2(_092_),
    .B1(_080_),
    .Y(_093_));
 sky130_fd_sc_hd__o22ai_1 _342_ (.A1(_034_),
    .A2(_086_),
    .B1(_089_),
    .B2(_093_),
    .Y(_004_));
 sky130_fd_sc_hd__o21ai_0 _343_ (.A1(_052_),
    .A2(_083_),
    .B1(_030_),
    .Y(_094_));
 sky130_fd_sc_hd__mux2i_1 _344_ (.A0(_028_),
    .A1(_055_),
    .S(_206_),
    .Y(_095_));
 sky130_fd_sc_hd__a221oi_1 _345_ (.A1(_219_),
    .A2(_094_),
    .B1(_095_),
    .B2(_072_),
    .C1(_042_),
    .Y(_096_));
 sky130_fd_sc_hd__nor2_1 _346_ (.A(_080_),
    .B(net24),
    .Y(_097_));
 sky130_fd_sc_hd__a31oi_1 _347_ (.A1(_199_),
    .A2(_040_),
    .A3(_096_),
    .B1(_097_),
    .Y(_005_));
 sky130_fd_sc_hd__nand2_1 _348_ (.A(_064_),
    .B(_029_),
    .Y(_098_));
 sky130_fd_sc_hd__nand2_1 _349_ (.A(_220_),
    .B(_224_),
    .Y(_099_));
 sky130_fd_sc_hd__buf_2 _350_ (.A(_044_),
    .X(_100_));
 sky130_fd_sc_hd__a21o_1 _351_ (.A1(_098_),
    .A2(_099_),
    .B1(_100_),
    .X(_101_));
 sky130_fd_sc_hd__o21ai_0 _352_ (.A1(_082_),
    .A2(_226_),
    .B1(_101_),
    .Y(_102_));
 sky130_fd_sc_hd__nor2b_1 _353_ (.A(_207_),
    .B_N(_235_),
    .Y(_103_));
 sky130_fd_sc_hd__mux2i_1 _354_ (.A0(_103_),
    .A1(_202_),
    .S(_052_),
    .Y(_104_));
 sky130_fd_sc_hd__a21oi_1 _355_ (.A1(_069_),
    .A2(_104_),
    .B1(_022_),
    .Y(_105_));
 sky130_fd_sc_hd__o22ai_1 _356_ (.A1(_198_),
    .A2(net25),
    .B1(_075_),
    .B2(_105_),
    .Y(_106_));
 sky130_fd_sc_hd__a31oi_1 _357_ (.A1(_199_),
    .A2(_061_),
    .A3(_102_),
    .B1(_106_),
    .Y(_006_));
 sky130_fd_sc_hd__o21ai_0 _358_ (.A1(_220_),
    .A2(_227_),
    .B1(_100_),
    .Y(_107_));
 sky130_fd_sc_hd__nand3_1 _359_ (.A(_082_),
    .B(_028_),
    .C(_083_),
    .Y(_108_));
 sky130_fd_sc_hd__nand2_1 _360_ (.A(_107_),
    .B(_108_),
    .Y(_109_));
 sky130_fd_sc_hd__nor2b_1 _361_ (.A(_075_),
    .B_N(_040_),
    .Y(_110_));
 sky130_fd_sc_hd__nor2_1 _362_ (.A(_198_),
    .B(net32),
    .Y(_111_));
 sky130_fd_sc_hd__a311oi_1 _363_ (.A1(_080_),
    .A2(_061_),
    .A3(_109_),
    .B1(_110_),
    .C1(_111_),
    .Y(_007_));
 sky130_fd_sc_hd__nor2b_1 _364_ (.A(_210_),
    .B_N(_226_),
    .Y(_112_));
 sky130_fd_sc_hd__or2_1 _365_ (.A(_207_),
    .B(_226_),
    .X(_113_));
 sky130_fd_sc_hd__nand2_1 _366_ (.A(_045_),
    .B(net7),
    .Y(_114_));
 sky130_fd_sc_hd__nand3_1 _367_ (.A(_082_),
    .B(_113_),
    .C(_114_),
    .Y(_115_));
 sky130_fd_sc_hd__o31ai_1 _368_ (.A1(_206_),
    .A2(_202_),
    .A3(_112_),
    .B1(_115_),
    .Y(_116_));
 sky130_fd_sc_hd__nand3_1 _369_ (.A(_080_),
    .B(_061_),
    .C(_116_),
    .Y(_117_));
 sky130_fd_sc_hd__o221a_1 _370_ (.A1(_198_),
    .A2(net29),
    .B1(_075_),
    .B2(_088_),
    .C1(_117_),
    .X(_008_));
 sky130_fd_sc_hd__nor2_1 _371_ (.A(_045_),
    .B(_196_),
    .Y(_118_));
 sky130_fd_sc_hd__a211oi_1 _372_ (.A1(net7),
    .A2(_196_),
    .B1(_118_),
    .C1(_100_),
    .Y(_119_));
 sky130_fd_sc_hd__a31o_1 _373_ (.A1(_062_),
    .A2(_098_),
    .A3(_053_),
    .B1(_119_),
    .X(_120_));
 sky130_fd_sc_hd__nand4_1 _374_ (.A(_072_),
    .B(_041_),
    .C(_074_),
    .D(_078_),
    .Y(_121_));
 sky130_fd_sc_hd__mux2i_1 _375_ (.A0(net31),
    .A1(_121_),
    .S(_198_),
    .Y(_122_));
 sky130_fd_sc_hd__a31oi_1 _376_ (.A1(_199_),
    .A2(_061_),
    .A3(_120_),
    .B1(_122_),
    .Y(_009_));
 sky130_fd_sc_hd__inv_1 _377_ (.A(net23),
    .Y(_123_));
 sky130_fd_sc_hd__nor3_1 _378_ (.A(_043_),
    .B(_050_),
    .C(_073_),
    .Y(_124_));
 sky130_fd_sc_hd__a211oi_1 _379_ (.A1(_224_),
    .A2(_196_),
    .B1(_118_),
    .C1(_100_),
    .Y(_125_));
 sky130_fd_sc_hd__a31oi_1 _380_ (.A1(_062_),
    .A2(_209_),
    .A3(_114_),
    .B1(_125_),
    .Y(_126_));
 sky130_fd_sc_hd__o21ai_0 _381_ (.A1(_081_),
    .A2(_126_),
    .B1(_080_),
    .Y(_127_));
 sky130_fd_sc_hd__o22ai_1 _382_ (.A1(_034_),
    .A2(_123_),
    .B1(_124_),
    .B2(_127_),
    .Y(_010_));
 sky130_fd_sc_hd__inv_1 _383_ (.A(net34),
    .Y(_128_));
 sky130_fd_sc_hd__o21ai_1 _384_ (.A1(_231_),
    .A2(_064_),
    .B1(_065_),
    .Y(_129_));
 sky130_fd_sc_hd__o21ai_1 _385_ (.A1(_029_),
    .A2(_200_),
    .B1(_045_),
    .Y(_130_));
 sky130_fd_sc_hd__a21oi_1 _386_ (.A1(_082_),
    .A2(_029_),
    .B1(_208_),
    .Y(_131_));
 sky130_fd_sc_hd__o2111ai_1 _387_ (.A1(_211_),
    .A2(_200_),
    .B1(_072_),
    .C1(_130_),
    .D1(_131_),
    .Y(_132_));
 sky130_fd_sc_hd__o211ai_1 _388_ (.A1(_081_),
    .A2(_129_),
    .B1(_132_),
    .C1(_034_),
    .Y(_133_));
 sky130_fd_sc_hd__o21ai_0 _389_ (.A1(_034_),
    .A2(_128_),
    .B1(_133_),
    .Y(_011_));
 sky130_fd_sc_hd__o21ai_0 _390_ (.A1(_045_),
    .A2(_208_),
    .B1(_114_),
    .Y(_134_));
 sky130_fd_sc_hd__nor2_1 _391_ (.A(_100_),
    .B(_134_),
    .Y(_135_));
 sky130_fd_sc_hd__a31oi_1 _392_ (.A1(_062_),
    .A2(_099_),
    .A3(_113_),
    .B1(_135_),
    .Y(_136_));
 sky130_fd_sc_hd__nand2_1 _393_ (.A(_052_),
    .B(_211_),
    .Y(_137_));
 sky130_fd_sc_hd__nand4_1 _394_ (.A(_197_),
    .B(_072_),
    .C(_041_),
    .D(_137_),
    .Y(_138_));
 sky130_fd_sc_hd__a21oi_1 _395_ (.A1(_209_),
    .A2(_130_),
    .B1(_100_),
    .Y(_139_));
 sky130_fd_sc_hd__nor3b_1 _396_ (.A(_138_),
    .B(_139_),
    .C_N(_046_),
    .Y(_140_));
 sky130_fd_sc_hd__nor2_1 _397_ (.A(_198_),
    .B(net35),
    .Y(_141_));
 sky130_fd_sc_hd__a311oi_1 _398_ (.A1(_080_),
    .A2(_061_),
    .A3(_136_),
    .B1(_140_),
    .C1(_141_),
    .Y(_012_));
 sky130_fd_sc_hd__nand2_1 _399_ (.A(_052_),
    .B(_196_),
    .Y(_142_));
 sky130_fd_sc_hd__o21ai_1 _400_ (.A1(_208_),
    .A2(_202_),
    .B1(_052_),
    .Y(_143_));
 sky130_fd_sc_hd__and2_1 _401_ (.A(_218_),
    .B(_041_),
    .X(_144_));
 sky130_fd_sc_hd__mux2i_1 _402_ (.A0(_142_),
    .A1(_143_),
    .S(_144_),
    .Y(_145_));
 sky130_fd_sc_hd__o21ai_0 _403_ (.A1(_100_),
    .A2(_212_),
    .B1(_197_),
    .Y(_146_));
 sky130_fd_sc_hd__o32a_1 _404_ (.A1(_042_),
    .A2(_145_),
    .A3(_146_),
    .B1(net36),
    .B2(_034_),
    .X(_013_));
 sky130_fd_sc_hd__inv_1 _405_ (.A(net37),
    .Y(_147_));
 sky130_fd_sc_hd__nand2_1 _406_ (.A(_064_),
    .B(_227_),
    .Y(_148_));
 sky130_fd_sc_hd__o31ai_1 _407_ (.A1(_029_),
    .A2(_208_),
    .A3(_200_),
    .B1(_072_),
    .Y(_149_));
 sky130_fd_sc_hd__nor2_1 _408_ (.A(_029_),
    .B(_208_),
    .Y(_150_));
 sky130_fd_sc_hd__a21oi_1 _409_ (.A1(_212_),
    .A2(_150_),
    .B1(_022_),
    .Y(_151_));
 sky130_fd_sc_hd__a21oi_1 _410_ (.A1(_148_),
    .A2(_149_),
    .B1(_151_),
    .Y(_152_));
 sky130_fd_sc_hd__nand2_1 _411_ (.A(_082_),
    .B(_034_),
    .Y(_153_));
 sky130_fd_sc_hd__o22ai_1 _412_ (.A1(_034_),
    .A2(_147_),
    .B1(_152_),
    .B2(_153_),
    .Y(_014_));
 sky130_fd_sc_hd__nand2_1 _413_ (.A(_062_),
    .B(_069_),
    .Y(_154_));
 sky130_fd_sc_hd__o211ai_1 _414_ (.A1(_062_),
    .A2(_129_),
    .B1(_154_),
    .C1(_061_),
    .Y(_155_));
 sky130_fd_sc_hd__nand2_1 _415_ (.A(_220_),
    .B(_200_),
    .Y(_156_));
 sky130_fd_sc_hd__nor3_1 _416_ (.A(_044_),
    .B(_029_),
    .C(_208_),
    .Y(_157_));
 sky130_fd_sc_hd__a221o_1 _417_ (.A1(_100_),
    .A2(_069_),
    .B1(_156_),
    .B2(_157_),
    .C1(_022_),
    .X(_158_));
 sky130_fd_sc_hd__nor2_1 _418_ (.A(_080_),
    .B(net38),
    .Y(_159_));
 sky130_fd_sc_hd__a31oi_1 _419_ (.A1(_199_),
    .A2(_155_),
    .A3(_158_),
    .B1(_159_),
    .Y(_015_));
 sky130_fd_sc_hd__a21oi_1 _420_ (.A1(_036_),
    .A2(_130_),
    .B1(_082_),
    .Y(_160_));
 sky130_fd_sc_hd__a21oi_1 _421_ (.A1(_072_),
    .A2(_160_),
    .B1(_042_),
    .Y(_161_));
 sky130_fd_sc_hd__nand3b_1 _422_ (.A_N(_144_),
    .B(_148_),
    .C(_062_),
    .Y(_162_));
 sky130_fd_sc_hd__nor2_1 _423_ (.A(_080_),
    .B(net40),
    .Y(_163_));
 sky130_fd_sc_hd__a31oi_1 _424_ (.A1(_199_),
    .A2(_161_),
    .A3(_162_),
    .B1(_163_),
    .Y(_016_));
 sky130_fd_sc_hd__nor3_1 _425_ (.A(_206_),
    .B(_103_),
    .C(_202_),
    .Y(_164_));
 sky130_fd_sc_hd__nand2b_1 _426_ (.A_N(_235_),
    .B(_207_),
    .Y(_165_));
 sky130_fd_sc_hd__or3_1 _427_ (.A(_203_),
    .B(_207_),
    .C(_233_),
    .X(_166_));
 sky130_fd_sc_hd__o31ai_2 _428_ (.A1(_044_),
    .A2(_200_),
    .A3(_165_),
    .B1(_166_),
    .Y(_167_));
 sky130_fd_sc_hd__o21ai_0 _429_ (.A1(_164_),
    .A2(_167_),
    .B1(_069_),
    .Y(_168_));
 sky130_fd_sc_hd__nand2_1 _430_ (.A(_144_),
    .B(_168_),
    .Y(_169_));
 sky130_fd_sc_hd__nand2b_1 _431_ (.A_N(_202_),
    .B(_113_),
    .Y(_170_));
 sky130_fd_sc_hd__a21o_1 _432_ (.A1(_056_),
    .A2(_053_),
    .B1(_206_),
    .X(_171_));
 sky130_fd_sc_hd__o21ai_0 _433_ (.A1(_100_),
    .A2(_170_),
    .B1(_171_),
    .Y(_172_));
 sky130_fd_sc_hd__nand2_1 _434_ (.A(_061_),
    .B(_172_),
    .Y(_173_));
 sky130_fd_sc_hd__nor2_1 _435_ (.A(_080_),
    .B(net41),
    .Y(_174_));
 sky130_fd_sc_hd__a31oi_1 _436_ (.A1(_199_),
    .A2(_169_),
    .A3(_173_),
    .B1(_174_),
    .Y(_017_));
 sky130_fd_sc_hd__o21ai_0 _437_ (.A1(_164_),
    .A2(_167_),
    .B1(_137_),
    .Y(_175_));
 sky130_fd_sc_hd__o21ai_0 _438_ (.A1(_220_),
    .A2(_029_),
    .B1(_053_),
    .Y(_176_));
 sky130_fd_sc_hd__o21ai_0 _439_ (.A1(_100_),
    .A2(_176_),
    .B1(_171_),
    .Y(_177_));
 sky130_fd_sc_hd__a22oi_1 _440_ (.A1(_072_),
    .A2(_175_),
    .B1(_177_),
    .B2(_043_),
    .Y(_178_));
 sky130_fd_sc_hd__nor2_1 _441_ (.A(_034_),
    .B(net45),
    .Y(_179_));
 sky130_fd_sc_hd__a21oi_1 _442_ (.A1(_199_),
    .A2(_178_),
    .B1(_179_),
    .Y(_018_));
 sky130_fd_sc_hd__a21oi_1 _443_ (.A1(_082_),
    .A2(_170_),
    .B1(_164_),
    .Y(_180_));
 sky130_fd_sc_hd__a211oi_1 _444_ (.A1(_069_),
    .A2(_167_),
    .B1(_164_),
    .C1(_022_),
    .Y(_181_));
 sky130_fd_sc_hd__a21oi_1 _445_ (.A1(_061_),
    .A2(_180_),
    .B1(_181_),
    .Y(_182_));
 sky130_fd_sc_hd__nor2_1 _446_ (.A(_034_),
    .B(net47),
    .Y(_183_));
 sky130_fd_sc_hd__a21oi_1 _447_ (.A1(_199_),
    .A2(_182_),
    .B1(_183_),
    .Y(_019_));
 sky130_fd_sc_hd__o21ai_0 _448_ (.A1(_082_),
    .A2(_227_),
    .B1(_197_),
    .Y(_184_));
 sky130_fd_sc_hd__a31oi_1 _449_ (.A1(_082_),
    .A2(_220_),
    .A3(_200_),
    .B1(_184_),
    .Y(_185_));
 sky130_fd_sc_hd__o21ai_0 _450_ (.A1(_062_),
    .A2(_156_),
    .B1(_143_),
    .Y(_186_));
 sky130_fd_sc_hd__o22ai_1 _451_ (.A1(_198_),
    .A2(net48),
    .B1(_138_),
    .B2(_186_),
    .Y(_187_));
 sky130_fd_sc_hd__a21oi_1 _452_ (.A1(_061_),
    .A2(_185_),
    .B1(_187_),
    .Y(_020_));
 sky130_fd_sc_hd__o211ai_1 _453_ (.A1(_210_),
    .A2(_029_),
    .B1(_165_),
    .C1(_044_),
    .Y(_188_));
 sky130_fd_sc_hd__o211ai_1 _454_ (.A1(_210_),
    .A2(net7),
    .B1(_055_),
    .C1(_206_),
    .Y(_189_));
 sky130_fd_sc_hd__and3_1 _455_ (.A(_027_),
    .B(_188_),
    .C(_189_),
    .X(_190_));
 sky130_fd_sc_hd__nand2_1 _456_ (.A(_044_),
    .B(_208_),
    .Y(_191_));
 sky130_fd_sc_hd__o21ai_0 _457_ (.A1(_044_),
    .A2(_047_),
    .B1(_191_),
    .Y(_192_));
 sky130_fd_sc_hd__a21oi_1 _458_ (.A1(_069_),
    .A2(_209_),
    .B1(_052_),
    .Y(_193_));
 sky130_fd_sc_hd__a21oi_1 _459_ (.A1(_220_),
    .A2(_192_),
    .B1(_193_),
    .Y(_194_));
 sky130_fd_sc_hd__mux2i_1 _460_ (.A0(_190_),
    .A1(_194_),
    .S(_144_),
    .Y(_195_));
 sky130_fd_sc_hd__mux2_1 _461_ (.A0(net39),
    .A1(_195_),
    .S(_197_),
    .X(_021_));
 sky130_fd_sc_hd__ha_1 _462_ (.A(_223_),
    .B(_224_),
    .COUT(_225_),
    .SUM(_226_));
 sky130_fd_sc_hd__ha_1 _463_ (.A(_223_),
    .B(_224_),
    .COUT(_227_),
    .SUM(_228_));
 sky130_fd_sc_hd__ha_1 _464_ (.A(_223_),
    .B(net7),
    .COUT(_229_),
    .SUM(_230_));
 sky130_fd_sc_hd__ha_1 _465_ (.A(_223_),
    .B(net7),
    .COUT(_231_),
    .SUM(_232_));
 sky130_fd_sc_hd__ha_1 _466_ (.A(net6),
    .B(_224_),
    .COUT(_233_),
    .SUM(_234_));
 sky130_fd_sc_hd__ha_2 _467_ (.A(net6),
    .B(net7),
    .COUT(_235_),
    .SUM(_236_));
 sky130_fd_sc_hd__clkbuf_1 _468_ (.A(net32),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 _469_ (.A(net29),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 _470_ (.A(net29),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 _471_ (.A(net22),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 _472_ (.A(net23),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 _473_ (.A(net48),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 _474_ (.A(net45),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 _475_ (.A(net45),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 _476_ (.A(net38),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 _477_ (.A(net39),
    .X(net49));
 sky130_fd_sc_hd__dfrtp_1 \cosine_out[0]$_DFFE_PN0P_  (.D(_000_),
    .Q(net18),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \cosine_out[10]$_DFFE_PN0P_  (.D(_001_),
    .Q(net19),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \cosine_out[11]$_DFFE_PN0P_  (.D(_002_),
    .Q(net20),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \cosine_out[12]$_DFFE_PN0P_  (.D(_003_),
    .Q(net21),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \cosine_out[13]$_DFFE_PN0P_  (.D(_004_),
    .Q(net22),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \cosine_out[15]$_DFFE_PN0P_  (.D(_005_),
    .Q(net24),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \cosine_out[1]$_DFFE_PN0P_  (.D(_006_),
    .Q(net25),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \cosine_out[2]$_DFFE_PN0P_  (.D(_007_),
    .Q(net32),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \cosine_out[4]$_DFFE_PN0P_  (.D(_008_),
    .Q(net29),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \cosine_out[7]$_DFFE_PN0P_  (.D(_009_),
    .Q(net31),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \cosine_out[9]$_DFFE_PN0P_  (.D(_010_),
    .Q(net23),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \sine_out[0]$_DFFE_PN0P_  (.D(_011_),
    .Q(net34),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \sine_out[10]$_DFFE_PN0P_  (.D(_012_),
    .Q(net35),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \sine_out[11]$_DFFE_PN0P_  (.D(_013_),
    .Q(net36),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \sine_out[12]$_DFFE_PN0P_  (.D(_014_),
    .Q(net37),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \sine_out[13]$_DFFE_PN0P_  (.D(_015_),
    .Q(net38),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \sine_out[15]$_DFFE_PN0P_  (.D(_016_),
    .Q(net40),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \sine_out[1]$_DFFE_PN0P_  (.D(_017_),
    .Q(net41),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \sine_out[5]$_DFFE_PN0P_  (.D(_018_),
    .Q(net45),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \sine_out[7]$_DFFE_PN0P_  (.D(_019_),
    .Q(net47),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \sine_out[8]$_DFFE_PN0P_  (.D(_020_),
    .Q(net48),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \sine_out[9]$_DFFE_PN0P_  (.D(_021_),
    .Q(net39),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid_out$_DFF_PN0_  (.D(net2),
    .Q(net50),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__buf_8 hold1 (.A(net51),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_66 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(enable),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(phase_in[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(phase_in[10]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(phase_in[11]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(phase_in[12]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input6 (.A(phase_in[13]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(phase_in[14]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(phase_in[1]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(phase_in[2]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(phase_in[3]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(phase_in[4]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(phase_in[5]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(phase_in[6]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(phase_in[7]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(phase_in[8]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(phase_in[9]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net18),
    .X(cosine_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net19),
    .X(cosine_out[10]));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net20),
    .X(cosine_out[11]));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net21),
    .X(cosine_out[12]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net22),
    .X(cosine_out[13]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net23),
    .X(cosine_out[14]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net24),
    .X(cosine_out[15]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net25),
    .X(cosine_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net26),
    .X(cosine_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net27),
    .X(cosine_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net28),
    .X(cosine_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net29),
    .X(cosine_out[5]));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(net30),
    .X(cosine_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output30 (.A(net31),
    .X(cosine_out[7]));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(net32),
    .X(cosine_out[8]));
 sky130_fd_sc_hd__clkbuf_1 output32 (.A(net33),
    .X(cosine_out[9]));
 sky130_fd_sc_hd__clkbuf_1 output33 (.A(net34),
    .X(sine_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output34 (.A(net35),
    .X(sine_out[10]));
 sky130_fd_sc_hd__clkbuf_1 output35 (.A(net36),
    .X(sine_out[11]));
 sky130_fd_sc_hd__clkbuf_1 output36 (.A(net37),
    .X(sine_out[12]));
 sky130_fd_sc_hd__clkbuf_1 output37 (.A(net38),
    .X(sine_out[13]));
 sky130_fd_sc_hd__clkbuf_1 output38 (.A(net39),
    .X(sine_out[14]));
 sky130_fd_sc_hd__clkbuf_1 output39 (.A(net40),
    .X(sine_out[15]));
 sky130_fd_sc_hd__clkbuf_1 output40 (.A(net41),
    .X(sine_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output41 (.A(net42),
    .X(sine_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output42 (.A(net43),
    .X(sine_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output43 (.A(net44),
    .X(sine_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output44 (.A(net45),
    .X(sine_out[5]));
 sky130_fd_sc_hd__clkbuf_1 output45 (.A(net46),
    .X(sine_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output46 (.A(net47),
    .X(sine_out[7]));
 sky130_fd_sc_hd__clkbuf_1 output47 (.A(net48),
    .X(sine_out[8]));
 sky130_fd_sc_hd__clkbuf_1 output48 (.A(net49),
    .X(sine_out[9]));
 sky130_fd_sc_hd__clkbuf_1 output49 (.A(net50),
    .X(valid_out));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkinv_2 clkload0 (.A(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net51));
 sky130_fd_sc_hd__fill_4 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_54 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_62 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_143 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_53 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_66 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_102 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_13 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_64 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_102 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_81 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_60 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_90 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_42 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_94 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_153 ();
endmodule
