module shadow_register (clk,
    main_load_en,
    rst_n,
    shadow_capture_en,
    shadow_load_en,
    use_shadow_out,
    main_data_in,
    main_data_out,
    shadow_data_in,
    shadow_data_out);
 input clk;
 input main_load_en;
 input rst_n;
 input shadow_capture_en;
 input shadow_load_en;
 input use_shadow_out;
 input [31:0] main_data_in;
 output [31:0] main_data_out;
 input [31:0] shadow_data_in;
 output [31:0] shadow_data_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire \main_reg[0] ;
 wire \main_reg[10] ;
 wire \main_reg[11] ;
 wire \main_reg[12] ;
 wire \main_reg[13] ;
 wire \main_reg[14] ;
 wire \main_reg[15] ;
 wire \main_reg[16] ;
 wire \main_reg[17] ;
 wire \main_reg[18] ;
 wire \main_reg[19] ;
 wire \main_reg[1] ;
 wire \main_reg[20] ;
 wire \main_reg[21] ;
 wire \main_reg[22] ;
 wire \main_reg[23] ;
 wire \main_reg[24] ;
 wire \main_reg[25] ;
 wire \main_reg[26] ;
 wire \main_reg[27] ;
 wire \main_reg[28] ;
 wire \main_reg[29] ;
 wire \main_reg[2] ;
 wire \main_reg[30] ;
 wire \main_reg[31] ;
 wire \main_reg[3] ;
 wire \main_reg[4] ;
 wire \main_reg[5] ;
 wire \main_reg[6] ;
 wire \main_reg[7] ;
 wire \main_reg[8] ;
 wire \main_reg[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net134;

 gf180mcu_fd_sc_mcu9t5v0__buf_4 _108_ (.I(net34),
    .Z(_064_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _109_ (.I0(\main_reg[0] ),
    .I1(net2),
    .S(_064_),
    .Z(_000_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _110_ (.I0(\main_reg[10] ),
    .I1(net3),
    .S(_064_),
    .Z(_001_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _111_ (.I0(\main_reg[11] ),
    .I1(net4),
    .S(_064_),
    .Z(_002_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _112_ (.I0(\main_reg[12] ),
    .I1(net5),
    .S(_064_),
    .Z(_003_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _113_ (.I0(\main_reg[13] ),
    .I1(net6),
    .S(_064_),
    .Z(_004_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _114_ (.I0(\main_reg[14] ),
    .I1(net7),
    .S(_064_),
    .Z(_005_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _115_ (.I0(\main_reg[15] ),
    .I1(net8),
    .S(_064_),
    .Z(_006_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _116_ (.I0(\main_reg[16] ),
    .I1(net9),
    .S(_064_),
    .Z(_007_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _117_ (.I0(\main_reg[17] ),
    .I1(net10),
    .S(_064_),
    .Z(_008_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _118_ (.I0(\main_reg[18] ),
    .I1(net11),
    .S(_064_),
    .Z(_009_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _119_ (.I(net34),
    .Z(_065_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _120_ (.I0(\main_reg[19] ),
    .I1(net12),
    .S(_065_),
    .Z(_010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _121_ (.I0(\main_reg[1] ),
    .I1(net13),
    .S(_065_),
    .Z(_011_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _122_ (.I0(\main_reg[20] ),
    .I1(net14),
    .S(_065_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _123_ (.I0(\main_reg[21] ),
    .I1(net15),
    .S(_065_),
    .Z(_013_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _124_ (.I0(\main_reg[22] ),
    .I1(net16),
    .S(_065_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _125_ (.I0(\main_reg[23] ),
    .I1(net17),
    .S(_065_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _126_ (.I0(\main_reg[24] ),
    .I1(net18),
    .S(_065_),
    .Z(_016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _127_ (.I0(\main_reg[25] ),
    .I1(net19),
    .S(_065_),
    .Z(_017_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _128_ (.I0(\main_reg[26] ),
    .I1(net20),
    .S(_065_),
    .Z(_018_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _129_ (.I0(\main_reg[27] ),
    .I1(net21),
    .S(_065_),
    .Z(_019_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _130_ (.I(net34),
    .Z(_066_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _131_ (.I0(\main_reg[28] ),
    .I1(net22),
    .S(_066_),
    .Z(_020_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _132_ (.I0(\main_reg[29] ),
    .I1(net23),
    .S(_066_),
    .Z(_021_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _133_ (.I0(\main_reg[2] ),
    .I1(net24),
    .S(_066_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _134_ (.I0(\main_reg[30] ),
    .I1(net25),
    .S(_066_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _135_ (.I0(\main_reg[31] ),
    .I1(net26),
    .S(_066_),
    .Z(_024_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _136_ (.I0(\main_reg[3] ),
    .I1(net27),
    .S(_066_),
    .Z(_025_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _137_ (.I0(\main_reg[4] ),
    .I1(net28),
    .S(_066_),
    .Z(_026_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _138_ (.I0(\main_reg[5] ),
    .I1(net29),
    .S(_066_),
    .Z(_027_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _139_ (.I0(\main_reg[6] ),
    .I1(net30),
    .S(_066_),
    .Z(_028_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _140_ (.I0(\main_reg[7] ),
    .I1(net31),
    .S(_066_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _141_ (.I0(\main_reg[8] ),
    .I1(net32),
    .S(net34),
    .Z(_030_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _142_ (.I0(\main_reg[9] ),
    .I1(net33),
    .S(net34),
    .Z(_031_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _143_ (.I(net68),
    .Z(_067_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _144_ (.I0(net102),
    .I1(net36),
    .S(_067_),
    .Z(_068_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _145_ (.I(net35),
    .Z(_069_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _146_ (.I0(_068_),
    .I1(\main_reg[0] ),
    .S(_069_),
    .Z(_032_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _147_ (.I0(net103),
    .I1(net37),
    .S(_067_),
    .Z(_070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _148_ (.I0(_070_),
    .I1(\main_reg[10] ),
    .S(_069_),
    .Z(_033_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _149_ (.I0(net104),
    .I1(net38),
    .S(_067_),
    .Z(_071_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _150_ (.I0(_071_),
    .I1(\main_reg[11] ),
    .S(_069_),
    .Z(_034_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _151_ (.I0(net105),
    .I1(net39),
    .S(_067_),
    .Z(_072_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _152_ (.I0(_072_),
    .I1(\main_reg[12] ),
    .S(_069_),
    .Z(_035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _153_ (.I0(net106),
    .I1(net40),
    .S(_067_),
    .Z(_073_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _154_ (.I0(_073_),
    .I1(\main_reg[13] ),
    .S(_069_),
    .Z(_036_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _155_ (.I0(net107),
    .I1(net41),
    .S(_067_),
    .Z(_074_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _156_ (.I0(_074_),
    .I1(\main_reg[14] ),
    .S(_069_),
    .Z(_037_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _157_ (.I0(net108),
    .I1(net42),
    .S(_067_),
    .Z(_075_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _158_ (.I0(_075_),
    .I1(\main_reg[15] ),
    .S(_069_),
    .Z(_038_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _159_ (.I0(net109),
    .I1(net43),
    .S(_067_),
    .Z(_076_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _160_ (.I0(_076_),
    .I1(\main_reg[16] ),
    .S(_069_),
    .Z(_039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _161_ (.I0(net110),
    .I1(net44),
    .S(_067_),
    .Z(_077_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _162_ (.I0(_077_),
    .I1(\main_reg[17] ),
    .S(_069_),
    .Z(_040_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _163_ (.I0(net111),
    .I1(net45),
    .S(_067_),
    .Z(_078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _164_ (.I0(_078_),
    .I1(\main_reg[18] ),
    .S(_069_),
    .Z(_041_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _165_ (.I(net68),
    .Z(_079_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _166_ (.I0(net112),
    .I1(net46),
    .S(_079_),
    .Z(_080_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _167_ (.I(net35),
    .Z(_081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _168_ (.I0(_080_),
    .I1(\main_reg[19] ),
    .S(_081_),
    .Z(_042_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _169_ (.I0(net113),
    .I1(net47),
    .S(_079_),
    .Z(_082_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _170_ (.I0(_082_),
    .I1(\main_reg[1] ),
    .S(_081_),
    .Z(_043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _171_ (.I0(net114),
    .I1(net48),
    .S(_079_),
    .Z(_083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _172_ (.I0(_083_),
    .I1(\main_reg[20] ),
    .S(_081_),
    .Z(_044_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _173_ (.I0(net115),
    .I1(net49),
    .S(_079_),
    .Z(_084_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _174_ (.I0(_084_),
    .I1(\main_reg[21] ),
    .S(_081_),
    .Z(_045_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _175_ (.I0(net116),
    .I1(net50),
    .S(_079_),
    .Z(_085_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _176_ (.I0(_085_),
    .I1(\main_reg[22] ),
    .S(_081_),
    .Z(_046_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _177_ (.I0(net117),
    .I1(net51),
    .S(_079_),
    .Z(_086_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _178_ (.I0(_086_),
    .I1(\main_reg[23] ),
    .S(_081_),
    .Z(_047_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _179_ (.I0(net118),
    .I1(net52),
    .S(_079_),
    .Z(_087_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _180_ (.I0(_087_),
    .I1(\main_reg[24] ),
    .S(_081_),
    .Z(_048_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _181_ (.I0(net119),
    .I1(net53),
    .S(_079_),
    .Z(_088_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _182_ (.I0(_088_),
    .I1(\main_reg[25] ),
    .S(_081_),
    .Z(_049_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _183_ (.I0(net120),
    .I1(net54),
    .S(_079_),
    .Z(_089_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _184_ (.I0(_089_),
    .I1(\main_reg[26] ),
    .S(_081_),
    .Z(_050_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _185_ (.I0(net121),
    .I1(net55),
    .S(_079_),
    .Z(_090_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _186_ (.I0(_090_),
    .I1(\main_reg[27] ),
    .S(_081_),
    .Z(_051_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _187_ (.I(net68),
    .Z(_091_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _188_ (.I0(net122),
    .I1(net56),
    .S(_091_),
    .Z(_092_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _189_ (.I(net35),
    .Z(_093_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _190_ (.I0(_092_),
    .I1(\main_reg[28] ),
    .S(_093_),
    .Z(_052_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _191_ (.I0(net123),
    .I1(net57),
    .S(_091_),
    .Z(_094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _192_ (.I0(_094_),
    .I1(\main_reg[29] ),
    .S(_093_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _193_ (.I0(net124),
    .I1(net58),
    .S(_091_),
    .Z(_095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _194_ (.I0(_095_),
    .I1(\main_reg[2] ),
    .S(_093_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _195_ (.I0(net125),
    .I1(net59),
    .S(_091_),
    .Z(_096_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _196_ (.I0(_096_),
    .I1(\main_reg[30] ),
    .S(_093_),
    .Z(_055_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _197_ (.I0(net126),
    .I1(net60),
    .S(_091_),
    .Z(_097_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _198_ (.I0(_097_),
    .I1(\main_reg[31] ),
    .S(_093_),
    .Z(_056_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _199_ (.I0(net127),
    .I1(net61),
    .S(_091_),
    .Z(_098_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _200_ (.I0(_098_),
    .I1(\main_reg[3] ),
    .S(_093_),
    .Z(_057_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _201_ (.I0(net128),
    .I1(net62),
    .S(_091_),
    .Z(_099_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _202_ (.I0(_099_),
    .I1(\main_reg[4] ),
    .S(_093_),
    .Z(_058_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _203_ (.I0(net129),
    .I1(net63),
    .S(_091_),
    .Z(_100_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _204_ (.I0(_100_),
    .I1(\main_reg[5] ),
    .S(_093_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _205_ (.I0(net130),
    .I1(net64),
    .S(_091_),
    .Z(_101_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _206_ (.I0(_101_),
    .I1(\main_reg[6] ),
    .S(_093_),
    .Z(_060_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _207_ (.I0(net131),
    .I1(net65),
    .S(_091_),
    .Z(_102_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _208_ (.I0(_102_),
    .I1(\main_reg[7] ),
    .S(_093_),
    .Z(_061_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _209_ (.I0(net132),
    .I1(net66),
    .S(net68),
    .Z(_103_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _210_ (.I0(_103_),
    .I1(\main_reg[8] ),
    .S(net35),
    .Z(_062_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _211_ (.I0(net133),
    .I1(net67),
    .S(net68),
    .Z(_104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _212_ (.I0(_104_),
    .I1(\main_reg[9] ),
    .S(net35),
    .Z(_063_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _213_ (.I(net69),
    .Z(_105_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _214_ (.I0(\main_reg[0] ),
    .I1(net102),
    .S(_105_),
    .Z(net70));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _215_ (.I0(\main_reg[10] ),
    .I1(net103),
    .S(_105_),
    .Z(net71));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _216_ (.I0(\main_reg[11] ),
    .I1(net104),
    .S(_105_),
    .Z(net72));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _217_ (.I0(\main_reg[12] ),
    .I1(net105),
    .S(_105_),
    .Z(net73));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _218_ (.I0(\main_reg[13] ),
    .I1(net106),
    .S(_105_),
    .Z(net74));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _219_ (.I0(\main_reg[14] ),
    .I1(net107),
    .S(_105_),
    .Z(net75));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _220_ (.I0(\main_reg[15] ),
    .I1(net108),
    .S(_105_),
    .Z(net76));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _221_ (.I0(\main_reg[16] ),
    .I1(net109),
    .S(_105_),
    .Z(net77));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _222_ (.I0(\main_reg[17] ),
    .I1(net110),
    .S(_105_),
    .Z(net78));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _223_ (.I0(\main_reg[18] ),
    .I1(net111),
    .S(_105_),
    .Z(net79));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _224_ (.I(net69),
    .Z(_106_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _225_ (.I0(\main_reg[19] ),
    .I1(net112),
    .S(_106_),
    .Z(net80));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _226_ (.I0(\main_reg[1] ),
    .I1(net113),
    .S(_106_),
    .Z(net81));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _227_ (.I0(\main_reg[20] ),
    .I1(net114),
    .S(_106_),
    .Z(net82));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _228_ (.I0(\main_reg[21] ),
    .I1(net115),
    .S(_106_),
    .Z(net83));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _229_ (.I0(\main_reg[22] ),
    .I1(net116),
    .S(_106_),
    .Z(net84));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _230_ (.I0(\main_reg[23] ),
    .I1(net117),
    .S(_106_),
    .Z(net85));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _231_ (.I0(\main_reg[24] ),
    .I1(net118),
    .S(_106_),
    .Z(net86));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _232_ (.I0(\main_reg[25] ),
    .I1(net119),
    .S(_106_),
    .Z(net87));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _233_ (.I0(\main_reg[26] ),
    .I1(net120),
    .S(_106_),
    .Z(net88));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _234_ (.I0(\main_reg[27] ),
    .I1(net121),
    .S(_106_),
    .Z(net89));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _235_ (.I(net69),
    .Z(_107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _236_ (.I0(\main_reg[28] ),
    .I1(net122),
    .S(_107_),
    .Z(net90));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _237_ (.I0(\main_reg[29] ),
    .I1(net123),
    .S(_107_),
    .Z(net91));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _238_ (.I0(\main_reg[2] ),
    .I1(net124),
    .S(_107_),
    .Z(net92));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _239_ (.I0(\main_reg[30] ),
    .I1(net125),
    .S(_107_),
    .Z(net93));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _240_ (.I0(\main_reg[31] ),
    .I1(net126),
    .S(_107_),
    .Z(net94));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _241_ (.I0(\main_reg[3] ),
    .I1(net127),
    .S(_107_),
    .Z(net95));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _242_ (.I0(\main_reg[4] ),
    .I1(net128),
    .S(_107_),
    .Z(net96));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _243_ (.I0(\main_reg[5] ),
    .I1(net129),
    .S(_107_),
    .Z(net97));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _244_ (.I0(\main_reg[6] ),
    .I1(net130),
    .S(_107_),
    .Z(net98));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _245_ (.I0(\main_reg[7] ),
    .I1(net131),
    .S(_107_),
    .Z(net99));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _246_ (.I0(\main_reg[8] ),
    .I1(net132),
    .S(net69),
    .Z(net100));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _247_ (.I0(\main_reg[9] ),
    .I1(net133),
    .S(net69),
    .Z(net101));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[0]$_DFFE_PN0P_  (.D(_000_),
    .RN(net1),
    .CLK(clknet_3_2__leaf_clk),
    .Q(\main_reg[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[10]$_DFFE_PN0P_  (.D(_001_),
    .RN(net1),
    .CLK(clknet_3_3__leaf_clk),
    .Q(\main_reg[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[11]$_DFFE_PN0P_  (.D(_002_),
    .RN(net1),
    .CLK(clknet_3_2__leaf_clk),
    .Q(\main_reg[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[12]$_DFFE_PN0P_  (.D(_003_),
    .RN(net1),
    .CLK(clknet_3_3__leaf_clk),
    .Q(\main_reg[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[13]$_DFFE_PN0P_  (.D(_004_),
    .RN(net1),
    .CLK(clknet_3_3__leaf_clk),
    .Q(\main_reg[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[14]$_DFFE_PN0P_  (.D(_005_),
    .RN(net1),
    .CLK(clknet_3_2__leaf_clk),
    .Q(\main_reg[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[15]$_DFFE_PN0P_  (.D(_006_),
    .RN(net1),
    .CLK(clknet_3_3__leaf_clk),
    .Q(\main_reg[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[16]$_DFFE_PN0P_  (.D(_007_),
    .RN(net1),
    .CLK(clknet_3_6__leaf_clk),
    .Q(\main_reg[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[17]$_DFFE_PN0P_  (.D(_008_),
    .RN(net1),
    .CLK(clknet_3_3__leaf_clk),
    .Q(\main_reg[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[18]$_DFFE_PN0P_  (.D(_009_),
    .RN(net1),
    .CLK(clknet_3_2__leaf_clk),
    .Q(\main_reg[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[19]$_DFFE_PN0P_  (.D(_010_),
    .RN(net1),
    .CLK(clknet_3_1__leaf_clk),
    .Q(\main_reg[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[1]$_DFFE_PN0P_  (.D(_011_),
    .RN(net1),
    .CLK(clknet_3_3__leaf_clk),
    .Q(\main_reg[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[20]$_DFFE_PN0P_  (.D(_012_),
    .RN(net1),
    .CLK(clknet_3_0__leaf_clk),
    .Q(\main_reg[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[21]$_DFFE_PN0P_  (.D(_013_),
    .RN(net1),
    .CLK(clknet_3_0__leaf_clk),
    .Q(\main_reg[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[22]$_DFFE_PN0P_  (.D(_014_),
    .RN(net1),
    .CLK(clknet_3_1__leaf_clk),
    .Q(\main_reg[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[23]$_DFFE_PN0P_  (.D(_015_),
    .RN(net1),
    .CLK(clknet_3_1__leaf_clk),
    .Q(\main_reg[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[24]$_DFFE_PN0P_  (.D(_016_),
    .RN(net1),
    .CLK(clknet_3_1__leaf_clk),
    .Q(\main_reg[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[25]$_DFFE_PN0P_  (.D(_017_),
    .RN(net1),
    .CLK(clknet_3_0__leaf_clk),
    .Q(\main_reg[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[26]$_DFFE_PN0P_  (.D(_018_),
    .RN(net1),
    .CLK(clknet_3_0__leaf_clk),
    .Q(\main_reg[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[27]$_DFFE_PN0P_  (.D(_019_),
    .RN(net1),
    .CLK(clknet_3_3__leaf_clk),
    .Q(\main_reg[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[28]$_DFFE_PN0P_  (.D(_020_),
    .RN(net1),
    .CLK(clknet_3_7__leaf_clk),
    .Q(\main_reg[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[29]$_DFFE_PN0P_  (.D(_021_),
    .RN(net1),
    .CLK(clknet_3_5__leaf_clk),
    .Q(\main_reg[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[2]$_DFFE_PN0P_  (.D(_022_),
    .RN(net1),
    .CLK(clknet_3_4__leaf_clk),
    .Q(\main_reg[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[30]$_DFFE_PN0P_  (.D(_023_),
    .RN(net1),
    .CLK(clknet_3_6__leaf_clk),
    .Q(\main_reg[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[31]$_DFFE_PN0P_  (.D(_024_),
    .RN(net1),
    .CLK(clknet_3_4__leaf_clk),
    .Q(\main_reg[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[3]$_DFFE_PN0P_  (.D(_025_),
    .RN(net1),
    .CLK(clknet_3_6__leaf_clk),
    .Q(\main_reg[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[4]$_DFFE_PN0P_  (.D(_026_),
    .RN(net1),
    .CLK(clknet_3_7__leaf_clk),
    .Q(\main_reg[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[5]$_DFFE_PN0P_  (.D(_027_),
    .RN(net1),
    .CLK(clknet_3_5__leaf_clk),
    .Q(\main_reg[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[6]$_DFFE_PN0P_  (.D(_028_),
    .RN(net1),
    .CLK(clknet_3_4__leaf_clk),
    .Q(\main_reg[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[7]$_DFFE_PN0P_  (.D(_029_),
    .RN(net1),
    .CLK(clknet_3_5__leaf_clk),
    .Q(\main_reg[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[8]$_DFFE_PN0P_  (.D(_030_),
    .RN(net1),
    .CLK(clknet_3_5__leaf_clk),
    .Q(\main_reg[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \main_reg[9]$_DFFE_PN0P_  (.D(_031_),
    .RN(net1),
    .CLK(clknet_3_5__leaf_clk),
    .Q(\main_reg[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[0]$_DFFE_PN0P_  (.D(_032_),
    .RN(net1),
    .CLK(clknet_3_2__leaf_clk),
    .Q(net102));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[10]$_DFFE_PN0P_  (.D(_033_),
    .RN(net1),
    .CLK(clknet_3_3__leaf_clk),
    .Q(net103));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[11]$_DFFE_PN0P_  (.D(_034_),
    .RN(net1),
    .CLK(clknet_3_6__leaf_clk),
    .Q(net104));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[12]$_DFFE_PN0P_  (.D(_035_),
    .RN(net1),
    .CLK(clknet_3_2__leaf_clk),
    .Q(net105));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[13]$_DFFE_PN0P_  (.D(_036_),
    .RN(net1),
    .CLK(clknet_3_3__leaf_clk),
    .Q(net106));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[14]$_DFFE_PN0P_  (.D(_037_),
    .RN(net1),
    .CLK(clknet_3_2__leaf_clk),
    .Q(net107));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[15]$_DFFE_PN0P_  (.D(_038_),
    .RN(net1),
    .CLK(clknet_3_2__leaf_clk),
    .Q(net108));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[16]$_DFFE_PN0P_  (.D(_039_),
    .RN(net1),
    .CLK(clknet_3_2__leaf_clk),
    .Q(net109));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[17]$_DFFE_PN0P_  (.D(_040_),
    .RN(net1),
    .CLK(clknet_3_3__leaf_clk),
    .Q(net110));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[18]$_DFFE_PN0P_  (.D(_041_),
    .RN(net1),
    .CLK(clknet_3_3__leaf_clk),
    .Q(net111));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[19]$_DFFE_PN0P_  (.D(_042_),
    .RN(net1),
    .CLK(clknet_3_1__leaf_clk),
    .Q(net112));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[1]$_DFFE_PN0P_  (.D(_043_),
    .RN(net1),
    .CLK(clknet_3_3__leaf_clk),
    .Q(net113));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[20]$_DFFE_PN0P_  (.D(_044_),
    .RN(net1),
    .CLK(clknet_3_0__leaf_clk),
    .Q(net114));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[21]$_DFFE_PN0P_  (.D(_045_),
    .RN(net1),
    .CLK(clknet_3_0__leaf_clk),
    .Q(net115));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[22]$_DFFE_PN0P_  (.D(_046_),
    .RN(net1),
    .CLK(clknet_3_1__leaf_clk),
    .Q(net116));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[23]$_DFFE_PN0P_  (.D(_047_),
    .RN(net1),
    .CLK(clknet_3_1__leaf_clk),
    .Q(net117));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[24]$_DFFE_PN0P_  (.D(_048_),
    .RN(net1),
    .CLK(clknet_3_1__leaf_clk),
    .Q(net118));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[25]$_DFFE_PN0P_  (.D(_049_),
    .RN(net1),
    .CLK(clknet_3_1__leaf_clk),
    .Q(net119));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[26]$_DFFE_PN0P_  (.D(_050_),
    .RN(net1),
    .CLK(clknet_3_0__leaf_clk),
    .Q(net120));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[27]$_DFFE_PN0P_  (.D(_051_),
    .RN(net1),
    .CLK(clknet_3_3__leaf_clk),
    .Q(net121));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[28]$_DFFE_PN0P_  (.D(_052_),
    .RN(net1),
    .CLK(clknet_3_6__leaf_clk),
    .Q(net122));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[29]$_DFFE_PN0P_  (.D(_053_),
    .RN(net1),
    .CLK(clknet_3_4__leaf_clk),
    .Q(net123));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[2]$_DFFE_PN0P_  (.D(_054_),
    .RN(net1),
    .CLK(clknet_3_4__leaf_clk),
    .Q(net124));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[30]$_DFFE_PN0P_  (.D(_055_),
    .RN(net1),
    .CLK(clknet_3_6__leaf_clk),
    .Q(net125));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[31]$_DFFE_PN0P_  (.D(_056_),
    .RN(net1),
    .CLK(clknet_3_4__leaf_clk),
    .Q(net126));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[3]$_DFFE_PN0P_  (.D(_057_),
    .RN(net1),
    .CLK(clknet_3_6__leaf_clk),
    .Q(net127));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[4]$_DFFE_PN0P_  (.D(_058_),
    .RN(net1),
    .CLK(clknet_3_7__leaf_clk),
    .Q(net128));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[5]$_DFFE_PN0P_  (.D(_059_),
    .RN(net1),
    .CLK(clknet_3_5__leaf_clk),
    .Q(net129));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[6]$_DFFE_PN0P_  (.D(_060_),
    .RN(net1),
    .CLK(clknet_3_7__leaf_clk),
    .Q(net130));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[7]$_DFFE_PN0P_  (.D(_061_),
    .RN(net1),
    .CLK(clknet_3_5__leaf_clk),
    .Q(net131));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[8]$_DFFE_PN0P_  (.D(_062_),
    .RN(net1),
    .CLK(clknet_3_5__leaf_clk),
    .Q(net132));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \shadow_reg[9]$_DFFE_PN0P_  (.D(_063_),
    .RN(net1),
    .CLK(clknet_3_5__leaf_clk),
    .Q(net133));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 hold1 (.I(net134),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Right_145 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Right_146 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Right_147 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Right_148 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Right_149 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Right_150 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Right_151 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Right_152 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Right_153 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Right_154 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Right_155 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Right_156 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Right_157 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Right_158 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_159_Right_159 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_160_Right_160 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_161_Right_161 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_162_Right_162 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_163_Right_163 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_164_Right_164 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_165_Right_165 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_166_Right_166 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_167_Right_167 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_168_Right_168 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_169_Right_169 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_170_Right_170 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_171_Right_171 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_172_Right_172 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_173_Right_173 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_174_Right_174 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_175_Right_175 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_176_Right_176 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_177_Right_177 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_178_Right_178 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_179_Right_179 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_180_Right_180 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_181_Right_181 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_182_Right_182 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_183_Right_183 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_184_Right_184 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_185_Right_185 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_186_Right_186 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_187_Right_187 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_188_Right_188 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_189_Right_189 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_190_Right_190 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_191_Right_191 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_192_Right_192 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_193_Right_193 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_194_Right_194 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_195_Right_195 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_196_Right_196 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_197_Right_197 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_198_Right_198 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_199_Right_199 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_200_Right_200 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_201_Right_201 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_202_Right_202 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_203_Right_203 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_204_Right_204 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_205_Right_205 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_206_Right_206 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_207_Right_207 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_208_Right_208 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_209_Right_209 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_210_Right_210 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_211_Right_211 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_212_Right_212 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_213_Right_213 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_214_Right_214 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_215_Right_215 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_216_Right_216 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_217_Right_217 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_218_Right_218 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_219_Right_219 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_220_Right_220 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_221_Right_221 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_222_Right_222 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_223_Right_223 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_224_Right_224 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_225_Right_225 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_226_Right_226 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_227_Right_227 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_228_Right_228 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_229_Right_229 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_230_Right_230 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_231_Right_231 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_232_Right_232 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_233_Right_233 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_234_Right_234 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_235_Right_235 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_236_Right_236 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_237_Right_237 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_238_Right_238 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_239_Right_239 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_240_Right_240 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_241_Right_241 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_242_Right_242 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_243_Right_243 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_244_Right_244 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_245_Right_245 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_246_Right_246 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_247_Right_247 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_248_Right_248 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_249_Right_249 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_250_Right_250 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_251_Right_251 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_252_Right_252 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_253_Right_253 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_254_Right_254 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_255_Right_255 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_256_Right_256 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_257_Right_257 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_258_Right_258 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_259_Right_259 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_260_Right_260 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_261_Right_261 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_262_Right_262 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_263_Right_263 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_264_Right_264 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_265_Right_265 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_266_Right_266 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_267_Right_267 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_268_Right_268 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_269_Right_269 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_270_Right_270 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_271_Right_271 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_272_Right_272 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_273_Right_273 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_274_Right_274 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_275_Right_275 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_276_Right_276 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_277_Right_277 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_278_Right_278 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_279_Right_279 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_280_Right_280 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_281_Right_281 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_282_Right_282 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_283_Right_283 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_284_Right_284 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_285_Right_285 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_286_Right_286 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_287_Right_287 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_288_Right_288 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_289_Right_289 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_290_Right_290 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_291_Right_291 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_292_Right_292 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_293_Right_293 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_294 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_295 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_296 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_297 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_298 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_299 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_300 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_301 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_302 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_303 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_304 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_305 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_306 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_307 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_308 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_309 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_310 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_311 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_312 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_313 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_314 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_315 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_316 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_317 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_318 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_319 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_320 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_321 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_322 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_323 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_324 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_325 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_326 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_327 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_328 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_329 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_330 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_331 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_332 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_333 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_334 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_335 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_336 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Left_337 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Left_338 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Left_339 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Left_340 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Left_341 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Left_342 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Left_343 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Left_344 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Left_345 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Left_346 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Left_347 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Left_348 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Left_349 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Left_350 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Left_351 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Left_352 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Left_353 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Left_354 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Left_355 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Left_356 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Left_357 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Left_358 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Left_359 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Left_360 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Left_361 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Left_362 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Left_363 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Left_364 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Left_365 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Left_366 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Left_367 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Left_368 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Left_369 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Left_370 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Left_371 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Left_372 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Left_373 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Left_374 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Left_375 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Left_376 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Left_377 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Left_378 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Left_379 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Left_380 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Left_381 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Left_382 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Left_383 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Left_384 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Left_385 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Left_386 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Left_387 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Left_388 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Left_389 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Left_390 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Left_391 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Left_392 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Left_393 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Left_394 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Left_395 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Left_396 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Left_397 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Left_398 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Left_399 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Left_400 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Left_401 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Left_402 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Left_403 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Left_404 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Left_405 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Left_406 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Left_407 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Left_408 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Left_409 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Left_410 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Left_411 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Left_412 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Left_413 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Left_414 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Left_415 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Left_416 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Left_417 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Left_418 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Left_419 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Left_420 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Left_421 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Left_422 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Left_423 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Left_424 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Left_425 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Left_426 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Left_427 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Left_428 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Left_429 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Left_430 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Left_431 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Left_432 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Left_433 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Left_434 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Left_435 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Left_436 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Left_437 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Left_438 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Left_439 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Left_440 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Left_441 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Left_442 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Left_443 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Left_444 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Left_445 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Left_446 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Left_447 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Left_448 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Left_449 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Left_450 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Left_451 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Left_452 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_159_Left_453 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_160_Left_454 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_161_Left_455 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_162_Left_456 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_163_Left_457 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_164_Left_458 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_165_Left_459 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_166_Left_460 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_167_Left_461 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_168_Left_462 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_169_Left_463 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_170_Left_464 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_171_Left_465 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_172_Left_466 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_173_Left_467 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_174_Left_468 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_175_Left_469 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_176_Left_470 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_177_Left_471 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_178_Left_472 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_179_Left_473 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_180_Left_474 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_181_Left_475 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_182_Left_476 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_183_Left_477 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_184_Left_478 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_185_Left_479 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_186_Left_480 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_187_Left_481 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_188_Left_482 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_189_Left_483 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_190_Left_484 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_191_Left_485 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_192_Left_486 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_193_Left_487 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_194_Left_488 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_195_Left_489 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_196_Left_490 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_197_Left_491 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_198_Left_492 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_199_Left_493 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_200_Left_494 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_201_Left_495 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_202_Left_496 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_203_Left_497 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_204_Left_498 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_205_Left_499 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_206_Left_500 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_207_Left_501 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_208_Left_502 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_209_Left_503 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_210_Left_504 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_211_Left_505 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_212_Left_506 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_213_Left_507 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_214_Left_508 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_215_Left_509 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_216_Left_510 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_217_Left_511 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_218_Left_512 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_219_Left_513 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_220_Left_514 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_221_Left_515 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_222_Left_516 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_223_Left_517 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_224_Left_518 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_225_Left_519 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_226_Left_520 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_227_Left_521 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_228_Left_522 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_229_Left_523 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_230_Left_524 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_231_Left_525 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_232_Left_526 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_233_Left_527 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_234_Left_528 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_235_Left_529 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_236_Left_530 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_237_Left_531 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_238_Left_532 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_239_Left_533 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_240_Left_534 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_241_Left_535 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_242_Left_536 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_243_Left_537 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_244_Left_538 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_245_Left_539 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_246_Left_540 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_247_Left_541 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_248_Left_542 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_249_Left_543 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_250_Left_544 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_251_Left_545 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_252_Left_546 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_253_Left_547 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_254_Left_548 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_255_Left_549 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_256_Left_550 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_257_Left_551 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_258_Left_552 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_259_Left_553 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_260_Left_554 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_261_Left_555 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_262_Left_556 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_263_Left_557 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_264_Left_558 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_265_Left_559 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_266_Left_560 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_267_Left_561 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_268_Left_562 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_269_Left_563 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_270_Left_564 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_271_Left_565 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_272_Left_566 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_273_Left_567 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_274_Left_568 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_275_Left_569 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_276_Left_570 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_277_Left_571 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_278_Left_572 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_279_Left_573 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_280_Left_574 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_281_Left_575 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_282_Left_576 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_283_Left_577 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_284_Left_578 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_285_Left_579 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_286_Left_580 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_287_Left_581 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_288_Left_582 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_289_Left_583 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_290_Left_584 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_291_Left_585 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_292_Left_586 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_293_Left_587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_961 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_962 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_963 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_964 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_965 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_966 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_967 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_968 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_969 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_970 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_971 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_972 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_973 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_974 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_975 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_976 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_977 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_978 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_979 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_980 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_981 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_982 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_983 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_984 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_985 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_986 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_987 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_988 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_989 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_990 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_991 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_992 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_993 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_994 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_995 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_996 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_997 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_998 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_999 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_1961 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_1962 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_1963 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_1965 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_1966 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1967 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1969 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1971 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_1978 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1981 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1983 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1985 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1987 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_1988 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_1989 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_1991 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_1993 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_1995 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_1998 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_2001 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_2003 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_2004 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_2010 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_2014 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_2015 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_2017 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_2018 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_2019 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_2020 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_2023 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_2025 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_2027 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_2028 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_2029 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_2030 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_2031 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_2032 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_2033 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_2034 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_2035 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_2036 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_2037 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_2039 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_2041 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_2043 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_2044 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_2045 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_2047 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_2048 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_2051 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_2052 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_2053 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_2054 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_2059 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_2060 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_2061 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_2063 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_2065 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_2067 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_2069 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_2071 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_2072 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_2073 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_2074 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_2075 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_2076 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_2077 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_2078 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_2080 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_2082 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_2085 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_2086 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_2087 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_2089 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_2090 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_2091 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_2092 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_2093 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_2096 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_2098 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_2099 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_2100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_2107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_2112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_2121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_2123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_2125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_2127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_2128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_2136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_2137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_2139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_2140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_2141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_2142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_2143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_2144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_2145 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_2146 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_2147 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_2148 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_2149 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_2150 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_2151 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_2153 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_2155 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_2156 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_2157 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_2158 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_2159 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_2160 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_2161 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_2163 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_2164 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_2165 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_2166 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_2167 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_2168 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_2169 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_2170 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_2171 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_2172 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_2173 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_2174 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_2175 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_2176 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_2177 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_2178 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_2179 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_2180 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_2181 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_2182 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_2183 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_2184 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_2185 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_2186 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_2187 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_2188 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_2189 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_2190 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_2191 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_2192 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_2193 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_2194 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_2195 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_2196 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_2197 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_2198 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_2199 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_2200 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_2201 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_2203 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_2204 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_2205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_2206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_2207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_2208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_2209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_2210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_2211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_2212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_2213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_2217 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_2221 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_2222 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_2223 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_2224 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_2225 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_2226 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_2227 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_2228 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_2229 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_2230 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_2231 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_2232 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_2233 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_2234 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_2235 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_2236 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_2237 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_2238 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_2239 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_2240 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_2241 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_2242 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_2243 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_2244 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_2245 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_2246 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_2247 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_2248 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_2249 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_2250 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_2251 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_2252 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_2253 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_2254 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_2255 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_2256 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_2257 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_2258 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_2259 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_2260 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_2261 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_2262 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_2263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_2264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_2265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_2267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_2268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_2269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_2270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_2271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_2272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_2273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_2274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_2275 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_2276 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_2277 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_2278 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_2279 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_2281 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_2282 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_2283 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_2284 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_2285 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_2286 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_2287 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_2288 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_2289 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_2290 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_2291 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_2292 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_2293 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_2294 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_2295 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_2296 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_2297 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_2298 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_2299 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_2300 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_2301 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_2302 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_2303 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_2304 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_2305 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_2306 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_2307 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_2308 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_2309 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_2310 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_2311 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_2314 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_2315 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_2317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_2318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_2319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_2320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_2321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_2322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_2323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_2324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_2325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_2326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_2327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_2328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_2329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_2331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_2332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_2333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_2334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_2335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_2336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_2337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_2338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_2339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_2340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_2341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_2342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_2343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_2344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_2345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_2346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_2347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_2348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_2349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_2350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_2351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_2352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_2353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_2354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_2355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_2356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_2357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_2358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_2359 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_2360 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_2361 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_2362 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_2363 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_2364 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_2365 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_2366 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_2367 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_2368 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_2369 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_2370 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_2371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_2372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_2373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_2374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_2375 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_2376 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_2377 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_2378 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_2379 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_2381 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_2382 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_2383 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_2384 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_2385 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_2386 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_2387 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_2388 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_2389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_2390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_2391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_2392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_2393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_2395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_2396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_2397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_2398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_2399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_2400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_2401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_2402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_2403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_2404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_2405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_2406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_2407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_2408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_2409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_2410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_2411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_2412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_2413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_2414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_2415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_2416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_2417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_2418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_2419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_2420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_2421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_2422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_2423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_2424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_2425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_2426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_2427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_2428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_2429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_2430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_2431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_2432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_2433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_2434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_2435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_2436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_2437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_2438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_2439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_2440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_2441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_2442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_2443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_2445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_2446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_2447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_2448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_2449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_2450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_2451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_2452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_2453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_2454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_2455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_2456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_2457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_2459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_2460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_2461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_2462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_2463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_2464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_2465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_2466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_2467 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_2468 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_2469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_2470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_2471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_2472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_2473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_2474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_2475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_2476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_2477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_2478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_2479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_2480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_2481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_2482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_2483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_2484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_2485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_2486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_2487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_2488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_2489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_2492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_2493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_2495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_2496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_2497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_2498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_2499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_2500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_2501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_2502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_2503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_2504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_2505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_2506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_2507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_2509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_2510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_2511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_2512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_2513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_2514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_2515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_2516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_2517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_2518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_2519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_2520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_2521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_2522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_2523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_2524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_2525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_2526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_2527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_2528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_2529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_2530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_2531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_2532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_2533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_2534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_2535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_2536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_2537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_2538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_2539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_2540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_2541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_2542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_2543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_2544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_2545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_2546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_2547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_2548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_2549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_2550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_2551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_2552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_2553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_2554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_2555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_2556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_2557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_2559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_2560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_2561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_2562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_2563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_2564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_2565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_2566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_2567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_2568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_2569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_2570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_2571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_2573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_2574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_2575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_2576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_2577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_2578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_2579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_2580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_2581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_2582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_2583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_2584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_2585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_2586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_2587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_2588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_2589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_2590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_2591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_2592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_2593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_2594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_2595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_2596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_2597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_2598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_2599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_2600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_2601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_2602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_2603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_2604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_2605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_2606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_2607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_2608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_2609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_2610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_2611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_2612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_2613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_2614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_2615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_2616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_2617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_2618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_2619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_2620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_2621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_2623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_2624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_2625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_2626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_2627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_2628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_2629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_2630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_2631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_2632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_2633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_2634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_2635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_2637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_2639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_2640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_2641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_2642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_2643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_2644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_2645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_2647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_2648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_2649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_2651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_2652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_2653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_2654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_2655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_2656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_2657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_2658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_2659 ();
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input1 (.I(main_data_in[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(main_data_in[10]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(main_data_in[11]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(main_data_in[12]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(main_data_in[13]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(main_data_in[14]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(main_data_in[15]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(main_data_in[16]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(main_data_in[17]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(main_data_in[18]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input11 (.I(main_data_in[19]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input12 (.I(main_data_in[1]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input13 (.I(main_data_in[20]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input14 (.I(main_data_in[21]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input15 (.I(main_data_in[22]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input16 (.I(main_data_in[23]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input17 (.I(main_data_in[24]),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input18 (.I(main_data_in[25]),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input19 (.I(main_data_in[26]),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input20 (.I(main_data_in[27]),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input21 (.I(main_data_in[28]),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input22 (.I(main_data_in[29]),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input23 (.I(main_data_in[2]),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input24 (.I(main_data_in[30]),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input25 (.I(main_data_in[31]),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input26 (.I(main_data_in[3]),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input27 (.I(main_data_in[4]),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input28 (.I(main_data_in[5]),
    .Z(net29));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input29 (.I(main_data_in[6]),
    .Z(net30));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input30 (.I(main_data_in[7]),
    .Z(net31));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input31 (.I(main_data_in[8]),
    .Z(net32));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input32 (.I(main_data_in[9]),
    .Z(net33));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 input33 (.I(main_load_en),
    .Z(net34));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 input34 (.I(shadow_capture_en),
    .Z(net35));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input35 (.I(shadow_data_in[0]),
    .Z(net36));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input36 (.I(shadow_data_in[10]),
    .Z(net37));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input37 (.I(shadow_data_in[11]),
    .Z(net38));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input38 (.I(shadow_data_in[12]),
    .Z(net39));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input39 (.I(shadow_data_in[13]),
    .Z(net40));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input40 (.I(shadow_data_in[14]),
    .Z(net41));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input41 (.I(shadow_data_in[15]),
    .Z(net42));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input42 (.I(shadow_data_in[16]),
    .Z(net43));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input43 (.I(shadow_data_in[17]),
    .Z(net44));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input44 (.I(shadow_data_in[18]),
    .Z(net45));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input45 (.I(shadow_data_in[19]),
    .Z(net46));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input46 (.I(shadow_data_in[1]),
    .Z(net47));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input47 (.I(shadow_data_in[20]),
    .Z(net48));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input48 (.I(shadow_data_in[21]),
    .Z(net49));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input49 (.I(shadow_data_in[22]),
    .Z(net50));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input50 (.I(shadow_data_in[23]),
    .Z(net51));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input51 (.I(shadow_data_in[24]),
    .Z(net52));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input52 (.I(shadow_data_in[25]),
    .Z(net53));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input53 (.I(shadow_data_in[26]),
    .Z(net54));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input54 (.I(shadow_data_in[27]),
    .Z(net55));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input55 (.I(shadow_data_in[28]),
    .Z(net56));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input56 (.I(shadow_data_in[29]),
    .Z(net57));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input57 (.I(shadow_data_in[2]),
    .Z(net58));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input58 (.I(shadow_data_in[30]),
    .Z(net59));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input59 (.I(shadow_data_in[31]),
    .Z(net60));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input60 (.I(shadow_data_in[3]),
    .Z(net61));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input61 (.I(shadow_data_in[4]),
    .Z(net62));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input62 (.I(shadow_data_in[5]),
    .Z(net63));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input63 (.I(shadow_data_in[6]),
    .Z(net64));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input64 (.I(shadow_data_in[7]),
    .Z(net65));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input65 (.I(shadow_data_in[8]),
    .Z(net66));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input66 (.I(shadow_data_in[9]),
    .Z(net67));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input67 (.I(shadow_load_en),
    .Z(net68));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 input68 (.I(use_shadow_out),
    .Z(net69));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output69 (.I(net70),
    .Z(main_data_out[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output70 (.I(net71),
    .Z(main_data_out[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output71 (.I(net72),
    .Z(main_data_out[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output72 (.I(net73),
    .Z(main_data_out[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output73 (.I(net74),
    .Z(main_data_out[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output74 (.I(net75),
    .Z(main_data_out[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output75 (.I(net76),
    .Z(main_data_out[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output76 (.I(net77),
    .Z(main_data_out[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output77 (.I(net78),
    .Z(main_data_out[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output78 (.I(net79),
    .Z(main_data_out[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output79 (.I(net80),
    .Z(main_data_out[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output80 (.I(net81),
    .Z(main_data_out[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output81 (.I(net82),
    .Z(main_data_out[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output82 (.I(net83),
    .Z(main_data_out[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output83 (.I(net84),
    .Z(main_data_out[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output84 (.I(net85),
    .Z(main_data_out[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output85 (.I(net86),
    .Z(main_data_out[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output86 (.I(net87),
    .Z(main_data_out[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output87 (.I(net88),
    .Z(main_data_out[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output88 (.I(net89),
    .Z(main_data_out[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output89 (.I(net90),
    .Z(main_data_out[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output90 (.I(net91),
    .Z(main_data_out[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output91 (.I(net92),
    .Z(main_data_out[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output92 (.I(net93),
    .Z(main_data_out[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output93 (.I(net94),
    .Z(main_data_out[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output94 (.I(net95),
    .Z(main_data_out[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output95 (.I(net96),
    .Z(main_data_out[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output96 (.I(net97),
    .Z(main_data_out[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output97 (.I(net98),
    .Z(main_data_out[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output98 (.I(net99),
    .Z(main_data_out[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output99 (.I(net100),
    .Z(main_data_out[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output100 (.I(net101),
    .Z(main_data_out[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output101 (.I(net102),
    .Z(shadow_data_out[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output102 (.I(net103),
    .Z(shadow_data_out[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output103 (.I(net104),
    .Z(shadow_data_out[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output104 (.I(net105),
    .Z(shadow_data_out[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output105 (.I(net106),
    .Z(shadow_data_out[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output106 (.I(net107),
    .Z(shadow_data_out[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output107 (.I(net108),
    .Z(shadow_data_out[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output108 (.I(net109),
    .Z(shadow_data_out[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output109 (.I(net110),
    .Z(shadow_data_out[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output110 (.I(net111),
    .Z(shadow_data_out[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output111 (.I(net112),
    .Z(shadow_data_out[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output112 (.I(net113),
    .Z(shadow_data_out[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output113 (.I(net114),
    .Z(shadow_data_out[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output114 (.I(net115),
    .Z(shadow_data_out[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output115 (.I(net116),
    .Z(shadow_data_out[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output116 (.I(net117),
    .Z(shadow_data_out[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output117 (.I(net118),
    .Z(shadow_data_out[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output118 (.I(net119),
    .Z(shadow_data_out[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output119 (.I(net120),
    .Z(shadow_data_out[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output120 (.I(net121),
    .Z(shadow_data_out[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output121 (.I(net122),
    .Z(shadow_data_out[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output122 (.I(net123),
    .Z(shadow_data_out[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output123 (.I(net124),
    .Z(shadow_data_out[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output124 (.I(net125),
    .Z(shadow_data_out[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output125 (.I(net126),
    .Z(shadow_data_out[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output126 (.I(net127),
    .Z(shadow_data_out[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output127 (.I(net128),
    .Z(shadow_data_out[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output128 (.I(net129),
    .Z(shadow_data_out[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output129 (.I(net130),
    .Z(shadow_data_out[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output130 (.I(net131),
    .Z(shadow_data_out[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output131 (.I(net132),
    .Z(shadow_data_out[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output132 (.I(net133),
    .Z(shadow_data_out[9]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_2_0_0_clk (.I(clknet_0_clk),
    .Z(clknet_2_0_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_2_1_0_clk (.I(clknet_0_clk),
    .Z(clknet_2_1_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_2_2_0_clk (.I(clknet_0_clk),
    .Z(clknet_2_2_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_2_3_0_clk (.I(clknet_0_clk),
    .Z(clknet_2_3_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_3_0__f_clk (.I(clknet_2_0_0_clk),
    .Z(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_3_1__f_clk (.I(clknet_2_0_0_clk),
    .Z(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_3_2__f_clk (.I(clknet_2_1_0_clk),
    .Z(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_3_3__f_clk (.I(clknet_2_1_0_clk),
    .Z(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_3_4__f_clk (.I(clknet_2_2_0_clk),
    .Z(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_3_5__f_clk (.I(clknet_2_2_0_clk),
    .Z(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_3_6__f_clk (.I(clknet_2_3_0_clk),
    .Z(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_3_7__f_clk (.I(clknet_2_3_0_clk),
    .Z(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload0 (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload1 (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload2 (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload3 (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net134));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_1 (.I(net1));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_2 (.I(net1));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_2048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_2052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_2308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_2604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_2606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_2590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_2594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_2625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_2633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_2588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_2592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_2594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_2644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_2590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_2594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_2645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_2649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_2651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_2588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_2592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_2643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_2651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_2590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_2643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_2651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_2588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_2596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_2600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_2647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_2651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_2590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_2606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_2614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_2616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_2647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_2651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_2590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_2647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_2651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_2588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_2596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_2590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_2606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_2608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_2624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_2632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_2634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_2604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_2606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_2630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_2634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_191_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_197_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_199_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_201_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_203_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_205_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_207_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_208_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_208_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_209_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_210_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_210_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_211_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_213_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_214_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_214_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_215_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_215_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_216_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_216_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_217_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_218_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_218_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_219_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_219_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_220_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_220_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_221_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_221_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_222_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_222_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_223_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_223_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_223_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_224_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_224_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_225_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_227_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_227_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_228_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_228_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_229_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_229_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_230_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_230_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_231_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_231_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_232_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_232_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_233_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_233_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_233_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_233_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_235_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_235_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_235_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_236_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_236_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_237_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_237_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_237_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_238_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_238_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_239_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_239_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_239_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_240_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_240_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_241_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_241_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_241_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_242_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_242_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_243_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_243_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_243_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_244_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_244_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_245_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_245_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_246_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_246_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_247_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_247_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_247_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_248_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_248_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_249_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_249_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_249_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_250_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_250_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_251_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_251_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_251_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_252_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_252_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_253_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_253_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_253_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_254_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_254_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_255_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_255_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_255_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_256_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_256_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_257_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_257_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_257_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_258_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_258_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_259_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_259_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_259_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_260_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_260_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_261_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_261_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_261_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_262_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_262_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_263_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_263_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_263_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_264_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_264_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_265_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_265_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_265_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_266_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_266_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_267_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_267_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_267_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_268_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_268_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_269_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_269_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_269_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_270_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_270_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_271_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_271_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_271_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_272_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_272_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_273_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_273_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_273_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_274_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_274_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_275_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_275_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_275_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_276_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_276_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_277_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_277_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_277_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_277_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_277_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_277_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_277_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_277_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_277_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_277_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_277_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_278_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_278_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_278_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_278_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_278_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_278_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_278_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_278_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_278_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_278_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_279_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_279_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_279_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_279_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_279_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_279_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_280_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_280_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_280_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_280_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_280_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_280_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_280_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_281_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_281_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_281_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_281_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_281_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_281_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_282_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_282_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_282_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_282_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_282_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_282_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_283_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_283_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_283_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_283_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_283_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_283_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_283_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_283_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_283_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_284_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_284_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_284_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_284_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_284_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_284_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_285_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_285_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_285_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_285_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_285_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_285_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_285_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_285_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_286_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_286_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_286_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_286_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_286_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_286_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_286_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_286_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_286_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_287_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_287_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_287_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_287_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_287_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_287_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_287_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_287_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_287_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_287_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_287_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_288_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_288_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_288_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_288_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_288_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_288_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_288_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_288_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_288_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_288_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_288_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_289_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_289_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_289_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_289_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_289_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_289_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_289_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_289_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_289_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_289_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_289_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_290_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_290_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_290_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_290_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_290_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_290_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_290_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_290_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_290_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_290_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_290_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_290_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_291_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_291_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_291_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_291_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_291_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_291_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_291_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_291_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_291_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_292_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_292_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_292_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_292_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_292_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_292_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_292_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_292_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_292_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_293_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_293_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_293_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_293_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_293_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_293_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_293_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_293_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_293_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_293_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_293_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_293_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_293_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_293_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_293_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_293_2298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_293_2476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_293_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_293_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_293_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_2650 ();
endmodule
