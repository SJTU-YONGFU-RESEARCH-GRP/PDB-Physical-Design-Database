module constant(
    output y
);

assign y = 0;
endmodule