
* cell smart_fifo
.SUBCKT smart_fifo
* net 1 wr_data[31]
* net 2 wr_data[2]
* net 3 wr_data[30]
* net 4 wr_data[3]
* net 5 wr_data[4]
* net 6 wr_data[5]
* net 7 wr_data[6]
* net 8 wr_data[7]
* net 9 wr_data[8]
* net 10 wr_data[9]
* net 11 wr_data[10]
* net 12 wr_data[11]
* net 13 wr_data[12]
* net 23 PWELL
* net 37 clk
* net 38 NWELL
* net 160 wr_data[13]
* net 625 wr_data[29]
* net 626 wr_data[28]
* net 842 wr_data[14]
* net 1010 wr_data[0]
* net 1113 wr_data[15]
* net 1167 rd_data[28]
* net 1200 rd_data[31]
* net 1201 rd_data[4]
* net 1258 rd_data[29]
* net 1259 rd_data[3]
* net 1260 rd_data[6]
* net 1274 rd_data[9]
* net 1275 rd_data[8]
* net 1276 rd_data[13]
* net 1290 rd_data[5]
* net 1308 rd_data[7]
* net 1322 wr_data[27]
* net 1323 rd_data[30]
* net 1341 rd_data[11]
* net 1342 rd_data[10]
* net 1360 rd_data[2]
* net 1381 wr_data[16]
* net 1382 rd_data[12]
* net 1395 rd_data[27]
* net 1421 data_count[4]
* net 1422 rd_data[0]
* net 1464 rd_data[14]
* net 1465 rd_valid
* net 1466 rd_data[15]
* net 1555 wr_data[26]
* net 1569 rd_data[16]
* net 1653 rd_data[17]
* net 1688 rd_data[26]
* net 1867 wr_data[25]
* net 1889 wr_data[18]
* net 1921 wr_data[17]
* net 2028 error_detected
* net 2070 underflow_detected
* net 2071 clear_errors
* net 2122 error_count[1]
* net 2162 error_count[4]
* net 2163 error_count[3]
* net 2164 error_count[0]
* net 2256 error_count[6]
* net 2294 error_count[8]
* net 2295 error_count[7]
* net 2374 error_count[10]
* net 2417 error_count[5]
* net 2454 rd_en
* net 2515 wr_data[24]
* net 2516 wr_data[23]
* net 2517 wr_data[22]
* net 2518 rd_data[24]
* net 2519 rd_data[23]
* net 2520 rd_data[25]
* net 2522 rd_data[22]
* net 2523 wr_data[21]
* net 2525 rd_data[21]
* net 2526 wr_data[19]
* net 2527 rd_data[20]
* net 2528 rd_data[19]
* net 2529 rd_data[1]
* net 2530 wr_data[1]
* net 2532 wr_data[20]
* net 2533 wr_en
* net 2534 rd_data[18]
* net 2535 overflow_detected
* net 2537 wr_ready
* net 2538 full
* net 2539 rst_n
* net 2540 empty
* net 2541 data_count[1]
* net 2542 data_count[2]
* net 2543 data_count[0]
* net 2544 almost_empty
* net 2545 almost_full
* net 2547 data_count[3]
* net 2548 error_count[15]
* net 2551 error_count[9]
* net 2552 error_count[12]
* net 2553 error_count[2]
* net 2554 error_count[13]
* net 2555 error_count[11]
* net 2556 error_count[14]
* cell instance $1 r0 *1 10.175,0.35
X$1 1 VIA_via5_0
* cell instance $2 r0 *1 18.905,0.07
X$2 1 VIA_via2_5
* cell instance $3 r0 *1 18.905,2.03
X$3 1 VIA_via1_4
* cell instance $4 r0 *1 18.81,1.4
X$4 1 23 38 26 CLKBUF_X2
* cell instance $5 r0 *1 19.135,0.07
X$5 1 VIA_via3_2
* cell instance $6 r0 *1 19.135,0.07
X$6 1 VIA_via4_0
* cell instance $7 r0 *1 8.455,2.03
X$7 2 VIA_via1_4
* cell instance $8 r0 *1 8.36,1.4
X$8 2 23 38 27 CLKBUF_X2
* cell instance $9 r0 *1 8.455,2.03
X$9 2 VIA_via2_5
* cell instance $10 r0 *1 8.495,2.03
X$10 2 VIA_via3_2
* cell instance $11 r0 *1 8.495,2.03
X$11 2 VIA_via4_0
* cell instance $12 r0 *1 8.495,2.03
X$12 2 VIA_via5_0
* cell instance $13 r0 *1 9.615,2.03
X$13 3 VIA_via3_2
* cell instance $14 r0 *1 9.595,2.03
X$14 3 VIA_via2_5
* cell instance $15 r0 *1 9.615,2.03
X$15 3 VIA_via4_0
* cell instance $16 r0 *1 9.615,2.03
X$16 3 VIA_via5_0
* cell instance $17 r0 *1 9.595,2.03
X$17 3 VIA_via1_4
* cell instance $18 r0 *1 9.5,1.4
X$18 3 23 38 24 CLKBUF_X2
* cell instance $19 r0 *1 28.025,2.03
X$19 4 VIA_via1_4
* cell instance $20 r0 *1 27.93,1.4
X$20 4 23 38 29 BUF_X1
* cell instance $21 r0 *1 28.025,2.03
X$21 4 VIA_via2_5
* cell instance $22 r0 *1 28.095,2.03
X$22 4 VIA_via3_2
* cell instance $23 r0 *1 28.095,2.03
X$23 4 VIA_via4_0
* cell instance $24 r0 *1 28.095,2.03
X$24 4 VIA_via5_0
* cell instance $25 r0 *1 32.965,2.03
X$25 5 VIA_via1_4
* cell instance $26 r0 *1 32.87,1.4
X$26 5 23 38 25 CLKBUF_X2
* cell instance $27 r0 *1 32.965,2.03
X$27 5 VIA_via2_5
* cell instance $28 r0 *1 33.135,2.03
X$28 5 VIA_via4_0
* cell instance $29 r0 *1 33.135,2.03
X$29 5 VIA_via3_2
* cell instance $30 r0 *1 33.135,2.03
X$30 5 VIA_via5_0
* cell instance $31 r0 *1 38.095,2.03
X$31 6 VIA_via1_4
* cell instance $32 r0 *1 38,1.4
X$32 6 23 38 98 CLKBUF_X2
* cell instance $33 r0 *1 38.095,2.03
X$33 6 VIA_via2_5
* cell instance $34 r0 *1 38.175,2.03
X$34 6 VIA_via3_2
* cell instance $35 r0 *1 38.175,2.03
X$35 6 VIA_via4_0
* cell instance $36 r0 *1 38.175,2.03
X$36 6 VIA_via5_0
* cell instance $37 r0 *1 45.315,2.03
X$37 7 VIA_via1_4
* cell instance $38 r0 *1 45.22,1.4
X$38 7 23 38 75 CLKBUF_X2
* cell instance $39 r0 *1 45.315,2.03
X$39 7 VIA_via2_5
* cell instance $40 r0 *1 45.455,2.03
X$40 7 VIA_via3_2
* cell instance $41 r0 *1 45.455,2.03
X$41 7 VIA_via4_0
* cell instance $42 r0 *1 45.455,2.03
X$42 7 VIA_via5_0
* cell instance $43 r0 *1 51.965,2.03
X$43 8 VIA_via1_4
* cell instance $44 r0 *1 51.87,1.4
X$44 8 23 38 66 CLKBUF_X2
* cell instance $45 r0 *1 51.965,2.03
X$45 8 VIA_via2_5
* cell instance $46 r0 *1 52.175,2.03
X$46 8 VIA_via4_0
* cell instance $47 r0 *1 52.175,2.03
X$47 8 VIA_via3_2
* cell instance $48 r0 *1 52.175,2.03
X$48 8 VIA_via5_0
* cell instance $49 r0 *1 53.855,2.03
X$49 9 VIA_via5_0
* cell instance $50 r0 *1 53.855,2.03
X$50 9 VIA_via4_0
* cell instance $51 r0 *1 53.855,2.03
X$51 9 VIA_via3_2
* cell instance $52 r0 *1 54.055,2.03
X$52 9 VIA_via1_4
* cell instance $53 r0 *1 53.96,1.4
X$53 9 23 38 112 CLKBUF_X2
* cell instance $54 r0 *1 54.055,2.03
X$54 9 VIA_via2_5
* cell instance $55 r0 *1 59.565,2.03
X$55 10 VIA_via1_4
* cell instance $56 r0 *1 59.47,1.4
X$56 10 23 38 121 CLKBUF_X2
* cell instance $57 r0 *1 59.565,2.03
X$57 10 VIA_via2_5
* cell instance $58 r0 *1 60.015,2.03
X$58 10 VIA_via4_0
* cell instance $59 r0 *1 60.015,2.03
X$59 10 VIA_via3_2
* cell instance $60 r0 *1 60.015,2.03
X$60 10 VIA_via5_0
* cell instance $61 r0 *1 71.725,2.03
X$61 11 VIA_via1_4
* cell instance $62 r0 *1 71.63,1.4
X$62 11 23 38 77 BUF_X1
* cell instance $63 r0 *1 71.725,2.03
X$63 11 VIA_via2_5
* cell instance $64 r0 *1 71.775,2.03
X$64 11 VIA_via3_2
* cell instance $65 r0 *1 71.775,2.03
X$65 11 VIA_via4_0
* cell instance $66 r0 *1 71.775,2.03
X$66 11 VIA_via5_0
* cell instance $67 r0 *1 79.615,1.75
X$67 12 VIA_via5_0
* cell instance $68 r0 *1 79.615,1.75
X$68 12 VIA_via4_0
* cell instance $69 r0 *1 79.895,3.57
X$69 12 VIA_via1_4
* cell instance $70 m0 *1 79.8,4.2
X$70 12 23 38 49 CLKBUF_X2
* cell instance $71 r0 *1 79.895,3.57
X$71 12 VIA_via2_5
* cell instance $72 r0 *1 79.615,3.57
X$72 12 VIA_via3_2
* cell instance $73 r0 *1 92.435,2.03
X$73 13 VIA_via1_4
* cell instance $74 r0 *1 92.34,1.4
X$74 13 23 38 53 CLKBUF_X2
* cell instance $75 r0 *1 92.435,2.03
X$75 13 VIA_via2_5
* cell instance $76 r0 *1 92.495,2.03
X$76 13 VIA_via3_2
* cell instance $77 r0 *1 92.495,2.03
X$77 13 VIA_via4_0
* cell instance $78 r0 *1 92.495,2.03
X$78 13 VIA_via5_0
* cell instance $79 r0 *1 16.625,10.43
X$79 14 VIA_via2_5
* cell instance $80 r0 *1 25.935,9.17
X$80 14 VIA_via2_5
* cell instance $81 r0 *1 26.125,9.17
X$81 14 VIA_via2_5
* cell instance $82 r0 *1 21.755,10.43
X$82 14 VIA_via2_5
* cell instance $83 r0 *1 23.655,9.17
X$83 14 VIA_via2_5
* cell instance $84 r0 *1 19.665,10.43
X$84 14 VIA_via1_4
* cell instance $85 r0 *1 18.05,9.8
X$85 23 3031 250 205 14 38 DFF_X1
* cell instance $86 r0 *1 19.665,10.43
X$86 14 VIA_via2_5
* cell instance $87 r0 *1 23.655,8.05
X$87 14 VIA_via1_4
* cell instance $88 r0 *1 23.18,7
X$88 149 23 38 14 CLKBUF_X3
* cell instance $89 r0 *1 16.625,11.97
X$89 14 VIA_via1_4
* cell instance $90 m0 *1 15.01,12.6
X$90 23 2785 270 271 14 38 DFF_X1
* cell instance $91 r0 *1 21.755,11.97
X$91 14 VIA_via1_4
* cell instance $92 m0 *1 20.14,12.6
X$92 23 2774 273 167 14 38 DFF_X1
* cell instance $93 r0 *1 22.135,9.17
X$93 14 VIA_via1_4
* cell instance $94 m0 *1 22.04,9.8
X$94 14 23 38 CLKBUF_X1
* cell instance $95 r0 *1 22.135,9.17
X$95 14 VIA_via2_5
* cell instance $96 r0 *1 25.555,9.17
X$96 14 VIA_via1_4
* cell instance $97 m0 *1 23.94,9.8
X$97 23 2802 165 193 14 38 DFF_X1
* cell instance $98 r0 *1 25.555,9.17
X$98 14 VIA_via2_5
* cell instance $99 r0 *1 25.935,10.43
X$99 14 VIA_via1_4
* cell instance $100 r0 *1 24.32,9.8
X$100 23 2996 206 168 14 38 DFF_X1
* cell instance $101 r0 *1 26.125,2.03
X$101 14 VIA_via1_4
* cell instance $102 r0 *1 24.51,1.4
X$102 23 2991 21 39 14 38 DFF_X1
* cell instance $103 r0 *1 25.935,4.83
X$103 14 VIA_via1_4
* cell instance $104 r0 *1 24.32,4.2
X$104 23 2947 115 72 14 38 DFF_X1
* cell instance $105 r0 *1 69.065,2.45
X$105 15 VIA_via2_5
* cell instance $106 r0 *1 70.585,2.45
X$106 15 VIA_via2_5
* cell instance $107 r0 *1 70.775,2.03
X$107 15 VIA_via1_4
* cell instance $108 r0 *1 67.64,1.4
X$108 23 2866 15 22 32 38 DFF_X1
* cell instance $109 r0 *1 70.205,4.83
X$109 15 VIA_via1_4
* cell instance $110 r0 *1 69.92,4.2
X$110 15 80 33 23 38 262 MUX2_X1
* cell instance $111 r0 *1 69.065,3.57
X$111 15 VIA_via1_4
* cell instance $112 m0 *1 68.21,4.2
X$112 78 51 15 23 38 22 MUX2_X1
* cell instance $113 r0 *1 78.375,2.03
X$113 16 VIA_via2_5
* cell instance $114 r0 *1 80.465,2.03
X$114 16 VIA_via1_4
* cell instance $115 r0 *1 79.61,1.4
X$115 53 17 16 23 38 20 MUX2_X1
* cell instance $116 r0 *1 80.465,2.03
X$116 16 VIA_via2_5
* cell instance $117 r0 *1 79.135,2.03
X$117 16 VIA_via1_4
* cell instance $118 r0 *1 76,1.4
X$118 23 3109 16 20 34 38 DFF_X1
* cell instance $119 r0 *1 79.135,2.03
X$119 16 VIA_via2_5
* cell instance $120 r0 *1 78.185,4.83
X$120 16 VIA_via1_4
* cell instance $121 r0 *1 77.33,4.2
X$121 50 80 16 23 38 110 MUX2_X1
* cell instance $122 r0 *1 80.655,72.17
X$122 17 VIA_via1_7
* cell instance $123 r0 *1 80.56,71.4
X$123 1111 17 1916 23 38 1886 MUX2_X1
* cell instance $124 r0 *1 75.715,37.03
X$124 17 VIA_via1_7
* cell instance $125 m0 *1 75.62,37.8
X$125 710 17 866 23 38 921 MUX2_X1
* cell instance $126 r0 *1 75.715,37.03
X$126 17 VIA_via2_5
* cell instance $127 r0 *1 66.975,3.43
X$127 17 VIA_via1_7
* cell instance $128 m0 *1 66.88,4.2
X$128 77 17 47 23 38 65 MUX2_X1
* cell instance $129 r0 *1 66.975,3.43
X$129 17 VIA_via2_5
* cell instance $130 r0 *1 79.705,2.17
X$130 17 VIA_via1_7
* cell instance $131 r0 *1 79.705,2.31
X$131 17 VIA_via2_5
* cell instance $132 r0 *1 70.205,3.43
X$132 17 VIA_via1_7
* cell instance $133 m0 *1 70.11,4.2
X$133 49 17 33 23 38 63 MUX2_X1
* cell instance $134 r0 *1 70.205,3.43
X$134 17 VIA_via2_5
* cell instance $135 r0 *1 76.665,58.17
X$135 17 VIA_via1_7
* cell instance $136 r0 *1 76.57,57.4
X$136 1073 17 1498 23 38 1548 MUX2_X1
* cell instance $137 r0 *1 76.665,58.31
X$137 17 VIA_via2_5
* cell instance $138 r0 *1 81.605,45.43
X$138 17 VIA_via1_7
* cell instance $139 m0 *1 81.51,46.2
X$139 806 17 1109 23 38 1110 MUX2_X1
* cell instance $140 r0 *1 81.605,45.43
X$140 17 VIA_via2_5
* cell instance $141 r0 *1 66.975,72.17
X$141 17 VIA_via1_7
* cell instance $142 r0 *1 66.88,71.4
X$142 1335 17 1914 23 38 1896 MUX2_X1
* cell instance $143 r0 *1 81.795,2.31
X$143 17 VIA_via2_5
* cell instance $144 r0 *1 78.375,16.17
X$144 17 VIA_via2_5
* cell instance $145 r0 *1 81.795,16.03
X$145 17 VIA_via2_5
* cell instance $146 r0 *1 69.445,55.79
X$146 17 VIA_via2_5
* cell instance $147 r0 *1 66.975,72.59
X$147 17 VIA_via2_5
* cell instance $148 r0 *1 80.655,72.59
X$148 17 VIA_via2_5
* cell instance $149 r0 *1 70.205,2.31
X$149 17 VIA_via2_5
* cell instance $150 r0 *1 70.585,50.75
X$150 17 VIA_via2_5
* cell instance $151 r0 *1 69.635,50.75
X$151 17 VIA_via2_5
* cell instance $152 r0 *1 81.225,45.43
X$152 17 VIA_via2_5
* cell instance $153 r0 *1 81.225,43.75
X$153 17 VIA_via2_5
* cell instance $154 r0 *1 77.805,34.23
X$154 17 VIA_via2_5
* cell instance $155 r0 *1 77.995,34.09
X$155 17 VIA_via2_5
* cell instance $156 r0 *1 75.715,43.75
X$156 17 VIA_via2_5
* cell instance $157 r0 *1 77.805,37.03
X$157 17 VIA_via2_5
* cell instance $158 r0 *1 75.715,42.77
X$158 17 VIA_via2_5
* cell instance $159 r0 *1 82.365,16.03
X$159 17 VIA_via1_4
* cell instance $160 r0 *1 82.27,15.4
X$160 377 17 378 23 38 409 MUX2_X1
* cell instance $161 r0 *1 82.365,16.03
X$161 17 VIA_via2_5
* cell instance $162 r0 *1 69.635,42.77
X$162 17 VIA_via1_4
* cell instance $163 m0 *1 69.54,43.4
X$163 675 17 1040 23 38 1090 MUX2_X1
* cell instance $164 r0 *1 69.635,42.77
X$164 17 VIA_via2_5
* cell instance $165 r0 *1 66.025,55.65
X$165 17 VIA_via1_4
* cell instance $166 r0 *1 64.98,54.6
X$166 821 38 17 23 BUF_X4
* cell instance $167 r0 *1 66.025,55.79
X$167 17 VIA_via2_5
* cell instance $168 r0 *1 67.855,72.59
X$168 17 VIA_via3_2
* cell instance $169 r0 *1 67.855,58.31
X$169 17 VIA_via3_2
* cell instance $170 r0 *1 67.855,55.79
X$170 17 VIA_via3_2
* cell instance $171 r0 *1 12.065,11.97
X$171 18 VIA_via2_5
* cell instance $172 r0 *1 11.305,6.37
X$172 18 VIA_via2_5
* cell instance $173 r0 *1 10.735,6.37
X$173 18 VIA_via2_5
* cell instance $174 r0 *1 11.115,11.97
X$174 18 VIA_via2_5
* cell instance $175 r0 *1 11.495,2.03
X$175 18 VIA_via2_5
* cell instance $176 r0 *1 5.035,11.97
X$176 18 VIA_via2_5
* cell instance $177 r0 *1 10.735,8.75
X$177 18 VIA_via1_4
* cell instance $178 m0 *1 10.26,9.8
X$178 149 23 38 18 CLKBUF_X3
* cell instance $179 r0 *1 11.115,9.59
X$179 18 VIA_via1_7
* cell instance $180 r0 *1 11.305,9.17
X$180 18 VIA_via1_4
* cell instance $181 m0 *1 11.21,9.8
X$181 18 23 38 3143 INV_X1
* cell instance $182 r0 *1 9.785,11.97
X$182 18 VIA_via1_4
* cell instance $183 m0 *1 8.17,12.6
X$183 23 2784 201 200 18 38 DFF_X1
* cell instance $184 r0 *1 9.785,11.97
X$184 18 VIA_via2_5
* cell instance $185 r0 *1 11.495,3.57
X$185 18 VIA_via1_4
* cell instance $186 m0 *1 9.88,4.2
X$186 23 2738 69 55 18 38 DFF_X1
* cell instance $187 r0 *1 13.775,2.03
X$187 18 VIA_via1_4
* cell instance $188 r0 *1 12.16,1.4
X$188 23 3043 56 19 18 38 DFF_X1
* cell instance $189 r0 *1 13.775,2.03
X$189 18 VIA_via2_5
* cell instance $190 r0 *1 9.215,6.37
X$190 18 VIA_via1_4
* cell instance $191 m0 *1 7.6,7
X$191 23 2754 106 129 18 38 DFF_X1
* cell instance $192 r0 *1 9.215,6.37
X$192 18 VIA_via2_5
* cell instance $193 r0 *1 12.255,13.23
X$193 18 VIA_via1_4
* cell instance $194 r0 *1 10.64,12.6
X$194 23 3045 246 269 18 38 DFF_X1
* cell instance $195 r0 *1 5.035,13.23
X$195 18 VIA_via1_4
* cell instance $196 r0 *1 3.42,12.6
X$196 23 3038 294 268 18 38 DFF_X1
* cell instance $197 r0 *1 14.725,3.01
X$197 19 VIA_via1_7
* cell instance $198 m0 *1 13.49,4.2
X$198 27 40 56 23 38 19 MUX2_X1
* cell instance $199 r0 *1 14.725,1.89
X$199 19 VIA_via2_5
* cell instance $200 r0 *1 13.015,2.03
X$200 19 VIA_via1_4
* cell instance $201 r0 *1 13.015,1.89
X$201 19 VIA_via2_5
* cell instance $202 r0 *1 80.845,2.17
X$202 20 VIA_via1_4
* cell instance $203 r0 *1 80.845,2.17
X$203 20 VIA_via2_5
* cell instance $204 r0 *1 76.855,2.03
X$204 20 VIA_via1_4
* cell instance $205 r0 *1 76.855,2.17
X$205 20 VIA_via2_5
* cell instance $206 r0 *1 25.745,2.03
X$206 21 VIA_via2_5
* cell instance $207 r0 *1 25.935,6.37
X$207 21 VIA_via1_4
* cell instance $208 m0 *1 25.65,7
X$208 21 70 115 23 38 95 MUX2_X1
* cell instance $209 r0 *1 27.645,2.03
X$209 21 VIA_via1_4
* cell instance $210 r0 *1 27.645,2.03
X$210 21 VIA_via2_5
* cell instance $211 r0 *1 25.745,3.57
X$211 21 VIA_via1_4
* cell instance $212 m0 *1 24.89,4.2
X$212 26 42 21 23 38 39 MUX2_X1
* cell instance $213 r0 *1 69.445,3.01
X$213 22 VIA_via1_7
* cell instance $214 r0 *1 69.445,2.03
X$214 22 VIA_via2_5
* cell instance $215 r0 *1 68.495,2.03
X$215 22 VIA_via1_4
* cell instance $216 r0 *1 68.495,2.03
X$216 22 VIA_via2_5
* cell instance $217 m0 *1 28.88,74.2
X$217 1905 1927 1511 1787 38 23 1928 OAI22_X2
* cell instance $218 m0 *1 28.69,74.2
X$218 23 38 FILLCELL_X1
* cell instance $219 m0 *1 30.59,74.2
X$219 1905 1927 1629 1157 1727 38 23 1906 OAI221_X1
* cell instance $220 m0 *1 31.73,74.2
X$220 23 38 FILLCELL_X4
* cell instance $221 m0 *1 32.49,74.2
X$221 1823 1728 23 38 1908 NAND2_X1
* cell instance $222 m0 *1 33.06,74.2
X$222 23 38 FILLCELL_X2
* cell instance $223 r0 *1 28.69,74.2
X$223 1971 1972 1629 1157 1727 38 23 1942 OAI221_X1
* cell instance $224 r0 *1 29.83,74.2
X$224 1636 1963 23 38 1907 NAND2_X1
* cell instance $225 r0 *1 30.4,74.2
X$225 23 38 FILLCELL_X4
* cell instance $226 r0 *1 31.16,74.2
X$226 1743 1907 1942 1804 1943 38 23 2038 OAI221_X1
* cell instance $227 r0 *1 32.3,74.2
X$227 1928 1765 1908 38 23 1973 OAI21_X2
* cell instance $228 m0 *1 33.63,74.2
X$228 1909 23 38 1795 CLKBUF_X3
* cell instance $229 m0 *1 33.44,74.2
X$229 23 38 FILLCELL_X1
* cell instance $230 m0 *1 34.58,74.2
X$230 23 38 FILLCELL_X16
* cell instance $231 m0 *1 37.62,74.2
X$231 23 38 FILLCELL_X8
* cell instance $232 m0 *1 39.14,74.2
X$232 23 2618 1912 1930 1933 38 DFF_X1
* cell instance $233 m0 *1 42.37,74.2
X$233 1912 1184 1964 23 38 1932 MUX2_X1
* cell instance $234 m0 *1 43.7,74.2
X$234 23 38 FILLCELL_X8
* cell instance $235 m0 *1 45.22,74.2
X$235 23 38 FILLCELL_X2
* cell instance $236 r0 *1 33.63,74.2
X$236 1963 1638 23 38 1943 NAND2_X1
* cell instance $237 r0 *1 34.2,74.2
X$237 23 3055 1944 1966 1933 38 DFF_X1
* cell instance $238 r0 *1 37.43,74.2
X$238 1636 1944 23 38 1999 NAND2_X1
* cell instance $239 r0 *1 38,74.2
X$239 23 38 FILLCELL_X4
* cell instance $240 r0 *1 38.76,74.2
X$240 23 38 FILLCELL_X2
* cell instance $241 r0 *1 39.14,74.2
X$241 23 3062 1964 1965 1933 38 DFF_X1
* cell instance $242 r0 *1 42.37,74.2
X$242 1636 1945 23 38 1975 NAND2_X1
* cell instance $243 r0 *1 42.94,74.2
X$243 1945 1638 23 38 2042 NAND2_X1
* cell instance $244 r0 *1 43.51,74.2
X$244 1964 1434 1813 23 38 1965 MUX2_X1
* cell instance $245 r0 *1 44.84,74.2
X$245 23 38 FILLCELL_X4
* cell instance $246 r0 *1 45.6,74.2
X$246 23 38 FILLCELL_X1
* cell instance $247 m0 *1 45.79,74.2
X$247 23 2701 1961 1962 1933 38 DFF_X1
* cell instance $248 m0 *1 45.6,74.2
X$248 23 38 FILLCELL_X1
* cell instance $249 m0 *1 49.02,74.2
X$249 23 38 FILLCELL_X16
* cell instance $250 m0 *1 52.06,74.2
X$250 23 38 FILLCELL_X8
* cell instance $251 m0 *1 53.58,74.2
X$251 23 2853 1948 1958 1960 38 DFF_X1
* cell instance $252 m0 *1 56.81,74.2
X$252 23 38 FILLCELL_X16
* cell instance $253 m0 *1 59.85,74.2
X$253 23 38 FILLCELL_X4
* cell instance $254 m0 *1 60.61,74.2
X$254 23 38 FILLCELL_X2
* cell instance $255 r0 *1 45.79,74.2
X$255 1932 1177 23 38 1996 NOR2_X1
* cell instance $256 r0 *1 46.36,74.2
X$256 23 38 FILLCELL_X4
* cell instance $257 r0 *1 47.12,74.2
X$257 23 38 FILLCELL_X1
* cell instance $258 r0 *1 47.31,74.2
X$258 1813 1492 1961 23 38 1962 MUX2_X1
* cell instance $259 r0 *1 48.64,74.2
X$259 1961 414 1946 23 38 1994 MUX2_X1
* cell instance $260 r0 *1 49.97,74.2
X$260 23 38 FILLCELL_X2
* cell instance $261 r0 *1 50.35,74.2
X$261 23 38 FILLCELL_X1
* cell instance $262 r0 *1 50.54,74.2
X$262 23 2876 1977 1993 1960 38 DFF_X1
* cell instance $263 r0 *1 53.77,74.2
X$263 1485 1879 1934 1142 1956 1978 23 38 1947 OAI33_X1
* cell instance $264 r0 *1 55.1,74.2
X$264 23 38 FILLCELL_X2
* cell instance $265 r0 *1 55.48,74.2
X$265 1743 1989 1990 1804 1957 38 23 1958 OAI221_X1
* cell instance $266 r0 *1 56.62,74.2
X$266 23 38 FILLCELL_X1
* cell instance $267 r0 *1 56.81,74.2
X$267 1948 1638 23 38 1957 NAND2_X1
* cell instance $268 r0 *1 57.38,74.2
X$268 1979 414 2020 23 38 1987 MUX2_X1
* cell instance $269 r0 *1 58.71,74.2
X$269 23 38 FILLCELL_X2
* cell instance $270 r0 *1 59.14,74.2
X$270 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $271 r0 *1 59.14,74.2
X$271 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $272 r0 *1 59.14,74.2
X$272 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $273 r0 *1 59.09,74.2
X$273 23 38 FILLCELL_X1
* cell instance $274 r0 *1 59.28,74.2
X$274 1198 23 38 1787 CLKBUF_X3
* cell instance $275 r0 *1 60.23,74.2
X$275 23 38 FILLCELL_X8
* cell instance $276 m0 *1 61.18,74.2
X$276 1880 373 1561 23 38 1901 MUX2_X1
* cell instance $277 m0 *1 60.99,74.2
X$277 23 38 FILLCELL_X1
* cell instance $278 m0 *1 62.51,74.2
X$278 23 38 FILLCELL_X4
* cell instance $279 m0 *1 63.27,74.2
X$279 23 38 FILLCELL_X2
* cell instance $280 r0 *1 61.75,74.2
X$280 1951 23 38 1157 CLKBUF_X3
* cell instance $281 r0 *1 62.7,74.2
X$281 23 38 FILLCELL_X16
* cell instance $282 m0 *1 66.88,74.2
X$282 1913 1099 1914 23 38 1897 MUX2_X1
* cell instance $283 m0 *1 63.65,74.2
X$283 23 2834 1913 1931 1915 38 DFF_X1
* cell instance $284 m0 *1 68.21,74.2
X$284 23 38 FILLCELL_X2
* cell instance $285 r0 *1 65.74,74.2
X$285 23 38 FILLCELL_X2
* cell instance $286 r0 *1 66.12,74.2
X$286 1686 23 38 1727 CLKBUF_X3
* cell instance $287 r0 *1 67.07,74.2
X$287 23 38 FILLCELL_X16
* cell instance $288 m0 *1 71.82,74.2
X$288 23 38 FILLCELL_X2
* cell instance $289 m0 *1 68.59,74.2
X$289 23 2835 1914 1896 1915 38 DFF_X1
* cell instance $290 r0 *1 70.11,74.2
X$290 1594 23 38 1206 CLKBUF_X3
* cell instance $291 r0 *1 71.06,74.2
X$291 23 38 FILLCELL_X8
* cell instance $292 m0 *1 75.43,74.2
X$292 1829 441 1770 23 38 1929 MUX2_X1
* cell instance $293 m0 *1 72.2,74.2
X$293 23 2850 1829 1929 1648 38 DFF_X1
* cell instance $294 m0 *1 76.76,74.2
X$294 23 38 FILLCELL_X4
* cell instance $295 m0 *1 77.52,74.2
X$295 23 38 FILLCELL_X2
* cell instance $296 r0 *1 72.58,74.2
X$296 23 38 FILLCELL_X4
* cell instance $297 r0 *1 73.34,74.2
X$297 23 38 FILLCELL_X1
* cell instance $298 r0 *1 73.53,74.2
X$298 1953 23 38 1594 INV_X8
* cell instance $299 r0 *1 75.24,74.2
X$299 23 1594 1331 38 BUF_X32
* cell instance $300 m0 *1 81.13,74.2
X$300 23 2836 1916 1886 1917 38 DFF_X1
* cell instance $301 m0 *1 77.9,74.2
X$301 23 2838 1885 1884 1917 38 DFF_X1
* cell instance $302 m0 *1 84.36,74.2
X$302 23 38 FILLCELL_X8
* cell instance $303 m0 *1 85.88,74.2
X$303 23 38 FILLCELL_X2
* cell instance $304 r0 *1 84.55,74.2
X$304 1951 23 38 1506 CLKBUF_X3
* cell instance $305 r0 *1 85.5,74.2
X$305 23 38 FILLCELL_X2
* cell instance $306 r0 *1 85.88,74.2
X$306 1949 23 38 1804 CLKBUF_X3
* cell instance $307 m0 *1 86.45,74.2
X$307 1230 23 38 1918 INV_X1
* cell instance $308 m0 *1 86.26,74.2
X$308 23 38 FILLCELL_X1
* cell instance $309 m0 *1 86.83,74.2
X$309 23 2832 1920 1919 1917 38 DFF_X1
* cell instance $310 m0 *1 90.06,74.2
X$310 23 1743 38 1332 BUF_X8
* cell instance $311 m0 *1 92.53,74.2
X$311 23 38 FILLCELL_X16
* cell instance $312 m0 *1 95.57,74.2
X$312 23 38 FILLCELL_X8
* cell instance $313 r180 *1 97.28,74.2
X$313 23 38 23 38 TAPCELL_X1
* cell instance $314 r0 *1 86.83,74.2
X$314 1226 1918 1984 23 1919 38 AOI21_X1
* cell instance $315 r0 *1 87.59,74.2
X$315 1949 23 38 1226 CLKBUF_X3
* cell instance $316 r0 *1 88.54,74.2
X$316 23 38 FILLCELL_X16
* cell instance $317 r0 *1 91.58,74.2
X$317 23 38 FILLCELL_X8
* cell instance $318 r0 *1 93.1,74.2
X$318 23 38 FILLCELL_X2
* cell instance $319 r0 *1 93.48,74.2
X$319 23 3104 1985 1986 2026 38 DFF_X1
* cell instance $320 r0 *1 96.71,74.2
X$320 23 38 FILLCELL_X2
* cell instance $321 m90 *1 97.28,74.2
X$321 23 38 23 38 TAPCELL_X1
* cell instance $322 m0 *1 16.53,37.8
X$322 875 831 23 38 970 NOR2_X1
* cell instance $323 m0 *1 15.96,37.8
X$323 873 831 23 38 917 NOR2_X1
* cell instance $324 m0 *1 17.1,37.8
X$324 871 831 23 38 918 NOR2_X1
* cell instance $325 m0 *1 17.67,37.8
X$325 857 829 23 38 877 NOR2_X1
* cell instance $326 m0 *1 18.24,37.8
X$326 23 38 FILLCELL_X2
* cell instance $327 r0 *1 15.96,37.8
X$327 967 937 23 38 920 NOR2_X1
* cell instance $328 r0 *1 16.53,37.8
X$328 915 831 23 38 931 NOR2_X1
* cell instance $329 r0 *1 17.1,37.8
X$329 932 920 888 891 917 889 23 38 890 OAI33_X1
* cell instance $330 r0 *1 18.43,37.8
X$330 23 38 FILLCELL_X2
* cell instance $331 m0 *1 19.19,37.8
X$331 878 829 23 38 892 NOR2_X1
* cell instance $332 m0 *1 18.62,37.8
X$332 827 829 23 38 922 NOR2_X1
* cell instance $333 m0 *1 19.76,37.8
X$333 23 38 FILLCELL_X8
* cell instance $334 m0 *1 21.28,37.8
X$334 23 2695 894 924 763 38 DFF_X1
* cell instance $335 m0 *1 24.51,37.8
X$335 23 38 FILLCELL_X4
* cell instance $336 m0 *1 25.27,37.8
X$336 23 38 FILLCELL_X2
* cell instance $337 r0 *1 18.81,37.8
X$337 23 38 FILLCELL_X1
* cell instance $338 r0 *1 19,37.8
X$338 933 893 23 38 972 NOR2_X1
* cell instance $339 r0 *1 19.57,37.8
X$339 23 38 FILLCELL_X8
* cell instance $340 r0 *1 21.09,37.8
X$340 23 38 FILLCELL_X2
* cell instance $341 r0 *1 21.47,37.8
X$341 23 38 FILLCELL_X1
* cell instance $342 r0 *1 21.66,37.8
X$342 894 929 358 23 38 924 MUX2_X1
* cell instance $343 r0 *1 22.99,37.8
X$343 851 900 894 23 38 973 MUX2_X1
* cell instance $344 r0 *1 24.32,37.8
X$344 973 893 23 38 975 NOR2_X1
* cell instance $345 r0 *1 24.89,37.8
X$345 23 38 FILLCELL_X4
* cell instance $346 r0 *1 25.65,37.8
X$346 932 935 975 891 896 895 23 38 897 OAI33_X1
* cell instance $347 m0 *1 25.84,37.8
X$347 698 829 23 38 895 NOR2_X1
* cell instance $348 m0 *1 25.65,37.8
X$348 23 38 FILLCELL_X1
* cell instance $349 m0 *1 26.41,37.8
X$349 23 38 FILLCELL_X2
* cell instance $350 m0 *1 27.36,37.8
X$350 898 858 421 23 38 880 MUX2_X1
* cell instance $351 m0 *1 26.79,37.8
X$351 852 831 23 38 896 NOR2_X1
* cell instance $352 m0 *1 28.69,37.8
X$352 23 2848 898 880 763 38 DFF_X1
* cell instance $353 m0 *1 31.92,37.8
X$353 23 38 FILLCELL_X16
* cell instance $354 m0 *1 34.96,37.8
X$354 23 2697 947 926 942 38 DFF_X1
* cell instance $355 m0 *1 38.19,37.8
X$355 23 38 FILLCELL_X8
* cell instance $356 m0 *1 39.71,37.8
X$356 23 2837 834 860 636 38 DFF_X1
* cell instance $357 m0 *1 42.94,37.8
X$357 23 38 FILLCELL_X4
* cell instance $358 m0 *1 43.7,37.8
X$358 23 38 FILLCELL_X1
* cell instance $359 m0 *1 43.89,37.8
X$359 834 900 836 23 38 885 MUX2_X1
* cell instance $360 m0 *1 45.22,37.8
X$360 23 38 FILLCELL_X2
* cell instance $361 r0 *1 26.98,37.8
X$361 23 38 FILLCELL_X1
* cell instance $362 r0 *1 27.17,37.8
X$362 939 929 421 23 38 938 MUX2_X1
* cell instance $363 r0 *1 28.5,37.8
X$363 23 38 FILLCELL_X2
* cell instance $364 r0 *1 28.88,37.8
X$364 898 900 939 23 38 940 MUX2_X1
* cell instance $365 r0 *1 30.21,37.8
X$365 23 38 FILLCELL_X4
* cell instance $366 r0 *1 30.97,37.8
X$366 23 38 FILLCELL_X1
* cell instance $367 r0 *1 31.16,37.8
X$367 943 941 510 23 38 1019 MUX2_X1
* cell instance $368 r0 *1 32.49,37.8
X$368 945 992 510 23 38 944 MUX2_X1
* cell instance $369 r0 *1 33.82,37.8
X$369 23 38 FILLCELL_X2
* cell instance $370 r0 *1 34.2,37.8
X$370 947 929 510 23 38 926 MUX2_X1
* cell instance $371 r0 *1 35.53,37.8
X$371 899 858 510 23 38 980 MUX2_X1
* cell instance $372 r0 *1 36.86,37.8
X$372 899 900 947 23 38 948 MUX2_X1
* cell instance $373 r0 *1 38.19,37.8
X$373 23 38 FILLCELL_X2
* cell instance $374 r0 *1 38.57,37.8
X$374 23 38 FILLCELL_X1
* cell instance $375 r0 *1 38.76,37.8
X$375 23 2961 899 980 636 38 DFF_X1
* cell instance $376 r0 *1 41.99,37.8
X$376 23 38 FILLCELL_X8
* cell instance $377 r0 *1 43.51,37.8
X$377 836 929 398 23 38 835 MUX2_X1
* cell instance $378 r0 *1 44.84,37.8
X$378 23 38 FILLCELL_X1
* cell instance $379 r0 *1 45.03,37.8
X$379 932 982 927 891 983 837 23 38 901 OAI33_X1
* cell instance $380 m0 *1 46.17,37.8
X$380 23 38 FILLCELL_X8
* cell instance $381 m0 *1 45.6,37.8
X$381 885 840 23 38 927 NOR2_X1
* cell instance $382 m0 *1 47.69,37.8
X$382 23 38 FILLCELL_X1
* cell instance $383 m0 *1 47.88,37.8
X$383 770 190 23 38 983 NOR2_X1
* cell instance $384 m0 *1 48.45,37.8
X$384 23 38 FILLCELL_X2
* cell instance $385 r0 *1 46.36,37.8
X$385 23 38 FILLCELL_X1
* cell instance $386 r0 *1 46.55,37.8
X$386 984 929 301 23 38 986 MUX2_X1
* cell instance $387 r0 *1 47.88,37.8
X$387 23 3124 984 986 839 38 DFF_X1
* cell instance $388 m0 *1 49.78,37.8
X$388 23 38 FILLCELL_X8
* cell instance $389 m0 *1 48.83,37.8
X$389 863 23 38 762 CLKBUF_X3
* cell instance $390 m0 *1 51.3,37.8
X$390 23 38 FILLCELL_X4
* cell instance $391 m0 *1 52.06,37.8
X$391 795 190 23 38 903 NOR2_X1
* cell instance $392 m0 *1 52.63,37.8
X$392 744 23 38 839 CLKBUF_X3
* cell instance $393 m0 *1 53.58,37.8
X$393 556 863 904 23 38 985 MUX2_X1
* cell instance $394 m0 *1 54.91,37.8
X$394 23 2821 905 886 839 38 DFF_X1
* cell instance $395 m0 *1 58.14,37.8
X$395 23 2820 856 884 839 38 DFF_X1
* cell instance $396 m0 *1 61.37,37.8
X$396 620 38 438 23 BUF_X4
* cell instance $397 m0 *1 62.7,37.8
X$397 23 38 FILLCELL_X1
* cell instance $398 m0 *1 62.89,37.8
X$398 599 38 174 23 BUF_X4
* cell instance $399 m0 *1 64.22,37.8
X$399 23 38 FILLCELL_X32
* cell instance $400 m0 *1 70.3,37.8
X$400 23 38 FILLCELL_X4
* cell instance $401 m0 *1 71.06,37.8
X$401 800 438 866 23 38 883 MUX2_X1
* cell instance $402 m0 *1 72.39,37.8
X$402 23 2710 866 921 801 38 DFF_X1
* cell instance $403 m0 *1 76.95,37.8
X$403 23 38 FILLCELL_X2
* cell instance $404 r0 *1 51.11,37.8
X$404 1027 840 23 38 987 NOR2_X1
* cell instance $405 r0 *1 51.68,37.8
X$405 932 902 987 891 903 861 23 38 925 OAI33_X1
* cell instance $406 r0 *1 53.01,37.8
X$406 23 38 FILLCELL_X2
* cell instance $407 r0 *1 53.39,37.8
X$407 23 2873 904 985 839 38 DFF_X1
* cell instance $408 r0 *1 56.62,37.8
X$408 904 144 905 23 38 950 MUX2_X1
* cell instance $409 r0 *1 57.95,37.8
X$409 23 38 FILLCELL_X4
* cell instance $410 r0 *1 58.71,37.8
X$410 23 38 FILLCELL_X2
* cell instance $411 r0 *1 59.14,37.8
X$411 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $412 r0 *1 59.14,37.8
X$412 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $413 r0 *1 59.14,37.8
X$413 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $414 r0 *1 59.09,37.8
X$414 640 863 951 23 38 952 MUX2_X1
* cell instance $415 r0 *1 60.42,37.8
X$415 951 144 856 23 38 953 MUX2_X1
* cell instance $416 r0 *1 61.75,37.8
X$416 23 38 FILLCELL_X4
* cell instance $417 r0 *1 62.51,37.8
X$417 23 38 FILLCELL_X2
* cell instance $418 r0 *1 62.89,37.8
X$418 23 38 FILLCELL_X1
* cell instance $419 r0 *1 63.08,37.8
X$419 23 2868 906 923 954 38 DFF_X1
* cell instance $420 r0 *1 66.31,37.8
X$420 906 520 799 23 38 923 MUX2_X1
* cell instance $421 r0 *1 67.64,37.8
X$421 23 38 FILLCELL_X16
* cell instance $422 r0 *1 70.68,37.8
X$422 23 38 FILLCELL_X8
* cell instance $423 r0 *1 72.2,37.8
X$423 862 38 263 23 BUF_X4
* cell instance $424 r0 *1 73.53,37.8
X$424 23 38 FILLCELL_X8
* cell instance $425 r0 *1 75.05,37.8
X$425 23 38 FILLCELL_X4
* cell instance $426 r0 *1 75.81,37.8
X$426 23 38 FILLCELL_X1
* cell instance $427 r0 *1 76,37.8
X$427 974 88 907 23 38 976 MUX2_X1
* cell instance $428 r0 *1 77.33,37.8
X$428 744 23 38 801 CLKBUF_X3
* cell instance $429 m0 *1 77.52,37.8
X$429 919 881 23 38 882 NOR2_X1
* cell instance $430 m0 *1 77.33,37.8
X$430 23 38 FILLCELL_X1
* cell instance $431 m0 *1 78.09,37.8
X$431 868 862 867 23 38 919 MUX2_X1
* cell instance $432 m0 *1 79.42,37.8
X$432 23 38 FILLCELL_X2
* cell instance $433 r0 *1 78.28,37.8
X$433 23 38 FILLCELL_X8
* cell instance $434 m0 *1 81.13,37.8
X$434 23 38 FILLCELL_X8
* cell instance $435 m0 *1 79.8,37.8
X$435 710 79 867 23 38 908 MUX2_X1
* cell instance $436 m0 *1 82.65,37.8
X$436 23 38 FILLCELL_X2
* cell instance $437 r0 *1 79.8,37.8
X$437 23 2929 867 908 801 38 DFF_X1
* cell instance $438 m0 *1 84.36,37.8
X$438 23 38 FILLCELL_X8
* cell instance $439 m0 *1 83.03,37.8
X$439 710 133 868 23 38 909 MUX2_X1
* cell instance $440 m0 *1 85.88,37.8
X$440 23 38 FILLCELL_X2
* cell instance $441 r0 *1 83.03,37.8
X$441 23 2883 868 909 1042 38 DFF_X1
* cell instance $442 r0 *1 86.26,37.8
X$442 910 174 907 23 38 869 MUX2_X1
* cell instance $443 m0 *1 89.49,37.8
X$443 23 38 FILLCELL_X4
* cell instance $444 m0 *1 86.26,37.8
X$444 23 2842 910 869 876 38 DFF_X1
* cell instance $445 m0 *1 90.25,37.8
X$445 23 38 FILLCELL_X1
* cell instance $446 m0 *1 90.44,37.8
X$446 912 261 23 38 913 NOR2_X1
* cell instance $447 m0 *1 91.01,37.8
X$447 23 38 FILLCELL_X4
* cell instance $448 m0 *1 91.77,37.8
X$448 23 38 FILLCELL_X2
* cell instance $449 r0 *1 87.59,37.8
X$449 911 223 907 23 38 956 MUX2_X1
* cell instance $450 r0 *1 88.92,37.8
X$450 23 38 FILLCELL_X2
* cell instance $451 r0 *1 89.3,37.8
X$451 23 38 FILLCELL_X1
* cell instance $452 r0 *1 89.49,37.8
X$452 911 188 910 23 38 912 MUX2_X1
* cell instance $453 r0 *1 90.82,37.8
X$453 227 913 966 225 963 964 23 38 914 OAI33_X1
* cell instance $454 r0 *1 92.15,37.8
X$454 23 38 FILLCELL_X2
* cell instance $455 m0 *1 92.72,37.8
X$455 23 38 FILLCELL_X16
* cell instance $456 m0 *1 92.15,37.8
X$456 872 177 23 38 964 NOR2_X1
* cell instance $457 m0 *1 95.76,37.8
X$457 23 38 FILLCELL_X4
* cell instance $458 m0 *1 96.52,37.8
X$458 23 38 FILLCELL_X2
* cell instance $459 r0 *1 92.53,37.8
X$459 957 274 23 38 963 NOR2_X1
* cell instance $460 r0 *1 93.1,37.8
X$460 23 38 FILLCELL_X2
* cell instance $461 r0 *1 93.48,37.8
X$461 23 2902 958 959 876 38 DFF_X1
* cell instance $462 r0 *1 96.71,37.8
X$462 23 38 FILLCELL_X2
* cell instance $463 r180 *1 97.28,37.8
X$463 23 38 23 38 TAPCELL_X1
* cell instance $464 m0 *1 96.9,37.8
X$464 23 38 FILLCELL_X1
* cell instance $465 m90 *1 97.28,37.8
X$465 23 38 23 38 TAPCELL_X1
* cell instance $466 m0 *1 7.98,60.2
X$466 1486 23 38 1292 CLKBUF_X3
* cell instance $467 m0 *1 4.75,60.2
X$467 23 2611 1481 1571 1292 38 DFF_X1
* cell instance $468 m0 *1 8.93,60.2
X$468 23 2613 1507 1545 1292 38 DFF_X1
* cell instance $469 m0 *1 12.16,60.2
X$469 1598 1530 1531 23 38 1574 MUX2_X1
* cell instance $470 m0 *1 13.49,60.2
X$470 23 2594 1531 1574 1326 38 DFF_X1
* cell instance $471 m0 *1 16.72,60.2
X$471 1532 1492 1533 23 38 1546 MUX2_X1
* cell instance $472 m0 *1 18.05,60.2
X$472 1533 792 1531 23 38 1575 MUX2_X1
* cell instance $473 m0 *1 19.38,60.2
X$473 23 38 FILLCELL_X8
* cell instance $474 m0 *1 20.9,60.2
X$474 23 38 FILLCELL_X1
* cell instance $475 m0 *1 21.09,60.2
X$475 1486 23 38 1399 CLKBUF_X3
* cell instance $476 m0 *1 22.04,60.2
X$476 1399 23 38 CLKBUF_X1
* cell instance $477 m0 *1 22.61,60.2
X$477 1575 829 23 38 1625 NOR2_X1
* cell instance $478 m0 *1 23.18,60.2
X$478 23 38 FILLCELL_X4
* cell instance $479 m0 *1 23.94,60.2
X$479 23 38 FILLCELL_X2
* cell instance $480 m0 *1 1.33,60.2
X$480 23 38 FILLCELL_X16
* cell instance $481 m0 *1 1.14,60.2
X$481 23 38 23 38 TAPCELL_X1
* cell instance $482 m0 *1 4.37,60.2
X$482 23 38 FILLCELL_X2
* cell instance $483 r0 *1 1.14,60.2
X$483 23 38 23 38 TAPCELL_X1
* cell instance $484 r0 *1 1.33,60.2
X$484 23 38 FILLCELL_X4
* cell instance $485 r0 *1 2.09,60.2
X$485 23 38 FILLCELL_X2
* cell instance $486 r0 *1 2.47,60.2
X$486 23 38 FILLCELL_X1
* cell instance $487 r0 *1 2.66,60.2
X$487 1555 23 38 1598 BUF_X1
* cell instance $488 r0 *1 3.14,60.2
X$488 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $489 r0 *1 3.14,60.2
X$489 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $490 r0 *1 3.14,60.2
X$490 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $491 r0 *1 3.23,60.2
X$491 23 2946 1654 1614 1556 38 DFF_X1
* cell instance $492 r0 *1 6.46,60.2
X$492 23 38 FILLCELL_X8
* cell instance $493 r0 *1 7.98,60.2
X$493 23 38 FILLCELL_X4
* cell instance $494 r0 *1 8.74,60.2
X$494 23 38 FILLCELL_X2
* cell instance $495 r0 *1 9.12,60.2
X$495 23 2954 1599 1618 1292 38 DFF_X1
* cell instance $496 r0 *1 12.35,60.2
X$496 23 38 FILLCELL_X16
* cell instance $497 r0 *1 15.39,60.2
X$497 23 38 FILLCELL_X8
* cell instance $498 r0 *1 16.91,60.2
X$498 23 38 FILLCELL_X1
* cell instance $499 r0 *1 17.1,60.2
X$499 23 2944 1600 1622 1399 38 DFF_X1
* cell instance $500 r0 *1 20.33,60.2
X$500 23 38 FILLCELL_X8
* cell instance $501 r0 *1 21.85,60.2
X$501 1576 937 23 38 1626 NOR2_X1
* cell instance $502 r0 *1 22.42,60.2
X$502 23 38 FILLCELL_X4
* cell instance $503 r0 *1 23.18,60.2
X$503 23 38 FILLCELL_X1
* cell instance $504 r0 *1 23.37,60.2
X$504 1601 994 1666 23 38 1576 MUX2_X1
* cell instance $505 m0 *1 27.55,60.2
X$505 23 38 FILLCELL_X8
* cell instance $506 m0 *1 24.32,60.2
X$506 23 2630 1534 1547 1399 38 DFF_X1
* cell instance $507 m0 *1 29.07,60.2
X$507 23 38 FILLCELL_X1
* cell instance $508 m0 *1 29.26,60.2
X$508 1513 1426 1629 1157 1139 38 23 1604 OAI221_X1
* cell instance $509 m0 *1 30.4,60.2
X$509 23 38 FILLCELL_X4
* cell instance $510 m0 *1 31.16,60.2
X$510 988 23 38 893 CLKBUF_X3
* cell instance $511 m0 *1 32.11,60.2
X$511 23 38 FILLCELL_X4
* cell instance $512 m0 *1 32.87,60.2
X$512 23 38 FILLCELL_X1
* cell instance $513 m0 *1 33.06,60.2
X$513 403 23 38 937 CLKBUF_X3
* cell instance $514 m0 *1 34.01,60.2
X$514 403 38 1537 23 BUF_X4
* cell instance $515 m0 *1 35.34,60.2
X$515 23 38 FILLCELL_X2
* cell instance $516 r0 *1 24.7,60.2
X$516 23 38 FILLCELL_X16
* cell instance $517 r0 *1 27.74,60.2
X$517 23 38 FILLCELL_X4
* cell instance $518 r0 *1 28.5,60.2
X$518 23 38 FILLCELL_X1
* cell instance $519 r0 *1 28.69,60.2
X$519 23 2989 1450 1603 1262 38 DFF_X1
* cell instance $520 r0 *1 31.92,60.2
X$520 23 38 FILLCELL_X32
* cell instance $521 m0 *1 37.05,60.2
X$521 23 38 FILLCELL_X2
* cell instance $522 m0 *1 35.72,60.2
X$522 403 38 1579 23 BUF_X4
* cell instance $523 m0 *1 38.38,60.2
X$523 840 38 1535 23 BUF_X4
* cell instance $524 m0 *1 37.43,60.2
X$524 988 23 38 831 CLKBUF_X3
* cell instance $525 m0 *1 39.71,60.2
X$525 1583 1487 1490 23 38 1549 MUX2_X1
* cell instance $526 m0 *1 41.04,60.2
X$526 23 38 FILLCELL_X4
* cell instance $527 m0 *1 41.8,60.2
X$527 23 38 FILLCELL_X1
* cell instance $528 m0 *1 41.99,60.2
X$528 1583 1454 1489 23 38 1585 MUX2_X1
* cell instance $529 m0 *1 43.32,60.2
X$529 23 38 FILLCELL_X1
* cell instance $530 m0 *1 43.51,60.2
X$530 1585 1105 23 38 1550 NOR2_X1
* cell instance $531 m0 *1 44.08,60.2
X$531 1298 1140 23 38 1552 NAND2_X1
* cell instance $532 m0 *1 44.65,60.2
X$532 23 2793 1536 1554 1404 38 DFF_X1
* cell instance $533 m0 *1 47.88,60.2
X$533 23 38 FILLCELL_X1
* cell instance $534 m0 *1 48.07,60.2
X$534 1175 38 1487 23 BUF_X4
* cell instance $535 m0 *1 49.4,60.2
X$535 23 2566 1525 1553 1404 38 DFF_X1
* cell instance $536 m0 *1 52.63,60.2
X$536 23 38 FILLCELL_X2
* cell instance $537 r0 *1 38,60.2
X$537 23 38 FILLCELL_X4
* cell instance $538 r0 *1 38.76,60.2
X$538 23 2988 1557 1580 1404 38 DFF_X1
* cell instance $539 r0 *1 41.99,60.2
X$539 1557 1383 1490 23 38 1580 MUX2_X1
* cell instance $540 r0 *1 43.32,60.2
X$540 23 38 FILLCELL_X8
* cell instance $541 r0 *1 44.84,60.2
X$541 23 38 FILLCELL_X2
* cell instance $542 r0 *1 45.22,60.2
X$542 23 38 FILLCELL_X1
* cell instance $543 r0 *1 45.41,60.2
X$543 1490 1544 1558 23 38 1632 MUX2_X1
* cell instance $544 r0 *1 46.74,60.2
X$544 1486 23 38 1404 CLKBUF_X3
* cell instance $545 r0 *1 47.69,60.2
X$545 23 38 FILLCELL_X1
* cell instance $546 r0 *1 47.88,60.2
X$546 1491 541 1536 23 38 1551 MUX2_X1
* cell instance $547 r0 *1 49.21,60.2
X$547 1587 23 38 1490 CLKBUF_X2
* cell instance $548 r0 *1 49.97,60.2
X$548 23 38 FILLCELL_X1
* cell instance $549 r0 *1 50.16,60.2
X$549 1587 1530 1559 23 38 1631 MUX2_X1
* cell instance $550 r0 *1 51.49,60.2
X$550 23 38 FILLCELL_X4
* cell instance $551 r0 *1 52.25,60.2
X$551 1525 414 1559 23 38 1589 MUX2_X1
* cell instance $552 m0 *1 53.2,60.2
X$552 1551 1177 23 38 1560 NOR2_X1
* cell instance $553 m0 *1 53.01,60.2
X$553 23 38 FILLCELL_X1
* cell instance $554 m0 *1 53.77,60.2
X$554 23 38 FILLCELL_X2
* cell instance $555 r0 *1 53.58,60.2
X$555 23 38 FILLCELL_X1
* cell instance $556 r0 *1 53.77,60.2
X$556 1485 1550 1560 476 1628 1590 23 38 1641 OAI33_X1
* cell instance $557 m0 *1 54.72,60.2
X$557 23 38 FILLCELL_X8
* cell instance $558 m0 *1 54.15,60.2
X$558 1589 1537 23 38 1590 NOR2_X1
* cell instance $559 m0 *1 56.24,60.2
X$559 23 38 FILLCELL_X4
* cell instance $560 m0 *1 57,60.2
X$560 1494 38 988 23 BUF_X4
* cell instance $561 m0 *1 58.33,60.2
X$561 403 38 374 23 BUF_X4
* cell instance $562 m0 *1 59.66,60.2
X$562 1495 1442 38 23 1408 AND2_X1
* cell instance $563 m0 *1 60.42,60.2
X$563 23 38 FILLCELL_X8
* cell instance $564 m0 *1 61.94,60.2
X$564 23 38 FILLCELL_X1
* cell instance $565 m0 *1 62.13,60.2
X$565 1494 38 840 23 BUF_X4
* cell instance $566 m0 *1 63.46,60.2
X$566 23 38 FILLCELL_X4
* cell instance $567 m0 *1 64.22,60.2
X$567 23 38 FILLCELL_X2
* cell instance $568 r0 *1 55.1,60.2
X$568 23 38 FILLCELL_X1
* cell instance $569 r0 *1 55.29,60.2
X$569 1587 1346 1606 23 38 1682 MUX2_X1
* cell instance $570 r0 *1 56.62,60.2
X$570 23 38 FILLCELL_X16
* cell instance $571 r0 *1 59.14,60.2
X$571 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $572 r0 *1 59.14,60.2
X$572 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $573 r0 *1 59.14,60.2
X$573 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $574 r0 *1 59.66,60.2
X$574 23 38 FILLCELL_X8
* cell instance $575 r0 *1 61.18,60.2
X$575 23 38 FILLCELL_X1
* cell instance $576 r0 *1 61.37,60.2
X$576 23 2895 1608 1595 1644 38 DFF_X1
* cell instance $577 r0 *1 64.6,60.2
X$577 1608 174 1561 23 38 1595 MUX2_X1
* cell instance $578 m0 *1 65.17,60.2
X$578 23 38 FILLCELL_X8
* cell instance $579 m0 *1 64.6,60.2
X$579 1597 23 38 1495 BUF_X1
* cell instance $580 m0 *1 66.69,60.2
X$580 23 38 FILLCELL_X2
* cell instance $581 r0 *1 65.93,60.2
X$581 23 38 FILLCELL_X2
* cell instance $582 r0 *1 66.31,60.2
X$582 227 1627 1593 225 1596 1562 23 38 1563 OAI33_X1
* cell instance $583 m0 *1 67.64,60.2
X$583 23 38 FILLCELL_X8
* cell instance $584 m0 *1 67.07,60.2
X$584 1371 1535 23 38 1596 NOR2_X1
* cell instance $585 m0 *1 69.16,60.2
X$585 23 2569 1538 1592 1301 38 DFF_X1
* cell instance $586 m0 *1 72.39,60.2
X$586 1538 559 1497 23 38 1592 MUX2_X1
* cell instance $587 m0 *1 73.72,60.2
X$587 23 38 FILLCELL_X4
* cell instance $588 m0 *1 74.48,60.2
X$588 23 2674 1498 1548 1336 38 DFF_X1
* cell instance $589 m0 *1 77.71,60.2
X$589 23 38 FILLCELL_X8
* cell instance $590 m0 *1 79.23,60.2
X$590 1073 240 1540 23 38 1565 MUX2_X1
* cell instance $591 m0 *1 80.56,60.2
X$591 23 38 FILLCELL_X16
* cell instance $592 m0 *1 83.6,60.2
X$592 23 38 FILLCELL_X1
* cell instance $593 m0 *1 83.79,60.2
X$593 1198 23 38 1304 CLKBUF_X3
* cell instance $594 m0 *1 84.74,60.2
X$594 1577 223 1497 23 38 1581 MUX2_X1
* cell instance $595 m0 *1 86.07,60.2
X$595 23 2669 1577 1581 1227 38 DFF_X1
* cell instance $596 m0 *1 89.3,60.2
X$596 23 38 FILLCELL_X8
* cell instance $597 m0 *1 90.82,60.2
X$597 23 38 FILLCELL_X4
* cell instance $598 m0 *1 91.58,60.2
X$598 23 38 FILLCELL_X1
* cell instance $599 m0 *1 91.77,60.2
X$599 1228 1570 23 38 1567 NAND2_X1
* cell instance $600 m0 *1 92.34,60.2
X$600 1225 1573 1462 1226 1543 38 23 1541 OAI221_X1
* cell instance $601 m0 *1 93.48,60.2
X$601 1228 1502 23 38 1573 NAND2_X1
* cell instance $602 m0 *1 94.05,60.2
X$602 1502 1239 23 38 1543 NAND2_X1
* cell instance $603 m0 *1 94.62,60.2
X$603 1570 1230 23 38 1542 NAND2_X1
* cell instance $604 m0 *1 95.19,60.2
X$604 23 38 FILLCELL_X8
* cell instance $605 m0 *1 96.71,60.2
X$605 23 38 FILLCELL_X2
* cell instance $606 r0 *1 67.64,60.2
X$606 23 1594 1332 38 BUF_X16
* cell instance $607 r0 *1 72.39,60.2
X$607 1564 520 1497 23 38 1624 MUX2_X1
* cell instance $608 r0 *1 73.72,60.2
X$608 1538 541 1564 23 38 1588 MUX2_X1
* cell instance $609 r0 *1 75.05,60.2
X$609 23 38 FILLCELL_X4
* cell instance $610 r0 *1 75.81,60.2
X$610 23 38 FILLCELL_X2
* cell instance $611 r0 *1 76.19,60.2
X$611 1392 23 38 1336 CLKBUF_X3
* cell instance $612 r0 *1 77.14,60.2
X$612 1588 1177 23 38 1621 NOR2_X1
* cell instance $613 r0 *1 77.71,60.2
X$613 23 38 FILLCELL_X4
* cell instance $614 r0 *1 78.47,60.2
X$614 23 38 FILLCELL_X1
* cell instance $615 r0 *1 78.66,60.2
X$615 1620 374 23 38 1678 NOR2_X1
* cell instance $616 r0 *1 79.23,60.2
X$616 23 2889 1540 1565 1336 38 DFF_X1
* cell instance $617 r0 *1 82.46,60.2
X$617 1586 88 1497 23 38 1619 MUX2_X1
* cell instance $618 r0 *1 83.79,60.2
X$618 1582 174 1497 23 38 1584 MUX2_X1
* cell instance $619 r0 *1 85.12,60.2
X$619 23 2856 1582 1584 1227 38 DFF_X1
* cell instance $620 r0 *1 88.35,60.2
X$620 227 1616 1578 225 1152 1471 23 38 1566 OAI33_X1
* cell instance $621 r0 *1 89.68,60.2
X$621 1331 38 1306 23 BUF_X4
* cell instance $622 r0 *1 91.01,60.2
X$622 23 38 FILLCELL_X2
* cell instance $623 r0 *1 91.39,60.2
X$623 1225 1567 1461 1226 1568 38 23 1572 OAI221_X1
* cell instance $624 r0 *1 92.53,60.2
X$624 1570 1239 23 38 1568 NAND2_X1
* cell instance $625 r0 *1 93.1,60.2
X$625 23 38 FILLCELL_X1
* cell instance $626 r0 *1 93.29,60.2
X$626 23 2879 1570 1572 1227 38 DFF_X1
* cell instance $627 r0 *1 96.52,60.2
X$627 23 38 FILLCELL_X2
* cell instance $628 r0 *1 96.9,60.2
X$628 23 38 FILLCELL_X1
* cell instance $629 m90 *1 97.28,60.2
X$629 23 38 23 38 TAPCELL_X1
* cell instance $630 r180 *1 97.28,60.2
X$630 23 38 23 38 TAPCELL_X1
* cell instance $631 r0 *1 3.14,3.4
X$631 23 VIA_via5_6_960_2800_5_2_600_600
* cell instance $632 r0 *1 3.14,3.4
X$632 23 VIA_via4_5_960_2800_5_2_600_600
* cell instance $633 r0 *1 3.14,3.4
X$633 23 VIA_via6_7_960_2800_4_1_600_600
* cell instance $634 r0 *1 59.14,33.4
X$634 23 VIA_via5_6_960_2800_5_2_600_600
* cell instance $635 r0 *1 59.14,33.4
X$635 23 VIA_via4_5_960_2800_5_2_600_600
* cell instance $636 r0 *1 59.14,33.4
X$636 23 VIA_via6_7_960_2800_4_1_600_600
* cell instance $637 r0 *1 3.14,33.4
X$637 23 VIA_via5_6_960_2800_5_2_600_600
* cell instance $638 r0 *1 3.14,33.4
X$638 23 VIA_via4_5_960_2800_5_2_600_600
* cell instance $639 r0 *1 3.14,33.4
X$639 23 VIA_via6_7_960_2800_4_1_600_600
* cell instance $640 r0 *1 59.14,3.4
X$640 23 VIA_via5_6_960_2800_5_2_600_600
* cell instance $641 r0 *1 59.14,3.4
X$641 23 VIA_via4_5_960_2800_5_2_600_600
* cell instance $642 r0 *1 59.14,3.4
X$642 23 VIA_via6_7_960_2800_4_1_600_600
* cell instance $643 m0 *1 36.86,96.6
X$643 2220 1346 2524 23 38 2514 MUX2_X1
* cell instance $644 m0 *1 36.67,96.6
X$644 23 38 FILLCELL_X1
* cell instance $645 m0 *1 38.19,96.6
X$645 2523 23 38 2220 BUF_X1
* cell instance $646 m0 *1 38.76,96.6
X$646 2147 23 38 2522 BUF_X1
* cell instance $647 m0 *1 39.33,96.6
X$647 23 38 FILLCELL_X2
* cell instance $648 m0 *1 10.07,40.6
X$648 928 941 453 23 38 962 MUX2_X1
* cell instance $649 m0 *1 6.84,40.6
X$649 23 2709 1012 965 789 38 DFF_X1
* cell instance $650 m0 *1 11.4,40.6
X$650 23 38 FILLCELL_X4
* cell instance $651 m0 *1 12.16,40.6
X$651 23 38 FILLCELL_X1
* cell instance $652 m0 *1 12.35,40.6
X$652 968 929 295 23 38 989 MUX2_X1
* cell instance $653 m0 *1 13.68,40.6
X$653 23 38 FILLCELL_X4
* cell instance $654 m0 *1 14.44,40.6
X$654 23 38 FILLCELL_X1
* cell instance $655 m0 *1 14.63,40.6
X$655 930 900 968 23 38 969 MUX2_X1
* cell instance $656 m0 *1 15.96,40.6
X$656 23 38 FILLCELL_X1
* cell instance $657 m0 *1 16.15,40.6
X$657 969 893 23 38 888 NOR2_X1
* cell instance $658 m0 *1 16.72,40.6
X$658 23 38 FILLCELL_X1
* cell instance $659 m0 *1 16.91,40.6
X$659 932 1013 972 891 970 892 23 38 1017 OAI33_X1
* cell instance $660 m0 *1 18.24,40.6
X$660 1016 900 934 23 38 933 MUX2_X1
* cell instance $661 m0 *1 19.57,40.6
X$661 934 929 453 23 38 1018 MUX2_X1
* cell instance $662 m0 *1 20.9,40.6
X$662 23 38 FILLCELL_X16
* cell instance $663 m0 *1 23.94,40.6
X$663 23 38 FILLCELL_X8
* cell instance $664 m0 *1 25.46,40.6
X$664 23 38 FILLCELL_X2
* cell instance $665 m0 *1 1.33,40.6
X$665 23 38 FILLCELL_X4
* cell instance $666 m0 *1 1.14,40.6
X$666 23 38 23 38 TAPCELL_X1
* cell instance $667 m0 *1 2.09,40.6
X$667 23 38 FILLCELL_X2
* cell instance $668 r0 *1 1.14,40.6
X$668 23 38 23 38 TAPCELL_X1
* cell instance $669 r0 *1 1.33,40.6
X$669 23 38 FILLCELL_X16
* cell instance $670 m0 *1 5.7,40.6
X$670 23 38 FILLCELL_X4
* cell instance $671 m0 *1 2.47,40.6
X$671 23 2708 1011 961 789 38 DFF_X1
* cell instance $672 m0 *1 6.46,40.6
X$672 23 38 FILLCELL_X2
* cell instance $673 r0 *1 3.14,40.6
X$673 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $674 r0 *1 3.14,40.6
X$674 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $675 r0 *1 3.14,40.6
X$675 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $676 r0 *1 4.37,40.6
X$676 23 38 FILLCELL_X4
* cell instance $677 r0 *1 5.13,40.6
X$677 1011 941 295 23 38 961 MUX2_X1
* cell instance $678 r0 *1 6.46,40.6
X$678 1011 994 887 23 38 967 MUX2_X1
* cell instance $679 r0 *1 7.79,40.6
X$679 1012 992 453 23 38 965 MUX2_X1
* cell instance $680 r0 *1 9.12,40.6
X$680 928 994 1012 23 38 1015 MUX2_X1
* cell instance $681 r0 *1 10.45,40.6
X$681 23 38 FILLCELL_X8
* cell instance $682 r0 *1 11.97,40.6
X$682 23 38 FILLCELL_X2
* cell instance $683 r0 *1 12.35,40.6
X$683 23 3077 968 989 991 38 DFF_X1
* cell instance $684 r0 *1 15.58,40.6
X$684 23 38 FILLCELL_X1
* cell instance $685 r0 *1 15.77,40.6
X$685 1015 937 23 38 1013 NOR2_X1
* cell instance $686 r0 *1 16.34,40.6
X$686 23 38 FILLCELL_X2
* cell instance $687 r0 *1 16.72,40.6
X$687 1016 858 453 23 38 990 MUX2_X1
* cell instance $688 r0 *1 18.05,40.6
X$688 23 38 FILLCELL_X2
* cell instance $689 r0 *1 18.43,40.6
X$689 23 3072 934 1018 991 38 DFF_X1
* cell instance $690 r0 *1 21.66,40.6
X$690 23 38 FILLCELL_X2
* cell instance $691 r0 *1 22.04,40.6
X$691 23 2949 1031 1029 991 38 DFF_X1
* cell instance $692 r0 *1 25.27,40.6
X$692 23 38 FILLCELL_X16
* cell instance $693 m0 *1 26.41,40.6
X$693 23 2847 939 938 942 38 DFF_X1
* cell instance $694 m0 *1 25.84,40.6
X$694 936 937 23 38 935 NOR2_X1
* cell instance $695 m0 *1 29.64,40.6
X$695 940 893 23 38 1020 NOR2_X1
* cell instance $696 m0 *1 30.21,40.6
X$696 23 2736 943 1019 942 38 DFF_X1
* cell instance $697 m0 *1 33.44,40.6
X$697 943 994 945 23 38 995 MUX2_X1
* cell instance $698 m0 *1 34.77,40.6
X$698 932 996 981 891 946 859 23 38 997 OAI33_X1
* cell instance $699 m0 *1 36.1,40.6
X$699 23 38 FILLCELL_X8
* cell instance $700 m0 *1 37.62,40.6
X$700 23 38 FILLCELL_X1
* cell instance $701 m0 *1 37.81,40.6
X$701 948 840 23 38 981 NOR2_X1
* cell instance $702 m0 *1 38.38,40.6
X$702 23 38 FILLCELL_X8
* cell instance $703 m0 *1 39.9,40.6
X$703 23 38 FILLCELL_X2
* cell instance $704 r0 *1 28.31,40.6
X$704 23 38 FILLCELL_X8
* cell instance $705 r0 *1 29.83,40.6
X$705 23 38 FILLCELL_X2
* cell instance $706 r0 *1 30.21,40.6
X$706 23 38 FILLCELL_X1
* cell instance $707 r0 *1 30.4,40.6
X$707 932 1022 1020 891 1023 993 23 38 1021 OAI33_X1
* cell instance $708 r0 *1 31.73,40.6
X$708 23 3063 945 944 942 38 DFF_X1
* cell instance $709 r0 *1 34.96,40.6
X$709 995 881 23 38 996 NOR2_X1
* cell instance $710 r0 *1 35.53,40.6
X$710 23 38 FILLCELL_X16
* cell instance $711 r0 *1 38.57,40.6
X$711 23 38 FILLCELL_X2
* cell instance $712 r0 *1 38.95,40.6
X$712 794 829 23 38 1086 NOR2_X1
* cell instance $713 r0 *1 39.52,40.6
X$713 998 941 398 23 38 949 MUX2_X1
* cell instance $714 m0 *1 43.51,40.6
X$714 23 38 FILLCELL_X4
* cell instance $715 m0 *1 40.28,40.6
X$715 23 2717 998 949 1035 38 DFF_X1
* cell instance $716 m0 *1 44.27,40.6
X$716 23 38 FILLCELL_X2
* cell instance $717 r0 *1 40.85,40.6
X$717 23 38 FILLCELL_X4
* cell instance $718 r0 *1 41.61,40.6
X$718 23 38 FILLCELL_X2
* cell instance $719 r0 *1 41.99,40.6
X$719 999 992 398 23 38 1034 MUX2_X1
* cell instance $720 r0 *1 43.32,40.6
X$720 998 862 999 23 38 1000 MUX2_X1
* cell instance $721 r0 *1 44.65,40.6
X$721 23 38 FILLCELL_X16
* cell instance $722 m0 *1 44.84,40.6
X$722 1000 881 23 38 982 NOR2_X1
* cell instance $723 m0 *1 44.65,40.6
X$723 23 38 FILLCELL_X1
* cell instance $724 m0 *1 45.41,40.6
X$724 23 38 FILLCELL_X16
* cell instance $725 m0 *1 48.45,40.6
X$725 23 2728 1002 1001 839 38 DFF_X1
* cell instance $726 m0 *1 51.68,40.6
X$726 23 38 FILLCELL_X8
* cell instance $727 m0 *1 53.2,40.6
X$727 23 38 FILLCELL_X1
* cell instance $728 m0 *1 53.39,40.6
X$728 988 38 190 23 BUF_X4
* cell instance $729 m0 *1 54.72,40.6
X$729 23 38 FILLCELL_X1
* cell instance $730 m0 *1 54.91,40.6
X$730 988 23 38 367 CLKBUF_X3
* cell instance $731 m0 *1 55.86,40.6
X$731 23 38 FILLCELL_X8
* cell instance $732 m0 *1 57.38,40.6
X$732 950 190 23 38 1003 NOR2_X1
* cell instance $733 m0 *1 57.95,40.6
X$733 23 38 FILLCELL_X4
* cell instance $734 m0 *1 58.71,40.6
X$734 23 2817 951 952 1038 38 DFF_X1
* cell instance $735 m0 *1 61.94,40.6
X$735 23 38 FILLCELL_X1
* cell instance $736 m0 *1 62.13,40.6
X$736 953 190 23 38 1004 NOR2_X1
* cell instance $737 m0 *1 62.7,40.6
X$737 23 38 FILLCELL_X4
* cell instance $738 m0 *1 63.46,40.6
X$738 955 559 799 23 38 1026 MUX2_X1
* cell instance $739 m0 *1 64.79,40.6
X$739 23 38 FILLCELL_X4
* cell instance $740 m0 *1 65.55,40.6
X$740 23 38 FILLCELL_X2
* cell instance $741 r0 *1 47.69,40.6
X$741 23 38 FILLCELL_X2
* cell instance $742 r0 *1 48.07,40.6
X$742 23 38 FILLCELL_X1
* cell instance $743 r0 *1 48.26,40.6
X$743 1002 858 301 23 38 1001 MUX2_X1
* cell instance $744 r0 *1 49.59,40.6
X$744 23 38 FILLCELL_X2
* cell instance $745 r0 *1 49.97,40.6
X$745 1002 900 984 23 38 1027 MUX2_X1
* cell instance $746 r0 *1 51.3,40.6
X$746 23 38 FILLCELL_X16
* cell instance $747 r0 *1 54.34,40.6
X$747 23 38 FILLCELL_X8
* cell instance $748 r0 *1 55.86,40.6
X$748 988 38 372 23 BUF_X4
* cell instance $749 r0 *1 57.19,40.6
X$749 23 38 FILLCELL_X16
* cell instance $750 r0 *1 59.14,40.6
X$750 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $751 r0 *1 59.14,40.6
X$751 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $752 r0 *1 59.14,40.6
X$752 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $753 r0 *1 60.23,40.6
X$753 23 38 FILLCELL_X4
* cell instance $754 r0 *1 60.99,40.6
X$754 23 38 FILLCELL_X1
* cell instance $755 r0 *1 61.18,40.6
X$755 598 38 223 23 BUF_X4
* cell instance $756 r0 *1 62.51,40.6
X$756 23 38 FILLCELL_X4
* cell instance $757 r0 *1 63.27,40.6
X$757 23 38 FILLCELL_X2
* cell instance $758 r0 *1 63.65,40.6
X$758 23 38 FILLCELL_X1
* cell instance $759 r0 *1 63.84,40.6
X$759 23 2927 955 1026 954 38 DFF_X1
* cell instance $760 m0 *1 67.26,40.6
X$760 23 38 FILLCELL_X4
* cell instance $761 m0 *1 65.93,40.6
X$761 955 541 906 23 38 979 MUX2_X1
* cell instance $762 m0 *1 68.02,40.6
X$762 979 367 23 38 978 NOR2_X1
* cell instance $763 m0 *1 68.59,40.6
X$763 799 260 1005 23 38 1025 MUX2_X1
* cell instance $764 m0 *1 69.92,40.6
X$764 23 38 FILLCELL_X4
* cell instance $765 m0 *1 70.68,40.6
X$765 675 240 977 23 38 1024 MUX2_X1
* cell instance $766 m0 *1 72.01,40.6
X$766 23 2734 977 1024 801 38 DFF_X1
* cell instance $767 m0 *1 75.24,40.6
X$767 23 38 FILLCELL_X4
* cell instance $768 m0 *1 76,40.6
X$768 23 2800 974 976 801 38 DFF_X1
* cell instance $769 m0 *1 79.23,40.6
X$769 23 38 FILLCELL_X2
* cell instance $770 r0 *1 67.07,40.6
X$770 23 38 FILLCELL_X2
* cell instance $771 r0 *1 67.45,40.6
X$771 23 38 FILLCELL_X1
* cell instance $772 r0 *1 67.64,40.6
X$772 23 2892 1005 1025 954 38 DFF_X1
* cell instance $773 r0 *1 70.87,40.6
X$773 1005 414 977 23 38 1006 MUX2_X1
* cell instance $774 r0 *1 72.2,40.6
X$774 23 38 FILLCELL_X16
* cell instance $775 r0 *1 75.24,40.6
X$775 23 38 FILLCELL_X4
* cell instance $776 r0 *1 76,40.6
X$776 23 2899 1047 1046 801 38 DFF_X1
* cell instance $777 r0 *1 79.23,40.6
X$777 23 38 FILLCELL_X4
* cell instance $778 m0 *1 79.8,40.6
X$778 1008 130 907 23 38 1007 MUX2_X1
* cell instance $779 m0 *1 79.61,40.6
X$779 23 38 FILLCELL_X1
* cell instance $780 m0 *1 81.13,40.6
X$780 23 38 FILLCELL_X4
* cell instance $781 m0 *1 81.89,40.6
X$781 23 38 FILLCELL_X1
* cell instance $782 m0 *1 82.08,40.6
X$782 974 724 1008 23 38 971 MUX2_X1
* cell instance $783 m0 *1 83.41,40.6
X$783 23 38 FILLCELL_X8
* cell instance $784 m0 *1 84.93,40.6
X$784 23 38 FILLCELL_X4
* cell instance $785 m0 *1 85.69,40.6
X$785 23 38 FILLCELL_X2
* cell instance $786 r0 *1 79.99,40.6
X$786 23 2896 1008 1007 1042 38 DFF_X1
* cell instance $787 r0 *1 83.22,40.6
X$787 23 38 FILLCELL_X4
* cell instance $788 r0 *1 83.98,40.6
X$788 23 38 FILLCELL_X2
* cell instance $789 r0 *1 84.36,40.6
X$789 675 23 38 799 BUF_X2
* cell instance $790 r0 *1 85.12,40.6
X$790 23 38 FILLCELL_X4
* cell instance $791 r0 *1 85.88,40.6
X$791 23 38 FILLCELL_X2
* cell instance $792 m0 *1 86.64,40.6
X$792 23 38 FILLCELL_X4
* cell instance $793 m0 *1 86.07,40.6
X$793 971 190 23 38 966 NOR2_X1
* cell instance $794 m0 *1 87.4,40.6
X$794 23 38 FILLCELL_X1
* cell instance $795 m0 *1 87.59,40.6
X$795 23 2804 911 956 876 38 DFF_X1
* cell instance $796 m0 *1 90.82,40.6
X$796 23 38 FILLCELL_X2
* cell instance $797 r0 *1 86.26,40.6
X$797 806 23 38 907 BUF_X2
* cell instance $798 r0 *1 87.02,40.6
X$798 23 38 FILLCELL_X2
* cell instance $799 r0 *1 87.4,40.6
X$799 23 38 FILLCELL_X1
* cell instance $800 r0 *1 87.59,40.6
X$800 1010 23 38 710 CLKBUF_X2
* cell instance $801 r0 *1 88.35,40.6
X$801 23 38 FILLCELL_X16
* cell instance $802 m0 *1 92.53,40.6
X$802 23 38 FILLCELL_X2
* cell instance $803 m0 *1 91.2,40.6
X$803 1009 263 958 23 38 957 MUX2_X1
* cell instance $804 r0 *1 91.39,40.6
X$804 23 38 FILLCELL_X2
* cell instance $805 r0 *1 91.77,40.6
X$805 806 191 1009 23 38 1014 MUX2_X1
* cell instance $806 m0 *1 93.1,40.6
X$806 806 187 958 23 38 959 MUX2_X1
* cell instance $807 m0 *1 92.91,40.6
X$807 23 38 FILLCELL_X1
* cell instance $808 m0 *1 94.43,40.6
X$808 23 38 FILLCELL_X8
* cell instance $809 m0 *1 95.95,40.6
X$809 23 38 FILLCELL_X4
* cell instance $810 m0 *1 96.71,40.6
X$810 23 38 FILLCELL_X2
* cell instance $811 r0 *1 93.1,40.6
X$811 23 2861 1009 1014 876 38 DFF_X1
* cell instance $812 r0 *1 96.33,40.6
X$812 23 38 FILLCELL_X4
* cell instance $813 r180 *1 97.28,40.6
X$813 23 38 23 38 TAPCELL_X1
* cell instance $814 m90 *1 97.28,40.6
X$814 23 38 23 38 TAPCELL_X1
* cell instance $815 m0 *1 91.77,15.4
X$815 377 191 313 23 38 335 MUX2_X1
* cell instance $816 m0 *1 91.58,15.4
X$816 23 38 FILLCELL_X1
* cell instance $817 m0 *1 93.1,15.4
X$817 23 38 FILLCELL_X2
* cell instance $818 r0 *1 91.58,15.4
X$818 23 2908 313 335 310 38 DFF_X1
* cell instance $819 m0 *1 96.71,15.4
X$819 23 38 FILLCELL_X2
* cell instance $820 m0 *1 93.48,15.4
X$820 23 2609 336 311 310 38 DFF_X1
* cell instance $821 r0 *1 94.81,15.4
X$821 377 187 336 23 38 311 MUX2_X1
* cell instance $822 r0 *1 96.14,15.4
X$822 23 38 FILLCELL_X4
* cell instance $823 r0 *1 96.9,15.4
X$823 23 38 FILLCELL_X1
* cell instance $824 r180 *1 97.28,15.4
X$824 23 38 23 38 TAPCELL_X1
* cell instance $825 m90 *1 97.28,15.4
X$825 23 38 23 38 TAPCELL_X1
* cell instance $826 m0 *1 10.45,51.8
X$826 1327 212 1294 23 38 1311 MUX2_X1
* cell instance $827 m0 *1 7.22,51.8
X$827 23 2606 1294 1293 1326 38 DFF_X1
* cell instance $828 m0 *1 11.78,51.8
X$828 1311 254 23 38 1295 NOR2_X1
* cell instance $829 m0 *1 12.35,51.8
X$829 23 38 FILLCELL_X16
* cell instance $830 m0 *1 15.39,51.8
X$830 890 340 1136 1137 38 23 1312 OAI22_X2
* cell instance $831 m0 *1 17.1,51.8
X$831 1312 1210 1296 38 23 1343 OAI21_X4
* cell instance $832 m0 *1 19.57,51.8
X$832 1017 433 1136 1137 38 23 1261 OAI22_X2
* cell instance $833 m0 *1 21.28,51.8
X$833 1017 433 1138 1157 1139 38 23 1297 OAI221_X1
* cell instance $834 m0 *1 22.42,51.8
X$834 1330 1122 23 38 1314 NAND2_X1
* cell instance $835 m0 *1 22.99,51.8
X$835 23 38 FILLCELL_X4
* cell instance $836 m0 *1 23.75,51.8
X$836 23 2628 1170 1315 1326 38 DFF_X1
* cell instance $837 m0 *1 26.98,51.8
X$837 23 38 FILLCELL_X1
* cell instance $838 m0 *1 27.17,51.8
X$838 1158 1170 23 38 1281 NAND2_X1
* cell instance $839 m0 *1 27.74,51.8
X$839 1170 1140 23 38 1243 NAND2_X1
* cell instance $840 m0 *1 28.31,51.8
X$840 23 38 FILLCELL_X16
* cell instance $841 m0 *1 31.35,51.8
X$841 1171 1140 23 38 1263 NAND2_X1
* cell instance $842 m0 *1 31.92,51.8
X$842 23 38 FILLCELL_X4
* cell instance $843 m0 *1 32.68,51.8
X$843 23 38 FILLCELL_X2
* cell instance $844 m0 *1 1.33,51.8
X$844 23 38 FILLCELL_X4
* cell instance $845 m0 *1 1.14,51.8
X$845 23 38 23 38 TAPCELL_X1
* cell instance $846 m0 *1 2.09,51.8
X$846 23 2614 1362 1291 1292 38 DFF_X1
* cell instance $847 m0 *1 5.32,51.8
X$847 23 38 FILLCELL_X8
* cell instance $848 m0 *1 6.84,51.8
X$848 23 38 FILLCELL_X2
* cell instance $849 r0 *1 1.14,51.8
X$849 23 38 23 38 TAPCELL_X1
* cell instance $850 r0 *1 1.33,51.8
X$850 1343 23 38 1360 BUF_X1
* cell instance $851 r0 *1 1.9,51.8
X$851 23 38 FILLCELL_X1
* cell instance $852 r0 *1 2.09,51.8
X$852 1285 23 38 1290 BUF_X1
* cell instance $853 r0 *1 2.66,51.8
X$853 1324 23 38 1323 BUF_X1
* cell instance $854 r0 *1 3.14,51.8
X$854 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $855 r0 *1 3.14,51.8
X$855 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $856 r0 *1 3.14,51.8
X$856 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $857 r0 *1 3.23,51.8
X$857 1322 23 38 1325 CLKBUF_X2
* cell instance $858 r0 *1 3.99,51.8
X$858 23 3007 1423 1345 1292 38 DFF_X1
* cell instance $859 r0 *1 7.22,51.8
X$859 1325 1346 1294 23 38 1293 MUX2_X1
* cell instance $860 r0 *1 8.55,51.8
X$860 23 38 FILLCELL_X2
* cell instance $861 r0 *1 8.93,51.8
X$861 23 2976 1327 1385 1326 38 DFF_X1
* cell instance $862 r0 *1 12.16,51.8
X$862 23 38 FILLCELL_X4
* cell instance $863 r0 *1 12.92,51.8
X$863 23 2987 1387 1328 1326 38 DFF_X1
* cell instance $864 r0 *1 16.15,51.8
X$864 23 38 FILLCELL_X8
* cell instance $865 r0 *1 17.67,51.8
X$865 23 38 FILLCELL_X4
* cell instance $866 r0 *1 18.43,51.8
X$866 1261 1210 1314 38 23 1324 OAI21_X4
* cell instance $867 r0 *1 20.9,51.8
X$867 23 38 FILLCELL_X2
* cell instance $868 r0 *1 21.28,51.8
X$868 1158 1330 23 38 1329 NAND2_X1
* cell instance $869 r0 *1 21.85,51.8
X$869 1206 1329 1297 1208 1349 38 23 1400 OAI221_X1
* cell instance $870 r0 *1 22.99,51.8
X$870 1330 1140 23 38 1349 NAND2_X1
* cell instance $871 r0 *1 23.56,51.8
X$871 23 38 FILLCELL_X32
* cell instance $872 r0 *1 29.64,51.8
X$872 23 38 FILLCELL_X16
* cell instance $873 r0 *1 32.68,51.8
X$873 23 38 FILLCELL_X4
* cell instance $874 m0 *1 33.63,51.8
X$874 23 2811 1143 1264 1262 38 DFF_X1
* cell instance $875 m0 *1 33.06,51.8
X$875 1158 1143 23 38 1249 NAND2_X1
* cell instance $876 m0 *1 36.86,51.8
X$876 1143 1140 23 38 1251 NAND2_X1
* cell instance $877 m0 *1 37.43,51.8
X$877 23 38 FILLCELL_X1
* cell instance $878 m0 *1 37.62,51.8
X$878 1368 1122 23 38 1265 NAND2_X1
* cell instance $879 m0 *1 38.19,51.8
X$879 1298 1122 23 38 1287 NAND2_X1
* cell instance $880 m0 *1 38.76,51.8
X$880 23 1063 428 1136 1286 1137 38 OAI22_X4
* cell instance $881 m0 *1 41.99,51.8
X$881 1158 1298 23 38 1353 NAND2_X1
* cell instance $882 m0 *1 42.56,51.8
X$882 620 38 1454 23 BUF_X4
* cell instance $883 m0 *1 43.89,51.8
X$883 1299 38 634 23 BUF_X4
* cell instance $884 m0 *1 45.22,51.8
X$884 1299 38 620 23 BUF_X4
* cell instance $885 m0 *1 46.55,51.8
X$885 23 38 FILLCELL_X1
* cell instance $886 m0 *1 46.74,51.8
X$886 599 38 1289 23 BUF_X4
* cell instance $887 m0 *1 48.07,51.8
X$887 620 38 541 23 BUF_X4
* cell instance $888 m0 *1 49.4,51.8
X$888 23 38 FILLCELL_X8
* cell instance $889 m0 *1 50.92,51.8
X$889 23 38 FILLCELL_X2
* cell instance $890 r0 *1 33.44,51.8
X$890 23 38 FILLCELL_X2
* cell instance $891 r0 *1 33.82,51.8
X$891 988 38 1177 23 BUF_X4
* cell instance $892 r0 *1 35.15,51.8
X$892 23 1331 1213 38 BUF_X32
* cell instance $893 r0 *1 44.46,51.8
X$893 23 3009 1298 1394 1174 38 DFF_X1
* cell instance $894 r0 *1 47.69,51.8
X$894 1332 1353 1191 1319 1552 38 23 1394 OAI221_X1
* cell instance $895 r0 *1 48.83,51.8
X$895 597 38 1383 23 BUF_X4
* cell instance $896 r0 *1 50.16,51.8
X$896 557 38 1369 23 BUF_X4
* cell instance $897 m0 *1 52.63,51.8
X$897 23 38 FILLCELL_X1
* cell instance $898 m0 *1 51.3,51.8
X$898 1299 38 862 23 BUF_X4
* cell instance $899 m0 *1 52.82,51.8
X$899 1318 23 38 1138 CLKBUF_X3
* cell instance $900 m0 *1 53.77,51.8
X$900 925 426 1138 1198 1300 38 23 1266 OAI221_X1
* cell instance $901 m0 *1 54.91,51.8
X$901 23 1136 38 1300 BUF_X8
* cell instance $902 m0 *1 57.38,51.8
X$902 23 38 FILLCELL_X2
* cell instance $903 r0 *1 51.49,51.8
X$903 23 38 FILLCELL_X1
* cell instance $904 r0 *1 51.68,51.8
X$904 1145 23 38 1485 CLKBUF_X3
* cell instance $905 r0 *1 52.63,51.8
X$905 620 38 188 23 BUF_X4
* cell instance $906 r0 *1 53.96,51.8
X$906 23 38 FILLCELL_X1
* cell instance $907 r0 *1 54.15,51.8
X$907 1158 1333 23 38 1334 NAND2_X1
* cell instance $908 r0 *1 54.72,51.8
X$908 1332 1334 1266 1319 1357 38 23 1440 OAI221_X1
* cell instance $909 r0 *1 55.86,51.8
X$909 925 426 1136 1240 38 23 1352 OAI22_X2
* cell instance $910 r0 *1 57.57,51.8
X$910 1333 1140 23 38 1357 NAND2_X1
* cell instance $911 m0 *1 60.99,51.8
X$911 1214 38 373 23 BUF_X4
* cell instance $912 m0 *1 57.76,51.8
X$912 23 2567 1217 1288 1301 38 DFF_X1
* cell instance $913 m0 *1 62.32,51.8
X$913 23 38 FILLCELL_X4
* cell instance $914 m0 *1 63.08,51.8
X$914 23 38 FILLCELL_X2
* cell instance $915 r0 *1 58.14,51.8
X$915 1333 1268 23 38 1351 NAND2_X1
* cell instance $916 r0 *1 58.71,51.8
X$916 23 38 FILLCELL_X8
* cell instance $917 r0 *1 59.14,51.8
X$917 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $918 r0 *1 59.14,51.8
X$918 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $919 r0 *1 59.14,51.8
X$919 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $920 r0 *1 60.23,51.8
X$920 23 38 FILLCELL_X1
* cell instance $921 r0 *1 60.42,51.8
X$921 1130 38 559 23 BUF_X4
* cell instance $922 r0 *1 61.75,51.8
X$922 1065 38 520 23 BUF_X4
* cell instance $923 r0 *1 63.08,51.8
X$923 23 38 FILLCELL_X8
* cell instance $924 m0 *1 63.65,51.8
X$924 23 2570 1267 1359 1301 38 DFF_X1
* cell instance $925 m0 *1 63.46,51.8
X$925 23 38 FILLCELL_X1
* cell instance $926 m0 *1 66.88,51.8
X$926 1335 187 1302 23 38 1284 MUX2_X1
* cell instance $927 m0 *1 68.21,51.8
X$927 1321 23 38 1145 CLKBUF_X2
* cell instance $928 m0 *1 68.97,51.8
X$928 23 38 FILLCELL_X4
* cell instance $929 m0 *1 69.73,51.8
X$929 1220 1219 23 38 1321 OR2_X1
* cell instance $930 m0 *1 70.49,51.8
X$930 1355 23 38 1220 INV_X1
* cell instance $931 m0 *1 70.87,51.8
X$931 23 38 FILLCELL_X32
* cell instance $932 m0 *1 76.95,51.8
X$932 23 38 FILLCELL_X2
* cell instance $933 r0 *1 64.6,51.8
X$933 23 38 FILLCELL_X1
* cell instance $934 r0 *1 64.79,51.8
X$934 1335 191 1267 23 38 1359 MUX2_X1
* cell instance $935 r0 *1 66.12,51.8
X$935 1267 1358 1302 23 38 1371 MUX2_X1
* cell instance $936 r0 *1 67.45,51.8
X$936 1145 23 38 475 CLKBUF_X3
* cell instance $937 r0 *1 68.4,51.8
X$937 23 38 FILLCELL_X2
* cell instance $938 r0 *1 68.78,51.8
X$938 23 38 FILLCELL_X1
* cell instance $939 r0 *1 68.97,51.8
X$939 1356 23 38 515 BUF_X2
* cell instance $940 r0 *1 69.73,51.8
X$940 1355 1219 23 38 1356 OR2_X1
* cell instance $941 r0 *1 70.49,51.8
X$941 23 38 FILLCELL_X16
* cell instance $942 r0 *1 73.53,51.8
X$942 23 3116 1337 1354 1336 38 DFF_X1
* cell instance $943 r0 *1 76.76,51.8
X$943 1073 79 1337 23 38 1354 MUX2_X1
* cell instance $944 m0 *1 80.56,51.8
X$944 1111 133 1269 23 38 1320 MUX2_X1
* cell instance $945 m0 *1 77.33,51.8
X$945 23 2675 1269 1320 1223 38 DFF_X1
* cell instance $946 m0 *1 81.89,51.8
X$946 1218 624 1318 1198 1300 38 23 1376 OAI221_X1
* cell instance $947 m0 *1 83.03,51.8
X$947 23 38 FILLCELL_X1
* cell instance $948 m0 *1 83.22,51.8
X$948 1218 624 1240 1224 38 23 1317 OAI22_X1
* cell instance $949 m0 *1 84.17,51.8
X$949 1225 1303 1317 38 1278 23 OAI21_X1
* cell instance $950 m0 *1 84.93,51.8
X$950 474 285 1304 1305 38 23 1316 OAI22_X1
* cell instance $951 m0 *1 85.88,51.8
X$951 23 38 FILLCELL_X16
* cell instance $952 m0 *1 88.92,51.8
X$952 1306 1270 1316 38 1384 23 OAI21_X1
* cell instance $953 m0 *1 89.68,51.8
X$953 483 265 1304 1305 38 23 1273 OAI22_X1
* cell instance $954 m0 *1 90.63,51.8
X$954 23 38 FILLCELL_X1
* cell instance $955 m0 *1 90.82,51.8
X$955 1225 1307 1279 1226 1313 38 23 1271 OAI221_X1
* cell instance $956 m0 *1 91.96,51.8
X$956 649 608 1304 1305 38 23 1277 OAI22_X1
* cell instance $957 m0 *1 92.91,51.8
X$957 1228 1272 23 38 1307 NAND2_X1
* cell instance $958 m0 *1 93.48,51.8
X$958 23 38 FILLCELL_X1
* cell instance $959 m0 *1 93.67,51.8
X$959 1272 1239 23 38 1313 NAND2_X1
* cell instance $960 m0 *1 94.24,51.8
X$960 23 38 FILLCELL_X1
* cell instance $961 m0 *1 94.43,51.8
X$961 1272 1230 23 38 1309 NAND2_X1
* cell instance $962 m0 *1 95,51.8
X$962 1306 1309 1273 38 1310 23 OAI21_X1
* cell instance $963 m0 *1 95.76,51.8
X$963 1340 23 38 1275 BUF_X1
* cell instance $964 m0 *1 96.33,51.8
X$964 1306 1231 1277 38 1344 23 OAI21_X1
* cell instance $965 r180 *1 97.28,51.8
X$965 23 38 23 38 TAPCELL_X1
* cell instance $966 r0 *1 78.09,51.8
X$966 23 38 FILLCELL_X8
* cell instance $967 r0 *1 79.61,51.8
X$967 1162 522 1318 1198 1300 38 23 1375 OAI221_X1
* cell instance $968 r0 *1 80.75,51.8
X$968 1269 1373 1283 23 38 1391 MUX2_X1
* cell instance $969 r0 *1 82.08,51.8
X$969 1392 23 38 1223 CLKBUF_X3
* cell instance $970 r0 *1 83.03,51.8
X$970 1162 522 1240 1224 38 23 1350 OAI22_X1
* cell instance $971 r0 *1 83.98,51.8
X$971 1225 1351 1352 38 1339 23 OAI21_X1
* cell instance $972 r0 *1 84.74,51.8
X$972 1225 1338 1350 38 1340 23 OAI21_X1
* cell instance $973 r0 *1 85.5,51.8
X$973 1377 1268 23 38 1338 NAND2_X1
* cell instance $974 r0 *1 86.07,51.8
X$974 23 38 FILLCELL_X16
* cell instance $975 r0 *1 89.11,51.8
X$975 23 38 FILLCELL_X2
* cell instance $976 r0 *1 89.49,51.8
X$976 23 38 FILLCELL_X1
* cell instance $977 r0 *1 89.68,51.8
X$977 534 277 1304 1305 38 23 1348 OAI22_X1
* cell instance $978 r0 *1 90.63,51.8
X$978 534 277 1241 1240 1224 38 23 1379 OAI221_X1
* cell instance $979 r0 *1 91.77,51.8
X$979 23 38 FILLCELL_X4
* cell instance $980 r0 *1 92.53,51.8
X$980 23 38 FILLCELL_X2
* cell instance $981 r0 *1 92.91,51.8
X$981 23 38 FILLCELL_X1
* cell instance $982 r0 *1 93.1,51.8
X$982 1306 1380 1348 38 1347 23 OAI21_X1
* cell instance $983 r0 *1 93.86,51.8
X$983 23 38 FILLCELL_X8
* cell instance $984 r0 *1 95.38,51.8
X$984 1339 23 38 1308 BUF_X1
* cell instance $985 r0 *1 95.95,51.8
X$985 1310 23 38 1341 BUF_X1
* cell instance $986 r0 *1 96.52,51.8
X$986 1344 23 38 1276 BUF_X1
* cell instance $987 m90 *1 97.28,51.8
X$987 23 38 23 38 TAPCELL_X1
* cell instance $988 m0 *1 69.92,4.2
X$988 23 38 FILLCELL_X1
* cell instance $989 m0 *1 71.44,4.2
X$989 23 2692 33 63 34 38 DFF_X1
* cell instance $990 m0 *1 74.67,4.2
X$990 23 2596 50 60 34 38 DFF_X1
* cell instance $991 m0 *1 77.9,4.2
X$991 52 51 50 23 38 60 MUX2_X1
* cell instance $992 m0 *1 79.23,4.2
X$992 23 38 FILLCELL_X2
* cell instance $993 r0 *1 71.25,4.2
X$993 23 38 FILLCELL_X8
* cell instance $994 r0 *1 72.77,4.2
X$994 23 38 FILLCELL_X2
* cell instance $995 r0 *1 73.15,4.2
X$995 77 79 81 23 38 125 MUX2_X1
* cell instance $996 r0 *1 74.48,4.2
X$996 23 38 FILLCELL_X4
* cell instance $997 r0 *1 75.24,4.2
X$997 23 38 FILLCELL_X2
* cell instance $998 r0 *1 75.62,4.2
X$998 23 38 FILLCELL_X1
* cell instance $999 r0 *1 75.81,4.2
X$999 49 23 38 78 BUF_X2
* cell instance $1000 r0 *1 76.57,4.2
X$1000 23 38 FILLCELL_X4
* cell instance $1001 r0 *1 78.66,4.2
X$1001 23 38 FILLCELL_X4
* cell instance $1002 r0 *1 79.42,4.2
X$1002 23 38 FILLCELL_X2
* cell instance $1003 m0 *1 79.61,4.2
X$1003 23 38 FILLCELL_X1
* cell instance $1004 m0 *1 80.56,4.2
X$1004 23 38 FILLCELL_X8
* cell instance $1005 m0 *1 82.08,4.2
X$1005 23 38 FILLCELL_X1
* cell instance $1006 m0 *1 82.27,4.2
X$1006 23 2801 86 35 36 38 DFF_X1
* cell instance $1007 m0 *1 85.5,4.2
X$1007 53 23 38 52 BUF_X2
* cell instance $1008 m0 *1 86.26,4.2
X$1008 23 38 FILLCELL_X32
* cell instance $1009 m0 *1 92.34,4.2
X$1009 23 38 FILLCELL_X16
* cell instance $1010 m0 *1 95.38,4.2
X$1010 23 38 FILLCELL_X8
* cell instance $1011 m0 *1 96.9,4.2
X$1011 23 38 FILLCELL_X1
* cell instance $1012 r180 *1 97.28,4.2
X$1012 23 38 23 38 TAPCELL_X1
* cell instance $1013 r0 *1 79.8,4.2
X$1013 82 88 52 23 38 132 MUX2_X1
* cell instance $1014 r0 *1 81.13,4.2
X$1014 23 38 FILLCELL_X1
* cell instance $1015 r0 *1 81.32,4.2
X$1015 86 88 78 23 38 35 MUX2_X1
* cell instance $1016 r0 *1 82.65,4.2
X$1016 23 2898 145 109 83 38 DFF_X1
* cell instance $1017 r0 *1 85.88,4.2
X$1017 23 38 FILLCELL_X4
* cell instance $1018 r0 *1 86.64,4.2
X$1018 23 38 FILLCELL_X1
* cell instance $1019 r0 *1 86.83,4.2
X$1019 23 3084 54 108 83 38 DFF_X1
* cell instance $1020 r0 *1 90.06,4.2
X$1020 49 79 85 23 38 84 MUX2_X1
* cell instance $1021 r0 *1 91.39,4.2
X$1021 23 3129 85 84 83 38 DFF_X1
* cell instance $1022 r0 *1 94.62,4.2
X$1022 23 38 FILLCELL_X8
* cell instance $1023 r0 *1 96.14,4.2
X$1023 23 38 FILLCELL_X4
* cell instance $1024 r0 *1 96.9,4.2
X$1024 23 38 FILLCELL_X1
* cell instance $1025 m90 *1 97.28,4.2
X$1025 23 38 23 38 TAPCELL_X1
* cell instance $1026 m0 *1 73.53,23.8
X$1026 580 541 477 23 38 478 MUX2_X1
* cell instance $1027 m0 *1 72.2,23.8
X$1027 580 559 52 23 38 537 MUX2_X1
* cell instance $1028 m0 *1 74.86,23.8
X$1028 23 38 FILLCELL_X1
* cell instance $1029 m0 *1 75.05,23.8
X$1029 607 367 23 38 577 NOR2_X1
* cell instance $1030 m0 *1 75.62,23.8
X$1030 23 38 FILLCELL_X1
* cell instance $1031 m0 *1 75.81,23.8
X$1031 562 373 524 23 38 523 MUX2_X1
* cell instance $1032 m0 *1 77.14,23.8
X$1032 23 38 FILLCELL_X1
* cell instance $1033 m0 *1 77.33,23.8
X$1033 616 438 562 23 38 618 MUX2_X1
* cell instance $1034 m0 *1 78.66,23.8
X$1034 475 617 577 476 563 564 23 38 649 OAI33_X1
* cell instance $1035 m0 *1 79.99,23.8
X$1035 565 374 23 38 564 NOR2_X1
* cell instance $1036 m0 *1 80.56,23.8
X$1036 23 38 FILLCELL_X2
* cell instance $1037 r0 *1 72.2,23.8
X$1037 606 559 524 23 38 605 MUX2_X1
* cell instance $1038 r0 *1 73.53,23.8
X$1038 606 541 642 23 38 607 MUX2_X1
* cell instance $1039 r0 *1 74.86,23.8
X$1039 23 38 FILLCELL_X1
* cell instance $1040 r0 *1 75.05,23.8
X$1040 616 441 524 23 38 619 MUX2_X1
* cell instance $1041 r0 *1 76.38,23.8
X$1041 23 2911 616 619 445 38 DFF_X1
* cell instance $1042 r0 *1 79.61,23.8
X$1042 618 370 23 38 617 NOR2_X1
* cell instance $1043 r0 *1 80.18,23.8
X$1043 23 38 FILLCELL_X32
* cell instance $1044 m0 *1 81.89,23.8
X$1044 524 260 525 23 38 575 MUX2_X1
* cell instance $1045 m0 *1 80.94,23.8
X$1045 139 23 38 445 CLKBUF_X3
* cell instance $1046 m0 *1 83.22,23.8
X$1046 23 2580 525 575 445 38 DFF_X1
* cell instance $1047 m0 *1 86.45,23.8
X$1047 573 223 524 23 38 566 MUX2_X1
* cell instance $1048 m0 *1 87.78,23.8
X$1048 23 38 FILLCELL_X4
* cell instance $1049 m0 *1 88.54,23.8
X$1049 23 38 FILLCELL_X2
* cell instance $1050 r0 *1 86.26,23.8
X$1050 23 38 FILLCELL_X1
* cell instance $1051 r0 *1 86.45,23.8
X$1051 650 190 23 38 613 NOR2_X1
* cell instance $1052 r0 *1 87.02,23.8
X$1052 23 38 FILLCELL_X16
* cell instance $1053 m0 *1 89.11,23.8
X$1053 573 188 529 23 38 572 MUX2_X1
* cell instance $1054 m0 *1 88.92,23.8
X$1054 23 38 FILLCELL_X1
* cell instance $1055 m0 *1 90.44,23.8
X$1055 572 261 23 38 612 NOR2_X1
* cell instance $1056 m0 *1 91.01,23.8
X$1056 23 38 FILLCELL_X4
* cell instance $1057 m0 *1 91.77,23.8
X$1057 23 38 FILLCELL_X2
* cell instance $1058 r0 *1 90.06,23.8
X$1058 23 38 FILLCELL_X4
* cell instance $1059 r0 *1 90.82,23.8
X$1059 23 38 FILLCELL_X2
* cell instance $1060 r0 *1 91.2,23.8
X$1060 227 612 613 225 567 609 23 38 608 OAI33_X1
* cell instance $1061 m0 *1 92.34,23.8
X$1061 570 177 23 38 609 NOR2_X1
* cell instance $1062 m0 *1 92.15,23.8
X$1062 23 38 FILLCELL_X1
* cell instance $1063 m0 *1 92.91,23.8
X$1063 23 38 FILLCELL_X2
* cell instance $1064 r0 *1 92.53,23.8
X$1064 23 38 FILLCELL_X16
* cell instance $1065 m0 *1 93.48,23.8
X$1065 568 126 480 23 38 570 MUX2_X1
* cell instance $1066 m0 *1 93.29,23.8
X$1066 23 38 FILLCELL_X1
* cell instance $1067 m0 *1 94.81,23.8
X$1067 377 133 568 23 38 527 MUX2_X1
* cell instance $1068 m0 *1 96.14,23.8
X$1068 23 38 FILLCELL_X4
* cell instance $1069 m0 *1 96.9,23.8
X$1069 23 38 FILLCELL_X1
* cell instance $1070 r180 *1 97.28,23.8
X$1070 23 38 23 38 TAPCELL_X1
* cell instance $1071 r0 *1 95.57,23.8
X$1071 23 38 FILLCELL_X8
* cell instance $1072 m90 *1 97.28,23.8
X$1072 23 38 23 38 TAPCELL_X1
* cell instance $1073 m0 *1 54.53,46.2
X$1073 1101 1065 556 23 38 1131 MUX2_X1
* cell instance $1074 m0 *1 51.3,46.2
X$1074 23 2780 1100 1165 1038 38 DFF_X1
* cell instance $1075 m0 *1 55.86,46.2
X$1075 23 38 FILLCELL_X8
* cell instance $1076 m0 *1 57.38,46.2
X$1076 23 38 FILLCELL_X1
* cell instance $1077 m0 *1 57.57,46.2
X$1077 1128 1130 640 23 38 1129 MUX2_X1
* cell instance $1078 m0 *1 58.9,46.2
X$1078 1038 23 38 CLKBUF_X1
* cell instance $1079 m0 *1 59.47,46.2
X$1079 1128 900 1092 23 38 1127 MUX2_X1
* cell instance $1080 m0 *1 60.8,46.2
X$1080 23 38 FILLCELL_X2
* cell instance $1081 r0 *1 51.3,46.2
X$1081 1145 23 38 932 CLKBUF_X3
* cell instance $1082 r0 *1 52.25,46.2
X$1082 1100 1130 556 23 38 1165 MUX2_X1
* cell instance $1083 r0 *1 53.58,46.2
X$1083 1100 900 1101 23 38 1166 MUX2_X1
* cell instance $1084 r0 *1 54.91,46.2
X$1084 23 38 FILLCELL_X4
* cell instance $1085 r0 *1 55.67,46.2
X$1085 1166 840 23 38 1189 NOR2_X1
* cell instance $1086 r0 *1 56.24,46.2
X$1086 1145 1190 1189 891 1003 798 23 38 1162 OAI33_X1
* cell instance $1087 r0 *1 57.57,46.2
X$1087 23 38 FILLCELL_X4
* cell instance $1088 r0 *1 58.33,46.2
X$1088 744 23 38 1038 CLKBUF_X3
* cell instance $1089 r0 *1 59.14,46.2
X$1089 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $1090 r0 *1 59.14,46.2
X$1090 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $1091 r0 *1 59.14,46.2
X$1091 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $1092 r0 *1 59.28,46.2
X$1092 23 38 FILLCELL_X4
* cell instance $1093 r0 *1 60.04,46.2
X$1093 23 38 FILLCELL_X1
* cell instance $1094 r0 *1 60.23,46.2
X$1094 600 38 225 23 BUF_X4
* cell instance $1095 m0 *1 61.37,46.2
X$1095 1127 840 23 38 1102 NOR2_X1
* cell instance $1096 m0 *1 61.18,46.2
X$1096 23 38 FILLCELL_X1
* cell instance $1097 m0 *1 61.94,46.2
X$1097 23 38 FILLCELL_X16
* cell instance $1098 m0 *1 64.98,46.2
X$1098 23 38 FILLCELL_X8
* cell instance $1099 m0 *1 66.5,46.2
X$1099 954 23 38 CLKBUF_X1
* cell instance $1100 m0 *1 67.07,46.2
X$1100 1067 1105 23 38 1159 NOR2_X1
* cell instance $1101 m0 *1 67.64,46.2
X$1101 799 51 1103 23 38 1161 MUX2_X1
* cell instance $1102 m0 *1 68.97,46.2
X$1102 23 38 FILLCELL_X1
* cell instance $1103 m0 *1 69.16,46.2
X$1103 1103 1099 1040 23 38 1123 MUX2_X1
* cell instance $1104 m0 *1 70.49,46.2
X$1104 23 38 FILLCELL_X1
* cell instance $1105 m0 *1 70.68,46.2
X$1105 1123 372 23 38 1104 NOR2_X1
* cell instance $1106 m0 *1 71.25,46.2
X$1106 23 38 FILLCELL_X16
* cell instance $1107 m0 *1 74.29,46.2
X$1107 23 38 FILLCELL_X4
* cell instance $1108 m0 *1 75.05,46.2
X$1108 23 38 FILLCELL_X2
* cell instance $1109 r0 *1 61.56,46.2
X$1109 1145 1176 1102 864 1004 1163 23 38 1218 OAI33_X1
* cell instance $1110 r0 *1 62.89,46.2
X$1110 23 38 FILLCELL_X16
* cell instance $1111 r0 *1 65.93,46.2
X$1111 23 38 FILLCELL_X4
* cell instance $1112 r0 *1 66.69,46.2
X$1112 23 38 FILLCELL_X1
* cell instance $1113 r0 *1 66.88,46.2
X$1113 23 2875 1103 1161 954 38 DFF_X1
* cell instance $1114 r0 *1 70.11,46.2
X$1114 475 1159 978 476 1104 1147 23 38 1146 OAI33_X1
* cell instance $1115 r0 *1 71.44,46.2
X$1115 23 38 FILLCELL_X4
* cell instance $1116 r0 *1 72.2,46.2
X$1116 23 38 FILLCELL_X1
* cell instance $1117 r0 *1 72.39,46.2
X$1117 1221 559 907 23 38 1186 MUX2_X1
* cell instance $1118 r0 *1 73.72,46.2
X$1118 23 38 FILLCELL_X8
* cell instance $1119 r0 *1 75.24,46.2
X$1119 23 2900 1107 1106 1042 38 DFF_X1
* cell instance $1120 m0 *1 76,46.2
X$1120 907 51 1107 23 38 1106 MUX2_X1
* cell instance $1121 m0 *1 75.43,46.2
X$1121 1089 1105 23 38 1156 NOR2_X1
* cell instance $1122 m0 *1 77.33,46.2
X$1122 23 38 FILLCELL_X2
* cell instance $1123 m0 *1 79.04,46.2
X$1123 1120 372 23 38 1108 NOR2_X1
* cell instance $1124 m0 *1 77.71,46.2
X$1124 1107 1099 1109 23 38 1120 MUX2_X1
* cell instance $1125 m0 *1 79.61,46.2
X$1125 23 38 FILLCELL_X8
* cell instance $1126 m0 *1 81.13,46.2
X$1126 23 38 FILLCELL_X2
* cell instance $1127 r0 *1 78.47,46.2
X$1127 475 1156 1183 476 1108 1148 23 38 1154 OAI33_X1
* cell instance $1128 r0 *1 79.8,46.2
X$1128 23 38 FILLCELL_X4
* cell instance $1129 r0 *1 80.56,46.2
X$1129 23 38 FILLCELL_X2
* cell instance $1130 r0 *1 80.94,46.2
X$1130 23 38 FILLCELL_X1
* cell instance $1131 r0 *1 81.13,46.2
X$1131 23 2910 1109 1110 1042 38 DFF_X1
* cell instance $1132 m0 *1 82.84,46.2
X$1132 23 38 FILLCELL_X4
* cell instance $1133 m0 *1 83.6,46.2
X$1133 744 23 38 1042 CLKBUF_X3
* cell instance $1134 m0 *1 84.55,46.2
X$1134 23 38 FILLCELL_X8
* cell instance $1135 m0 *1 86.07,46.2
X$1135 1111 191 1069 23 38 1118 MUX2_X1
* cell instance $1136 m0 *1 87.4,46.2
X$1136 1111 187 1070 23 38 1116 MUX2_X1
* cell instance $1137 m0 *1 88.73,46.2
X$1137 23 38 FILLCELL_X4
* cell instance $1138 m0 *1 89.49,46.2
X$1138 23 38 FILLCELL_X2
* cell instance $1139 r0 *1 84.36,46.2
X$1139 23 38 FILLCELL_X32
* cell instance $1140 m0 *1 90.06,46.2
X$1140 1112 274 23 38 1153 NOR2_X1
* cell instance $1141 m0 *1 89.87,46.2
X$1141 23 38 FILLCELL_X1
* cell instance $1142 m0 *1 90.63,46.2
X$1142 23 38 FILLCELL_X4
* cell instance $1143 m0 *1 91.39,46.2
X$1143 1071 274 23 38 1152 NOR2_X1
* cell instance $1144 m0 *1 91.96,46.2
X$1144 23 38 FILLCELL_X1
* cell instance $1145 m0 *1 92.15,46.2
X$1145 23 2807 1072 1114 876 38 DFF_X1
* cell instance $1146 m0 *1 95.38,46.2
X$1146 23 38 FILLCELL_X4
* cell instance $1147 m0 *1 96.14,46.2
X$1147 1113 23 38 806 CLKBUF_X2
* cell instance $1148 m0 *1 96.9,46.2
X$1148 23 38 FILLCELL_X1
* cell instance $1149 r180 *1 97.28,46.2
X$1149 23 38 23 38 TAPCELL_X1
* cell instance $1150 r0 *1 90.44,46.2
X$1150 23 38 FILLCELL_X32
* cell instance $1151 r0 *1 96.52,46.2
X$1151 23 38 FILLCELL_X2
* cell instance $1152 r0 *1 96.9,46.2
X$1152 23 38 FILLCELL_X1
* cell instance $1153 m90 *1 97.28,46.2
X$1153 23 38 23 38 TAPCELL_X1
* cell instance $1154 m0 *1 5.7,71.4
X$1154 1789 412 1819 23 38 1840 MUX2_X1
* cell instance $1155 m0 *1 2.47,71.4
X$1155 23 2615 1819 1835 1556 38 DFF_X1
* cell instance $1156 m0 *1 7.03,71.4
X$1156 1819 1369 1791 23 38 1835 MUX2_X1
* cell instance $1157 m0 *1 8.36,71.4
X$1157 23 38 FILLCELL_X16
* cell instance $1158 m0 *1 11.4,71.4
X$1158 1840 354 23 38 1869 NOR2_X1
* cell instance $1159 m0 *1 11.97,71.4
X$1159 23 38 FILLCELL_X8
* cell instance $1160 m0 *1 13.49,71.4
X$1160 23 38 FILLCELL_X2
* cell instance $1161 m0 *1 1.33,71.4
X$1161 23 38 FILLCELL_X4
* cell instance $1162 m0 *1 1.14,71.4
X$1162 23 38 23 38 TAPCELL_X1
* cell instance $1163 m0 *1 2.09,71.4
X$1163 23 38 FILLCELL_X2
* cell instance $1164 r0 *1 1.14,71.4
X$1164 23 38 23 38 TAPCELL_X1
* cell instance $1165 r0 *1 1.33,71.4
X$1165 23 38 FILLCELL_X1
* cell instance $1166 r0 *1 1.52,71.4
X$1166 1867 23 38 1935 BUF_X1
* cell instance $1167 r0 *1 2.09,71.4
X$1167 23 38 FILLCELL_X16
* cell instance $1168 r0 *1 3.14,71.4
X$1168 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $1169 r0 *1 3.14,71.4
X$1169 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $1170 r0 *1 3.14,71.4
X$1170 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $1171 r0 *1 5.13,71.4
X$1171 23 38 FILLCELL_X8
* cell instance $1172 r0 *1 6.65,71.4
X$1172 23 38 FILLCELL_X4
* cell instance $1173 r0 *1 7.41,71.4
X$1173 23 3001 1868 1890 1635 38 DFF_X1
* cell instance $1174 r0 *1 10.64,71.4
X$1174 1868 1289 1791 23 38 1890 MUX2_X1
* cell instance $1175 r0 *1 11.97,71.4
X$1175 23 38 FILLCELL_X4
* cell instance $1176 r0 *1 12.73,71.4
X$1176 23 2951 1870 1923 1635 38 DFF_X1
* cell instance $1177 m0 *1 14.06,71.4
X$1177 23 2572 1842 1841 1635 38 DFF_X1
* cell instance $1178 m0 *1 13.87,71.4
X$1178 23 38 FILLCELL_X1
* cell instance $1179 m0 *1 17.29,71.4
X$1179 23 38 FILLCELL_X2
* cell instance $1180 r0 *1 15.96,71.4
X$1180 23 38 FILLCELL_X2
* cell instance $1181 r0 *1 16.34,71.4
X$1181 1870 1184 1842 23 38 1891 MUX2_X1
* cell instance $1182 m0 *1 17.86,71.4
X$1182 1843 1488 1820 23 38 1792 MUX2_X1
* cell instance $1183 m0 *1 17.67,71.4
X$1183 23 38 FILLCELL_X1
* cell instance $1184 m0 *1 19.19,71.4
X$1184 23 2573 1871 1845 1848 38 DFF_X1
* cell instance $1185 m0 *1 22.42,71.4
X$1185 23 2620 1821 1847 1848 38 DFF_X1
* cell instance $1186 m0 *1 25.65,71.4
X$1186 1821 1488 1822 23 38 1847 MUX2_X1
* cell instance $1187 m0 *1 26.98,71.4
X$1187 23 38 FILLCELL_X16
* cell instance $1188 m0 *1 30.02,71.4
X$1188 23 38 FILLCELL_X1
* cell instance $1189 m0 *1 30.21,71.4
X$1189 1206 1824 1906 1804 1852 38 23 1850 OAI221_X1
* cell instance $1190 m0 *1 31.35,71.4
X$1190 1636 1823 23 38 1824 NAND2_X1
* cell instance $1191 m0 *1 31.92,71.4
X$1191 23 38 FILLCELL_X1
* cell instance $1192 m0 *1 32.11,71.4
X$1192 1823 1638 23 38 1852 NAND2_X1
* cell instance $1193 m0 *1 32.68,71.4
X$1193 1855 1488 1725 23 38 1894 MUX2_X1
* cell instance $1194 m0 *1 34.01,71.4
X$1194 1851 1177 23 38 1911 NOR2_X1
* cell instance $1195 m0 *1 34.58,71.4
X$1195 23 38 FILLCELL_X4
* cell instance $1196 m0 *1 35.34,71.4
X$1196 23 38 FILLCELL_X1
* cell instance $1197 m0 *1 35.53,71.4
X$1197 1810 1454 1855 23 38 1873 MUX2_X1
* cell instance $1198 m0 *1 36.86,71.4
X$1198 23 38 FILLCELL_X8
* cell instance $1199 m0 *1 38.38,71.4
X$1199 23 38 FILLCELL_X4
* cell instance $1200 m0 *1 39.14,71.4
X$1200 1856 1487 1730 23 38 1895 MUX2_X1
* cell instance $1201 m0 *1 40.47,71.4
X$1201 1856 1454 1825 23 38 1874 MUX2_X1
* cell instance $1202 m0 *1 41.8,71.4
X$1202 23 38 FILLCELL_X8
* cell instance $1203 m0 *1 43.32,71.4
X$1203 23 38 FILLCELL_X4
* cell instance $1204 m0 *1 44.08,71.4
X$1204 23 38 FILLCELL_X1
* cell instance $1205 m0 *1 44.27,71.4
X$1205 1268 23 38 1728 CLKBUF_X3
* cell instance $1206 m0 *1 45.22,71.4
X$1206 23 38 FILLCELL_X8
* cell instance $1207 m0 *1 46.74,71.4
X$1207 23 38 FILLCELL_X2
* cell instance $1208 r0 *1 17.67,71.4
X$1208 23 38 FILLCELL_X4
* cell instance $1209 r0 *1 18.43,71.4
X$1209 23 38 FILLCELL_X1
* cell instance $1210 r0 *1 18.62,71.4
X$1210 1891 893 23 38 1904 NOR2_X1
* cell instance $1211 r0 *1 19.19,71.4
X$1211 1871 1487 1820 23 38 1845 MUX2_X1
* cell instance $1212 r0 *1 20.52,71.4
X$1212 1871 1454 1843 23 38 1872 MUX2_X1
* cell instance $1213 r0 *1 21.85,71.4
X$1213 23 38 FILLCELL_X16
* cell instance $1214 r0 *1 24.89,71.4
X$1214 23 38 FILLCELL_X1
* cell instance $1215 r0 *1 25.08,71.4
X$1215 1794 1454 1821 23 38 1926 MUX2_X1
* cell instance $1216 r0 *1 26.41,71.4
X$1216 23 38 FILLCELL_X8
* cell instance $1217 r0 *1 27.93,71.4
X$1217 23 38 FILLCELL_X4
* cell instance $1218 r0 *1 28.69,71.4
X$1218 23 38 FILLCELL_X1
* cell instance $1219 r0 *1 28.88,71.4
X$1219 23 2979 1823 1850 1795 38 DFF_X1
* cell instance $1220 r0 *1 32.11,71.4
X$1220 23 38 FILLCELL_X2
* cell instance $1221 r0 *1 32.49,71.4
X$1221 23 38 FILLCELL_X1
* cell instance $1222 r0 *1 32.68,71.4
X$1222 1795 23 38 3149 INV_X1
* cell instance $1223 r0 *1 33.06,71.4
X$1223 23 2975 1855 1894 1795 38 DFF_X1
* cell instance $1224 r0 *1 36.29,71.4
X$1224 23 38 FILLCELL_X2
* cell instance $1225 r0 *1 36.67,71.4
X$1225 23 38 FILLCELL_X1
* cell instance $1226 r0 *1 36.86,71.4
X$1226 1873 1105 23 38 1910 NOR2_X1
* cell instance $1227 r0 *1 37.43,71.4
X$1227 23 38 FILLCELL_X1
* cell instance $1228 r0 *1 37.62,71.4
X$1228 23 2982 1856 1895 1639 38 DFF_X1
* cell instance $1229 r0 *1 40.85,71.4
X$1229 23 38 FILLCELL_X1
* cell instance $1230 r0 *1 41.04,71.4
X$1230 1874 1105 23 38 1998 NOR2_X1
* cell instance $1231 r0 *1 41.61,71.4
X$1231 23 38 FILLCELL_X1
* cell instance $1232 r0 *1 41.8,71.4
X$1232 1912 1446 1813 23 38 1930 MUX2_X1
* cell instance $1233 r0 *1 43.13,71.4
X$1233 23 38 FILLCELL_X16
* cell instance $1234 r0 *1 46.17,71.4
X$1234 23 38 FILLCELL_X1
* cell instance $1235 r0 *1 46.36,71.4
X$1235 1949 23 38 1208 CLKBUF_X3
* cell instance $1236 m0 *1 47.31,71.4
X$1236 1859 1105 23 38 1875 NOR2_X1
* cell instance $1237 m0 *1 47.12,71.4
X$1237 23 38 FILLCELL_X1
* cell instance $1238 m0 *1 47.88,71.4
X$1238 23 2726 1876 1877 1735 38 DFF_X1
* cell instance $1239 m0 *1 51.11,71.4
X$1239 23 38 FILLCELL_X2
* cell instance $1240 r0 *1 47.31,71.4
X$1240 23 38 FILLCELL_X4
* cell instance $1241 r0 *1 48.07,71.4
X$1241 1876 1487 1767 23 38 1877 MUX2_X1
* cell instance $1242 r0 *1 49.4,71.4
X$1242 23 2886 1878 1898 1735 38 DFF_X1
* cell instance $1243 m0 *1 52.82,71.4
X$1243 1786 1177 23 38 1934 NOR2_X1
* cell instance $1244 m0 *1 51.49,71.4
X$1244 1878 1488 1767 23 38 1898 MUX2_X1
* cell instance $1245 m0 *1 53.39,71.4
X$1245 1863 1765 1862 38 23 1866 OAI21_X2
* cell instance $1246 m0 *1 54.72,71.4
X$1246 1743 1865 1864 1804 1860 38 23 1861 OAI221_X1
* cell instance $1247 m0 *1 55.86,71.4
X$1247 1797 1728 23 38 1862 NAND2_X1
* cell instance $1248 m0 *1 56.43,71.4
X$1248 1797 1638 23 38 1860 NAND2_X1
* cell instance $1249 m0 *1 57,71.4
X$1249 23 38 FILLCELL_X8
* cell instance $1250 m0 *1 58.52,71.4
X$1250 23 38 FILLCELL_X4
* cell instance $1251 m0 *1 59.28,71.4
X$1251 23 38 FILLCELL_X2
* cell instance $1252 r0 *1 52.63,71.4
X$1252 1876 1454 1878 23 38 1899 MUX2_X1
* cell instance $1253 r0 *1 53.96,71.4
X$1253 1899 1105 23 38 1879 NOR2_X1
* cell instance $1254 r0 *1 54.53,71.4
X$1254 1318 23 38 1629 CLKBUF_X3
* cell instance $1255 r0 *1 55.48,71.4
X$1255 1478 23 38 1636 CLKBUF_X3
* cell instance $1256 r0 *1 56.43,71.4
X$1256 23 38 FILLCELL_X16
* cell instance $1257 r0 *1 59.14,71.4
X$1257 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $1258 r0 *1 59.14,71.4
X$1258 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $1259 r0 *1 59.14,71.4
X$1259 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $1260 r0 *1 59.47,71.4
X$1260 23 2914 1880 1901 1684 38 DFF_X1
* cell instance $1261 m0 *1 59.85,71.4
X$1261 23 2585 1826 1858 1684 38 DFF_X1
* cell instance $1262 m0 *1 59.66,71.4
X$1262 23 38 FILLCELL_X1
* cell instance $1263 m0 *1 63.08,71.4
X$1263 1826 441 1561 23 38 1858 MUX2_X1
* cell instance $1264 m0 *1 64.41,71.4
X$1264 23 38 FILLCELL_X2
* cell instance $1265 r0 *1 62.7,71.4
X$1265 1826 1454 1880 23 38 1900 MUX2_X1
* cell instance $1266 r0 *1 64.03,71.4
X$1266 1561 51 1913 23 38 1931 MUX2_X1
* cell instance $1267 m0 *1 68.02,71.4
X$1267 1561 260 1853 23 38 1827 MUX2_X1
* cell instance $1268 m0 *1 64.79,71.4
X$1268 23 2582 1853 1827 1684 38 DFF_X1
* cell instance $1269 m0 *1 69.35,71.4
X$1269 23 38 FILLCELL_X4
* cell instance $1270 m0 *1 70.11,71.4
X$1270 23 38 FILLCELL_X1
* cell instance $1271 m0 *1 70.3,71.4
X$1271 1335 240 1828 23 38 1814 MUX2_X1
* cell instance $1272 m0 *1 71.63,71.4
X$1272 23 38 FILLCELL_X16
* cell instance $1273 m0 *1 74.67,71.4
X$1273 1829 1454 1883 23 38 1830 MUX2_X1
* cell instance $1274 m0 *1 76,71.4
X$1274 23 38 FILLCELL_X8
* cell instance $1275 m0 *1 77.52,71.4
X$1275 23 38 FILLCELL_X1
* cell instance $1276 m0 *1 77.71,71.4
X$1276 1892 1605 23 38 1844 NOR2_X1
* cell instance $1277 m0 *1 78.28,71.4
X$1277 23 38 FILLCELL_X4
* cell instance $1278 m0 *1 79.04,71.4
X$1278 23 38 FILLCELL_X2
* cell instance $1279 r0 *1 65.36,71.4
X$1279 23 38 FILLCELL_X1
* cell instance $1280 r0 *1 65.55,71.4
X$1280 1900 1105 23 38 1881 NOR2_X1
* cell instance $1281 r0 *1 66.12,71.4
X$1281 23 38 FILLCELL_X1
* cell instance $1282 r0 *1 66.31,71.4
X$1282 1897 1605 23 38 1882 NOR2_X1
* cell instance $1283 r0 *1 68.21,71.4
X$1283 23 38 FILLCELL_X2
* cell instance $1284 r0 *1 68.59,71.4
X$1284 1853 414 1828 23 38 1800 MUX2_X1
* cell instance $1285 r0 *1 69.92,71.4
X$1285 23 38 FILLCELL_X8
* cell instance $1286 r0 *1 71.44,71.4
X$1286 23 38 FILLCELL_X4
* cell instance $1287 r0 *1 72.2,71.4
X$1287 23 38 FILLCELL_X1
* cell instance $1288 r0 *1 72.39,71.4
X$1288 23 3102 1883 1893 1648 38 DFF_X1
* cell instance $1289 r0 *1 75.62,71.4
X$1289 1883 373 1770 23 38 1893 MUX2_X1
* cell instance $1290 r0 *1 76.95,71.4
X$1290 23 38 FILLCELL_X4
* cell instance $1291 r0 *1 77.71,71.4
X$1291 1770 51 1885 23 38 1884 MUX2_X1
* cell instance $1292 r0 *1 79.04,71.4
X$1292 23 38 FILLCELL_X1
* cell instance $1293 r0 *1 79.23,71.4
X$1293 1885 1099 1916 23 38 1892 MUX2_X1
* cell instance $1294 m0 *1 79.61,71.4
X$1294 1770 260 1833 23 38 1839 MUX2_X1
* cell instance $1295 m0 *1 79.42,71.4
X$1295 23 38 FILLCELL_X1
* cell instance $1296 m0 *1 80.94,71.4
X$1296 23 2676 1833 1839 1648 38 DFF_X1
* cell instance $1297 m0 *1 84.17,71.4
X$1297 23 38 FILLCELL_X2
* cell instance $1298 r0 *1 81.89,71.4
X$1298 23 38 FILLCELL_X2
* cell instance $1299 r0 *1 82.27,71.4
X$1299 1833 414 1887 23 38 1837 MUX2_X1
* cell instance $1300 r0 *1 83.6,71.4
X$1300 23 38 FILLCELL_X4
* cell instance $1301 r0 *1 84.36,71.4
X$1301 23 38 FILLCELL_X2
* cell instance $1302 m0 *1 85.88,71.4
X$1302 23 38 FILLCELL_X2
* cell instance $1303 m0 *1 84.55,71.4
X$1303 1111 240 1887 23 38 1888 MUX2_X1
* cell instance $1304 r0 *1 84.74,71.4
X$1304 23 2858 1887 1888 1714 38 DFF_X1
* cell instance $1305 m0 *1 87.02,71.4
X$1305 23 38 FILLCELL_X32
* cell instance $1306 m0 *1 86.26,71.4
X$1306 1111 23 38 1770 BUF_X2
* cell instance $1307 m0 *1 93.1,71.4
X$1307 23 38 FILLCELL_X16
* cell instance $1308 m0 *1 96.14,71.4
X$1308 23 38 FILLCELL_X4
* cell instance $1309 m0 *1 96.9,71.4
X$1309 23 38 FILLCELL_X1
* cell instance $1310 r180 *1 97.28,71.4
X$1310 23 38 23 38 TAPCELL_X1
* cell instance $1311 r0 *1 87.97,71.4
X$1311 1268 23 38 1230 CLKBUF_X3
* cell instance $1312 r0 *1 88.92,71.4
X$1312 1920 23 38 1268 BUF_X2
* cell instance $1313 r0 *1 89.68,71.4
X$1313 23 38 FILLCELL_X16
* cell instance $1314 r0 *1 92.72,71.4
X$1314 23 38 FILLCELL_X4
* cell instance $1315 r0 *1 93.48,71.4
X$1315 23 38 FILLCELL_X2
* cell instance $1316 r0 *1 93.86,71.4
X$1316 23 38 FILLCELL_X1
* cell instance $1317 r0 *1 94.05,71.4
X$1317 1889 23 38 1335 BUF_X2
* cell instance $1318 r0 *1 94.81,71.4
X$1318 1921 23 38 1111 BUF_X2
* cell instance $1319 r0 *1 95.57,71.4
X$1319 23 38 FILLCELL_X8
* cell instance $1320 m90 *1 97.28,71.4
X$1320 23 38 23 38 TAPCELL_X1
* cell instance $1321 m0 *1 83.98,93.8
X$1321 2456 2483 2457 23 38 2484 MUX2_X1
* cell instance $1322 m0 *1 83.79,93.8
X$1322 23 38 FILLCELL_X1
* cell instance $1323 m0 *1 85.31,93.8
X$1323 23 38 FILLCELL_X1
* cell instance $1324 m0 *1 85.5,93.8
X$1324 2412 2057 38 23 2485 AND2_X1
* cell instance $1325 m0 *1 86.26,93.8
X$1325 2058 23 38 2373 CLKBUF_X3
* cell instance $1326 m0 *1 87.21,93.8
X$1326 2485 2379 2487 23 38 2486 MUX2_X1
* cell instance $1327 m0 *1 88.54,93.8
X$1327 1319 2412 23 38 2487 NOR2_X1
* cell instance $1328 m0 *1 89.11,93.8
X$1328 23 38 FILLCELL_X1
* cell instance $1329 m0 *1 89.3,93.8
X$1329 23 2828 2414 2459 2373 38 DFF_X1
* cell instance $1330 m0 *1 92.53,93.8
X$1330 23 38 FILLCELL_X16
* cell instance $1331 m0 *1 95.57,93.8
X$1331 23 38 FILLCELL_X8
* cell instance $1332 r180 *1 97.28,93.8
X$1332 23 38 23 38 TAPCELL_X1
* cell instance $1333 r0 *1 83.79,93.8
X$1333 23 3123 2411 2484 2373 38 DFF_X1
* cell instance $1334 r0 *1 87.02,93.8
X$1334 23 38 FILLCELL_X2
* cell instance $1335 r0 *1 87.4,93.8
X$1335 23 3125 2412 2486 2373 38 DFF_X1
* cell instance $1336 r0 *1 90.63,93.8
X$1336 23 38 FILLCELL_X32
* cell instance $1337 r0 *1 96.71,93.8
X$1337 23 38 FILLCELL_X2
* cell instance $1338 m90 *1 97.28,93.8
X$1338 23 38 23 38 TAPCELL_X1
* cell instance $1339 m0 *1 4.94,65.8
X$1339 1598 1346 1746 23 38 1709 MUX2_X1
* cell instance $1340 m0 *1 1.71,65.8
X$1340 23 2607 1689 1710 1556 38 DFF_X1
* cell instance $1341 m0 *1 6.27,65.8
X$1341 23 38 FILLCELL_X1
* cell instance $1342 m0 *1 6.46,65.8
X$1342 1689 1358 1746 23 38 1712 MUX2_X1
* cell instance $1343 m0 *1 7.79,65.8
X$1343 1718 23 38 1688 BUF_X1
* cell instance $1344 m0 *1 8.36,65.8
X$1344 23 38 FILLCELL_X8
* cell instance $1345 m0 *1 9.88,65.8
X$1345 23 38 FILLCELL_X2
* cell instance $1346 m0 *1 1.33,65.8
X$1346 23 38 FILLCELL_X2
* cell instance $1347 m0 *1 1.14,65.8
X$1347 23 38 23 38 TAPCELL_X1
* cell instance $1348 r0 *1 1.14,65.8
X$1348 23 38 23 38 TAPCELL_X1
* cell instance $1349 r0 *1 1.33,65.8
X$1349 23 38 FILLCELL_X4
* cell instance $1350 r0 *1 2.09,65.8
X$1350 23 38 FILLCELL_X2
* cell instance $1351 r0 *1 2.47,65.8
X$1351 23 38 FILLCELL_X1
* cell instance $1352 r0 *1 2.66,65.8
X$1352 23 3003 1746 1709 1556 38 DFF_X1
* cell instance $1353 r0 *1 3.14,65.8
X$1353 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $1354 r0 *1 3.14,65.8
X$1354 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $1355 r0 *1 3.14,65.8
X$1355 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $1356 r0 *1 5.89,65.8
X$1356 1486 23 38 1556 CLKBUF_X3
* cell instance $1357 r0 *1 6.84,65.8
X$1357 23 38 FILLCELL_X1
* cell instance $1358 r0 *1 7.03,65.8
X$1358 23 3004 1717 1747 1556 38 DFF_X1
* cell instance $1359 r0 *1 10.26,65.8
X$1359 23 2943 1762 1779 1635 38 DFF_X1
* cell instance $1360 m0 *1 10.45,65.8
X$1360 1712 1535 23 38 1691 NOR2_X1
* cell instance $1361 m0 *1 10.26,65.8
X$1361 23 38 FILLCELL_X1
* cell instance $1362 m0 *1 11.02,65.8
X$1362 1425 1749 1778 548 1691 1690 23 38 1720 OAI33_X1
* cell instance $1363 m0 *1 12.35,65.8
X$1363 23 38 FILLCELL_X1
* cell instance $1364 m0 *1 12.54,65.8
X$1364 1762 627 1692 23 38 1719 MUX2_X1
* cell instance $1365 m0 *1 13.87,65.8
X$1365 1692 1289 1532 23 38 1721 MUX2_X1
* cell instance $1366 m0 *1 15.2,65.8
X$1366 23 38 FILLCELL_X8
* cell instance $1367 m0 *1 16.72,65.8
X$1367 23 38 FILLCELL_X4
* cell instance $1368 m0 *1 17.48,65.8
X$1368 23 38 FILLCELL_X2
* cell instance $1369 r0 *1 13.49,65.8
X$1369 1719 381 23 38 1749 NOR2_X1
* cell instance $1370 r0 *1 14.06,65.8
X$1370 23 2952 1692 1721 1635 38 DFF_X1
* cell instance $1371 r0 *1 17.29,65.8
X$1371 23 38 FILLCELL_X4
* cell instance $1372 m0 *1 18.05,65.8
X$1372 23 2574 1724 1722 1693 38 DFF_X1
* cell instance $1373 m0 *1 17.86,65.8
X$1373 23 38 FILLCELL_X1
* cell instance $1374 m0 *1 21.28,65.8
X$1374 23 38 FILLCELL_X4
* cell instance $1375 m0 *1 22.04,65.8
X$1375 23 38 FILLCELL_X1
* cell instance $1376 m0 *1 22.23,65.8
X$1376 23 2626 1666 1716 1693 38 DFF_X1
* cell instance $1377 m0 *1 25.46,65.8
X$1377 23 2788 1694 1752 1693 38 DFF_X1
* cell instance $1378 m0 *1 28.69,65.8
X$1378 23 38 FILLCELL_X8
* cell instance $1379 m0 *1 30.21,65.8
X$1379 23 38 FILLCELL_X1
* cell instance $1380 m0 *1 30.4,65.8
X$1380 23 2823 1637 1696 1262 38 DFF_X1
* cell instance $1381 m0 *1 33.63,65.8
X$1381 23 38 FILLCELL_X8
* cell instance $1382 m0 *1 35.15,65.8
X$1382 23 2812 1729 1758 1795 38 DFF_X1
* cell instance $1383 m0 *1 38.38,65.8
X$1383 23 2829 1731 1697 1639 38 DFF_X1
* cell instance $1384 m0 *1 41.61,65.8
X$1384 23 38 FILLCELL_X8
* cell instance $1385 m0 *1 43.13,65.8
X$1385 23 38 FILLCELL_X2
* cell instance $1386 r0 *1 18.05,65.8
X$1386 1724 1488 1791 23 38 1722 MUX2_X1
* cell instance $1387 r0 *1 19.38,65.8
X$1387 23 38 FILLCELL_X2
* cell instance $1388 r0 *1 19.76,65.8
X$1388 23 38 FILLCELL_X1
* cell instance $1389 r0 *1 19.95,65.8
X$1389 1723 994 1724 23 38 1780 MUX2_X1
* cell instance $1390 r0 *1 21.28,65.8
X$1390 23 2994 1723 1781 1693 38 DFF_X1
* cell instance $1391 r0 *1 24.51,65.8
X$1391 1486 23 38 1693 CLKBUF_X3
* cell instance $1392 r0 *1 25.46,65.8
X$1392 23 38 FILLCELL_X2
* cell instance $1393 r0 *1 25.84,65.8
X$1393 1764 1434 1725 23 38 1763 MUX2_X1
* cell instance $1394 r0 *1 27.17,65.8
X$1394 23 38 FILLCELL_X1
* cell instance $1395 r0 *1 27.36,65.8
X$1395 1694 1446 1725 23 38 1752 MUX2_X1
* cell instance $1396 r0 *1 28.69,65.8
X$1396 23 38 FILLCELL_X2
* cell instance $1397 r0 *1 29.07,65.8
X$1397 23 38 FILLCELL_X1
* cell instance $1398 r0 *1 29.26,65.8
X$1398 1726 1720 1629 1157 1727 38 23 1695 OAI221_X1
* cell instance $1399 r0 *1 30.4,65.8
X$1399 1726 1720 1511 1787 38 23 1754 OAI22_X2
* cell instance $1400 r0 *1 32.11,65.8
X$1400 1754 1765 1757 38 23 1718 OAI21_X2
* cell instance $1401 r0 *1 33.44,65.8
X$1401 1637 1728 23 38 1757 NAND2_X1
* cell instance $1402 r0 *1 34.01,65.8
X$1402 23 38 FILLCELL_X8
* cell instance $1403 r0 *1 35.53,65.8
X$1403 23 38 FILLCELL_X4
* cell instance $1404 r0 *1 36.29,65.8
X$1404 1729 1434 1730 23 38 1758 MUX2_X1
* cell instance $1405 r0 *1 37.62,65.8
X$1405 1731 1446 1730 23 38 1697 MUX2_X1
* cell instance $1406 r0 *1 38.95,65.8
X$1406 1731 1184 1729 23 38 1732 MUX2_X1
* cell instance $1407 r0 *1 40.28,65.8
X$1407 23 38 FILLCELL_X8
* cell instance $1408 r0 *1 41.8,65.8
X$1408 23 38 FILLCELL_X2
* cell instance $1409 r0 *1 42.18,65.8
X$1409 23 2984 1733 1766 1639 38 DFF_X1
* cell instance $1410 m0 *1 44.08,65.8
X$1410 23 38 FILLCELL_X16
* cell instance $1411 m0 *1 43.51,65.8
X$1411 1639 23 38 CLKBUF_X1
* cell instance $1412 m0 *1 47.12,65.8
X$1412 23 38 FILLCELL_X4
* cell instance $1413 m0 *1 47.88,65.8
X$1413 1734 1446 1767 23 38 1698 MUX2_X1
* cell instance $1414 m0 *1 49.21,65.8
X$1414 23 38 FILLCELL_X8
* cell instance $1415 m0 *1 50.73,65.8
X$1415 23 38 FILLCELL_X4
* cell instance $1416 m0 *1 51.49,65.8
X$1416 23 2601 1677 1760 1735 38 DFF_X1
* cell instance $1417 m0 *1 54.72,65.8
X$1417 1425 1679 1761 225 1699 1700 23 38 1736 OAI33_X1
* cell instance $1418 m0 *1 56.05,65.8
X$1418 1701 1483 23 38 1700 NOR2_X1
* cell instance $1419 m0 *1 56.62,65.8
X$1419 1587 1480 1702 23 38 1642 MUX2_X1
* cell instance $1420 m0 *1 57.95,65.8
X$1420 23 38 FILLCELL_X1
* cell instance $1421 m0 *1 58.14,65.8
X$1421 1737 1373 1702 23 38 1701 MUX2_X1
* cell instance $1422 m0 *1 59.47,65.8
X$1422 23 38 FILLCELL_X2
* cell instance $1423 r0 *1 45.41,65.8
X$1423 23 38 FILLCELL_X4
* cell instance $1424 r0 *1 46.17,65.8
X$1424 1733 1454 1782 23 38 1859 MUX2_X1
* cell instance $1425 r0 *1 47.5,65.8
X$1425 23 38 FILLCELL_X1
* cell instance $1426 r0 *1 47.69,65.8
X$1426 23 3121 1734 1698 1639 38 DFF_X1
* cell instance $1427 r0 *1 50.92,65.8
X$1427 1734 541 1784 23 38 1786 MUX2_X1
* cell instance $1428 r0 *1 52.25,65.8
X$1428 23 38 FILLCELL_X1
* cell instance $1429 r0 *1 52.44,65.8
X$1429 1392 23 38 1735 CLKBUF_X3
* cell instance $1430 r0 *1 53.39,65.8
X$1430 23 38 FILLCELL_X4
* cell instance $1431 r0 *1 54.15,65.8
X$1431 23 38 FILLCELL_X1
* cell instance $1432 r0 *1 54.34,65.8
X$1432 1641 1736 1629 1506 1727 38 23 1864 OAI221_X1
* cell instance $1433 r0 *1 55.48,65.8
X$1433 23 38 FILLCELL_X2
* cell instance $1434 r0 *1 55.86,65.8
X$1434 23 38 FILLCELL_X1
* cell instance $1435 r0 *1 56.05,65.8
X$1435 1587 1493 1737 23 38 1768 MUX2_X1
* cell instance $1436 r0 *1 57.38,65.8
X$1436 23 38 FILLCELL_X8
* cell instance $1437 r0 *1 58.9,65.8
X$1437 23 38 FILLCELL_X4
* cell instance $1438 r0 *1 59.14,65.8
X$1438 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $1439 r0 *1 59.14,65.8
X$1439 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $1440 r0 *1 59.14,65.8
X$1440 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $1441 r0 *1 59.66,65.8
X$1441 23 38 FILLCELL_X1
* cell instance $1442 m0 *1 60.04,65.8
X$1442 23 2584 1739 1703 1684 38 DFF_X1
* cell instance $1443 m0 *1 59.85,65.8
X$1443 23 38 FILLCELL_X1
* cell instance $1444 m0 *1 63.27,65.8
X$1444 1739 520 1561 23 38 1703 MUX2_X1
* cell instance $1445 m0 *1 64.6,65.8
X$1445 23 38 FILLCELL_X8
* cell instance $1446 m0 *1 66.12,65.8
X$1446 23 38 FILLCELL_X4
* cell instance $1447 m0 *1 66.88,65.8
X$1447 1704 88 1561 23 38 1759 MUX2_X1
* cell instance $1448 m0 *1 68.21,65.8
X$1448 23 38 FILLCELL_X4
* cell instance $1449 m0 *1 68.97,65.8
X$1449 1392 23 38 1644 CLKBUF_X3
* cell instance $1450 m0 *1 69.92,65.8
X$1450 1644 23 38 3141 INV_X1
* cell instance $1451 m0 *1 70.3,65.8
X$1451 23 38 FILLCELL_X8
* cell instance $1452 m0 *1 71.82,65.8
X$1452 23 38 FILLCELL_X2
* cell instance $1453 r0 *1 59.85,65.8
X$1453 23 2925 1738 1788 1684 38 DFF_X1
* cell instance $1454 r0 *1 63.08,65.8
X$1454 1738 541 1739 23 38 1769 MUX2_X1
* cell instance $1455 r0 *1 64.41,65.8
X$1455 23 38 FILLCELL_X8
* cell instance $1456 r0 *1 65.93,65.8
X$1456 23 2906 1704 1759 1644 38 DFF_X1
* cell instance $1457 r0 *1 69.16,65.8
X$1457 23 38 FILLCELL_X8
* cell instance $1458 r0 *1 70.68,65.8
X$1458 23 38 FILLCELL_X1
* cell instance $1459 r0 *1 70.87,65.8
X$1459 1300 38 1305 23 BUF_X4
* cell instance $1460 r0 *1 72.2,65.8
X$1460 23 38 FILLCELL_X4
* cell instance $1461 m0 *1 73.15,65.8
X$1461 23 38 FILLCELL_X8
* cell instance $1462 m0 *1 72.2,65.8
X$1462 1318 23 38 1241 CLKBUF_X3
* cell instance $1463 m0 *1 74.67,65.8
X$1463 23 38 FILLCELL_X1
* cell instance $1464 m0 *1 74.86,65.8
X$1464 23 2681 1610 1715 1336 38 DFF_X1
* cell instance $1465 m0 *1 78.09,65.8
X$1465 23 2623 1611 1753 1648 38 DFF_X1
* cell instance $1466 m0 *1 81.32,65.8
X$1466 1519 23 38 1239 CLKBUF_X3
* cell instance $1467 m0 *1 82.27,65.8
X$1467 23 38 FILLCELL_X16
* cell instance $1468 m0 *1 85.31,65.8
X$1468 23 38 FILLCELL_X2
* cell instance $1469 r0 *1 72.96,65.8
X$1469 23 38 FILLCELL_X1
* cell instance $1470 r0 *1 73.15,65.8
X$1470 1392 23 38 3138 INV_X2
* cell instance $1471 r0 *1 73.72,65.8
X$1471 1802 520 1770 23 38 1771 MUX2_X1
* cell instance $1472 r0 *1 75.05,65.8
X$1472 434 23 38 1392 CLKBUF_X3
* cell instance $1473 r0 *1 76,65.8
X$1473 23 38 FILLCELL_X2
* cell instance $1474 r0 *1 76.38,65.8
X$1474 23 38 FILLCELL_X1
* cell instance $1475 r0 *1 76.57,65.8
X$1475 23 2903 1755 1756 1336 38 DFF_X1
* cell instance $1476 r0 *1 79.8,65.8
X$1476 1478 23 38 1228 CLKBUF_X3
* cell instance $1477 r0 *1 80.75,65.8
X$1477 23 38 FILLCELL_X4
* cell instance $1478 r0 *1 81.51,65.8
X$1478 23 38 FILLCELL_X2
* cell instance $1479 r0 *1 81.89,65.8
X$1479 23 2880 1740 1751 1648 38 DFF_X1
* cell instance $1480 r0 *1 85.12,65.8
X$1480 23 38 FILLCELL_X2
* cell instance $1481 r0 *1 85.5,65.8
X$1481 1740 130 1770 23 38 1751 MUX2_X1
* cell instance $1482 m0 *1 85.88,65.8
X$1482 1773 1650 23 38 1713 NOR2_X1
* cell instance $1483 m0 *1 85.69,65.8
X$1483 23 38 FILLCELL_X1
* cell instance $1484 m0 *1 86.45,65.8
X$1484 23 38 FILLCELL_X8
* cell instance $1485 m0 *1 87.97,65.8
X$1485 23 38 FILLCELL_X2
* cell instance $1486 r0 *1 86.83,65.8
X$1486 23 38 FILLCELL_X2
* cell instance $1487 r0 *1 87.21,65.8
X$1487 23 38 FILLCELL_X1
* cell instance $1488 r0 *1 87.4,65.8
X$1488 1741 188 1750 23 38 1705 MUX2_X1
* cell instance $1489 m0 *1 88.92,65.8
X$1489 23 38 FILLCELL_X2
* cell instance $1490 m0 *1 88.35,65.8
X$1490 1705 1579 23 38 1651 NOR2_X1
* cell instance $1491 r0 *1 88.73,65.8
X$1491 23 2912 1750 1774 1714 38 DFF_X1
* cell instance $1492 m0 *1 90.44,65.8
X$1492 23 38 FILLCELL_X16
* cell instance $1493 m0 *1 89.3,65.8
X$1493 1706 1652 1241 1506 1224 38 23 1711 OAI221_X1
* cell instance $1494 m0 *1 93.48,65.8
X$1494 23 38 FILLCELL_X2
* cell instance $1495 r0 *1 91.96,65.8
X$1495 1228 1742 23 38 1777 NAND2_X1
* cell instance $1496 r0 *1 92.53,65.8
X$1496 23 38 FILLCELL_X2
* cell instance $1497 r0 *1 92.91,65.8
X$1497 1743 1748 1707 1226 1744 38 23 1775 OAI221_X1
* cell instance $1498 m0 *1 94.05,65.8
X$1498 1745 1239 23 38 1744 NAND2_X1
* cell instance $1499 m0 *1 93.86,65.8
X$1499 23 38 FILLCELL_X1
* cell instance $1500 m0 *1 94.62,65.8
X$1500 1742 1230 23 38 1708 NAND2_X1
* cell instance $1501 m0 *1 95.19,65.8
X$1501 23 38 FILLCELL_X2
* cell instance $1502 r0 *1 94.05,65.8
X$1502 1228 1745 23 38 1748 NAND2_X1
* cell instance $1503 r0 *1 94.62,65.8
X$1503 23 38 FILLCELL_X8
* cell instance $1504 m0 *1 96.14,65.8
X$1504 23 38 FILLCELL_X4
* cell instance $1505 m0 *1 95.57,65.8
X$1505 1745 1230 23 38 1612 NAND2_X1
* cell instance $1506 m0 *1 96.9,65.8
X$1506 23 38 FILLCELL_X1
* cell instance $1507 r180 *1 97.28,65.8
X$1507 23 38 23 38 TAPCELL_X1
* cell instance $1508 r0 *1 96.14,65.8
X$1508 23 38 FILLCELL_X4
* cell instance $1509 r0 *1 96.9,65.8
X$1509 23 38 FILLCELL_X1
* cell instance $1510 m90 *1 97.28,65.8
X$1510 23 38 23 38 TAPCELL_X1
* cell instance $1511 m0 *1 64.98,96.6
X$1511 2536 23 38 2535 BUF_X1
* cell instance $1512 m0 *1 64.79,96.6
X$1512 23 38 FILLCELL_X1
* cell instance $1513 m0 *1 65.55,96.6
X$1513 23 38 FILLCELL_X2
* cell instance $1514 m0 *1 75.05,96.6
X$1514 2481 23 38 2541 BUF_X1
* cell instance $1515 m0 *1 74.48,96.6
X$1515 1953 23 38 2540 BUF_X1
* cell instance $1516 m0 *1 75.62,96.6
X$1516 2452 23 38 2542 BUF_X1
* cell instance $1517 m0 *1 76.19,96.6
X$1517 2451 23 38 2543 BUF_X1
* cell instance $1518 m0 *1 76.76,96.6
X$1518 2563 23 38 2544 BUF_X1
* cell instance $1519 m0 *1 77.33,96.6
X$1519 23 38 FILLCELL_X1
* cell instance $1520 m0 *1 77.52,96.6
X$1520 2452 2409 23 38 2494 NAND2_X1
* cell instance $1521 m0 *1 78.09,96.6
X$1521 2493 23 38 2545 BUF_X1
* cell instance $1522 m0 *1 78.66,96.6
X$1522 2546 23 38 2547 BUF_X1
* cell instance $1523 m0 *1 79.23,96.6
X$1523 23 38 FILLCELL_X1
* cell instance $1524 m0 *1 79.42,96.6
X$1524 2512 23 38 2548 BUF_X1
* cell instance $1525 m0 *1 79.99,96.6
X$1525 2510 23 38 2546 INV_X1
* cell instance $1526 m0 *1 80.37,96.6
X$1526 23 38 FILLCELL_X1
* cell instance $1527 m0 *1 80.56,96.6
X$1527 1319 2512 23 38 2550 NOR2_X1
* cell instance $1528 m0 *1 81.13,96.6
X$1528 23 38 FILLCELL_X8
* cell instance $1529 m0 *1 82.65,96.6
X$1529 23 38 FILLCELL_X2
* cell instance $1530 m0 *1 66.12,96.6
X$1530 2561 23 38 2538 BUF_X1
* cell instance $1531 m0 *1 65.93,96.6
X$1531 23 38 FILLCELL_X1
* cell instance $1532 m0 *1 66.69,96.6
X$1532 23 38 FILLCELL_X4
* cell instance $1533 m0 *1 67.45,96.6
X$1533 23 38 FILLCELL_X2
* cell instance $1534 m0 *1 88.54,96.6
X$1534 2412 23 38 2555 BUF_X1
* cell instance $1535 m0 *1 87.97,96.6
X$1535 2373 23 38 CLKBUF_X1
* cell instance $1536 m0 *1 89.11,96.6
X$1536 23 38 FILLCELL_X8
* cell instance $1537 m0 *1 90.63,96.6
X$1537 23 38 FILLCELL_X4
* cell instance $1538 m0 *1 91.39,96.6
X$1538 2414 23 38 2556 BUF_X1
* cell instance $1539 m0 *1 91.96,96.6
X$1539 23 38 FILLCELL_X16
* cell instance $1540 m0 *1 95,96.6
X$1540 23 38 FILLCELL_X8
* cell instance $1541 m0 *1 96.52,96.6
X$1541 23 38 FILLCELL_X2
* cell instance $1542 m0 *1 53.58,96.6
X$1542 1866 23 38 2528 BUF_X1
* cell instance $1543 m0 *1 53.39,96.6
X$1543 23 38 FILLCELL_X1
* cell instance $1544 m0 *1 54.15,96.6
X$1544 23 38 FILLCELL_X4
* cell instance $1545 m0 *1 54.91,96.6
X$1545 23 38 FILLCELL_X1
* cell instance $1546 m0 *1 55.1,96.6
X$1546 2110 23 38 2529 BUF_X1
* cell instance $1547 m0 *1 55.67,96.6
X$1547 23 38 FILLCELL_X4
* cell instance $1548 m0 *1 56.43,96.6
X$1548 23 38 FILLCELL_X2
* cell instance $1549 m0 *1 83.6,96.6
X$1549 2411 23 38 2552 BUF_X1
* cell instance $1550 m0 *1 83.03,96.6
X$1550 2192 23 38 2551 BUF_X1
* cell instance $1551 m0 *1 84.17,96.6
X$1551 2059 23 38 2553 BUF_X1
* cell instance $1552 m0 *1 84.74,96.6
X$1552 2369 23 38 2554 BUF_X1
* cell instance $1553 m0 *1 85.31,96.6
X$1553 23 38 FILLCELL_X8
* cell instance $1554 m0 *1 86.83,96.6
X$1554 23 38 FILLCELL_X4
* cell instance $1555 m0 *1 87.59,96.6
X$1555 23 38 FILLCELL_X2
* cell instance $1556 m0 *1 57,96.6
X$1556 2530 23 38 2151 BUF_X1
* cell instance $1557 m0 *1 56.81,96.6
X$1557 23 38 FILLCELL_X1
* cell instance $1558 m0 *1 57.57,96.6
X$1558 23 38 FILLCELL_X4
* cell instance $1559 m0 *1 58.33,96.6
X$1559 23 38 FILLCELL_X2
* cell instance $1560 m0 *1 13.3,96.6
X$1560 2515 23 38 2199 BUF_X1
* cell instance $1561 m0 *1 13.11,96.6
X$1561 23 38 FILLCELL_X1
* cell instance $1562 m0 *1 13.87,96.6
X$1562 23 38 FILLCELL_X4
* cell instance $1563 m0 *1 14.63,96.6
X$1563 2516 23 38 2217 BUF_X1
* cell instance $1564 m0 *1 15.2,96.6
X$1564 23 38 FILLCELL_X32
* cell instance $1565 m0 *1 21.28,96.6
X$1565 23 38 FILLCELL_X32
* cell instance $1566 m0 *1 27.36,96.6
X$1566 23 38 FILLCELL_X8
* cell instance $1567 m0 *1 28.88,96.6
X$1567 23 38 FILLCELL_X4
* cell instance $1568 m0 *1 29.64,96.6
X$1568 2517 23 38 2218 BUF_X1
* cell instance $1569 m0 *1 30.21,96.6
X$1569 2169 23 38 2518 BUF_X1
* cell instance $1570 m0 *1 30.78,96.6
X$1570 2304 23 38 2519 BUF_X1
* cell instance $1571 m0 *1 31.35,96.6
X$1571 1973 23 38 2520 BUF_X1
* cell instance $1572 m0 *1 31.92,96.6
X$1572 1909 23 38 2355 CLKBUF_X3
* cell instance $1573 m0 *1 32.87,96.6
X$1573 23 38 FILLCELL_X1
* cell instance $1574 m0 *1 33.06,96.6
X$1574 23 2643 2505 2521 2355 38 DFF_X1
* cell instance $1575 m0 *1 36.29,96.6
X$1575 23 38 FILLCELL_X2
* cell instance $1576 r0 *1 15.39,1.4
X$1576 23 38 FILLCELL_X16
* cell instance $1577 r0 *1 18.43,1.4
X$1577 23 38 FILLCELL_X2
* cell instance $1578 m0 *1 39.9,96.6
X$1578 23 2638 2558 2557 2333 38 DFF_X1
* cell instance $1579 m0 *1 39.71,96.6
X$1579 23 38 FILLCELL_X1
* cell instance $1580 m0 *1 43.13,96.6
X$1580 23 38 FILLCELL_X16
* cell instance $1581 m0 *1 46.17,96.6
X$1581 23 38 FILLCELL_X8
* cell instance $1582 m0 *1 47.69,96.6
X$1582 23 38 FILLCELL_X4
* cell instance $1583 m0 *1 48.45,96.6
X$1583 23 2721 2506 2559 2316 38 DFF_X1
* cell instance $1584 m0 *1 51.68,96.6
X$1584 2183 23 38 2527 BUF_X1
* cell instance $1585 m0 *1 52.25,96.6
X$1585 23 38 FILLCELL_X4
* cell instance $1586 m0 *1 53.01,96.6
X$1586 23 38 FILLCELL_X2
* cell instance $1587 m0 *1 28.12,91
X$1587 23 2650 2356 2354 2355 38 DFF_X1
* cell instance $1588 m0 *1 27.93,91
X$1588 23 38 FILLCELL_X1
* cell instance $1589 m0 *1 31.35,91
X$1589 23 38 FILLCELL_X16
* cell instance $1590 m0 *1 34.39,91
X$1590 23 38 FILLCELL_X4
* cell instance $1591 m0 *1 35.15,91
X$1591 23 38 FILLCELL_X2
* cell instance $1592 r0 *1 27.93,91
X$1592 2441 1373 2440 23 38 2467 MUX2_X1
* cell instance $1593 r0 *1 29.26,91
X$1593 23 38 FILLCELL_X8
* cell instance $1594 r0 *1 30.78,91
X$1594 23 38 FILLCELL_X2
* cell instance $1595 r0 *1 31.16,91
X$1595 2467 1483 23 38 2468 NOR2_X1
* cell instance $1596 r0 *1 31.73,91
X$1596 23 38 FILLCELL_X4
* cell instance $1597 r0 *1 32.49,91
X$1597 23 38 FILLCELL_X2
* cell instance $1598 r0 *1 32.87,91
X$1598 2442 1535 23 38 2357 NOR2_X1
* cell instance $1599 r0 *1 33.44,91
X$1599 23 38 FILLCELL_X16
* cell instance $1600 m0 *1 36.86,91
X$1600 2358 627 2331 23 38 2424 MUX2_X1
* cell instance $1601 m0 *1 35.53,91
X$1601 2358 1403 1730 23 38 2386 MUX2_X1
* cell instance $1602 m0 *1 38.19,91
X$1602 2424 1579 23 38 2390 NOR2_X1
* cell instance $1603 m0 *1 38.76,91
X$1603 23 38 FILLCELL_X4
* cell instance $1604 m0 *1 39.52,91
X$1604 2359 1535 23 38 2360 NOR2_X1
* cell instance $1605 m0 *1 40.09,91
X$1605 23 38 FILLCELL_X1
* cell instance $1606 m0 *1 40.28,91
X$1606 1425 2390 2425 548 2360 2399 23 38 2013 OAI33_X1
* cell instance $1607 m0 *1 41.61,91
X$1607 2426 1483 23 38 2399 NOR2_X1
* cell instance $1608 m0 *1 42.18,91
X$1608 23 38 FILLCELL_X4
* cell instance $1609 m0 *1 42.94,91
X$1609 23 38 FILLCELL_X2
* cell instance $1610 r0 *1 36.48,91
X$1610 23 38 FILLCELL_X8
* cell instance $1611 r0 *1 38,91
X$1611 23 38 FILLCELL_X4
* cell instance $1612 r0 *1 38.76,91
X$1612 23 38 FILLCELL_X2
* cell instance $1613 r0 *1 39.14,91
X$1613 23 3070 2443 2469 2333 38 DFF_X1
* cell instance $1614 r0 *1 42.37,91
X$1614 1909 23 38 2333 CLKBUF_X3
* cell instance $1615 r0 *1 43.32,91
X$1615 23 38 FILLCELL_X8
* cell instance $1616 m0 *1 43.89,91
X$1616 23 38 FILLCELL_X8
* cell instance $1617 m0 *1 43.32,91
X$1617 2361 1650 23 38 2425 NOR2_X1
* cell instance $1618 m0 *1 45.41,91
X$1618 23 38 FILLCELL_X1
* cell instance $1619 m0 *1 45.6,91
X$1619 2401 1289 1813 23 38 2400 MUX2_X1
* cell instance $1620 m0 *1 46.93,91
X$1620 23 38 FILLCELL_X2
* cell instance $1621 r0 *1 44.84,91
X$1621 23 38 FILLCELL_X4
* cell instance $1622 r0 *1 45.6,91
X$1622 23 3067 2401 2400 2333 38 DFF_X1
* cell instance $1623 m0 *1 47.5,91
X$1623 2334 627 2401 23 38 2427 MUX2_X1
* cell instance $1624 m0 *1 47.31,91
X$1624 23 38 FILLCELL_X1
* cell instance $1625 m0 *1 48.83,91
X$1625 23 38 FILLCELL_X1
* cell instance $1626 m0 *1 49.02,91
X$1626 2362 1369 1813 23 38 2393 MUX2_X1
* cell instance $1627 m0 *1 50.35,91
X$1627 23 2588 2362 2393 2316 38 DFF_X1
* cell instance $1628 m0 *1 53.58,91
X$1628 2397 724 2362 23 38 2431 MUX2_X1
* cell instance $1629 m0 *1 54.91,91
X$1629 2431 1650 23 38 2430 NOR2_X1
* cell instance $1630 m0 *1 55.48,91
X$1630 2316 23 38 CLKBUF_X1
* cell instance $1631 m0 *1 56.05,91
X$1631 23 38 FILLCELL_X1
* cell instance $1632 m0 *1 56.24,91
X$1632 2363 1373 2402 23 38 2398 MUX2_X1
* cell instance $1633 m0 *1 57.57,91
X$1633 23 38 FILLCELL_X2
* cell instance $1634 r0 *1 48.83,91
X$1634 23 38 FILLCELL_X4
* cell instance $1635 r0 *1 49.59,91
X$1635 23 38 FILLCELL_X1
* cell instance $1636 r0 *1 49.78,91
X$1636 2427 1579 23 38 2444 NOR2_X1
* cell instance $1637 r0 *1 50.35,91
X$1637 1425 2444 2430 548 2470 2471 23 38 2016 OAI33_X1
* cell instance $1638 r0 *1 51.68,91
X$1638 2445 1535 23 38 2470 NOR2_X1
* cell instance $1639 r0 *1 52.25,91
X$1639 23 38 FILLCELL_X4
* cell instance $1640 r0 *1 53.01,91
X$1640 2446 1483 23 38 2471 NOR2_X1
* cell instance $1641 r0 *1 53.58,91
X$1641 23 38 FILLCELL_X2
* cell instance $1642 r0 *1 53.96,91
X$1642 2058 23 38 2316 CLKBUF_X3
* cell instance $1643 r0 *1 54.91,91
X$1643 23 3127 2363 2447 2316 38 DFF_X1
* cell instance $1644 m0 *1 59.28,91
X$1644 23 38 FILLCELL_X8
* cell instance $1645 m0 *1 57.95,91
X$1645 2151 1480 2402 23 38 2403 MUX2_X1
* cell instance $1646 m0 *1 60.8,91
X$1646 23 38 FILLCELL_X2
* cell instance $1647 r0 *1 58.14,91
X$1647 23 3089 2402 2403 2316 38 DFF_X1
* cell instance $1648 r0 *1 59.14,91
X$1648 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $1649 r0 *1 59.14,91
X$1649 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $1650 r0 *1 59.14,91
X$1650 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $1651 m0 *1 64.41,91
X$1651 23 2579 2364 2396 2246 38 DFF_X1
* cell instance $1652 m0 *1 61.18,91
X$1652 23 2657 1370 2404 2246 38 DFF_X1
* cell instance $1653 m0 *1 67.64,91
X$1653 23 38 FILLCELL_X2
* cell instance $1654 r0 *1 61.37,91
X$1654 23 38 FILLCELL_X8
* cell instance $1655 r0 *1 62.89,91
X$1655 23 38 FILLCELL_X2
* cell instance $1656 r0 *1 63.27,91
X$1656 23 38 FILLCELL_X1
* cell instance $1657 r0 *1 63.46,91
X$1657 2236 23 38 2155 INV_X2
* cell instance $1658 r0 *1 64.03,91
X$1658 2246 23 38 CLKBUF_X1
* cell instance $1659 r0 *1 64.6,91
X$1659 23 2473 2284 2404 2246 38 DFF_X1
* cell instance $1660 r0 *1 67.83,91
X$1660 23 38 FILLCELL_X1
* cell instance $1661 m0 *1 68.78,91
X$1661 2405 2391 2365 23 38 2404 MUX2_X1
* cell instance $1662 m0 *1 68.02,91
X$1662 2284 2057 38 23 2405 AND2_X1
* cell instance $1663 m0 *1 70.11,91
X$1663 1319 2284 23 38 2365 NOR2_X1
* cell instance $1664 m0 *1 70.68,91
X$1664 23 38 FILLCELL_X4
* cell instance $1665 m0 *1 71.44,91
X$1665 23 38 FILLCELL_X1
* cell instance $1666 m0 *1 71.63,91
X$1666 2187 2186 2450 38 23 2406 HA_X1
* cell instance $1667 m0 *1 73.53,91
X$1667 2366 2190 2232 23 2391 38 AOI21_X1
* cell instance $1668 m0 *1 74.29,91
X$1668 23 38 FILLCELL_X4
* cell instance $1669 m0 *1 75.05,91
X$1669 23 38 FILLCELL_X1
* cell instance $1670 m0 *1 75.24,91
X$1670 2367 23 38 2407 INV_X1
* cell instance $1671 m0 *1 75.62,91
X$1671 2189 2428 38 2190 23 XOR2_X2
* cell instance $1672 m0 *1 77.33,91
X$1672 23 38 FILLCELL_X4
* cell instance $1673 m0 *1 78.09,91
X$1673 23 38 FILLCELL_X1
* cell instance $1674 m0 *1 78.28,91
X$1674 2454 23 38 2160 CLKBUF_X3
* cell instance $1675 m0 *1 79.23,91
X$1675 23 38 FILLCELL_X4
* cell instance $1676 m0 *1 79.99,91
X$1676 2387 1686 2065 23 38 2410 NOR3_X1
* cell instance $1677 m0 *1 80.75,91
X$1677 23 2677 2369 2389 2373 38 DFF_X1
* cell instance $1678 m0 *1 83.98,91
X$1678 2423 1300 2065 23 38 2483 NOR3_X1
* cell instance $1679 m0 *1 84.74,91
X$1679 2422 2370 2369 23 38 2387 NAND3_X1
* cell instance $1680 m0 *1 85.5,91
X$1680 2193 2337 2412 2338 23 38 2423 NAND4_X1
* cell instance $1681 m0 *1 86.45,91
X$1681 2193 2337 2232 2190 23 38 2376 NAND4_X1
* cell instance $1682 m0 *1 87.4,91
X$1682 23 38 FILLCELL_X1
* cell instance $1683 m0 *1 87.59,91
X$1683 2414 2063 2161 38 23 2422 AND3_X1
* cell instance $1684 m0 *1 88.54,91
X$1684 2378 1686 2065 23 38 2458 NOR3_X1
* cell instance $1685 m0 *1 89.3,91
X$1685 2377 2376 2371 23 38 2372 MUX2_X1
* cell instance $1686 m0 *1 90.63,91
X$1686 23 2826 2416 2372 2373 38 DFF_X1
* cell instance $1687 m0 *1 93.86,91
X$1687 23 38 FILLCELL_X2
* cell instance $1688 r0 *1 68.02,91
X$1688 2473 2364 2504 38 23 2449 HA_X1
* cell instance $1689 r0 *1 69.92,91
X$1689 2472 2154 2503 38 23 2501 HA_X1
* cell instance $1690 r0 *1 71.82,91
X$1690 2449 2478 2480 23 2429 38 AOI21_X1
* cell instance $1691 r0 *1 72.58,91
X$1691 23 38 FILLCELL_X1
* cell instance $1692 r0 *1 72.77,91
X$1692 2406 23 38 2562 BUF_X1
* cell instance $1693 r0 *1 73.34,91
X$1693 2406 23 38 2500 INV_X1
* cell instance $1694 r0 *1 73.72,91
X$1694 2450 23 38 2451 INV_X1
* cell instance $1695 r0 *1 74.1,91
X$1695 2408 2429 2407 38 2428 23 OAI21_X1
* cell instance $1696 r0 *1 74.86,91
X$1696 2452 2409 2451 2408 23 38 2498 NOR4_X1
* cell instance $1697 r0 *1 75.81,91
X$1697 2336 23 38 2408 INV_X1
* cell instance $1698 r0 *1 76.19,91
X$1698 23 38 FILLCELL_X1
* cell instance $1699 r0 *1 76.38,91
X$1699 2452 2451 2409 2408 38 2453 23 OR4_X2
* cell instance $1700 r0 *1 77.71,91
X$1700 2450 2409 23 38 2455 XOR2_X1
* cell instance $1701 r0 *1 78.85,91
X$1701 23 38 FILLCELL_X4
* cell instance $1702 r0 *1 79.61,91
X$1702 23 38 FILLCELL_X2
* cell instance $1703 r0 *1 79.99,91
X$1703 2156 23 38 2232 CLKBUF_X3
* cell instance $1704 r0 *1 80.94,91
X$1704 23 38 FILLCELL_X8
* cell instance $1705 r0 *1 82.46,91
X$1705 23 38 FILLCELL_X4
* cell instance $1706 r0 *1 83.22,91
X$1706 23 38 FILLCELL_X1
* cell instance $1707 r0 *1 83.41,91
X$1707 2411 2057 38 23 2456 AND2_X1
* cell instance $1708 r0 *1 84.17,91
X$1708 23 38 FILLCELL_X2
* cell instance $1709 r0 *1 84.55,91
X$1709 23 38 FILLCELL_X1
* cell instance $1710 r0 *1 84.74,91
X$1710 1319 2411 23 38 2457 NOR2_X1
* cell instance $1711 r0 *1 85.31,91
X$1711 23 38 FILLCELL_X1
* cell instance $1712 r0 *1 85.5,91
X$1712 2411 2412 2338 2192 23 38 2413 NAND4_X1
* cell instance $1713 r0 *1 86.45,91
X$1713 2413 2289 23 38 2370 NOR2_X1
* cell instance $1714 r0 *1 87.02,91
X$1714 23 38 FILLCELL_X2
* cell instance $1715 r0 *1 87.4,91
X$1715 1319 2414 23 38 2462 NOR2_X1
* cell instance $1716 r0 *1 87.97,91
X$1716 2414 2057 38 23 2415 AND2_X1
* cell instance $1717 r0 *1 88.73,91
X$1717 2415 2458 2462 23 38 2459 MUX2_X1
* cell instance $1718 r0 *1 90.06,91
X$1718 23 38 FILLCELL_X32
* cell instance $1719 m0 *1 94.81,91
X$1719 2416 23 38 2374 BUF_X1
* cell instance $1720 m0 *1 94.24,91
X$1720 2416 23 38 2338 BUF_X1
* cell instance $1721 m0 *1 95.38,91
X$1721 2293 23 38 2417 BUF_X1
* cell instance $1722 m0 *1 95.95,91
X$1722 23 38 FILLCELL_X4
* cell instance $1723 m0 *1 96.71,91
X$1723 23 38 FILLCELL_X2
* cell instance $1724 r0 *1 96.14,91
X$1724 23 38 FILLCELL_X4
* cell instance $1725 r0 *1 96.9,91
X$1725 23 38 FILLCELL_X1
* cell instance $1726 m90 *1 97.28,91
X$1726 23 38 23 38 TAPCELL_X1
* cell instance $1727 r180 *1 97.28,91
X$1727 23 38 23 38 TAPCELL_X1
* cell instance $1728 m0 *1 59.85,96.6
X$1728 23 2653 2507 2531 2246 38 DFF_X1
* cell instance $1729 m0 *1 59.66,96.6
X$1729 23 38 FILLCELL_X1
* cell instance $1730 m0 *1 63.08,96.6
X$1730 23 38 FILLCELL_X4
* cell instance $1731 m0 *1 63.84,96.6
X$1731 2533 23 38 2236 BUF_X1
* cell instance $1732 m0 *1 64.41,96.6
X$1732 23 38 FILLCELL_X2
* cell instance $1733 m0 *1 4.18,43.4
X$1733 23 2705 1028 1043 1094 38 DFF_X1
* cell instance $1734 m0 *1 3.99,43.4
X$1734 23 38 FILLCELL_X1
* cell instance $1735 m0 *1 7.41,43.4
X$1735 1028 941 502 23 38 1043 MUX2_X1
* cell instance $1736 m0 *1 8.74,43.4
X$1736 23 38 FILLCELL_X32
* cell instance $1737 m0 *1 14.82,43.4
X$1737 23 38 FILLCELL_X8
* cell instance $1738 m0 *1 16.34,43.4
X$1738 23 38 FILLCELL_X4
* cell instance $1739 m0 *1 17.1,43.4
X$1739 23 38 FILLCELL_X1
* cell instance $1740 m0 *1 17.29,43.4
X$1740 23 2699 1016 990 991 38 DFF_X1
* cell instance $1741 m0 *1 20.52,43.4
X$1741 23 38 FILLCELL_X2
* cell instance $1742 m0 *1 1.33,43.4
X$1742 23 38 FILLCELL_X8
* cell instance $1743 m0 *1 1.14,43.4
X$1743 23 38 23 38 TAPCELL_X1
* cell instance $1744 m0 *1 2.85,43.4
X$1744 23 38 FILLCELL_X4
* cell instance $1745 m0 *1 3.61,43.4
X$1745 23 38 FILLCELL_X2
* cell instance $1746 r0 *1 1.14,43.4
X$1746 23 38 23 38 TAPCELL_X1
* cell instance $1747 r0 *1 1.33,43.4
X$1747 23 38 FILLCELL_X16
* cell instance $1748 r0 *1 3.14,43.4
X$1748 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $1749 r0 *1 3.14,43.4
X$1749 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $1750 r0 *1 3.14,43.4
X$1750 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $1751 r0 *1 4.37,43.4
X$1751 23 38 FILLCELL_X8
* cell instance $1752 r0 *1 5.89,43.4
X$1752 23 38 FILLCELL_X2
* cell instance $1753 r0 *1 6.27,43.4
X$1753 23 38 FILLCELL_X1
* cell instance $1754 r0 *1 6.46,43.4
X$1754 1056 992 502 23 38 1075 MUX2_X1
* cell instance $1755 r0 *1 7.79,43.4
X$1755 1028 994 1056 23 38 1078 MUX2_X1
* cell instance $1756 r0 *1 9.12,43.4
X$1756 23 38 FILLCELL_X8
* cell instance $1757 r0 *1 10.64,43.4
X$1757 23 38 FILLCELL_X4
* cell instance $1758 r0 *1 11.4,43.4
X$1758 23 38 FILLCELL_X1
* cell instance $1759 r0 *1 11.59,43.4
X$1759 23 3078 1057 1077 1094 38 DFF_X1
* cell instance $1760 r0 *1 14.82,43.4
X$1760 1057 929 502 23 38 1077 MUX2_X1
* cell instance $1761 r0 *1 16.15,43.4
X$1761 1078 937 23 38 1079 NOR2_X1
* cell instance $1762 r0 *1 16.72,43.4
X$1762 23 38 FILLCELL_X1
* cell instance $1763 r0 *1 16.91,43.4
X$1763 932 1079 1096 891 918 922 23 38 1058 OAI33_X1
* cell instance $1764 r0 *1 18.24,43.4
X$1764 23 38 FILLCELL_X8
* cell instance $1765 r0 *1 19.76,43.4
X$1765 23 38 FILLCELL_X4
* cell instance $1766 r0 *1 20.52,43.4
X$1766 23 38 FILLCELL_X2
* cell instance $1767 m0 *1 1.9,21
X$1767 23 2747 465 526 447 38 DFF_X1
* cell instance $1768 m0 *1 1.71,21
X$1768 23 38 FILLCELL_X1
* cell instance $1769 m0 *1 5.13,21
X$1769 465 412 448 23 38 485 MUX2_X1
* cell instance $1770 m0 *1 6.46,21
X$1770 149 23 38 447 CLKBUF_X3
* cell instance $1771 m0 *1 7.41,21
X$1771 447 23 38 CLKBUF_X1
* cell instance $1772 m0 *1 7.98,21
X$1772 23 38 FILLCELL_X2
* cell instance $1773 m0 *1 1.33,21
X$1773 23 38 FILLCELL_X2
* cell instance $1774 m0 *1 1.14,21
X$1774 23 38 23 38 TAPCELL_X1
* cell instance $1775 r0 *1 1.14,21
X$1775 23 38 23 38 TAPCELL_X1
* cell instance $1776 r0 *1 1.33,21
X$1776 23 38 FILLCELL_X8
* cell instance $1777 r0 *1 2.85,21
X$1777 23 38 FILLCELL_X4
* cell instance $1778 r0 *1 3.14,21
X$1778 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $1779 r0 *1 3.14,21
X$1779 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $1780 r0 *1 3.14,21
X$1780 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $1781 r0 *1 3.61,21
X$1781 465 318 502 23 38 526 MUX2_X1
* cell instance $1782 r0 *1 4.94,21
X$1782 448 257 502 23 38 446 MUX2_X1
* cell instance $1783 r0 *1 6.27,21
X$1783 23 38 FILLCELL_X16
* cell instance $1784 m0 *1 8.55,21
X$1784 411 318 453 23 38 450 MUX2_X1
* cell instance $1785 m0 *1 8.36,21
X$1785 23 38 FILLCELL_X1
* cell instance $1786 m0 *1 9.88,21
X$1786 485 354 23 38 490 NOR2_X1
* cell instance $1787 m0 *1 10.45,21
X$1787 23 38 FILLCELL_X8
* cell instance $1788 m0 *1 11.97,21
X$1788 23 38 FILLCELL_X2
* cell instance $1789 r0 *1 9.31,21
X$1789 23 38 FILLCELL_X8
* cell instance $1790 r0 *1 10.83,21
X$1790 528 354 23 38 547 NOR2_X1
* cell instance $1791 r0 *1 11.4,21
X$1791 23 38 FILLCELL_X16
* cell instance $1792 m0 *1 12.54,21
X$1792 23 2737 451 488 503 38 DFF_X1
* cell instance $1793 m0 *1 12.35,21
X$1793 23 38 FILLCELL_X1
* cell instance $1794 m0 *1 15.77,21
X$1794 356 492 490 360 322 338 23 38 531 OAI33_X1
* cell instance $1795 m0 *1 17.1,21
X$1795 530 381 23 38 492 NOR2_X1
* cell instance $1796 m0 *1 17.67,21
X$1796 23 38 FILLCELL_X4
* cell instance $1797 m0 *1 18.43,21
X$1797 23 38 FILLCELL_X2
* cell instance $1798 r0 *1 14.44,21
X$1798 23 38 FILLCELL_X1
* cell instance $1799 r0 *1 14.63,21
X$1799 503 23 38 3148 INV_X1
* cell instance $1800 r0 *1 15.01,21
X$1800 149 23 38 503 CLKBUF_X3
* cell instance $1801 r0 *1 15.96,21
X$1801 549 472 504 23 38 530 MUX2_X1
* cell instance $1802 r0 *1 17.29,21
X$1802 504 437 502 23 38 550 MUX2_X1
* cell instance $1803 r0 *1 18.62,21
X$1803 23 38 FILLCELL_X4
* cell instance $1804 m0 *1 19,21
X$1804 466 437 453 23 38 493 MUX2_X1
* cell instance $1805 m0 *1 18.81,21
X$1805 23 38 FILLCELL_X1
* cell instance $1806 m0 *1 20.33,21
X$1806 23 2742 466 493 324 38 DFF_X1
* cell instance $1807 m0 *1 23.56,21
X$1807 23 38 FILLCELL_X4
* cell instance $1808 m0 *1 24.32,21
X$1808 149 23 38 324 CLKBUF_X3
* cell instance $1809 m0 *1 25.27,21
X$1809 324 23 38 3144 INV_X1
* cell instance $1810 m0 *1 25.65,21
X$1810 23 38 FILLCELL_X2
* cell instance $1811 r0 *1 19.38,21
X$1811 23 38 FILLCELL_X1
* cell instance $1812 r0 *1 19.57,21
X$1812 505 393 358 23 38 533 MUX2_X1
* cell instance $1813 r0 *1 20.9,21
X$1813 23 3042 505 533 324 38 DFF_X1
* cell instance $1814 r0 *1 24.13,21
X$1814 505 472 576 23 38 467 MUX2_X1
* cell instance $1815 r0 *1 25.46,21
X$1815 23 38 FILLCELL_X1
* cell instance $1816 r0 *1 25.65,21
X$1816 23 2923 507 506 324 38 DFF_X1
* cell instance $1817 m0 *1 29.26,21
X$1817 507 472 468 23 38 497 MUX2_X1
* cell instance $1818 m0 *1 26.03,21
X$1818 23 2773 468 495 324 38 DFF_X1
* cell instance $1819 m0 *1 30.59,21
X$1819 23 38 FILLCELL_X1
* cell instance $1820 m0 *1 30.78,21
X$1820 497 381 23 38 469 NOR2_X1
* cell instance $1821 m0 *1 31.35,21
X$1821 23 38 FILLCELL_X4
* cell instance $1822 m0 *1 32.11,21
X$1822 536 354 23 38 458 NOR2_X1
* cell instance $1823 m0 *1 32.68,21
X$1823 23 2776 470 511 329 38 DFF_X1
* cell instance $1824 m0 *1 35.91,21
X$1824 470 472 540 23 38 435 MUX2_X1
* cell instance $1825 m0 *1 37.24,21
X$1825 23 38 FILLCELL_X1
* cell instance $1826 m0 *1 37.43,21
X$1826 23 2786 554 553 329 38 DFF_X1
* cell instance $1827 m0 *1 40.66,21
X$1827 23 38 FILLCELL_X2
* cell instance $1828 r0 *1 28.88,21
X$1828 23 38 FILLCELL_X4
* cell instance $1829 r0 *1 29.64,21
X$1829 551 318 510 23 38 508 MUX2_X1
* cell instance $1830 r0 *1 30.97,21
X$1830 551 305 509 23 38 536 MUX2_X1
* cell instance $1831 r0 *1 32.3,21
X$1831 23 38 FILLCELL_X2
* cell instance $1832 r0 *1 32.68,21
X$1832 470 393 510 23 38 511 MUX2_X1
* cell instance $1833 r0 *1 34.01,21
X$1833 23 38 FILLCELL_X1
* cell instance $1834 r0 *1 34.2,21
X$1834 540 437 510 23 38 552 MUX2_X1
* cell instance $1835 r0 *1 35.53,21
X$1835 23 38 FILLCELL_X8
* cell instance $1836 r0 *1 37.05,21
X$1836 23 38 FILLCELL_X4
* cell instance $1837 r0 *1 37.81,21
X$1837 23 2860 578 542 329 38 DFF_X1
* cell instance $1838 r0 *1 41.04,21
X$1838 23 38 FILLCELL_X1
* cell instance $1839 m0 *1 41.23,21
X$1839 579 370 23 38 436 NOR2_X1
* cell instance $1840 m0 *1 41.04,21
X$1840 23 38 FILLCELL_X1
* cell instance $1841 m0 *1 41.8,21
X$1841 23 38 FILLCELL_X4
* cell instance $1842 m0 *1 42.56,21
X$1842 501 393 398 23 38 544 MUX2_X1
* cell instance $1843 m0 *1 43.89,21
X$1843 501 472 512 23 38 500 MUX2_X1
* cell instance $1844 m0 *1 45.22,21
X$1844 500 370 23 38 471 NOR2_X1
* cell instance $1845 m0 *1 45.79,21
X$1845 299 23 38 CLKBUF_X1
* cell instance $1846 m0 *1 46.36,21
X$1846 23 38 FILLCELL_X32
* cell instance $1847 m0 *1 52.44,21
X$1847 403 38 261 23 BUF_X4
* cell instance $1848 m0 *1 53.77,21
X$1848 23 2610 514 499 158 38 DFF_X1
* cell instance $1849 m0 *1 57,21
X$1849 23 38 FILLCELL_X4
* cell instance $1850 m0 *1 57.76,21
X$1850 588 367 23 38 516 NOR2_X1
* cell instance $1851 m0 *1 58.33,21
X$1851 23 38 FILLCELL_X2
* cell instance $1852 r0 *1 41.23,21
X$1852 23 2890 501 544 299 38 DFF_X1
* cell instance $1853 r0 *1 44.46,21
X$1853 23 38 FILLCELL_X2
* cell instance $1854 r0 *1 44.84,21
X$1854 23 38 FILLCELL_X1
* cell instance $1855 r0 *1 45.03,21
X$1855 512 437 398 23 38 581 MUX2_X1
* cell instance $1856 r0 *1 46.36,21
X$1856 23 38 FILLCELL_X4
* cell instance $1857 r0 *1 47.12,21
X$1857 23 38 FILLCELL_X2
* cell instance $1858 r0 *1 47.5,21
X$1858 23 38 FILLCELL_X1
* cell instance $1859 r0 *1 47.69,21
X$1859 23 3118 513 545 299 38 DFF_X1
* cell instance $1860 r0 *1 50.92,21
X$1860 513 472 555 23 38 546 MUX2_X1
* cell instance $1861 r0 *1 52.25,21
X$1861 23 38 FILLCELL_X1
* cell instance $1862 r0 *1 52.44,21
X$1862 515 23 38 356 CLKBUF_X3
* cell instance $1863 r0 *1 53.39,21
X$1863 23 3005 558 586 158 38 DFF_X1
* cell instance $1864 r0 *1 56.62,21
X$1864 546 370 23 38 587 NOR2_X1
* cell instance $1865 r0 *1 57.19,21
X$1865 23 38 FILLCELL_X4
* cell instance $1866 r0 *1 57.95,21
X$1866 515 587 516 360 517 518 23 38 522 OAI33_X1
* cell instance $1867 m0 *1 59.28,21
X$1867 23 38 FILLCELL_X2
* cell instance $1868 m0 *1 58.71,21
X$1868 134 374 23 38 518 NOR2_X1
* cell instance $1869 r0 *1 59.14,21
X$1869 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $1870 r0 *1 59.14,21
X$1870 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $1871 r0 *1 59.14,21
X$1871 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $1872 r0 *1 59.28,21
X$1872 23 38 FILLCELL_X1
* cell instance $1873 r0 *1 59.47,21
X$1873 23 2963 585 584 543 38 DFF_X1
* cell instance $1874 m0 *1 59.85,21
X$1874 23 2840 519 498 543 38 DFF_X1
* cell instance $1875 m0 *1 59.66,21
X$1875 23 38 FILLCELL_X1
* cell instance $1876 m0 *1 63.08,21
X$1876 123 374 23 38 603 NOR2_X1
* cell instance $1877 m0 *1 63.65,21
X$1877 23 38 FILLCELL_X4
* cell instance $1878 m0 *1 64.41,21
X$1878 23 38 FILLCELL_X2
* cell instance $1879 r0 *1 62.7,21
X$1879 519 520 48 23 38 498 MUX2_X1
* cell instance $1880 r0 *1 64.03,21
X$1880 23 38 FILLCELL_X8
* cell instance $1881 m0 *1 66.12,21
X$1881 23 2854 457 494 334 38 DFF_X1
* cell instance $1882 m0 *1 64.79,21
X$1882 475 440 560 476 496 406 23 38 474 OAI33_X1
* cell instance $1883 m0 *1 69.35,21
X$1883 23 38 FILLCELL_X2
* cell instance $1884 r0 *1 65.55,21
X$1884 23 38 FILLCELL_X4
* cell instance $1885 r0 *1 66.31,21
X$1885 23 38 FILLCELL_X1
* cell instance $1886 r0 *1 66.5,21
X$1886 538 520 78 23 38 582 MUX2_X1
* cell instance $1887 r0 *1 67.83,21
X$1887 23 38 FILLCELL_X2
* cell instance $1888 r0 *1 68.21,21
X$1888 23 38 FILLCELL_X1
* cell instance $1889 r0 *1 68.4,21
X$1889 561 541 538 23 38 539 MUX2_X1
* cell instance $1890 m0 *1 71.06,21
X$1890 23 38 FILLCELL_X1
* cell instance $1891 m0 *1 69.73,21
X$1891 475 442 521 476 407 419 23 38 483 OAI33_X1
* cell instance $1892 m0 *1 71.25,21
X$1892 23 2686 477 535 334 38 DFF_X1
* cell instance $1893 m0 *1 74.48,21
X$1893 139 23 38 334 CLKBUF_X3
* cell instance $1894 m0 *1 75.43,21
X$1894 478 367 23 38 489 NOR2_X1
* cell instance $1895 m0 *1 76,21
X$1895 23 38 FILLCELL_X2
* cell instance $1896 r0 *1 69.73,21
X$1896 539 367 23 38 521 NOR2_X1
* cell instance $1897 r0 *1 70.3,21
X$1897 23 38 FILLCELL_X2
* cell instance $1898 r0 *1 70.68,21
X$1898 23 2920 580 537 334 38 DFF_X1
* cell instance $1899 r0 *1 73.91,21
X$1899 23 38 FILLCELL_X2
* cell instance $1900 r0 *1 74.29,21
X$1900 477 520 52 23 38 535 MUX2_X1
* cell instance $1901 r0 *1 75.62,21
X$1901 23 38 FILLCELL_X4
* cell instance $1902 m0 *1 76.57,21
X$1902 475 491 489 476 443 486 23 38 534 OAI33_X1
* cell instance $1903 m0 *1 76.38,21
X$1903 23 38 FILLCELL_X1
* cell instance $1904 m0 *1 77.9,21
X$1904 524 51 444 23 38 487 MUX2_X1
* cell instance $1905 m0 *1 79.23,21
X$1905 23 38 FILLCELL_X2
* cell instance $1906 r0 *1 76.38,21
X$1906 23 2931 562 523 445 38 DFF_X1
* cell instance $1907 r0 *1 79.61,21
X$1907 532 372 23 38 563 NOR2_X1
* cell instance $1908 m0 *1 80.94,21
X$1908 23 38 FILLCELL_X4
* cell instance $1909 m0 *1 79.61,21
X$1909 444 80 378 23 38 532 MUX2_X1
* cell instance $1910 m0 *1 81.7,21
X$1910 23 38 FILLCELL_X2
* cell instance $1911 r0 *1 80.18,21
X$1911 23 38 FILLCELL_X8
* cell instance $1912 r0 *1 81.7,21
X$1912 23 38 FILLCELL_X1
* cell instance $1913 r0 *1 81.89,21
X$1913 525 414 479 23 38 565 MUX2_X1
* cell instance $1914 m0 *1 83.41,21
X$1914 23 2666 479 484 445 38 DFF_X1
* cell instance $1915 m0 *1 82.08,21
X$1915 377 240 479 23 38 484 MUX2_X1
* cell instance $1916 m0 *1 86.64,21
X$1916 23 38 FILLCELL_X8
* cell instance $1917 m0 *1 88.16,21
X$1917 23 2565 529 482 310 38 DFF_X1
* cell instance $1918 m0 *1 91.39,21
X$1918 23 38 FILLCELL_X8
* cell instance $1919 m0 *1 92.91,21
X$1919 23 38 FILLCELL_X2
* cell instance $1920 r0 *1 83.22,21
X$1920 23 38 FILLCELL_X8
* cell instance $1921 r0 *1 84.74,21
X$1921 23 38 FILLCELL_X1
* cell instance $1922 r0 *1 84.93,21
X$1922 377 23 38 524 BUF_X2
* cell instance $1923 r0 *1 85.69,21
X$1923 23 2930 573 566 445 38 DFF_X1
* cell instance $1924 r0 *1 88.92,21
X$1924 529 174 524 23 38 482 MUX2_X1
* cell instance $1925 r0 *1 90.25,21
X$1925 23 38 FILLCELL_X8
* cell instance $1926 r0 *1 91.77,21
X$1926 23 38 FILLCELL_X2
* cell instance $1927 r0 *1 92.15,21
X$1927 410 274 23 38 567 NOR2_X1
* cell instance $1928 r0 *1 92.72,21
X$1928 23 38 FILLCELL_X2
* cell instance $1929 r0 *1 93.1,21
X$1929 23 2926 568 527 310 38 DFF_X1
* cell instance $1930 m0 *1 96.52,21
X$1930 23 38 FILLCELL_X2
* cell instance $1931 m0 *1 93.29,21
X$1931 23 2571 480 481 310 38 DFF_X1
* cell instance $1932 r0 *1 96.33,21
X$1932 23 38 FILLCELL_X4
* cell instance $1933 r180 *1 97.28,21
X$1933 23 38 23 38 TAPCELL_X1
* cell instance $1934 m0 *1 96.9,21
X$1934 23 38 FILLCELL_X1
* cell instance $1935 m90 *1 97.28,21
X$1935 23 38 23 38 TAPCELL_X1
* cell instance $1936 r0 *1 67.45,1.4
X$1936 23 38 FILLCELL_X1
* cell instance $1937 r0 *1 70.87,1.4
X$1937 23 38 FILLCELL_X4
* cell instance $1938 r0 *1 72.2,1.4
X$1938 23 38 FILLCELL_X16
* cell instance $1939 r0 *1 75.24,1.4
X$1939 23 38 FILLCELL_X4
* cell instance $1940 r0 *1 79.23,1.4
X$1940 23 38 FILLCELL_X2
* cell instance $1941 m0 *1 68.78,96.6
X$1941 23 38 FILLCELL_X16
* cell instance $1942 m0 *1 67.83,96.6
X$1942 2539 23 38 1478 CLKBUF_X3
* cell instance $1943 m0 *1 71.82,96.6
X$1943 23 38 FILLCELL_X8
* cell instance $1944 m0 *1 73.34,96.6
X$1944 23 38 FILLCELL_X4
* cell instance $1945 m0 *1 74.1,96.6
X$1945 23 38 FILLCELL_X2
* cell instance $1946 m0 *1 1.33,68.6
X$1946 23 38 FILLCELL_X16
* cell instance $1947 m0 *1 1.14,68.6
X$1947 23 38 23 38 TAPCELL_X1
* cell instance $1948 m0 *1 4.37,68.6
X$1948 23 38 FILLCELL_X8
* cell instance $1949 m0 *1 5.89,68.6
X$1949 23 38 FILLCELL_X4
* cell instance $1950 m0 *1 6.65,68.6
X$1950 23 38 FILLCELL_X2
* cell instance $1951 r0 *1 1.14,68.6
X$1951 23 38 23 38 TAPCELL_X1
* cell instance $1952 r0 *1 1.33,68.6
X$1952 23 38 FILLCELL_X2
* cell instance $1953 r0 *1 1.71,68.6
X$1953 23 38 FILLCELL_X1
* cell instance $1954 r0 *1 1.9,68.6
X$1954 23 3002 1789 1834 1556 38 DFF_X1
* cell instance $1955 r0 *1 3.14,68.6
X$1955 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $1956 r0 *1 3.14,68.6
X$1956 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $1957 r0 *1 3.14,68.6
X$1957 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $1958 r0 *1 5.13,68.6
X$1958 1789 1383 1791 23 38 1834 MUX2_X1
* cell instance $1959 r0 *1 6.46,68.6
X$1959 23 38 FILLCELL_X4
* cell instance $1960 m0 *1 7.22,68.6
X$1960 23 2605 1790 1838 1556 38 DFF_X1
* cell instance $1961 m0 *1 7.03,68.6
X$1961 23 38 FILLCELL_X1
* cell instance $1962 m0 *1 10.45,68.6
X$1962 23 38 FILLCELL_X1
* cell instance $1963 m0 *1 10.64,68.6
X$1963 1717 1369 1532 23 38 1747 MUX2_X1
* cell instance $1964 m0 *1 11.97,68.6
X$1964 23 38 FILLCELL_X2
* cell instance $1965 r0 *1 7.22,68.6
X$1965 23 38 FILLCELL_X2
* cell instance $1966 r0 *1 7.6,68.6
X$1966 1790 1383 1532 23 38 1838 MUX2_X1
* cell instance $1967 r0 *1 8.93,68.6
X$1967 1790 412 1717 23 38 1836 MUX2_X1
* cell instance $1968 r0 *1 10.26,68.6
X$1968 23 38 FILLCELL_X2
* cell instance $1969 r0 *1 10.64,68.6
X$1969 1836 354 23 38 1778 NOR2_X1
* cell instance $1970 r0 *1 11.21,68.6
X$1970 23 38 FILLCELL_X8
* cell instance $1971 m0 *1 12.54,68.6
X$1971 1762 1403 1532 23 38 1779 MUX2_X1
* cell instance $1972 m0 *1 12.35,68.6
X$1972 23 38 FILLCELL_X1
* cell instance $1973 m0 *1 13.87,68.6
X$1973 23 38 FILLCELL_X16
* cell instance $1974 m0 *1 16.91,68.6
X$1974 23 38 FILLCELL_X8
* cell instance $1975 m0 *1 18.43,68.6
X$1975 23 38 FILLCELL_X4
* cell instance $1976 m0 *1 19.19,68.6
X$1976 23 38 FILLCELL_X2
* cell instance $1977 r0 *1 12.73,68.6
X$1977 23 38 FILLCELL_X4
* cell instance $1978 r0 *1 13.49,68.6
X$1978 23 38 FILLCELL_X2
* cell instance $1979 r0 *1 13.87,68.6
X$1979 23 38 FILLCELL_X1
* cell instance $1980 r0 *1 14.06,68.6
X$1980 1486 23 38 1635 CLKBUF_X3
* cell instance $1981 r0 *1 15.01,68.6
X$1981 1635 23 38 CLKBUF_X1
* cell instance $1982 r0 *1 15.58,68.6
X$1982 23 38 FILLCELL_X2
* cell instance $1983 r0 *1 15.96,68.6
X$1983 1842 1434 1791 23 38 1841 MUX2_X1
* cell instance $1984 r0 *1 17.29,68.6
X$1984 23 38 FILLCELL_X4
* cell instance $1985 r0 *1 18.05,68.6
X$1985 23 2948 1843 1792 1635 38 DFF_X1
* cell instance $1986 m0 *1 19.76,68.6
X$1986 1723 1487 1791 23 38 1781 MUX2_X1
* cell instance $1987 m0 *1 19.57,68.6
X$1987 23 38 FILLCELL_X1
* cell instance $1988 m0 *1 21.09,68.6
X$1988 1780 937 23 38 1793 NOR2_X1
* cell instance $1989 m0 *1 21.66,68.6
X$1989 23 38 FILLCELL_X4
* cell instance $1990 m0 *1 22.42,68.6
X$1990 23 38 FILLCELL_X2
* cell instance $1991 r0 *1 21.28,68.6
X$1991 23 38 FILLCELL_X16
* cell instance $1992 m0 *1 22.99,68.6
X$1992 434 23 38 1486 CLKBUF_X3
* cell instance $1993 m0 *1 22.8,68.6
X$1993 23 38 FILLCELL_X1
* cell instance $1994 m0 *1 23.94,68.6
X$1994 1486 23 38 3153 CLKBUF_X3
* cell instance $1995 m0 *1 24.89,68.6
X$1995 1693 23 38 CLKBUF_X1
* cell instance $1996 m0 *1 25.46,68.6
X$1996 23 38 FILLCELL_X2
* cell instance $1997 r0 *1 24.32,68.6
X$1997 23 38 FILLCELL_X4
* cell instance $1998 r0 *1 25.08,68.6
X$1998 23 38 FILLCELL_X2
* cell instance $1999 r0 *1 25.46,68.6
X$1999 23 38 FILLCELL_X1
* cell instance $2000 r0 *1 25.65,68.6
X$2000 1794 1487 1822 23 38 1849 MUX2_X1
* cell instance $2001 m0 *1 29.07,68.6
X$2001 1694 1184 1764 23 38 1851 MUX2_X1
* cell instance $2002 m0 *1 25.84,68.6
X$2002 23 2824 1764 1763 1693 38 DFF_X1
* cell instance $2003 m0 *1 30.4,68.6
X$2003 23 38 FILLCELL_X8
* cell instance $2004 m0 *1 31.92,68.6
X$2004 23 38 FILLCELL_X4
* cell instance $2005 m0 *1 32.68,68.6
X$2005 23 38 FILLCELL_X2
* cell instance $2006 r0 *1 26.98,68.6
X$2006 23 2999 1794 1849 1693 38 DFF_X1
* cell instance $2007 r0 *1 30.21,68.6
X$2007 23 38 FILLCELL_X16
* cell instance $2008 m0 *1 34.39,68.6
X$2008 23 38 FILLCELL_X16
* cell instance $2009 m0 *1 33.06,68.6
X$2009 1810 1487 1725 23 38 1812 MUX2_X1
* cell instance $2010 m0 *1 37.43,68.6
X$2010 23 38 FILLCELL_X8
* cell instance $2011 m0 *1 38.95,68.6
X$2011 23 38 FILLCELL_X2
* cell instance $2012 r0 *1 33.25,68.6
X$2012 23 38 FILLCELL_X1
* cell instance $2013 r0 *1 33.44,68.6
X$2013 23 2973 1810 1812 1795 38 DFF_X1
* cell instance $2014 r0 *1 36.67,68.6
X$2014 23 38 FILLCELL_X4
* cell instance $2015 r0 *1 37.43,68.6
X$2015 23 2983 1825 1854 1639 38 DFF_X1
* cell instance $2016 m0 *1 39.52,68.6
X$2016 1732 1177 23 38 1796 NOR2_X1
* cell instance $2017 m0 *1 39.33,68.6
X$2017 23 38 FILLCELL_X1
* cell instance $2018 m0 *1 40.09,68.6
X$2018 23 38 FILLCELL_X2
* cell instance $2019 m0 *1 41.42,68.6
X$2019 1733 1487 1813 23 38 1766 MUX2_X1
* cell instance $2020 m0 *1 40.47,68.6
X$2020 1486 23 38 1639 CLKBUF_X3
* cell instance $2021 m0 *1 42.75,68.6
X$2021 1782 1488 1813 23 38 1783 MUX2_X1
* cell instance $2022 m0 *1 44.08,68.6
X$2022 23 2814 1782 1783 1639 38 DFF_X1
* cell instance $2023 m0 *1 47.31,68.6
X$2023 23 38 FILLCELL_X4
* cell instance $2024 m0 *1 48.07,68.6
X$2024 1784 1434 1767 23 38 1816 MUX2_X1
* cell instance $2025 m0 *1 49.4,68.6
X$2025 23 2602 1784 1816 1735 38 DFF_X1
* cell instance $2026 m0 *1 52.63,68.6
X$2026 23 38 FILLCELL_X4
* cell instance $2027 m0 *1 53.39,68.6
X$2027 1641 1736 1511 1787 38 23 1863 OAI22_X2
* cell instance $2028 m0 *1 55.1,68.6
X$2028 23 38 FILLCELL_X4
* cell instance $2029 m0 *1 55.86,68.6
X$2029 23 2603 1737 1768 1735 38 DFF_X1
* cell instance $2030 m0 *1 59.09,68.6
X$2030 23 38 FILLCELL_X8
* cell instance $2031 m0 *1 60.61,68.6
X$2031 23 38 FILLCELL_X2
* cell instance $2032 r0 *1 40.66,68.6
X$2032 1825 1488 1730 23 38 1854 MUX2_X1
* cell instance $2033 r0 *1 41.99,68.6
X$2033 23 1331 1765 38 BUF_X32
* cell instance $2034 r0 *1 51.3,68.6
X$2034 23 38 FILLCELL_X8
* cell instance $2035 r0 *1 52.82,68.6
X$2035 23 38 FILLCELL_X4
* cell instance $2036 r0 *1 53.58,68.6
X$2036 23 38 FILLCELL_X2
* cell instance $2037 r0 *1 53.96,68.6
X$2037 23 38 FILLCELL_X1
* cell instance $2038 r0 *1 54.15,68.6
X$2038 1636 1797 23 38 1865 NAND2_X1
* cell instance $2039 r0 *1 54.72,68.6
X$2039 23 2888 1797 1861 1735 38 DFF_X1
* cell instance $2040 r0 *1 57.95,68.6
X$2040 23 38 FILLCELL_X32
* cell instance $2041 r0 *1 59.14,68.6
X$2041 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $2042 r0 *1 59.14,68.6
X$2042 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $2043 r0 *1 59.14,68.6
X$2043 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $2044 m0 *1 61.18,68.6
X$2044 1738 559 1561 23 38 1788 MUX2_X1
* cell instance $2045 m0 *1 60.99,68.6
X$2045 23 38 FILLCELL_X1
* cell instance $2046 m0 *1 62.51,68.6
X$2046 1392 23 38 1684 CLKBUF_X3
* cell instance $2047 m0 *1 63.46,68.6
X$2047 1684 23 38 CLKBUF_X1
* cell instance $2048 m0 *1 64.03,68.6
X$2048 1755 1728 23 38 1798 NAND2_X1
* cell instance $2049 m0 *1 64.6,68.6
X$2049 1769 1177 23 38 1818 NOR2_X1
* cell instance $2050 m0 *1 65.17,68.6
X$2050 23 38 FILLCELL_X4
* cell instance $2051 m0 *1 65.93,68.6
X$2051 23 38 FILLCELL_X1
* cell instance $2052 m0 *1 66.12,68.6
X$2052 1335 23 38 1561 CLKBUF_X2
* cell instance $2053 m0 *1 66.88,68.6
X$2053 1785 1563 1787 1305 38 23 1817 OAI22_X1
* cell instance $2054 m0 *1 67.83,68.6
X$2054 23 38 FILLCELL_X1
* cell instance $2055 m0 *1 68.02,68.6
X$2055 1785 1563 1241 1506 1727 38 23 1772 OAI221_X1
* cell instance $2056 m0 *1 69.16,68.6
X$2056 23 38 FILLCELL_X2
* cell instance $2057 r0 *1 64.03,68.6
X$2057 1817 1765 1798 38 23 1857 OAI21_X2
* cell instance $2058 r0 *1 65.36,68.6
X$2058 23 38 FILLCELL_X2
* cell instance $2059 r0 *1 65.74,68.6
X$2059 475 1881 1818 476 1882 1799 23 38 1785 OAI33_X1
* cell instance $2060 r0 *1 67.07,68.6
X$2060 23 38 FILLCELL_X2
* cell instance $2061 r0 *1 67.45,68.6
X$2061 23 2870 1828 1814 1915 38 DFF_X1
* cell instance $2062 m0 *1 70.11,68.6
X$2062 23 38 FILLCELL_X8
* cell instance $2063 m0 *1 69.54,68.6
X$2063 1800 1537 23 38 1799 NOR2_X1
* cell instance $2064 m0 *1 71.63,68.6
X$2064 23 38 FILLCELL_X1
* cell instance $2065 m0 *1 71.82,68.6
X$2065 1801 559 1770 23 38 1815 MUX2_X1
* cell instance $2066 m0 *1 73.15,68.6
X$2066 23 38 FILLCELL_X2
* cell instance $2067 r0 *1 70.68,68.6
X$2067 23 38 FILLCELL_X1
* cell instance $2068 r0 *1 70.87,68.6
X$2068 23 3101 1801 1815 1644 38 DFF_X1
* cell instance $2069 m0 *1 73.72,68.6
X$2069 23 2667 1802 1771 1644 38 DFF_X1
* cell instance $2070 m0 *1 73.53,68.6
X$2070 23 38 FILLCELL_X1
* cell instance $2071 m0 *1 76.95,68.6
X$2071 23 38 FILLCELL_X4
* cell instance $2072 m0 *1 77.71,68.6
X$2072 1743 1811 1772 1804 1809 38 23 1756 OAI221_X1
* cell instance $2073 m0 *1 78.85,68.6
X$2073 23 38 FILLCELL_X2
* cell instance $2074 r0 *1 74.1,68.6
X$2074 1801 541 1802 23 38 1803 MUX2_X1
* cell instance $2075 r0 *1 75.43,68.6
X$2075 23 38 FILLCELL_X1
* cell instance $2076 r0 *1 75.62,68.6
X$2076 1803 1177 23 38 1846 NOR2_X1
* cell instance $2077 r0 *1 76.19,68.6
X$2077 1830 1105 23 38 1831 NOR2_X1
* cell instance $2078 r0 *1 76.76,68.6
X$2078 23 38 FILLCELL_X2
* cell instance $2079 r0 *1 77.14,68.6
X$2079 475 1831 1846 476 1844 1832 23 38 1706 OAI33_X1
* cell instance $2080 r0 *1 78.47,68.6
X$2080 1837 1537 23 38 1832 NOR2_X1
* cell instance $2081 r0 *1 79.04,68.6
X$2081 23 38 FILLCELL_X4
* cell instance $2082 m0 *1 79.8,68.6
X$2082 23 38 FILLCELL_X1
* cell instance $2083 m0 *1 79.23,68.6
X$2083 1228 1755 23 38 1811 NAND2_X1
* cell instance $2084 m0 *1 79.99,68.6
X$2084 1755 1239 23 38 1809 NAND2_X1
* cell instance $2085 m0 *1 80.56,68.6
X$2085 23 38 FILLCELL_X8
* cell instance $2086 m0 *1 82.08,68.6
X$2086 23 38 FILLCELL_X1
* cell instance $2087 m0 *1 82.27,68.6
X$2087 1805 88 1770 23 38 1808 MUX2_X1
* cell instance $2088 m0 *1 83.6,68.6
X$2088 23 38 FILLCELL_X4
* cell instance $2089 m0 *1 84.36,68.6
X$2089 1805 724 1740 23 38 1773 MUX2_X1
* cell instance $2090 m0 *1 85.69,68.6
X$2090 23 38 FILLCELL_X2
* cell instance $2091 r0 *1 79.8,68.6
X$2091 23 38 FILLCELL_X1
* cell instance $2092 r0 *1 79.99,68.6
X$2092 1392 23 38 1648 CLKBUF_X3
* cell instance $2093 r0 *1 80.94,68.6
X$2093 1648 23 38 CLKBUF_X1
* cell instance $2094 r0 *1 81.51,68.6
X$2094 23 38 FILLCELL_X1
* cell instance $2095 r0 *1 81.7,68.6
X$2095 23 2891 1805 1808 1648 38 DFF_X1
* cell instance $2096 r0 *1 84.93,68.6
X$2096 23 2884 1741 1807 1714 38 DFF_X1
* cell instance $2097 m0 *1 86.26,68.6
X$2097 1741 223 1770 23 38 1807 MUX2_X1
* cell instance $2098 m0 *1 86.07,68.6
X$2098 23 38 FILLCELL_X1
* cell instance $2099 m0 *1 87.59,68.6
X$2099 1750 174 1770 23 38 1774 MUX2_X1
* cell instance $2100 m0 *1 88.92,68.6
X$2100 1392 23 38 1714 CLKBUF_X3
* cell instance $2101 m0 *1 89.87,68.6
X$2101 1714 23 38 3142 INV_X1
* cell instance $2102 m0 *1 90.25,68.6
X$2102 1743 1777 1711 1804 1776 38 23 1806 OAI221_X1
* cell instance $2103 m0 *1 91.39,68.6
X$2103 23 38 FILLCELL_X2
* cell instance $2104 r0 *1 88.16,68.6
X$2104 23 38 FILLCELL_X8
* cell instance $2105 r0 *1 89.68,68.6
X$2105 23 38 FILLCELL_X1
* cell instance $2106 r0 *1 89.87,68.6
X$2106 23 2882 1742 1806 1714 38 DFF_X1
* cell instance $2107 m0 *1 92.34,68.6
X$2107 23 38 FILLCELL_X2
* cell instance $2108 m0 *1 91.77,68.6
X$2108 1742 1239 23 38 1776 NAND2_X1
* cell instance $2109 m0 *1 92.91,68.6
X$2109 23 2575 1745 1775 1714 38 DFF_X1
* cell instance $2110 m0 *1 92.72,68.6
X$2110 23 38 FILLCELL_X1
* cell instance $2111 m0 *1 96.14,68.6
X$2111 23 38 FILLCELL_X4
* cell instance $2112 m0 *1 96.9,68.6
X$2112 23 38 FILLCELL_X1
* cell instance $2113 r180 *1 97.28,68.6
X$2113 23 38 23 38 TAPCELL_X1
* cell instance $2114 r0 *1 93.1,68.6
X$2114 23 38 FILLCELL_X16
* cell instance $2115 r0 *1 96.14,68.6
X$2115 23 38 FILLCELL_X4
* cell instance $2116 r0 *1 96.9,68.6
X$2116 23 38 FILLCELL_X1
* cell instance $2117 m90 *1 97.28,68.6
X$2117 23 38 23 38 TAPCELL_X1
* cell instance $2118 m0 *1 1.33,93.8
X$2118 23 38 FILLCELL_X16
* cell instance $2119 m0 *1 1.14,93.8
X$2119 23 38 23 38 TAPCELL_X1
* cell instance $2120 m0 *1 4.37,93.8
X$2120 23 38 FILLCELL_X4
* cell instance $2121 m0 *1 5.13,93.8
X$2121 23 38 FILLCELL_X1
* cell instance $2122 m0 *1 5.32,93.8
X$2122 23 2651 2474 2511 2434 38 DFF_X1
* cell instance $2123 m0 *1 8.55,93.8
X$2123 23 38 FILLCELL_X4
* cell instance $2124 m0 *1 9.31,93.8
X$2124 23 38 FILLCELL_X1
* cell instance $2125 m0 *1 9.5,93.8
X$2125 23 2672 2433 2461 2434 38 DFF_X1
* cell instance $2126 m0 *1 12.73,93.8
X$2126 2199 1480 2463 23 38 2488 MUX2_X1
* cell instance $2127 m0 *1 14.06,93.8
X$2127 2434 23 38 CLKBUF_X1
* cell instance $2128 m0 *1 14.63,93.8
X$2128 2217 1346 2489 23 38 2435 MUX2_X1
* cell instance $2129 m0 *1 15.96,93.8
X$2129 2217 1406 2475 23 38 2465 MUX2_X1
* cell instance $2130 m0 *1 17.29,93.8
X$2130 2475 1358 2489 23 38 2466 MUX2_X1
* cell instance $2131 m0 *1 18.62,93.8
X$2131 23 2673 2437 2436 2434 38 DFF_X1
* cell instance $2132 m0 *1 21.85,93.8
X$2132 2217 1493 2438 23 38 2439 MUX2_X1
* cell instance $2133 m0 *1 23.18,93.8
X$2133 23 38 FILLCELL_X8
* cell instance $2134 m0 *1 24.7,93.8
X$2134 23 38 FILLCELL_X1
* cell instance $2135 m0 *1 24.89,93.8
X$2135 23 2644 2440 2490 2355 38 DFF_X1
* cell instance $2136 m0 *1 28.12,93.8
X$2136 2218 1493 2441 23 38 2491 MUX2_X1
* cell instance $2137 m0 *1 29.45,93.8
X$2137 2218 1406 2495 23 38 2492 MUX2_X1
* cell instance $2138 m0 *1 30.78,93.8
X$2138 23 38 FILLCELL_X4
* cell instance $2139 m0 *1 31.54,93.8
X$2139 23 38 FILLCELL_X2
* cell instance $2140 r0 *1 1.14,93.8
X$2140 23 38 23 38 TAPCELL_X1
* cell instance $2141 r0 *1 1.33,93.8
X$2141 23 38 FILLCELL_X16
* cell instance $2142 r0 *1 3.14,93.8
X$2142 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $2143 r0 *1 3.14,93.4
X$2143 23 VIA_via5_6_960_2800_5_2_600_600
* cell instance $2144 r0 *1 3.14,93.4
X$2144 23 VIA_via4_5_960_2800_5_2_600_600
* cell instance $2145 r0 *1 3.14,93.4
X$2145 23 VIA_via6_7_960_2800_4_1_600_600
* cell instance $2146 r0 *1 3.14,93.8
X$2146 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $2147 r0 *1 3.14,93.8
X$2147 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $2148 r0 *1 4.37,93.8
X$2148 23 38 FILLCELL_X8
* cell instance $2149 r0 *1 5.89,93.8
X$2149 23 38 FILLCELL_X2
* cell instance $2150 r0 *1 6.27,93.8
X$2150 23 38 FILLCELL_X1
* cell instance $2151 r0 *1 6.46,93.8
X$2151 2199 1346 2474 23 38 2511 MUX2_X1
* cell instance $2152 r0 *1 7.79,93.8
X$2152 23 38 FILLCELL_X2
* cell instance $2153 r0 *1 8.17,93.8
X$2153 23 38 FILLCELL_X1
* cell instance $2154 r0 *1 8.36,93.8
X$2154 2432 1358 2474 23 38 2418 MUX2_X1
* cell instance $2155 r0 *1 9.69,93.8
X$2155 23 38 FILLCELL_X4
* cell instance $2156 r0 *1 10.45,93.8
X$2156 23 38 FILLCELL_X2
* cell instance $2157 r0 *1 10.83,93.8
X$2157 23 2962 2463 2488 2434 38 DFF_X1
* cell instance $2158 r0 *1 14.06,93.8
X$2158 23 38 FILLCELL_X1
* cell instance $2159 r0 *1 14.25,93.8
X$2159 23 2965 2489 2435 2434 38 DFF_X1
* cell instance $2160 r0 *1 17.48,93.8
X$2160 23 38 FILLCELL_X32
* cell instance $2161 r0 *1 23.56,93.8
X$2161 23 38 FILLCELL_X8
* cell instance $2162 r0 *1 25.08,93.8
X$2162 23 3079 2441 2491 2355 38 DFF_X1
* cell instance $2163 r0 *1 28.31,93.8
X$2163 23 38 FILLCELL_X4
* cell instance $2164 r0 *1 29.07,93.8
X$2164 23 38 FILLCELL_X1
* cell instance $2165 r0 *1 29.26,93.8
X$2165 23 3075 2495 2492 2355 38 DFF_X1
* cell instance $2166 m0 *1 33.25,93.8
X$2166 23 38 FILLCELL_X8
* cell instance $2167 m0 *1 31.92,93.8
X$2167 2495 1358 2505 23 38 2442 MUX2_X1
* cell instance $2168 m0 *1 34.77,93.8
X$2168 23 38 FILLCELL_X4
* cell instance $2169 m0 *1 35.53,93.8
X$2169 23 2634 2497 2496 2355 38 DFF_X1
* cell instance $2170 m0 *1 38.76,93.8
X$2170 2220 1406 2497 23 38 2496 MUX2_X1
* cell instance $2171 m0 *1 40.09,93.8
X$2171 23 38 FILLCELL_X4
* cell instance $2172 m0 *1 40.85,93.8
X$2172 2220 1493 2443 23 38 2469 MUX2_X1
* cell instance $2173 m0 *1 42.18,93.8
X$2173 2443 1373 2558 23 38 2426 MUX2_X1
* cell instance $2174 m0 *1 43.51,93.8
X$2174 23 38 FILLCELL_X8
* cell instance $2175 m0 *1 45.03,93.8
X$2175 23 38 FILLCELL_X2
* cell instance $2176 r0 *1 32.49,93.8
X$2176 23 38 FILLCELL_X2
* cell instance $2177 r0 *1 32.87,93.8
X$2177 2218 1346 2505 23 38 2521 MUX2_X1
* cell instance $2178 r0 *1 34.2,93.8
X$2178 2355 23 38 CLKBUF_X1
* cell instance $2179 r0 *1 34.77,93.8
X$2179 23 38 FILLCELL_X4
* cell instance $2180 r0 *1 35.53,93.8
X$2180 23 38 FILLCELL_X1
* cell instance $2181 r0 *1 35.72,93.8
X$2181 23 3021 2524 2514 2355 38 DFF_X1
* cell instance $2182 r0 *1 38.95,93.8
X$2182 2497 1358 2524 23 38 2359 MUX2_X1
* cell instance $2183 r0 *1 40.28,93.8
X$2183 2220 1480 2558 23 38 2557 MUX2_X1
* cell instance $2184 r0 *1 41.61,93.8
X$2184 23 38 FILLCELL_X2
* cell instance $2185 r0 *1 41.99,93.8
X$2185 23 38 FILLCELL_X1
* cell instance $2186 r0 *1 42.18,93.8
X$2186 2052 23 38 2525 BUF_X1
* cell instance $2187 r0 *1 42.75,93.8
X$2187 23 38 FILLCELL_X16
* cell instance $2188 m0 *1 48.64,93.8
X$2188 2182 1406 2476 23 38 2499 MUX2_X1
* cell instance $2189 m0 *1 45.41,93.8
X$2189 23 2639 2476 2499 2333 38 DFF_X1
* cell instance $2190 m0 *1 49.97,93.8
X$2190 23 38 FILLCELL_X2
* cell instance $2191 r0 *1 45.79,93.8
X$2191 23 38 FILLCELL_X2
* cell instance $2192 r0 *1 46.17,93.8
X$2192 2526 23 38 1587 BUF_X2
* cell instance $2193 r0 *1 46.93,93.8
X$2193 23 38 FILLCELL_X16
* cell instance $2194 r0 *1 49.97,93.8
X$2194 23 38 FILLCELL_X1
* cell instance $2195 r0 *1 50.16,93.8
X$2195 2182 1346 2506 23 38 2559 MUX2_X1
* cell instance $2196 m0 *1 51.68,93.8
X$2196 23 38 FILLCELL_X4
* cell instance $2197 m0 *1 50.35,93.8
X$2197 2476 1358 2506 23 38 2445 MUX2_X1
* cell instance $2198 m0 *1 52.44,93.8
X$2198 23 38 FILLCELL_X2
* cell instance $2199 r0 *1 51.49,93.8
X$2199 23 38 FILLCELL_X4
* cell instance $2200 r0 *1 52.25,93.8
X$2200 23 38 FILLCELL_X2
* cell instance $2201 r0 *1 52.63,93.8
X$2201 23 38 FILLCELL_X1
* cell instance $2202 r0 *1 52.82,93.8
X$2202 23 3126 2502 2477 2316 38 DFF_X1
* cell instance $2203 m0 *1 53.01,93.8
X$2203 2182 1493 2502 23 38 2477 MUX2_X1
* cell instance $2204 m0 *1 52.82,93.8
X$2204 23 38 FILLCELL_X1
* cell instance $2205 m0 *1 54.34,93.8
X$2205 23 38 FILLCELL_X2
* cell instance $2206 m0 *1 54.91,93.8
X$2206 2151 1493 2363 23 38 2447 MUX2_X1
* cell instance $2207 m0 *1 54.72,93.8
X$2207 23 38 FILLCELL_X1
* cell instance $2208 m0 *1 56.24,93.8
X$2208 23 38 FILLCELL_X32
* cell instance $2209 m0 *1 62.32,93.8
X$2209 23 38 FILLCELL_X16
* cell instance $2210 m0 *1 65.36,93.8
X$2210 2232 1240 23 38 2508 NAND2_X1
* cell instance $2211 m0 *1 65.93,93.8
X$2211 23 38 FILLCELL_X8
* cell instance $2212 m0 *1 67.45,93.8
X$2212 23 38 FILLCELL_X2
* cell instance $2213 r0 *1 56.05,93.8
X$2213 2502 1373 2507 23 38 2446 MUX2_X1
* cell instance $2214 r0 *1 57.38,93.8
X$2214 23 38 FILLCELL_X4
* cell instance $2215 r0 *1 58.14,93.8
X$2215 23 38 FILLCELL_X1
* cell instance $2216 r0 *1 58.33,93.8
X$2216 2182 1480 2507 23 38 2531 MUX2_X1
* cell instance $2217 r0 *1 59.14,93.8
X$2217 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $2218 r0 *1 59.14,93.4
X$2218 23 VIA_via5_6_960_2800_5_2_600_600
* cell instance $2219 r0 *1 59.14,93.4
X$2219 23 VIA_via4_5_960_2800_5_2_600_600
* cell instance $2220 r0 *1 59.14,93.4
X$2220 23 VIA_via6_7_960_2800_4_1_600_600
* cell instance $2221 r0 *1 59.14,93.8
X$2221 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $2222 r0 *1 59.14,93.8
X$2222 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $2223 r0 *1 59.66,93.8
X$2223 23 38 FILLCELL_X16
* cell instance $2224 r0 *1 62.7,93.8
X$2224 23 38 FILLCELL_X8
* cell instance $2225 r0 *1 64.22,93.8
X$2225 1857 23 38 2534 BUF_X1
* cell instance $2226 r0 *1 64.79,93.8
X$2226 2508 2155 23 38 2536 NOR2_X1
* cell instance $2227 r0 *1 65.36,93.8
X$2227 2508 23 38 2537 BUF_X1
* cell instance $2228 r0 *1 65.93,93.8
X$2228 2508 23 38 2561 INV_X1
* cell instance $2229 r0 *1 66.31,93.8
X$2229 23 38 FILLCELL_X16
* cell instance $2230 m0 *1 68.02,93.8
X$2230 2504 38 2478 23 BUF_X4
* cell instance $2231 m0 *1 67.83,93.8
X$2231 23 38 FILLCELL_X1
* cell instance $2232 m0 *1 69.35,93.8
X$2232 23 38 FILLCELL_X4
* cell instance $2233 m0 *1 70.11,93.8
X$2233 2503 2478 23 38 2479 NAND2_X1
* cell instance $2234 m0 *1 70.68,93.8
X$2234 2449 2478 2501 23 2448 38 AOI21_X1
* cell instance $2235 m0 *1 71.44,93.8
X$2235 23 2154 2480 2481 2500 2472 38 FA_X1
* cell instance $2236 m0 *1 74.48,93.8
X$2236 23 38 FILLCELL_X2
* cell instance $2237 r0 *1 69.35,93.8
X$2237 23 38 FILLCELL_X2
* cell instance $2238 r0 *1 69.73,93.8
X$2238 23 38 FILLCELL_X1
* cell instance $2239 r0 *1 69.92,93.8
X$2239 2448 2562 2479 38 23 2482 OAI21_X2
* cell instance $2240 r0 *1 71.25,93.8
X$2240 2480 2478 38 2452 23 XOR2_X2
* cell instance $2241 r0 *1 72.96,93.8
X$2241 23 38 FILLCELL_X4
* cell instance $2242 r0 *1 73.72,93.8
X$2242 2481 23 38 2409 BUF_X1
* cell instance $2243 r0 *1 74.29,93.8
X$2243 2452 2409 2451 2336 23 38 2513 NOR4_X1
* cell instance $2244 m0 *1 74.86,93.8
X$2244 2513 2498 2482 38 23 2156 MUX2_X2
* cell instance $2245 m0 *1 76.57,93.8
X$2245 2509 2453 2482 38 23 2287 MUX2_X2
* cell instance $2246 m0 *1 78.28,93.8
X$2246 2510 2494 2190 38 2493 23 OAI21_X1
* cell instance $2247 m0 *1 79.04,93.8
X$2247 1478 23 38 2057 BUF_X2
* cell instance $2248 m0 *1 79.8,93.8
X$2248 2549 2410 2550 23 38 2560 MUX2_X1
* cell instance $2249 m0 *1 81.13,93.8
X$2249 23 38 FILLCELL_X8
* cell instance $2250 m0 *1 82.65,93.8
X$2250 23 38 FILLCELL_X4
* cell instance $2251 m0 *1 83.41,93.8
X$2251 23 38 FILLCELL_X2
* cell instance $2252 r0 *1 75.24,93.8
X$2252 2336 2452 2409 2451 38 2509 23 OR4_X2
* cell instance $2253 r0 *1 76.57,93.8
X$2253 2336 2482 38 23 2510 XNOR2_X1
* cell instance $2254 r0 *1 77.71,93.8
X$2254 23 38 FILLCELL_X2
* cell instance $2255 r0 *1 78.09,93.8
X$2255 2455 1240 2546 2452 23 38 2563 NOR4_X1
* cell instance $2256 r0 *1 79.04,93.8
X$2256 2512 2057 38 23 2549 AND2_X1
* cell instance $2257 r0 *1 79.8,93.8
X$2257 23 38 FILLCELL_X2
* cell instance $2258 r0 *1 80.18,93.8
X$2258 23 3115 2512 2560 2373 38 DFF_X1
* cell instance $2259 r0 *1 83.41,93.8
X$2259 23 38 FILLCELL_X2
* cell instance $2260 m0 *1 1.33,79.8
X$2260 23 38 FILLCELL_X16
* cell instance $2261 m0 *1 1.14,79.8
X$2261 23 38 23 38 TAPCELL_X1
* cell instance $2262 m0 *1 4.37,79.8
X$2262 23 38 FILLCELL_X8
* cell instance $2263 m0 *1 5.89,79.8
X$2263 23 38 FILLCELL_X4
* cell instance $2264 m0 *1 6.65,79.8
X$2264 1909 23 38 1902 CLKBUF_X3
* cell instance $2265 m0 *1 7.6,79.8
X$2265 23 2656 2046 2123 2045 38 DFF_X1
* cell instance $2266 m0 *1 10.83,79.8
X$2266 23 38 FILLCELL_X2
* cell instance $2267 r0 *1 1.14,79.8
X$2267 23 38 23 38 TAPCELL_X1
* cell instance $2268 r0 *1 1.33,79.8
X$2268 23 38 FILLCELL_X2
* cell instance $2269 r0 *1 1.71,79.8
X$2269 23 38 FILLCELL_X1
* cell instance $2270 r0 *1 1.9,79.8
X$2270 23 2971 2165 2197 1902 38 DFF_X1
* cell instance $2271 r0 *1 3.14,79.8
X$2271 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $2272 r0 *1 3.14,79.8
X$2272 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $2273 r0 *1 3.14,79.8
X$2273 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $2274 r0 *1 5.13,79.8
X$2274 23 38 FILLCELL_X16
* cell instance $2275 r0 *1 8.17,79.8
X$2275 23 38 FILLCELL_X8
* cell instance $2276 r0 *1 9.69,79.8
X$2276 23 38 FILLCELL_X2
* cell instance $2277 r0 *1 10.07,79.8
X$2277 1935 1482 2046 23 38 2123 MUX2_X1
* cell instance $2278 m0 *1 11.4,79.8
X$2278 23 2670 2047 2072 1902 38 DFF_X1
* cell instance $2279 m0 *1 11.21,79.8
X$2279 23 38 FILLCELL_X1
* cell instance $2280 m0 *1 14.63,79.8
X$2280 23 38 FILLCELL_X4
* cell instance $2281 m0 *1 15.39,79.8
X$2281 23 38 FILLCELL_X2
* cell instance $2282 r0 *1 11.4,79.8
X$2282 23 38 FILLCELL_X16
* cell instance $2283 r0 *1 14.44,79.8
X$2283 23 38 FILLCELL_X4
* cell instance $2284 r0 *1 15.2,79.8
X$2284 1820 1492 2105 23 38 2142 MUX2_X1
* cell instance $2285 m0 *1 15.96,79.8
X$2285 2033 792 2047 23 38 2048 MUX2_X1
* cell instance $2286 m0 *1 15.77,79.8
X$2286 23 38 FILLCELL_X1
* cell instance $2287 m0 *1 17.29,79.8
X$2287 23 38 FILLCELL_X8
* cell instance $2288 m0 *1 18.81,79.8
X$2288 23 38 FILLCELL_X2
* cell instance $2289 r0 *1 16.53,79.8
X$2289 2105 792 2176 23 38 2077 MUX2_X1
* cell instance $2290 r0 *1 17.86,79.8
X$2290 23 38 FILLCELL_X2
* cell instance $2291 r0 *1 18.24,79.8
X$2291 23 38 FILLCELL_X1
* cell instance $2292 r0 *1 18.43,79.8
X$2292 1822 1544 2127 23 38 2143 MUX2_X1
* cell instance $2293 m0 *1 19.76,79.8
X$2293 23 38 FILLCELL_X32
* cell instance $2294 m0 *1 19.19,79.8
X$2294 2077 1537 23 38 2035 NOR2_X1
* cell instance $2295 m0 *1 25.84,79.8
X$2295 23 38 FILLCELL_X16
* cell instance $2296 m0 *1 28.88,79.8
X$2296 23 38 FILLCELL_X4
* cell instance $2297 m0 *1 29.64,79.8
X$2297 23 38 FILLCELL_X2
* cell instance $2298 r0 *1 19.76,79.8
X$2298 23 38 FILLCELL_X4
* cell instance $2299 r0 *1 20.52,79.8
X$2299 23 38 FILLCELL_X2
* cell instance $2300 r0 *1 20.9,79.8
X$2300 2127 813 2177 23 38 2080 MUX2_X1
* cell instance $2301 r0 *1 22.23,79.8
X$2301 23 38 FILLCELL_X4
* cell instance $2302 r0 *1 22.99,79.8
X$2302 23 38 FILLCELL_X2
* cell instance $2303 r0 *1 23.37,79.8
X$2303 1822 1492 2128 23 38 2167 MUX2_X1
* cell instance $2304 r0 *1 24.7,79.8
X$2304 23 38 FILLCELL_X4
* cell instance $2305 r0 *1 25.46,79.8
X$2305 2128 792 2178 23 38 2049 MUX2_X1
* cell instance $2306 r0 *1 26.79,79.8
X$2306 23 38 FILLCELL_X4
* cell instance $2307 r0 *1 27.55,79.8
X$2307 23 38 FILLCELL_X2
* cell instance $2308 r0 *1 27.93,79.8
X$2308 23 38 FILLCELL_X1
* cell instance $2309 r0 *1 28.12,79.8
X$2309 1725 1492 2106 23 38 2205 MUX2_X1
* cell instance $2310 r0 *1 29.45,79.8
X$2310 2106 792 2206 23 38 2088 MUX2_X1
* cell instance $2311 m0 *1 30.59,79.8
X$2311 1743 2083 2039 1804 2087 38 23 2086 OAI221_X1
* cell instance $2312 m0 *1 30.02,79.8
X$2312 1636 2050 23 38 2083 NAND2_X1
* cell instance $2313 m0 *1 31.73,79.8
X$2313 2084 1765 2085 38 23 2304 OAI21_X2
* cell instance $2314 m0 *1 33.06,79.8
X$2314 23 38 FILLCELL_X1
* cell instance $2315 m0 *1 33.25,79.8
X$2315 2050 1638 23 38 2087 NAND2_X1
* cell instance $2316 m0 *1 33.82,79.8
X$2316 2050 1728 23 38 2130 NAND2_X1
* cell instance $2317 m0 *1 34.39,79.8
X$2317 23 38 FILLCELL_X16
* cell instance $2318 m0 *1 37.43,79.8
X$2318 23 38 FILLCELL_X4
* cell instance $2319 m0 *1 38.19,79.8
X$2319 23 38 FILLCELL_X2
* cell instance $2320 r0 *1 30.78,79.8
X$2320 23 38 FILLCELL_X4
* cell instance $2321 r0 *1 31.54,79.8
X$2321 2082 2010 2130 38 23 2169 OAI21_X2
* cell instance $2322 r0 *1 32.87,79.8
X$2322 23 38 FILLCELL_X8
* cell instance $2323 r0 *1 34.39,79.8
X$2323 2107 1099 2180 23 38 2051 MUX2_X1
* cell instance $2324 r0 *1 35.72,79.8
X$2324 23 38 FILLCELL_X1
* cell instance $2325 r0 *1 35.91,79.8
X$2325 23 3020 2146 2173 1933 38 DFF_X1
* cell instance $2326 m0 *1 38.76,79.8
X$2326 23 2629 1945 2014 1933 38 DFF_X1
* cell instance $2327 m0 *1 38.57,79.8
X$2327 23 38 FILLCELL_X1
* cell instance $2328 m0 *1 41.99,79.8
X$2328 2109 1605 23 38 1974 NOR2_X1
* cell instance $2329 m0 *1 42.56,79.8
X$2329 23 38 FILLCELL_X8
* cell instance $2330 m0 *1 44.08,79.8
X$2330 23 38 FILLCELL_X4
* cell instance $2331 m0 *1 44.84,79.8
X$2331 23 38 FILLCELL_X1
* cell instance $2332 m0 *1 45.03,79.8
X$2332 1813 1544 2095 23 38 2133 MUX2_X1
* cell instance $2333 m0 *1 46.36,79.8
X$2333 23 38 FILLCELL_X4
* cell instance $2334 m0 *1 47.12,79.8
X$2334 2095 1099 2181 23 38 2044 MUX2_X1
* cell instance $2335 m0 *1 48.45,79.8
X$2335 23 2729 1946 2135 1960 38 DFF_X1
* cell instance $2336 m0 *1 51.68,79.8
X$2336 23 38 FILLCELL_X16
* cell instance $2337 m0 *1 54.72,79.8
X$2337 23 38 FILLCELL_X1
* cell instance $2338 m0 *1 54.91,79.8
X$2338 2053 2010 2103 38 23 2110 OAI21_X2
* cell instance $2339 m0 *1 56.24,79.8
X$2339 23 38 FILLCELL_X32
* cell instance $2340 m0 *1 62.32,79.8
X$2340 23 38 FILLCELL_X4
* cell instance $2341 m0 *1 63.08,79.8
X$2341 23 38 FILLCELL_X1
* cell instance $2342 m0 *1 63.27,79.8
X$2342 2102 2153 3133 38 23 2104 HA_X1
* cell instance $2343 m0 *1 65.17,79.8
X$2343 23 38 FILLCELL_X4
* cell instance $2344 m0 *1 65.93,79.8
X$2344 2111 23 38 1411 BUF_X2
* cell instance $2345 m0 *1 66.69,79.8
X$2345 23 38 FILLCELL_X4
* cell instance $2346 m0 *1 67.45,79.8
X$2346 23 38 FILLCELL_X1
* cell instance $2347 m0 *1 67.64,79.8
X$2347 2055 2057 38 23 2112 AND2_X1
* cell instance $2348 m0 *1 68.4,79.8
X$2348 23 38 FILLCELL_X4
* cell instance $2349 m0 *1 69.16,79.8
X$2349 23 2598 1982 2101 1981 38 DFF_X1
* cell instance $2350 m0 *1 72.39,79.8
X$2350 23 38 FILLCELL_X4
* cell instance $2351 m0 *1 73.15,79.8
X$2351 23 38 FILLCELL_X1
* cell instance $2352 m0 *1 73.34,79.8
X$2352 2056 2113 38 23 2136 AND2_X1
* cell instance $2353 m0 *1 74.1,79.8
X$2353 23 38 FILLCELL_X16
* cell instance $2354 m0 *1 77.14,79.8
X$2354 23 38 FILLCELL_X8
* cell instance $2355 m0 *1 78.66,79.8
X$2355 23 38 FILLCELL_X2
* cell instance $2356 r0 *1 39.14,79.8
X$2356 23 38 FILLCELL_X4
* cell instance $2357 r0 *1 39.9,79.8
X$2357 23 38 FILLCELL_X2
* cell instance $2358 r0 *1 40.28,79.8
X$2358 23 38 FILLCELL_X1
* cell instance $2359 r0 *1 40.47,79.8
X$2359 1730 1544 2108 23 38 2148 MUX2_X1
* cell instance $2360 r0 *1 41.8,79.8
X$2360 2108 1099 2221 23 38 2109 MUX2_X1
* cell instance $2361 r0 *1 43.13,79.8
X$2361 23 38 FILLCELL_X4
* cell instance $2362 r0 *1 43.89,79.8
X$2362 23 38 FILLCELL_X2
* cell instance $2363 r0 *1 44.27,79.8
X$2363 23 3056 2095 2133 2149 38 DFF_X1
* cell instance $2364 r0 *1 47.5,79.8
X$2364 23 38 FILLCELL_X2
* cell instance $2365 r0 *1 47.88,79.8
X$2365 23 38 FILLCELL_X1
* cell instance $2366 r0 *1 48.07,79.8
X$2366 2182 1530 1946 23 38 2135 MUX2_X1
* cell instance $2367 r0 *1 49.4,79.8
X$2367 23 38 FILLCELL_X8
* cell instance $2368 r0 *1 50.92,79.8
X$2368 23 38 FILLCELL_X2
* cell instance $2369 r0 *1 51.3,79.8
X$2369 1767 1544 2138 23 38 2150 MUX2_X1
* cell instance $2370 r0 *1 52.63,79.8
X$2370 23 38 FILLCELL_X2
* cell instance $2371 r0 *1 53.01,79.8
X$2371 2058 23 38 1960 CLKBUF_X3
* cell instance $2372 r0 *1 53.96,79.8
X$2372 23 38 FILLCELL_X4
* cell instance $2373 r0 *1 54.72,79.8
X$2373 23 38 FILLCELL_X2
* cell instance $2374 r0 *1 55.1,79.8
X$2374 23 38 FILLCELL_X1
* cell instance $2375 r0 *1 55.29,79.8
X$2375 2138 1099 2211 23 38 2054 MUX2_X1
* cell instance $2376 r0 *1 56.62,79.8
X$2376 23 38 FILLCELL_X2
* cell instance $2377 r0 *1 57,79.8
X$2377 771 38 1530 23 BUF_X4
* cell instance $2378 r0 *1 58.33,79.8
X$2378 23 3088 2020 2152 1915 38 DFF_X1
* cell instance $2379 r0 *1 59.14,79.8
X$2379 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $2380 r0 *1 59.14,79.8
X$2380 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $2381 r0 *1 59.14,79.8
X$2381 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $2382 r0 *1 61.56,79.8
X$2382 23 2172 1915 2153 2154 38 DFF_X2
* cell instance $2383 r0 *1 65.17,79.8
X$2383 2186 2153 2055 38 23 2111 HA_X1
* cell instance $2384 r0 *1 67.07,79.8
X$2384 2102 2113 38 23 2171 AND2_X1
* cell instance $2385 r0 *1 67.83,79.8
X$2385 2139 2157 2112 23 38 2172 MUX2_X1
* cell instance $2386 r0 *1 69.16,79.8
X$2386 2154 2113 38 23 2139 AND2_X1
* cell instance $2387 r0 *1 69.92,79.8
X$2387 2137 1984 2170 23 38 2099 MUX2_X1
* cell instance $2388 r0 *1 71.25,79.8
X$2388 23 38 FILLCELL_X1
* cell instance $2389 r0 *1 71.44,79.8
X$2389 2058 23 38 3137 INV_X2
* cell instance $2390 r0 *1 72.01,79.8
X$2390 2136 1984 2170 23 38 2158 MUX2_X1
* cell instance $2391 r0 *1 73.34,79.8
X$2391 434 23 38 2058 CLKBUF_X3
* cell instance $2392 r0 *1 74.29,79.8
X$2392 23 38 FILLCELL_X2
* cell instance $2393 r0 *1 74.67,79.8
X$2393 2134 2114 2168 23 38 2212 MUX2_X1
* cell instance $2394 r0 *1 76,79.8
X$2394 23 38 FILLCELL_X2
* cell instance $2395 r0 *1 76.38,79.8
X$2395 2116 2115 23 38 2168 NOR2_X1
* cell instance $2396 r0 *1 76.95,79.8
X$2396 2115 1478 38 23 2134 AND2_X1
* cell instance $2397 r0 *1 77.71,79.8
X$2397 23 38 FILLCELL_X8
* cell instance $2398 m0 *1 79.99,79.8
X$2398 23 38 FILLCELL_X2
* cell instance $2399 m0 *1 79.04,79.8
X$2399 1983 23 38 2116 CLKBUF_X3
* cell instance $2400 r0 *1 79.23,79.8
X$2400 1478 23 38 2113 BUF_X2
* cell instance $2401 r0 *1 79.99,79.8
X$2401 1951 38 2065 23 BUF_X4
* cell instance $2402 m0 *1 80.94,79.8
X$2402 23 2625 2059 2096 1917 38 DFF_X1
* cell instance $2403 m0 *1 80.37,79.8
X$2403 2160 23 38 1519 INV_X2
* cell instance $2404 m0 *1 84.17,79.8
X$2404 23 2092 1917 2060 2022 38 DFF_X2
* cell instance $2405 m0 *1 87.78,79.8
X$2405 2022 2023 2061 38 23 2062 HA_X1
* cell instance $2406 m0 *1 89.68,79.8
X$2406 23 38 FILLCELL_X1
* cell instance $2407 m0 *1 89.87,79.8
X$2407 2063 2064 2062 23 38 2074 NAND3_X1
* cell instance $2408 m0 *1 90.63,79.8
X$2408 23 38 FILLCELL_X2
* cell instance $2409 r0 *1 81.32,79.8
X$2409 23 38 FILLCELL_X2
* cell instance $2410 r0 *1 81.7,79.8
X$2410 1949 2059 23 38 2117 NOR2_X1
* cell instance $2411 r0 *1 82.27,79.8
X$2411 2117 2159 2131 23 38 2096 MUX2_X1
* cell instance $2412 r0 *1 83.6,79.8
X$2412 2059 1460 38 23 2131 AND2_X1
* cell instance $2413 r0 *1 84.36,79.8
X$2413 2160 2059 38 23 2132 AND2_X1
* cell instance $2414 r0 *1 85.12,79.8
X$2414 2132 23 38 2063 BUF_X2
* cell instance $2415 r0 *1 85.88,79.8
X$2415 23 38 FILLCELL_X4
* cell instance $2416 r0 *1 86.64,79.8
X$2416 2060 2057 38 23 2089 AND2_X1
* cell instance $2417 r0 *1 87.4,79.8
X$2417 2061 2057 38 23 2118 AND2_X1
* cell instance $2418 r0 *1 88.16,79.8
X$2418 23 38 FILLCELL_X2
* cell instance $2419 r0 *1 88.54,79.8
X$2419 2023 2022 2064 2069 38 23 2161 AND4_X1
* cell instance $2420 r0 *1 89.68,79.8
X$2420 2063 2022 2023 23 38 2129 NAND3_X1
* cell instance $2421 r0 *1 90.44,79.8
X$2421 2129 1686 2065 23 38 2119 NOR3_X1
* cell instance $2422 m0 *1 91.01,79.8
X$2422 23 38 FILLCELL_X1
* cell instance $2423 m0 *1 91.2,79.8
X$2423 2074 1686 2065 23 38 2076 NOR3_X1
* cell instance $2424 m0 *1 91.96,79.8
X$2424 2120 2076 2066 23 38 2073 MUX2_X1
* cell instance $2425 m0 *1 93.29,79.8
X$2425 23 2633 2069 2073 2026 38 DFF_X1
* cell instance $2426 m0 *1 96.52,79.8
X$2426 2071 23 38 2068 BUF_X1
* cell instance $2427 r180 *1 97.28,79.8
X$2427 23 38 23 38 TAPCELL_X1
* cell instance $2428 r0 *1 91.2,79.8
X$2428 2064 2113 38 23 2121 AND2_X1
* cell instance $2429 r0 *1 91.96,79.8
X$2429 2121 2119 2125 23 38 2067 MUX2_X1
* cell instance $2430 r0 *1 93.29,79.8
X$2430 2116 2064 23 38 2125 NOR2_X1
* cell instance $2431 r0 *1 93.86,79.8
X$2431 2124 23 38 2070 BUF_X1
* cell instance $2432 r0 *1 94.43,79.8
X$2432 2025 23 38 2124 INV_X1
* cell instance $2433 r0 *1 94.81,79.8
X$2433 2023 23 38 2122 BUF_X1
* cell instance $2434 r0 *1 95.38,79.8
X$2434 23 38 FILLCELL_X2
* cell instance $2435 r0 *1 95.76,79.8
X$2435 23 38 FILLCELL_X1
* cell instance $2436 r0 *1 95.95,79.8
X$2436 2022 23 38 2164 BUF_X1
* cell instance $2437 r0 *1 96.52,79.8
X$2437 2064 23 38 2163 BUF_X1
* cell instance $2438 m90 *1 97.28,79.8
X$2438 23 38 23 38 TAPCELL_X1
* cell instance $2439 m0 *1 1.33,18.2
X$2439 23 38 FILLCELL_X16
* cell instance $2440 m0 *1 1.14,18.2
X$2440 23 38 23 38 TAPCELL_X1
* cell instance $2441 m0 *1 4.37,18.2
X$2441 23 38 FILLCELL_X8
* cell instance $2442 m0 *1 5.89,18.2
X$2442 23 38 FILLCELL_X2
* cell instance $2443 r0 *1 1.14,18.2
X$2443 23 38 23 38 TAPCELL_X1
* cell instance $2444 r0 *1 1.33,18.2
X$2444 23 38 FILLCELL_X4
* cell instance $2445 r0 *1 2.09,18.2
X$2445 23 3039 448 446 447 38 DFF_X1
* cell instance $2446 r0 *1 3.14,18.2
X$2446 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $2447 r0 *1 3.14,18.2
X$2447 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $2448 r0 *1 3.14,18.2
X$2448 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $2449 r0 *1 5.32,18.2
X$2449 23 3040 411 450 447 38 DFF_X1
* cell instance $2450 m0 *1 9.5,18.2
X$2450 411 412 391 23 38 416 MUX2_X1
* cell instance $2451 m0 *1 6.27,18.2
X$2451 23 2745 391 449 447 38 DFF_X1
* cell instance $2452 m0 *1 10.83,18.2
X$2452 23 2782 392 413 503 38 DFF_X1
* cell instance $2453 m0 *1 14.06,18.2
X$2453 392 393 295 23 38 413 MUX2_X1
* cell instance $2454 m0 *1 15.39,18.2
X$2454 23 38 FILLCELL_X2
* cell instance $2455 r0 *1 8.55,18.2
X$2455 391 257 453 23 38 449 MUX2_X1
* cell instance $2456 r0 *1 9.88,18.2
X$2456 23 38 FILLCELL_X8
* cell instance $2457 r0 *1 11.4,18.2
X$2457 23 38 FILLCELL_X4
* cell instance $2458 r0 *1 12.16,18.2
X$2458 23 38 FILLCELL_X2
* cell instance $2459 r0 *1 12.54,18.2
X$2459 23 38 FILLCELL_X1
* cell instance $2460 r0 *1 12.73,18.2
X$2460 451 437 295 23 38 488 MUX2_X1
* cell instance $2461 r0 *1 14.06,18.2
X$2461 23 38 FILLCELL_X4
* cell instance $2462 r0 *1 14.82,18.2
X$2462 392 472 451 23 38 355 MUX2_X1
* cell instance $2463 m0 *1 16.34,18.2
X$2463 23 2741 432 394 503 38 DFF_X1
* cell instance $2464 m0 *1 15.77,18.2
X$2464 416 354 23 38 380 NOR2_X1
* cell instance $2465 m0 *1 19.57,18.2
X$2465 23 38 FILLCELL_X2
* cell instance $2466 r0 *1 16.15,18.2
X$2466 432 393 453 23 38 394 MUX2_X1
* cell instance $2467 r0 *1 17.48,18.2
X$2467 23 38 FILLCELL_X4
* cell instance $2468 r0 *1 18.24,18.2
X$2468 23 38 FILLCELL_X1
* cell instance $2469 r0 *1 18.43,18.2
X$2469 432 472 466 23 38 395 MUX2_X1
* cell instance $2470 r0 *1 19.76,18.2
X$2470 23 38 FILLCELL_X16
* cell instance $2471 m0 *1 20.52,18.2
X$2471 356 359 380 360 417 396 23 38 433 OAI33_X1
* cell instance $2472 m0 *1 19.95,18.2
X$2472 395 381 23 38 359 NOR2_X1
* cell instance $2473 m0 *1 21.85,18.2
X$2473 23 38 FILLCELL_X16
* cell instance $2474 m0 *1 24.89,18.2
X$2474 356 455 418 360 361 327 23 38 397 OAI33_X1
* cell instance $2475 m0 *1 26.22,18.2
X$2475 23 38 FILLCELL_X2
* cell instance $2476 r0 *1 22.8,18.2
X$2476 23 38 FILLCELL_X8
* cell instance $2477 r0 *1 24.32,18.2
X$2477 23 38 FILLCELL_X2
* cell instance $2478 r0 *1 24.7,18.2
X$2478 23 38 FILLCELL_X1
* cell instance $2479 r0 *1 24.89,18.2
X$2479 467 381 23 38 455 NOR2_X1
* cell instance $2480 r0 *1 25.46,18.2
X$2480 23 38 FILLCELL_X1
* cell instance $2481 r0 *1 25.65,18.2
X$2481 434 23 38 149 CLKBUF_X3
* cell instance $2482 r0 *1 26.6,18.2
X$2482 23 38 FILLCELL_X8
* cell instance $2483 m0 *1 27.17,18.2
X$2483 23 38 FILLCELL_X8
* cell instance $2484 m0 *1 26.6,18.2
X$2484 362 354 23 38 418 NOR2_X1
* cell instance $2485 m0 *1 28.69,18.2
X$2485 23 38 FILLCELL_X4
* cell instance $2486 m0 *1 29.45,18.2
X$2486 23 38 FILLCELL_X2
* cell instance $2487 r0 *1 28.12,18.2
X$2487 468 437 421 23 38 495 MUX2_X1
* cell instance $2488 r0 *1 29.45,18.2
X$2488 23 38 FILLCELL_X16
* cell instance $2489 m0 *1 30.02,18.2
X$2489 328 257 421 23 38 387 MUX2_X1
* cell instance $2490 m0 *1 29.83,18.2
X$2490 23 38 FILLCELL_X1
* cell instance $2491 m0 *1 31.35,18.2
X$2491 356 469 363 360 364 365 23 38 422 OAI33_X1
* cell instance $2492 m0 *1 32.68,18.2
X$2492 23 38 FILLCELL_X16
* cell instance $2493 m0 *1 35.72,18.2
X$2493 23 38 FILLCELL_X8
* cell instance $2494 m0 *1 37.24,18.2
X$2494 23 38 FILLCELL_X1
* cell instance $2495 m0 *1 37.43,18.2
X$2495 366 318 319 23 38 389 MUX2_X1
* cell instance $2496 m0 *1 38.76,18.2
X$2496 23 38 FILLCELL_X2
* cell instance $2497 r0 *1 32.49,18.2
X$2497 23 38 FILLCELL_X8
* cell instance $2498 r0 *1 34.01,18.2
X$2498 356 459 458 360 253 388 23 38 423 OAI33_X1
* cell instance $2499 r0 *1 35.34,18.2
X$2499 435 381 23 38 459 NOR2_X1
* cell instance $2500 r0 *1 35.91,18.2
X$2500 23 38 FILLCELL_X32
* cell instance $2501 m0 *1 39.33,18.2
X$2501 98 23 38 319 BUF_X2
* cell instance $2502 m0 *1 39.14,18.2
X$2502 23 38 FILLCELL_X1
* cell instance $2503 m0 *1 40.09,18.2
X$2503 356 436 425 360 331 429 23 38 428 OAI33_X1
* cell instance $2504 m0 *1 41.42,18.2
X$2504 23 38 FILLCELL_X8
* cell instance $2505 m0 *1 42.94,18.2
X$2505 23 38 FILLCELL_X2
* cell instance $2506 r0 *1 41.99,18.2
X$2506 23 38 FILLCELL_X8
* cell instance $2507 m0 *1 43.51,18.2
X$2507 368 318 398 23 38 350 MUX2_X1
* cell instance $2508 m0 *1 43.32,18.2
X$2508 23 38 FILLCELL_X1
* cell instance $2509 m0 *1 44.84,18.2
X$2509 369 367 23 38 399 NOR2_X1
* cell instance $2510 m0 *1 45.41,18.2
X$2510 23 38 FILLCELL_X2
* cell instance $2511 r0 *1 43.51,18.2
X$2511 23 38 FILLCELL_X4
* cell instance $2512 r0 *1 44.27,18.2
X$2512 356 471 399 360 430 400 23 38 460 OAI33_X1
* cell instance $2513 r0 *1 45.6,18.2
X$2513 149 23 38 299 CLKBUF_X3
* cell instance $2514 m0 *1 46.74,18.2
X$2514 23 2727 402 401 299 38 DFF_X1
* cell instance $2515 m0 *1 45.79,18.2
X$2515 403 23 38 370 CLKBUF_X3
* cell instance $2516 m0 *1 49.97,18.2
X$2516 23 38 FILLCELL_X4
* cell instance $2517 m0 *1 50.73,18.2
X$2517 23 38 FILLCELL_X2
* cell instance $2518 r0 *1 46.55,18.2
X$2518 23 38 FILLCELL_X1
* cell instance $2519 r0 *1 46.74,18.2
X$2519 402 393 301 23 38 401 MUX2_X1
* cell instance $2520 r0 *1 48.07,18.2
X$2520 463 437 301 23 38 352 MUX2_X1
* cell instance $2521 r0 *1 49.4,18.2
X$2521 402 472 463 23 38 464 MUX2_X1
* cell instance $2522 r0 *1 50.73,18.2
X$2522 23 38 FILLCELL_X4
* cell instance $2523 m0 *1 52.06,18.2
X$2523 356 404 371 360 427 390 23 38 426 OAI33_X1
* cell instance $2524 m0 *1 51.11,18.2
X$2524 403 23 38 248 CLKBUF_X3
* cell instance $2525 m0 *1 53.39,18.2
X$2525 23 38 FILLCELL_X4
* cell instance $2526 m0 *1 54.15,18.2
X$2526 23 38 FILLCELL_X2
* cell instance $2527 r0 *1 51.49,18.2
X$2527 23 38 FILLCELL_X2
* cell instance $2528 r0 *1 51.87,18.2
X$2528 464 370 23 38 404 NOR2_X1
* cell instance $2529 r0 *1 52.44,18.2
X$2529 23 38 FILLCELL_X16
* cell instance $2530 m0 *1 55.1,18.2
X$2530 23 38 FILLCELL_X16
* cell instance $2531 m0 *1 54.53,18.2
X$2531 405 372 23 38 427 NOR2_X1
* cell instance $2532 m0 *1 58.14,18.2
X$2532 23 38 FILLCELL_X1
* cell instance $2533 m0 *1 58.33,18.2
X$2533 424 372 23 38 517 NOR2_X1
* cell instance $2534 m0 *1 58.9,18.2
X$2534 23 38 FILLCELL_X1
* cell instance $2535 m0 *1 59.09,18.2
X$2535 23 2714 439 462 158 38 DFF_X1
* cell instance $2536 m0 *1 62.32,18.2
X$2536 386 373 48 23 38 347 MUX2_X1
* cell instance $2537 m0 *1 63.65,18.2
X$2537 23 38 FILLCELL_X8
* cell instance $2538 m0 *1 65.17,18.2
X$2538 23 38 FILLCELL_X2
* cell instance $2539 r0 *1 55.48,18.2
X$2539 23 38 FILLCELL_X1
* cell instance $2540 r0 *1 55.67,18.2
X$2540 139 23 38 158 CLKBUF_X3
* cell instance $2541 r0 *1 56.62,18.2
X$2541 158 23 38 CLKBUF_X1
* cell instance $2542 r0 *1 57.19,18.2
X$2542 23 38 FILLCELL_X16
* cell instance $2543 r0 *1 59.14,18.2
X$2543 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $2544 r0 *1 59.14,18.2
X$2544 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $2545 r0 *1 59.14,18.2
X$2545 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $2546 r0 *1 60.23,18.2
X$2546 23 38 FILLCELL_X1
* cell instance $2547 r0 *1 60.42,18.2
X$2547 439 441 48 23 38 462 MUX2_X1
* cell instance $2548 r0 *1 61.75,18.2
X$2548 439 438 386 23 38 461 MUX2_X1
* cell instance $2549 r0 *1 63.08,18.2
X$2549 23 38 FILLCELL_X4
* cell instance $2550 r0 *1 63.84,18.2
X$2550 23 38 FILLCELL_X2
* cell instance $2551 r0 *1 64.22,18.2
X$2551 23 38 FILLCELL_X1
* cell instance $2552 r0 *1 64.41,18.2
X$2552 461 370 23 38 440 NOR2_X1
* cell instance $2553 r0 *1 64.98,18.2
X$2553 23 38 FILLCELL_X2
* cell instance $2554 r0 *1 65.36,18.2
X$2554 23 38 FILLCELL_X1
* cell instance $2555 m0 *1 65.74,18.2
X$2555 306 374 23 38 406 NOR2_X1
* cell instance $2556 m0 *1 65.55,18.2
X$2556 23 38 FILLCELL_X1
* cell instance $2557 m0 *1 66.31,18.2
X$2557 23 38 FILLCELL_X1
* cell instance $2558 m0 *1 66.5,18.2
X$2558 23 2851 384 385 153 38 DFF_X1
* cell instance $2559 m0 *1 69.73,18.2
X$2559 420 374 23 38 419 NOR2_X1
* cell instance $2560 m0 *1 70.3,18.2
X$2560 23 38 FILLCELL_X1
* cell instance $2561 m0 *1 70.49,18.2
X$2561 262 372 23 38 407 NOR2_X1
* cell instance $2562 m0 *1 71.06,18.2
X$2562 23 38 FILLCELL_X4
* cell instance $2563 m0 *1 71.82,18.2
X$2563 23 38 FILLCELL_X1
* cell instance $2564 m0 *1 72.01,18.2
X$2564 23 2688 454 408 334 38 DFF_X1
* cell instance $2565 m0 *1 75.24,18.2
X$2565 23 38 FILLCELL_X2
* cell instance $2566 r0 *1 65.55,18.2
X$2566 105 372 23 38 496 NOR2_X1
* cell instance $2567 r0 *1 66.12,18.2
X$2567 23 38 FILLCELL_X8
* cell instance $2568 r0 *1 67.64,18.2
X$2568 457 441 78 23 38 494 MUX2_X1
* cell instance $2569 r0 *1 68.97,18.2
X$2569 457 438 384 23 38 456 MUX2_X1
* cell instance $2570 r0 *1 70.3,18.2
X$2570 456 370 23 38 442 NOR2_X1
* cell instance $2571 r0 *1 70.87,18.2
X$2571 23 38 FILLCELL_X8
* cell instance $2572 r0 *1 72.39,18.2
X$2572 23 38 FILLCELL_X1
* cell instance $2573 r0 *1 72.58,18.2
X$2573 454 441 52 23 38 408 MUX2_X1
* cell instance $2574 r0 *1 73.91,18.2
X$2574 434 23 38 139 CLKBUF_X3
* cell instance $2575 r0 *1 74.86,18.2
X$2575 23 38 FILLCELL_X2
* cell instance $2576 r0 *1 75.24,18.2
X$2576 454 438 375 23 38 452 MUX2_X1
* cell instance $2577 m0 *1 75.81,18.2
X$2577 375 373 52 23 38 383 MUX2_X1
* cell instance $2578 m0 *1 75.62,18.2
X$2578 23 38 FILLCELL_X1
* cell instance $2579 m0 *1 77.14,18.2
X$2579 23 38 FILLCELL_X1
* cell instance $2580 m0 *1 77.33,18.2
X$2580 52 260 376 23 38 382 MUX2_X1
* cell instance $2581 m0 *1 78.66,18.2
X$2581 23 38 FILLCELL_X4
* cell instance $2582 m0 *1 79.42,18.2
X$2582 415 374 23 38 486 NOR2_X1
* cell instance $2583 m0 *1 79.99,18.2
X$2583 376 414 307 23 38 415 MUX2_X1
* cell instance $2584 m0 *1 81.32,18.2
X$2584 23 38 FILLCELL_X4
* cell instance $2585 m0 *1 82.08,18.2
X$2585 23 2668 378 409 445 38 DFF_X1
* cell instance $2586 m0 *1 85.31,18.2
X$2586 23 38 FILLCELL_X8
* cell instance $2587 m0 *1 86.83,18.2
X$2587 23 38 FILLCELL_X1
* cell instance $2588 m0 *1 87.02,18.2
X$2588 23 2581 309 379 310 38 DFF_X1
* cell instance $2589 m0 *1 90.25,18.2
X$2589 23 38 FILLCELL_X8
* cell instance $2590 m0 *1 91.77,18.2
X$2590 23 38 FILLCELL_X4
* cell instance $2591 m0 *1 92.53,18.2
X$2591 23 38 FILLCELL_X2
* cell instance $2592 r0 *1 76.57,18.2
X$2592 452 370 23 38 491 NOR2_X1
* cell instance $2593 r0 *1 77.14,18.2
X$2593 23 38 FILLCELL_X2
* cell instance $2594 r0 *1 77.52,18.2
X$2594 23 38 FILLCELL_X1
* cell instance $2595 r0 *1 77.71,18.2
X$2595 110 372 23 38 443 NOR2_X1
* cell instance $2596 r0 *1 78.28,18.2
X$2596 23 2933 444 487 445 38 DFF_X1
* cell instance $2597 r0 *1 81.51,18.2
X$2597 23 38 FILLCELL_X32
* cell instance $2598 r0 *1 87.59,18.2
X$2598 23 38 FILLCELL_X16
* cell instance $2599 r0 *1 90.63,18.2
X$2599 23 38 FILLCELL_X4
* cell instance $2600 r0 *1 91.39,18.2
X$2600 23 38 FILLCELL_X2
* cell instance $2601 r0 *1 91.77,18.2
X$2601 139 23 38 310 CLKBUF_X3
* cell instance $2602 r0 *1 92.72,18.2
X$2602 310 23 38 CLKBUF_X1
* cell instance $2603 m0 *1 94.24,18.2
X$2603 23 38 FILLCELL_X8
* cell instance $2604 m0 *1 92.91,18.2
X$2604 313 263 336 23 38 410 MUX2_X1
* cell instance $2605 m0 *1 95.76,18.2
X$2605 23 38 FILLCELL_X4
* cell instance $2606 m0 *1 96.52,18.2
X$2606 23 38 FILLCELL_X2
* cell instance $2607 r0 *1 93.29,18.2
X$2607 23 38 FILLCELL_X1
* cell instance $2608 r0 *1 93.48,18.2
X$2608 377 79 480 23 38 481 MUX2_X1
* cell instance $2609 r0 *1 94.81,18.2
X$2609 23 38 FILLCELL_X8
* cell instance $2610 r0 *1 96.33,18.2
X$2610 23 38 FILLCELL_X4
* cell instance $2611 r180 *1 97.28,18.2
X$2611 23 38 23 38 TAPCELL_X1
* cell instance $2612 m0 *1 96.9,18.2
X$2612 23 38 FILLCELL_X1
* cell instance $2613 m90 *1 97.28,18.2
X$2613 23 38 23 38 TAPCELL_X1
* cell instance $2614 r0 *1 45.98,1.4
X$2614 23 38 FILLCELL_X16
* cell instance $2615 r0 *1 49.02,1.4
X$2615 23 38 FILLCELL_X8
* cell instance $2616 r0 *1 50.54,1.4
X$2616 23 38 FILLCELL_X4
* cell instance $2617 r0 *1 51.3,1.4
X$2617 23 38 FILLCELL_X2
* cell instance $2618 r0 *1 19.57,1.4
X$2618 23 38 FILLCELL_X16
* cell instance $2619 r0 *1 22.61,1.4
X$2619 23 38 FILLCELL_X8
* cell instance $2620 r0 *1 24.13,1.4
X$2620 23 38 FILLCELL_X2
* cell instance $2621 m0 *1 1.33,54.6
X$2621 23 38 FILLCELL_X8
* cell instance $2622 m0 *1 1.14,54.6
X$2622 23 38 23 38 TAPCELL_X1
* cell instance $2623 m0 *1 2.85,54.6
X$2623 23 38 FILLCELL_X2
* cell instance $2624 r0 *1 1.14,54.6
X$2624 23 38 23 38 TAPCELL_X1
* cell instance $2625 r0 *1 1.33,54.6
X$2625 23 38 FILLCELL_X8
* cell instance $2626 r0 *1 2.85,54.6
X$2626 23 38 FILLCELL_X4
* cell instance $2627 r0 *1 3.14,54.6
X$2627 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $2628 r0 *1 3.14,54.6
X$2628 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $2629 r0 *1 3.14,54.6
X$2629 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $2630 m0 *1 3.42,54.6
X$2630 1362 1383 1361 23 38 1291 MUX2_X1
* cell instance $2631 m0 *1 3.23,54.6
X$2631 23 38 FILLCELL_X1
* cell instance $2632 m0 *1 4.75,54.6
X$2632 1423 1369 1361 23 38 1345 MUX2_X1
* cell instance $2633 m0 *1 6.08,54.6
X$2633 23 38 FILLCELL_X2
* cell instance $2634 r0 *1 3.61,54.6
X$2634 23 38 FILLCELL_X1
* cell instance $2635 r0 *1 3.8,54.6
X$2635 1397 23 38 1395 BUF_X1
* cell instance $2636 r0 *1 4.37,54.6
X$2636 23 38 FILLCELL_X8
* cell instance $2637 r0 *1 5.89,54.6
X$2637 23 38 FILLCELL_X4
* cell instance $2638 m0 *1 6.65,54.6
X$2638 1362 412 1423 23 38 1424 MUX2_X1
* cell instance $2639 m0 *1 6.46,54.6
X$2639 23 38 FILLCELL_X1
* cell instance $2640 m0 *1 7.98,54.6
X$2640 23 38 FILLCELL_X2
* cell instance $2641 r0 *1 6.65,54.6
X$2641 23 38 FILLCELL_X1
* cell instance $2642 r0 *1 6.84,54.6
X$2642 1325 23 38 1361 BUF_X2
* cell instance $2643 r0 *1 7.6,54.6
X$2643 23 38 FILLCELL_X16
* cell instance $2644 m0 *1 8.55,54.6
X$2644 1325 1406 1327 23 38 1385 MUX2_X1
* cell instance $2645 m0 *1 8.36,54.6
X$2645 23 38 FILLCELL_X1
* cell instance $2646 m0 *1 9.88,54.6
X$2646 23 38 FILLCELL_X4
* cell instance $2647 m0 *1 10.64,54.6
X$2647 23 38 FILLCELL_X1
* cell instance $2648 m0 *1 10.83,54.6
X$2648 1424 354 23 38 1363 NOR2_X1
* cell instance $2649 m0 *1 11.4,54.6
X$2649 23 38 FILLCELL_X4
* cell instance $2650 m0 *1 12.16,54.6
X$2650 23 38 FILLCELL_X1
* cell instance $2651 m0 *1 12.35,54.6
X$2651 1387 1289 1361 23 38 1328 MUX2_X1
* cell instance $2652 m0 *1 13.68,54.6
X$2652 1428 381 23 38 1427 NOR2_X1
* cell instance $2653 m0 *1 14.25,54.6
X$2653 1396 627 1387 23 38 1428 MUX2_X1
* cell instance $2654 m0 *1 15.58,54.6
X$2654 1486 23 38 1326 CLKBUF_X3
* cell instance $2655 m0 *1 16.53,54.6
X$2655 1326 23 38 CLKBUF_X1
* cell instance $2656 m0 *1 17.1,54.6
X$2656 23 38 FILLCELL_X2
* cell instance $2657 r0 *1 10.64,54.6
X$2657 23 38 FILLCELL_X4
* cell instance $2658 r0 *1 11.4,54.6
X$2658 1425 1427 1363 548 1295 1467 23 38 1426 OAI33_X1
* cell instance $2659 r0 *1 12.73,54.6
X$2659 23 38 FILLCELL_X4
* cell instance $2660 r0 *1 13.49,54.6
X$2660 23 38 FILLCELL_X2
* cell instance $2661 r0 *1 13.87,54.6
X$2661 23 38 FILLCELL_X1
* cell instance $2662 r0 *1 14.06,54.6
X$2662 1396 1403 1361 23 38 1430 MUX2_X1
* cell instance $2663 r0 *1 15.39,54.6
X$2663 23 2980 1396 1430 1326 38 DFF_X1
* cell instance $2664 m0 *1 18.05,54.6
X$2664 1158 1364 23 38 1398 NAND2_X1
* cell instance $2665 m0 *1 17.48,54.6
X$2665 1364 1122 23 38 1296 NAND2_X1
* cell instance $2666 m0 *1 18.62,54.6
X$2666 1206 1398 1365 1208 1431 38 23 1389 OAI221_X1
* cell instance $2667 m0 *1 19.76,54.6
X$2667 890 340 1138 1157 1139 38 23 1365 OAI221_X1
* cell instance $2668 m0 *1 20.9,54.6
X$2668 23 2597 1330 1400 1399 38 DFF_X1
* cell instance $2669 m0 *1 24.13,54.6
X$2669 23 38 FILLCELL_X4
* cell instance $2670 m0 *1 24.89,54.6
X$2670 23 38 FILLCELL_X1
* cell instance $2671 m0 *1 25.08,54.6
X$2671 23 2792 1401 1432 1262 38 DFF_X1
* cell instance $2672 m0 *1 28.31,54.6
X$2672 1366 1434 1361 23 38 1436 MUX2_X1
* cell instance $2673 m0 *1 29.64,54.6
X$2673 23 2791 1366 1436 1262 38 DFF_X1
* cell instance $2674 m0 *1 32.87,54.6
X$2674 23 38 FILLCELL_X8
* cell instance $2675 m0 *1 34.39,54.6
X$2675 23 38 FILLCELL_X1
* cell instance $2676 m0 *1 34.58,54.6
X$2676 403 38 381 23 BUF_X4
* cell instance $2677 m0 *1 35.91,54.6
X$2677 23 38 FILLCELL_X1
* cell instance $2678 m0 *1 36.1,54.6
X$2678 1332 1437 1438 1208 1367 38 23 1393 OAI221_X1
* cell instance $2679 m0 *1 37.24,54.6
X$2679 23 2798 1368 1393 1174 38 DFF_X1
* cell instance $2680 m0 *1 40.47,54.6
X$2680 1063 428 1138 1198 1139 38 23 1438 OAI221_X1
* cell instance $2681 m0 *1 41.61,54.6
X$2681 862 38 1358 23 BUF_X4
* cell instance $2682 m0 *1 42.94,54.6
X$2682 634 38 1373 23 BUF_X4
* cell instance $2683 m0 *1 44.27,54.6
X$2683 1268 23 38 1122 CLKBUF_X3
* cell instance $2684 m0 *1 45.22,54.6
X$2684 1065 38 1434 23 BUF_X4
* cell instance $2685 m0 *1 46.55,54.6
X$2685 598 38 1403 23 BUF_X4
* cell instance $2686 m0 *1 47.88,54.6
X$2686 23 38 FILLCELL_X1
* cell instance $2687 m0 *1 48.07,54.6
X$2687 23 2730 1405 1439 1404 38 DFF_X1
* cell instance $2688 m0 *1 51.3,54.6
X$2688 23 38 FILLCELL_X4
* cell instance $2689 m0 *1 52.06,54.6
X$2689 1370 23 38 1299 BUF_X2
* cell instance $2690 m0 *1 52.82,54.6
X$2690 515 38 1425 23 BUF_X4
* cell instance $2691 m0 *1 54.15,54.6
X$2691 23 38 FILLCELL_X2
* cell instance $2692 r0 *1 18.62,54.6
X$2692 23 38 FILLCELL_X4
* cell instance $2693 r0 *1 19.38,54.6
X$2693 23 38 FILLCELL_X1
* cell instance $2694 r0 *1 19.57,54.6
X$2694 23 2978 1364 1389 1399 38 DFF_X1
* cell instance $2695 r0 *1 22.8,54.6
X$2695 1364 1140 23 38 1431 NAND2_X1
* cell instance $2696 r0 *1 23.37,54.6
X$2696 23 38 FILLCELL_X8
* cell instance $2697 r0 *1 24.89,54.6
X$2697 23 38 FILLCELL_X4
* cell instance $2698 r0 *1 25.65,54.6
X$2698 1401 1446 1361 23 38 1432 MUX2_X1
* cell instance $2699 r0 *1 26.98,54.6
X$2699 23 38 FILLCELL_X1
* cell instance $2700 r0 *1 27.17,54.6
X$2700 1401 1184 1366 23 38 1447 MUX2_X1
* cell instance $2701 r0 *1 28.5,54.6
X$2701 23 38 FILLCELL_X2
* cell instance $2702 r0 *1 28.88,54.6
X$2702 1402 1213 1474 38 23 1397 OAI21_X4
* cell instance $2703 r0 *1 31.35,54.6
X$2703 1450 1122 23 38 1474 NAND2_X1
* cell instance $2704 r0 *1 31.92,54.6
X$2704 23 38 FILLCELL_X4
* cell instance $2705 r0 *1 32.68,54.6
X$2705 23 38 FILLCELL_X1
* cell instance $2706 r0 *1 32.87,54.6
X$2706 23 3006 1452 1453 1174 38 DFF_X1
* cell instance $2707 r0 *1 36.1,54.6
X$2707 1368 1140 23 38 1367 NAND2_X1
* cell instance $2708 r0 *1 36.67,54.6
X$2708 1198 23 38 1137 CLKBUF_X3
* cell instance $2709 r0 *1 37.62,54.6
X$2709 1486 23 38 1174 CLKBUF_X3
* cell instance $2710 r0 *1 38.57,54.6
X$2710 620 38 792 23 BUF_X4
* cell instance $2711 r0 *1 39.9,54.6
X$2711 23 38 FILLCELL_X2
* cell instance $2712 r0 *1 40.28,54.6
X$2712 23 1331 1210 38 BUF_X32
* cell instance $2713 r0 *1 49.59,54.6
X$2713 23 2887 1455 1477 1404 38 DFF_X1
* cell instance $2714 r0 *1 52.82,54.6
X$2714 1405 188 1455 23 38 1591 MUX2_X1
* cell instance $2715 r0 *1 54.15,54.6
X$2715 286 38 1406 23 BUF_X4
* cell instance $2716 m0 *1 54.72,54.6
X$2716 23 2564 1333 1440 1301 38 DFF_X1
* cell instance $2717 m0 *1 54.53,54.6
X$2717 23 38 FILLCELL_X1
* cell instance $2718 m0 *1 57.95,54.6
X$2718 23 38 FILLCELL_X8
* cell instance $2719 m0 *1 59.47,54.6
X$2719 23 38 FILLCELL_X2
* cell instance $2720 r0 *1 55.48,54.6
X$2720 1478 23 38 1158 CLKBUF_X3
* cell instance $2721 r0 *1 56.43,54.6
X$2721 23 38 FILLCELL_X1
* cell instance $2722 r0 *1 56.62,54.6
X$2722 1519 23 38 1140 CLKBUF_X3
* cell instance $2723 r0 *1 57.57,54.6
X$2723 1407 38 881 23 BUF_X4
* cell instance $2724 r0 *1 58.9,54.6
X$2724 1408 23 38 1130 BUF_X2
* cell instance $2725 r0 *1 59.14,54.6
X$2725 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $2726 r0 *1 59.14,54.6
X$2726 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $2727 r0 *1 59.14,54.6
X$2727 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $2728 r0 *1 59.66,54.6
X$2728 1456 1442 38 23 1409 AND2_X1
* cell instance $2729 m0 *1 60.61,54.6
X$2729 1175 38 441 23 BUF_X4
* cell instance $2730 m0 *1 59.85,54.6
X$2730 1409 23 38 598 BUF_X2
* cell instance $2731 m0 *1 61.94,54.6
X$2731 1411 1444 38 23 1443 AND2_X1
* cell instance $2732 m0 *1 62.7,54.6
X$2732 1443 23 38 557 CLKBUF_X3
* cell instance $2733 m0 *1 63.65,54.6
X$2733 23 38 FILLCELL_X1
* cell instance $2734 m0 *1 63.84,54.6
X$2734 1411 1442 38 23 1441 AND2_X1
* cell instance $2735 m0 *1 64.6,54.6
X$2735 1441 23 38 597 CLKBUF_X3
* cell instance $2736 m0 *1 65.55,54.6
X$2736 597 38 88 23 BUF_X4
* cell instance $2737 m0 *1 66.88,54.6
X$2737 1301 23 38 CLKBUF_X1
* cell instance $2738 m0 *1 67.45,54.6
X$2738 23 38 FILLCELL_X8
* cell instance $2739 m0 *1 68.97,54.6
X$2739 23 38 FILLCELL_X2
* cell instance $2740 r0 *1 60.42,54.6
X$2740 1410 23 38 1065 BUF_X2
* cell instance $2741 r0 *1 61.18,54.6
X$2741 1457 1411 23 286 38 NAND2_X4
* cell instance $2742 r0 *1 62.89,54.6
X$2742 1412 23 38 599 BUF_X2
* cell instance $2743 r0 *1 63.65,54.6
X$2743 557 38 130 23 BUF_X4
* cell instance $2744 r0 *1 66.31,54.6
X$2744 1335 133 1413 23 38 1476 MUX2_X1
* cell instance $2745 r0 *1 67.64,54.6
X$2745 1392 23 38 1301 CLKBUF_X3
* cell instance $2746 r0 *1 68.59,54.6
X$2746 23 38 FILLCELL_X4
* cell instance $2747 m0 *1 69.54,54.6
X$2747 1335 79 1372 23 38 1414 MUX2_X1
* cell instance $2748 m0 *1 69.35,54.6
X$2748 23 38 FILLCELL_X1
* cell instance $2749 m0 *1 70.87,54.6
X$2749 23 38 FILLCELL_X8
* cell instance $2750 m0 *1 72.39,54.6
X$2750 23 38 FILLCELL_X4
* cell instance $2751 m0 *1 73.15,54.6
X$2751 23 38 FILLCELL_X2
* cell instance $2752 r0 *1 69.35,54.6
X$2752 23 38 FILLCELL_X1
* cell instance $2753 r0 *1 69.54,54.6
X$2753 23 2917 1372 1414 1301 38 DFF_X1
* cell instance $2754 r0 *1 72.77,54.6
X$2754 23 38 FILLCELL_X2
* cell instance $2755 r0 *1 73.15,54.6
X$2755 23 38 FILLCELL_X1
* cell instance $2756 r0 *1 73.34,54.6
X$2756 23 3107 1374 1475 1336 38 DFF_X1
* cell instance $2757 m0 *1 73.72,54.6
X$2757 881 38 177 23 BUF_X4
* cell instance $2758 m0 *1 73.53,54.6
X$2758 23 38 FILLCELL_X1
* cell instance $2759 m0 *1 75.05,54.6
X$2759 23 38 FILLCELL_X8
* cell instance $2760 m0 *1 76.57,54.6
X$2760 23 38 FILLCELL_X2
* cell instance $2761 r0 *1 76.57,54.6
X$2761 1073 133 1374 23 38 1475 MUX2_X1
* cell instance $2762 m0 *1 78.28,54.6
X$2762 23 38 FILLCELL_X1
* cell instance $2763 m0 *1 76.95,54.6
X$2763 1374 1373 1337 23 38 1524 MUX2_X1
* cell instance $2764 m0 *1 78.47,54.6
X$2764 23 2678 1416 1390 1223 38 DFF_X1
* cell instance $2765 m0 *1 81.7,54.6
X$2765 23 38 FILLCELL_X1
* cell instance $2766 m0 *1 81.89,54.6
X$2766 1332 1415 1376 1319 1417 38 23 1390 OAI221_X1
* cell instance $2767 m0 *1 83.03,54.6
X$2767 1223 23 38 CLKBUF_X1
* cell instance $2768 m0 *1 83.6,54.6
X$2768 1416 1268 23 38 1303 NAND2_X1
* cell instance $2769 m0 *1 84.17,54.6
X$2769 23 38 FILLCELL_X1
* cell instance $2770 m0 *1 84.36,54.6
X$2770 841 1088 1304 1305 38 23 1388 OAI22_X1
* cell instance $2771 m0 *1 85.31,54.6
X$2771 1088 841 1241 1300 1240 38 23 1418 OAI221_X1
* cell instance $2772 m0 *1 86.45,54.6
X$2772 23 38 FILLCELL_X8
* cell instance $2773 m0 *1 87.97,54.6
X$2773 23 38 FILLCELL_X4
* cell instance $2774 m0 *1 88.73,54.6
X$2774 23 38 FILLCELL_X1
* cell instance $2775 m0 *1 88.92,54.6
X$2775 1306 1435 1388 38 1386 23 OAI21_X1
* cell instance $2776 m0 *1 89.68,54.6
X$2776 23 38 FILLCELL_X4
* cell instance $2777 m0 *1 90.44,54.6
X$2777 23 38 FILLCELL_X1
* cell instance $2778 m0 *1 90.63,54.6
X$2778 1225 1433 1379 1226 1429 38 23 1378 OAI221_X1
* cell instance $2779 m0 *1 91.77,54.6
X$2779 1228 1420 23 38 1433 NAND2_X1
* cell instance $2780 m0 *1 92.34,54.6
X$2780 1420 1239 23 38 1429 NAND2_X1
* cell instance $2781 m0 *1 92.91,54.6
X$2781 1420 1230 23 38 1380 NAND2_X1
* cell instance $2782 m0 *1 93.48,54.6
X$2782 23 38 FILLCELL_X2
* cell instance $2783 r0 *1 77.9,54.6
X$2783 23 38 FILLCELL_X4
* cell instance $2784 r0 *1 78.66,54.6
X$2784 23 38 FILLCELL_X1
* cell instance $2785 r0 *1 78.85,54.6
X$2785 23 2877 1377 1473 1223 38 DFF_X1
* cell instance $2786 r0 *1 82.08,54.6
X$2786 1460 1416 23 38 1415 NAND2_X1
* cell instance $2787 r0 *1 82.65,54.6
X$2787 23 38 FILLCELL_X1
* cell instance $2788 r0 *1 82.84,54.6
X$2788 1416 1519 23 38 1417 NAND2_X1
* cell instance $2789 r0 *1 83.41,54.6
X$2789 23 38 FILLCELL_X8
* cell instance $2790 r0 *1 84.93,54.6
X$2790 23 38 FILLCELL_X1
* cell instance $2791 r0 *1 85.12,54.6
X$2791 1391 177 23 38 1515 NOR2_X1
* cell instance $2792 r0 *1 85.69,54.6
X$2792 23 2867 1419 1472 1223 38 DFF_X1
* cell instance $2793 r0 *1 88.92,54.6
X$2793 1419 1230 23 38 1435 NAND2_X1
* cell instance $2794 r0 *1 89.49,54.6
X$2794 23 38 FILLCELL_X1
* cell instance $2795 r0 *1 89.68,54.6
X$2795 23 3035 1420 1378 1227 38 DFF_X1
* cell instance $2796 r0 *1 92.91,54.6
X$2796 23 38 FILLCELL_X1
* cell instance $2797 r0 *1 93.1,54.6
X$2797 1154 914 1304 1305 38 23 1463 OAI22_X1
* cell instance $2798 m0 *1 94.43,54.6
X$2798 1381 23 38 1073 CLKBUF_X2
* cell instance $2799 m0 *1 93.86,54.6
X$2799 1386 23 38 1422 BUF_X1
* cell instance $2800 m0 *1 95.19,54.6
X$2800 1347 23 38 1382 BUF_X1
* cell instance $2801 m0 *1 95.76,54.6
X$2801 23 38 FILLCELL_X1
* cell instance $2802 m0 *1 95.95,54.6
X$2802 1384 23 38 1342 BUF_X1
* cell instance $2803 m0 *1 96.52,54.6
X$2803 1304 23 38 1421 BUF_X1
* cell instance $2804 r180 *1 97.28,54.6
X$2804 23 38 23 38 TAPCELL_X1
* cell instance $2805 r0 *1 94.05,54.6
X$2805 23 38 FILLCELL_X4
* cell instance $2806 r0 *1 94.81,54.6
X$2806 23 38 FILLCELL_X2
* cell instance $2807 r0 *1 95.19,54.6
X$2807 1470 23 38 1464 BUF_X1
* cell instance $2808 r0 *1 95.76,54.6
X$2808 23 38 FILLCELL_X4
* cell instance $2809 r0 *1 96.52,54.6
X$2809 23 38 FILLCELL_X2
* cell instance $2810 r0 *1 96.9,54.6
X$2810 23 38 FILLCELL_X1
* cell instance $2811 m90 *1 97.28,54.6
X$2811 23 38 23 38 TAPCELL_X1
* cell instance $2812 m0 *1 1.33,63
X$2812 23 38 FILLCELL_X8
* cell instance $2813 m0 *1 1.14,63
X$2813 23 38 23 38 TAPCELL_X1
* cell instance $2814 m0 *1 2.85,63
X$2814 23 38 FILLCELL_X4
* cell instance $2815 m0 *1 3.61,63
X$2815 23 38 FILLCELL_X2
* cell instance $2816 r0 *1 1.14,63
X$2816 23 38 23 38 TAPCELL_X1
* cell instance $2817 r0 *1 1.33,63
X$2817 23 38 FILLCELL_X8
* cell instance $2818 r0 *1 2.85,63
X$2818 23 38 FILLCELL_X2
* cell instance $2819 r0 *1 3.14,63
X$2819 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $2820 r0 *1 3.14,63
X$2820 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $2821 r0 *1 3.14,63.4
X$2821 23 VIA_via4_5_960_2800_5_2_600_600
* cell instance $2822 r0 *1 3.14,63
X$2822 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $2823 r0 *1 3.14,63.4
X$2823 23 VIA_via5_6_960_2800_5_2_600_600
* cell instance $2824 r0 *1 3.14,63.4
X$2824 23 VIA_via6_7_960_2800_4_1_600_600
* cell instance $2825 r0 *1 3.23,63
X$2825 1598 1406 1689 23 38 1710 MUX2_X1
* cell instance $2826 m0 *1 5.32,63
X$2826 1598 1480 1633 23 38 1655 MUX2_X1
* cell instance $2827 m0 *1 3.99,63
X$2827 1598 1493 1654 23 38 1614 MUX2_X1
* cell instance $2828 m0 *1 6.65,63
X$2828 23 38 FILLCELL_X2
* cell instance $2829 r0 *1 4.56,63
X$2829 23 38 FILLCELL_X2
* cell instance $2830 r0 *1 4.94,63
X$2830 23 2998 1633 1655 1556 38 DFF_X1
* cell instance $2831 m0 *1 8.36,63
X$2831 23 38 FILLCELL_X1
* cell instance $2832 m0 *1 7.03,63
X$2832 1654 70 1633 23 38 1617 MUX2_X1
* cell instance $2833 m0 *1 8.55,63
X$2833 1598 23 38 1532 BUF_X2
* cell instance $2834 m0 *1 9.31,63
X$2834 23 38 FILLCELL_X2
* cell instance $2835 r0 *1 8.17,63
X$2835 23 38 FILLCELL_X8
* cell instance $2836 m0 *1 9.88,63
X$2836 1532 1544 1599 23 38 1618 MUX2_X1
* cell instance $2837 m0 *1 9.69,63
X$2837 23 38 FILLCELL_X1
* cell instance $2838 m0 *1 11.21,63
X$2838 1598 1482 1659 23 38 1634 MUX2_X1
* cell instance $2839 m0 *1 12.54,63
X$2839 23 38 FILLCELL_X4
* cell instance $2840 m0 *1 13.3,63
X$2840 23 38 FILLCELL_X1
* cell instance $2841 m0 *1 13.49,63
X$2841 1599 813 1659 23 38 1623 MUX2_X1
* cell instance $2842 m0 *1 14.82,63
X$2842 23 38 FILLCELL_X2
* cell instance $2843 r0 *1 9.69,63
X$2843 23 38 FILLCELL_X4
* cell instance $2844 r0 *1 10.45,63
X$2844 23 38 FILLCELL_X1
* cell instance $2845 r0 *1 10.64,63
X$2845 1617 1483 23 38 1690 NOR2_X1
* cell instance $2846 r0 *1 11.21,63
X$2846 23 2942 1659 1634 1635 38 DFF_X1
* cell instance $2847 r0 *1 14.44,63
X$2847 23 38 FILLCELL_X8
* cell instance $2848 m0 *1 15.39,63
X$2848 23 2576 1661 1660 1399 38 DFF_X1
* cell instance $2849 m0 *1 15.2,63
X$2849 23 38 FILLCELL_X1
* cell instance $2850 m0 *1 18.62,63
X$2850 1600 1434 1532 23 38 1622 MUX2_X1
* cell instance $2851 m0 *1 19.95,63
X$2851 1662 893 23 38 1663 NOR2_X1
* cell instance $2852 m0 *1 20.52,63
X$2852 1623 831 23 38 1664 NOR2_X1
* cell instance $2853 m0 *1 21.09,63
X$2853 1485 1626 1663 1142 1664 1625 23 38 1726 OAI33_X1
* cell instance $2854 m0 *1 22.42,63
X$2854 23 38 FILLCELL_X2
* cell instance $2855 r0 *1 15.96,63
X$2855 23 38 FILLCELL_X2
* cell instance $2856 r0 *1 16.34,63
X$2856 1661 1446 1532 23 38 1660 MUX2_X1
* cell instance $2857 r0 *1 17.67,63
X$2857 23 38 FILLCELL_X2
* cell instance $2858 r0 *1 18.05,63
X$2858 23 38 FILLCELL_X1
* cell instance $2859 r0 *1 18.24,63
X$2859 1661 1184 1600 23 38 1662 MUX2_X1
* cell instance $2860 r0 *1 19.57,63
X$2860 23 38 FILLCELL_X2
* cell instance $2861 r0 *1 19.95,63
X$2861 23 2953 1601 1665 1693 38 DFF_X1
* cell instance $2862 m0 *1 24.13,63
X$2862 23 38 FILLCELL_X16
* cell instance $2863 m0 *1 22.8,63
X$2863 1601 1487 1532 23 38 1665 MUX2_X1
* cell instance $2864 m0 *1 27.17,63
X$2864 23 38 FILLCELL_X8
* cell instance $2865 m0 *1 28.69,63
X$2865 23 38 FILLCELL_X2
* cell instance $2866 r0 *1 23.18,63
X$2866 1666 1488 1532 23 38 1716 MUX2_X1
* cell instance $2867 r0 *1 24.51,63
X$2867 23 38 FILLCELL_X32
* cell instance $2868 m0 *1 29.64,63
X$2868 1206 1602 1604 1208 1630 38 23 1603 OAI221_X1
* cell instance $2869 m0 *1 29.07,63
X$2869 1636 1450 23 38 1602 NAND2_X1
* cell instance $2870 m0 *1 30.78,63
X$2870 1450 1638 23 38 1630 NAND2_X1
* cell instance $2871 m0 *1 31.35,63
X$2871 988 38 354 23 BUF_X4
* cell instance $2872 m0 *1 32.68,63
X$2872 23 38 FILLCELL_X16
* cell instance $2873 m0 *1 35.72,63
X$2873 23 38 FILLCELL_X1
* cell instance $2874 m0 *1 35.91,63
X$2874 988 38 1650 23 BUF_X4
* cell instance $2875 m0 *1 37.24,63
X$2875 23 38 FILLCELL_X4
* cell instance $2876 m0 *1 38,63
X$2876 23 38 FILLCELL_X2
* cell instance $2877 r0 *1 30.59,63
X$2877 23 38 FILLCELL_X2
* cell instance $2878 r0 *1 30.97,63
X$2878 1206 1667 1695 1208 1668 38 23 1696 OAI221_X1
* cell instance $2879 r0 *1 32.11,63
X$2879 1636 1637 23 38 1667 NAND2_X1
* cell instance $2880 r0 *1 32.68,63
X$2880 23 38 FILLCELL_X2
* cell instance $2881 r0 *1 33.06,63
X$2881 1637 1638 23 38 1668 NAND2_X1
* cell instance $2882 r0 *1 33.63,63
X$2882 23 38 FILLCELL_X32
* cell instance $2883 m0 *1 38.57,63
X$2883 988 38 1605 23 BUF_X4
* cell instance $2884 m0 *1 38.38,63
X$2884 23 38 FILLCELL_X1
* cell instance $2885 m0 *1 39.9,63
X$2885 23 38 FILLCELL_X4
* cell instance $2886 m0 *1 40.66,63
X$2886 23 38 FILLCELL_X1
* cell instance $2887 m0 *1 40.85,63
X$2887 1671 1369 1490 23 38 1670 MUX2_X1
* cell instance $2888 m0 *1 42.18,63
X$2888 23 38 FILLCELL_X4
* cell instance $2889 m0 *1 42.94,63
X$2889 1557 724 1671 23 38 1673 MUX2_X1
* cell instance $2890 m0 *1 44.27,63
X$2890 23 38 FILLCELL_X2
* cell instance $2891 r0 *1 39.71,63
X$2891 23 38 FILLCELL_X4
* cell instance $2892 r0 *1 40.47,63
X$2892 23 38 FILLCELL_X1
* cell instance $2893 r0 *1 40.66,63
X$2893 23 2986 1671 1670 1404 38 DFF_X1
* cell instance $2894 r0 *1 43.89,63
X$2894 23 38 FILLCELL_X8
* cell instance $2895 m0 *1 47.88,63
X$2895 1558 1099 1640 23 38 1676 MUX2_X1
* cell instance $2896 m0 *1 44.65,63
X$2896 23 2819 1558 1632 1404 38 DFF_X1
* cell instance $2897 m0 *1 49.21,63
X$2897 23 38 FILLCELL_X1
* cell instance $2898 m0 *1 49.4,63
X$2898 23 2600 1559 1631 1735 38 DFF_X1
* cell instance $2899 m0 *1 52.63,63
X$2899 1676 1605 23 38 1628 NOR2_X1
* cell instance $2900 m0 *1 53.2,63
X$2900 23 38 FILLCELL_X4
* cell instance $2901 m0 *1 53.96,63
X$2901 23 38 FILLCELL_X1
* cell instance $2902 m0 *1 54.15,63
X$2902 1591 1579 23 38 1679 NOR2_X1
* cell instance $2903 m0 *1 54.72,63
X$2903 23 38 FILLCELL_X4
* cell instance $2904 m0 *1 55.48,63
X$2904 23 38 FILLCELL_X1
* cell instance $2905 m0 *1 55.67,63
X$2905 23 2599 1606 1682 1735 38 DFF_X1
* cell instance $2906 m0 *1 58.9,63
X$2906 23 38 FILLCELL_X8
* cell instance $2907 m0 *1 60.42,63
X$2907 23 38 FILLCELL_X2
* cell instance $2908 r0 *1 45.41,63
X$2908 23 2990 1640 1675 1639 38 DFF_X1
* cell instance $2909 r0 *1 48.64,63
X$2909 1587 1482 1640 23 38 1675 MUX2_X1
* cell instance $2910 r0 *1 49.97,63
X$2910 23 38 FILLCELL_X8
* cell instance $2911 r0 *1 51.49,63
X$2911 23 38 FILLCELL_X4
* cell instance $2912 r0 *1 52.25,63
X$2912 1587 1406 1677 23 38 1760 MUX2_X1
* cell instance $2913 r0 *1 53.58,63
X$2913 1673 1650 23 38 1761 NOR2_X1
* cell instance $2914 r0 *1 54.15,63
X$2914 23 38 FILLCELL_X1
* cell instance $2915 r0 *1 54.34,63
X$2915 1677 1358 1606 23 38 1680 MUX2_X1
* cell instance $2916 r0 *1 55.67,63
X$2916 1680 1535 23 38 1699 NOR2_X1
* cell instance $2917 r0 *1 56.24,63
X$2917 23 38 FILLCELL_X2
* cell instance $2918 r0 *1 56.62,63
X$2918 23 38 FILLCELL_X1
* cell instance $2919 r0 *1 56.81,63
X$2919 23 2874 1702 1642 1684 38 DFF_X1
* cell instance $2920 r0 *1 59.14,63
X$2920 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $2921 r0 *1 59.14,63
X$2921 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $2922 r0 *1 59.14,63.4
X$2922 23 VIA_via4_5_960_2800_5_2_600_600
* cell instance $2923 r0 *1 59.14,63
X$2923 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $2924 r0 *1 59.14,63.4
X$2924 23 VIA_via5_6_960_2800_5_2_600_600
* cell instance $2925 r0 *1 59.14,63.4
X$2925 23 VIA_via6_7_960_2800_4_1_600_600
* cell instance $2926 r0 *1 60.04,63
X$2926 23 38 FILLCELL_X8
* cell instance $2927 m0 *1 64.03,63
X$2927 1643 188 1608 23 38 1687 MUX2_X1
* cell instance $2928 m0 *1 60.8,63
X$2928 23 2583 1643 1607 1684 38 DFF_X1
* cell instance $2929 m0 *1 65.36,63
X$2929 1686 23 38 1139 CLKBUF_X3
* cell instance $2930 m0 *1 66.31,63
X$2930 1687 1579 23 38 1627 NOR2_X1
* cell instance $2931 m0 *1 66.88,63
X$2931 1704 724 1645 23 38 1646 MUX2_X1
* cell instance $2932 m0 *1 68.21,63
X$2932 23 38 FILLCELL_X2
* cell instance $2933 r0 *1 61.56,63
X$2933 23 38 FILLCELL_X2
* cell instance $2934 r0 *1 61.94,63
X$2934 1643 223 1561 23 38 1607 MUX2_X1
* cell instance $2935 r0 *1 63.27,63
X$2935 23 2855 1645 1685 1644 38 DFF_X1
* cell instance $2936 r0 *1 66.5,63
X$2936 1645 130 1561 23 38 1685 MUX2_X1
* cell instance $2937 r0 *1 67.83,63
X$2937 23 38 FILLCELL_X2
* cell instance $2938 r0 *1 68.21,63
X$2938 1646 1650 23 38 1593 NOR2_X1
* cell instance $2939 m0 *1 71.82,63
X$2939 23 38 FILLCELL_X4
* cell instance $2940 m0 *1 68.59,63
X$2940 23 2604 1564 1624 1644 38 DFF_X1
* cell instance $2941 m0 *1 72.58,63
X$2941 23 38 FILLCELL_X2
* cell instance $2942 r0 *1 68.78,63
X$2942 23 38 FILLCELL_X16
* cell instance $2943 r0 *1 71.82,63
X$2943 23 38 FILLCELL_X2
* cell instance $2944 r0 *1 72.2,63
X$2944 23 3110 1647 1609 1336 38 DFF_X1
* cell instance $2945 m0 *1 73.15,63
X$2945 1647 441 1497 23 38 1609 MUX2_X1
* cell instance $2946 m0 *1 72.96,63
X$2946 23 38 FILLCELL_X1
* cell instance $2947 m0 *1 74.48,63
X$2947 1647 1454 1610 23 38 1683 MUX2_X1
* cell instance $2948 m0 *1 75.81,63
X$2948 23 38 FILLCELL_X1
* cell instance $2949 m0 *1 76,63
X$2949 1683 1105 23 38 1681 NOR2_X1
* cell instance $2950 m0 *1 76.57,63
X$2950 23 38 FILLCELL_X4
* cell instance $2951 m0 *1 77.33,63
X$2951 23 38 FILLCELL_X2
* cell instance $2952 r0 *1 75.43,63
X$2952 1610 373 1497 23 38 1715 MUX2_X1
* cell instance $2953 r0 *1 76.76,63
X$2953 23 38 FILLCELL_X8
* cell instance $2954 m0 *1 79.04,63
X$2954 1611 414 1540 23 38 1620 MUX2_X1
* cell instance $2955 m0 *1 77.71,63
X$2955 475 1681 1621 476 1539 1678 23 38 1615 OAI33_X1
* cell instance $2956 m0 *1 80.37,63
X$2956 23 38 FILLCELL_X4
* cell instance $2957 m0 *1 81.13,63
X$2957 23 38 FILLCELL_X2
* cell instance $2958 r0 *1 78.28,63
X$2958 23 38 FILLCELL_X2
* cell instance $2959 r0 *1 78.66,63
X$2959 1497 260 1611 23 38 1753 MUX2_X1
* cell instance $2960 r0 *1 79.99,63
X$2960 23 38 FILLCELL_X8
* cell instance $2961 r0 *1 81.51,63
X$2961 23 38 FILLCELL_X2
* cell instance $2962 m0 *1 84.74,63
X$2962 1586 724 1649 23 38 1674 MUX2_X1
* cell instance $2963 m0 *1 81.51,63
X$2963 23 2679 1586 1619 1714 38 DFF_X1
* cell instance $2964 m0 *1 86.07,63
X$2964 1674 1650 23 38 1578 NOR2_X1
* cell instance $2965 m0 *1 86.64,63
X$2965 23 38 FILLCELL_X1
* cell instance $2966 m0 *1 86.83,63
X$2966 1577 188 1582 23 38 1669 MUX2_X1
* cell instance $2967 m0 *1 88.16,63
X$2967 1669 1579 23 38 1616 NOR2_X1
* cell instance $2968 m0 *1 88.73,63
X$2968 227 1651 1713 225 1153 1515 23 38 1652 OAI33_X1
* cell instance $2969 m0 *1 90.06,63
X$2969 23 1225 38 1331 BUF_X8
* cell instance $2970 m0 *1 92.53,63
X$2970 23 38 FILLCELL_X2
* cell instance $2971 r0 *1 81.89,63
X$2971 23 38 FILLCELL_X1
* cell instance $2972 r0 *1 82.08,63
X$2972 23 2881 1649 1672 1648 38 DFF_X1
* cell instance $2973 r0 *1 85.31,63
X$2973 1649 130 1497 23 38 1672 MUX2_X1
* cell instance $2974 r0 *1 86.64,63
X$2974 23 38 FILLCELL_X8
* cell instance $2975 r0 *1 88.16,63
X$2975 23 38 FILLCELL_X4
* cell instance $2976 r0 *1 88.92,63
X$2976 23 38 FILLCELL_X2
* cell instance $2977 r0 *1 89.3,63
X$2977 1706 1652 1304 1305 38 23 1656 OAI22_X1
* cell instance $2978 r0 *1 90.25,63
X$2978 1686 23 38 1224 BUF_X2
* cell instance $2979 r0 *1 91.01,63
X$2979 23 38 FILLCELL_X4
* cell instance $2980 r0 *1 91.77,63
X$2980 1615 1566 1241 1506 1224 38 23 1707 OAI221_X1
* cell instance $2981 r0 *1 92.91,63
X$2981 23 38 FILLCELL_X8
* cell instance $2982 m0 *1 93.1,63
X$2982 1615 1566 1304 1305 38 23 1658 OAI22_X1
* cell instance $2983 m0 *1 92.91,63
X$2983 23 38 FILLCELL_X1
* cell instance $2984 m0 *1 94.05,63
X$2984 23 38 FILLCELL_X8
* cell instance $2985 m0 *1 95.57,63
X$2985 1306 1612 1658 38 1613 23 OAI21_X1
* cell instance $2986 m0 *1 96.33,63
X$2986 1613 23 38 1569 BUF_X1
* cell instance $2987 m0 *1 96.9,63
X$2987 23 38 FILLCELL_X1
* cell instance $2988 r180 *1 97.28,63
X$2988 23 38 23 38 TAPCELL_X1
* cell instance $2989 r0 *1 94.43,63
X$2989 23 38 FILLCELL_X2
* cell instance $2990 r0 *1 94.81,63
X$2990 1306 1708 1656 38 1657 23 OAI21_X1
* cell instance $2991 r0 *1 95.57,63
X$2991 23 38 FILLCELL_X4
* cell instance $2992 r0 *1 96.33,63
X$2992 23 38 FILLCELL_X1
* cell instance $2993 r0 *1 96.52,63
X$2993 1657 23 38 1653 BUF_X1
* cell instance $2994 m90 *1 97.28,63
X$2994 23 38 23 38 TAPCELL_X1
* cell instance $2995 m0 *1 26.22,43.4
X$2995 23 38 FILLCELL_X8
* cell instance $2996 m0 *1 24.89,43.4
X$2996 1031 994 1045 23 38 936 MUX2_X1
* cell instance $2997 m0 *1 27.74,43.4
X$2997 1059 992 421 23 38 1080 MUX2_X1
* cell instance $2998 m0 *1 29.07,43.4
X$2998 23 38 FILLCELL_X1
* cell instance $2999 m0 *1 29.26,43.4
X$2999 1032 941 421 23 38 1081 MUX2_X1
* cell instance $3000 m0 *1 30.59,43.4
X$3000 1032 994 1059 23 38 1050 MUX2_X1
* cell instance $3001 m0 *1 31.92,43.4
X$3001 1050 881 23 38 1022 NOR2_X1
* cell instance $3002 m0 *1 32.49,43.4
X$3002 23 38 FILLCELL_X1
* cell instance $3003 m0 *1 32.68,43.4
X$3003 693 23 38 942 CLKBUF_X3
* cell instance $3004 m0 *1 33.63,43.4
X$3004 942 23 38 CLKBUF_X1
* cell instance $3005 m0 *1 34.2,43.4
X$3005 23 38 FILLCELL_X8
* cell instance $3006 m0 *1 35.72,43.4
X$3006 23 38 FILLCELL_X4
* cell instance $3007 m0 *1 36.48,43.4
X$3007 1083 900 1124 23 38 1052 MUX2_X1
* cell instance $3008 m0 *1 37.81,43.4
X$3008 23 38 FILLCELL_X1
* cell instance $3009 m0 *1 38,43.4
X$3009 1052 840 23 38 1061 NOR2_X1
* cell instance $3010 m0 *1 38.57,43.4
X$3010 23 38 FILLCELL_X1
* cell instance $3011 m0 *1 38.76,43.4
X$3011 1053 831 23 38 1033 NOR2_X1
* cell instance $3012 m0 *1 39.33,43.4
X$3012 23 38 FILLCELL_X8
* cell instance $3013 m0 *1 40.85,43.4
X$3013 23 38 FILLCELL_X4
* cell instance $3014 m0 *1 41.61,43.4
X$3014 23 38 FILLCELL_X1
* cell instance $3015 m0 *1 41.8,43.4
X$3015 23 2720 999 1034 1035 38 DFF_X1
* cell instance $3016 m0 *1 45.03,43.4
X$3016 23 2711 1036 1064 1035 38 DFF_X1
* cell instance $3017 m0 *1 48.26,43.4
X$3017 1055 941 301 23 38 1037 MUX2_X1
* cell instance $3018 m0 *1 49.59,43.4
X$3018 1055 862 1036 23 38 1054 MUX2_X1
* cell instance $3019 m0 *1 50.92,43.4
X$3019 1054 881 23 38 902 NOR2_X1
* cell instance $3020 m0 *1 51.49,43.4
X$3020 23 38 FILLCELL_X16
* cell instance $3021 m0 *1 54.53,43.4
X$3021 23 38 FILLCELL_X4
* cell instance $3022 m0 *1 55.29,43.4
X$3022 23 38 FILLCELL_X1
* cell instance $3023 m0 *1 55.48,43.4
X$3023 864 23 38 891 CLKBUF_X3
* cell instance $3024 m0 *1 56.43,43.4
X$3024 23 38 FILLCELL_X2
* cell instance $3025 m0 *1 21.09,43.4
X$3025 1031 941 358 23 38 1029 MUX2_X1
* cell instance $3026 m0 *1 20.9,43.4
X$3026 23 38 FILLCELL_X1
* cell instance $3027 m0 *1 22.42,43.4
X$3027 1045 992 358 23 38 1030 MUX2_X1
* cell instance $3028 m0 *1 23.75,43.4
X$3028 23 38 FILLCELL_X4
* cell instance $3029 m0 *1 24.51,43.4
X$3029 23 38 FILLCELL_X2
* cell instance $3030 r0 *1 20.9,43.4
X$3030 23 38 FILLCELL_X1
* cell instance $3031 r0 *1 21.09,43.4
X$3031 693 23 38 991 CLKBUF_X3
* cell instance $3032 r0 *1 22.04,43.4
X$3032 991 23 38 3146 INV_X1
* cell instance $3033 r0 *1 22.42,43.4
X$3033 23 38 FILLCELL_X2
* cell instance $3034 r0 *1 22.8,43.4
X$3034 23 38 FILLCELL_X1
* cell instance $3035 r0 *1 22.99,43.4
X$3035 23 2995 1045 1030 991 38 DFF_X1
* cell instance $3036 r0 *1 26.22,43.4
X$3036 23 2956 1059 1080 942 38 DFF_X1
* cell instance $3037 r0 *1 29.45,43.4
X$3037 23 38 FILLCELL_X1
* cell instance $3038 r0 *1 29.64,43.4
X$3038 23 2958 1032 1081 942 38 DFF_X1
* cell instance $3039 r0 *1 32.87,43.4
X$3039 23 38 FILLCELL_X8
* cell instance $3040 r0 *1 34.39,43.4
X$3040 23 38 FILLCELL_X2
* cell instance $3041 r0 *1 34.77,43.4
X$3041 23 38 FILLCELL_X1
* cell instance $3042 r0 *1 34.96,43.4
X$3042 23 2966 1083 1060 942 38 DFF_X1
* cell instance $3043 r0 *1 38.19,43.4
X$3043 932 1062 1061 891 1033 1086 23 38 1063 OAI33_X1
* cell instance $3044 r0 *1 39.52,43.4
X$3044 1085 881 23 38 1062 NOR2_X1
* cell instance $3045 r0 *1 40.09,43.4
X$3045 23 38 FILLCELL_X1
* cell instance $3046 r0 *1 40.28,43.4
X$3046 1087 862 1098 23 38 1085 MUX2_X1
* cell instance $3047 r0 *1 41.61,43.4
X$3047 23 38 FILLCELL_X16
* cell instance $3048 r0 *1 44.65,43.4
X$3048 23 38 FILLCELL_X4
* cell instance $3049 r0 *1 45.41,43.4
X$3049 23 38 FILLCELL_X2
* cell instance $3050 r0 *1 45.79,43.4
X$3050 23 38 FILLCELL_X1
* cell instance $3051 r0 *1 45.98,43.4
X$3051 693 23 38 1035 CLKBUF_X3
* cell instance $3052 r0 *1 46.93,43.4
X$3052 1036 992 301 23 38 1064 MUX2_X1
* cell instance $3053 r0 *1 48.26,43.4
X$3053 23 3096 1055 1037 1035 38 DFF_X1
* cell instance $3054 r0 *1 51.49,43.4
X$3054 23 38 FILLCELL_X2
* cell instance $3055 r0 *1 51.87,43.4
X$3055 23 2878 1101 1131 1035 38 DFF_X1
* cell instance $3056 r0 *1 55.1,43.4
X$3056 23 38 FILLCELL_X8
* cell instance $3057 r0 *1 56.62,43.4
X$3057 23 2857 1128 1129 1038 38 DFF_X1
* cell instance $3058 m0 *1 57,43.4
X$3058 864 38 476 23 BUF_X4
* cell instance $3059 m0 *1 56.81,43.4
X$3059 23 38 FILLCELL_X1
* cell instance $3060 m0 *1 58.33,43.4
X$3060 23 38 FILLCELL_X2
* cell instance $3061 m0 *1 58.9,43.4
X$3061 620 38 900 23 BUF_X4
* cell instance $3062 m0 *1 58.71,43.4
X$3062 23 38 FILLCELL_X1
* cell instance $3063 m0 *1 60.23,43.4
X$3063 23 2816 1092 1091 1038 38 DFF_X1
* cell instance $3064 m0 *1 63.46,43.4
X$3064 23 38 FILLCELL_X1
* cell instance $3065 m0 *1 63.65,43.4
X$3065 1066 441 799 23 38 1093 MUX2_X1
* cell instance $3066 m0 *1 64.98,43.4
X$3066 23 2810 1051 1039 954 38 DFF_X1
* cell instance $3067 m0 *1 68.21,43.4
X$3067 744 23 38 954 CLKBUF_X3
* cell instance $3068 m0 *1 69.16,43.4
X$3068 23 38 FILLCELL_X2
* cell instance $3069 r0 *1 59.14,43.4
X$3069 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $3070 r0 *1 59.14,43.4
X$3070 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $3071 r0 *1 59.14,43.4
X$3071 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $3072 r0 *1 59.85,43.4
X$3072 1092 1065 640 23 38 1091 MUX2_X1
* cell instance $3073 r0 *1 61.18,43.4
X$3073 23 38 FILLCELL_X8
* cell instance $3074 r0 *1 62.7,43.4
X$3074 23 2863 1066 1093 1038 38 DFF_X1
* cell instance $3075 r0 *1 65.93,43.4
X$3075 23 38 FILLCELL_X1
* cell instance $3076 r0 *1 66.12,43.4
X$3076 1066 438 1051 23 38 1067 MUX2_X1
* cell instance $3077 r0 *1 67.45,43.4
X$3077 1051 373 799 23 38 1039 MUX2_X1
* cell instance $3078 r0 *1 68.78,43.4
X$3078 23 2945 1040 1090 954 38 DFF_X1
* cell instance $3079 m0 *1 70.87,43.4
X$3079 23 38 FILLCELL_X2
* cell instance $3080 m0 *1 71.44,43.4
X$3080 1006 374 23 38 1147 NOR2_X1
* cell instance $3081 m0 *1 71.25,43.4
X$3081 23 38 FILLCELL_X1
* cell instance $3082 m0 *1 72.01,43.4
X$3082 23 38 FILLCELL_X4
* cell instance $3083 m0 *1 72.77,43.4
X$3083 23 38 FILLCELL_X1
* cell instance $3084 m0 *1 72.96,43.4
X$3084 23 2687 1048 1049 801 38 DFF_X1
* cell instance $3085 m0 *1 76.19,43.4
X$3085 1047 373 907 23 38 1046 MUX2_X1
* cell instance $3086 m0 *1 77.52,43.4
X$3086 23 38 FILLCELL_X16
* cell instance $3087 m0 *1 80.56,43.4
X$3087 23 38 FILLCELL_X2
* cell instance $3088 r0 *1 72.01,43.4
X$3088 23 38 FILLCELL_X8
* cell instance $3089 r0 *1 73.53,43.4
X$3089 23 38 FILLCELL_X2
* cell instance $3090 r0 *1 73.91,43.4
X$3090 1048 441 907 23 38 1049 MUX2_X1
* cell instance $3091 r0 *1 75.24,43.4
X$3091 1048 438 1047 23 38 1089 MUX2_X1
* cell instance $3092 r0 *1 76.57,43.4
X$3092 23 38 FILLCELL_X8
* cell instance $3093 r0 *1 78.09,43.4
X$3093 23 38 FILLCELL_X4
* cell instance $3094 r0 *1 78.85,43.4
X$3094 23 38 FILLCELL_X2
* cell instance $3095 r0 *1 79.23,43.4
X$3095 23 38 FILLCELL_X1
* cell instance $3096 r0 *1 79.42,43.4
X$3096 1082 374 23 38 1148 NOR2_X1
* cell instance $3097 r0 *1 79.99,43.4
X$3097 23 38 FILLCELL_X1
* cell instance $3098 r0 *1 80.18,43.4
X$3098 23 2904 1041 1084 1042 38 DFF_X1
* cell instance $3099 m0 *1 82.27,43.4
X$3099 1041 414 1068 23 38 1082 MUX2_X1
* cell instance $3100 m0 *1 80.94,43.4
X$3100 907 260 1041 23 38 1084 MUX2_X1
* cell instance $3101 m0 *1 83.6,43.4
X$3101 23 2833 1068 1044 1042 38 DFF_X1
* cell instance $3102 m0 *1 86.83,43.4
X$3102 23 38 FILLCELL_X1
* cell instance $3103 m0 *1 87.02,43.4
X$3103 23 2830 1070 1116 1042 38 DFF_X1
* cell instance $3104 m0 *1 90.25,43.4
X$3104 23 38 FILLCELL_X8
* cell instance $3105 m0 *1 91.77,43.4
X$3105 876 23 38 CLKBUF_X1
* cell instance $3106 m0 *1 92.34,43.4
X$3106 744 23 38 876 CLKBUF_X3
* cell instance $3107 m0 *1 93.29,43.4
X$3107 23 2852 1074 1076 876 38 DFF_X1
* cell instance $3108 m0 *1 96.52,43.4
X$3108 23 38 FILLCELL_X2
* cell instance $3109 r0 *1 83.41,43.4
X$3109 806 240 1068 23 38 1044 MUX2_X1
* cell instance $3110 r0 *1 84.74,43.4
X$3110 23 38 FILLCELL_X2
* cell instance $3111 r0 *1 85.12,43.4
X$3111 23 38 FILLCELL_X1
* cell instance $3112 r0 *1 85.31,43.4
X$3112 23 2918 1069 1118 1042 38 DFF_X1
* cell instance $3113 r0 *1 88.54,43.4
X$3113 1069 263 1070 23 38 1112 MUX2_X1
* cell instance $3114 r0 *1 89.87,43.4
X$3114 23 38 FILLCELL_X2
* cell instance $3115 r0 *1 90.25,43.4
X$3115 23 38 FILLCELL_X1
* cell instance $3116 r0 *1 90.44,43.4
X$3116 1072 263 1074 23 38 1071 MUX2_X1
* cell instance $3117 r0 *1 91.77,43.4
X$3117 1073 191 1072 23 38 1114 MUX2_X1
* cell instance $3118 r0 *1 93.1,43.4
X$3118 23 38 FILLCELL_X4
* cell instance $3119 r0 *1 93.86,43.4
X$3119 23 38 FILLCELL_X2
* cell instance $3120 r0 *1 94.24,43.4
X$3120 1073 187 1074 23 38 1076 MUX2_X1
* cell instance $3121 r0 *1 95.57,43.4
X$3121 23 38 FILLCELL_X8
* cell instance $3122 r180 *1 97.28,43.4
X$3122 23 38 23 38 TAPCELL_X1
* cell instance $3123 m0 *1 96.9,43.4
X$3123 23 38 FILLCELL_X1
* cell instance $3124 m90 *1 97.28,43.4
X$3124 23 38 23 38 TAPCELL_X1
* cell instance $3125 m0 *1 1.33,37.8
X$3125 23 38 FILLCELL_X8
* cell instance $3126 m0 *1 1.14,37.8
X$3126 23 38 23 38 TAPCELL_X1
* cell instance $3127 m0 *1 2.85,37.8
X$3127 23 38 FILLCELL_X2
* cell instance $3128 r0 *1 1.14,37.8
X$3128 23 38 23 38 TAPCELL_X1
* cell instance $3129 r0 *1 1.33,37.8
X$3129 23 38 FILLCELL_X2
* cell instance $3130 r0 *1 1.71,37.8
X$3130 23 3025 887 960 789 38 DFF_X1
* cell instance $3131 r0 *1 3.14,37.8
X$3131 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $3132 r0 *1 3.14,37.8
X$3132 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $3133 r0 *1 3.14,37.8
X$3133 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $3134 m0 *1 6.46,37.8
X$3134 845 813 691 23 38 915 MUX2_X1
* cell instance $3135 m0 *1 3.23,37.8
X$3135 23 2694 845 870 789 38 DFF_X1
* cell instance $3136 m0 *1 7.79,37.8
X$3136 693 23 38 789 CLKBUF_X3
* cell instance $3137 m0 *1 8.74,37.8
X$3137 23 38 FILLCELL_X32
* cell instance $3138 m0 *1 14.82,37.8
X$3138 23 38 FILLCELL_X4
* cell instance $3139 m0 *1 15.58,37.8
X$3139 23 38 FILLCELL_X2
* cell instance $3140 r0 *1 4.94,37.8
X$3140 887 992 295 23 38 960 MUX2_X1
* cell instance $3141 r0 *1 6.27,37.8
X$3141 23 3065 928 962 789 38 DFF_X1
* cell instance $3142 r0 *1 9.5,37.8
X$3142 23 38 FILLCELL_X8
* cell instance $3143 r0 *1 11.02,37.8
X$3143 23 3073 930 916 789 38 DFF_X1
* cell instance $3144 r0 *1 14.25,37.8
X$3144 930 858 295 23 38 916 MUX2_X1
* cell instance $3145 r0 *1 15.58,37.8
X$3145 23 38 FILLCELL_X2
* cell instance $3146 m0 *1 1.33,46.2
X$3146 23 38 FILLCELL_X8
* cell instance $3147 m0 *1 1.14,46.2
X$3147 23 38 23 38 TAPCELL_X1
* cell instance $3148 m0 *1 2.85,46.2
X$3148 23 38 FILLCELL_X2
* cell instance $3149 r0 *1 1.14,46.2
X$3149 23 38 23 38 TAPCELL_X1
* cell instance $3150 r0 *1 1.33,46.2
X$3150 23 38 FILLCELL_X2
* cell instance $3151 r0 *1 1.71,46.2
X$3151 23 3026 1132 1149 1094 38 DFF_X1
* cell instance $3152 r0 *1 3.14,46.2
X$3152 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $3153 r0 *1 3.14,46.2
X$3153 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $3154 r0 *1 3.14,46.2
X$3154 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $3155 m0 *1 3.42,46.2
X$3155 1132 941 591 23 38 1149 MUX2_X1
* cell instance $3156 m0 *1 3.23,46.2
X$3156 23 38 FILLCELL_X1
* cell instance $3157 m0 *1 4.75,46.2
X$3157 23 38 FILLCELL_X2
* cell instance $3158 r0 *1 4.94,46.2
X$3158 1150 992 591 23 38 1168 MUX2_X1
* cell instance $3159 m0 *1 8.36,46.2
X$3159 23 38 FILLCELL_X8
* cell instance $3160 m0 *1 5.13,46.2
X$3160 23 2706 1056 1075 1094 38 DFF_X1
* cell instance $3161 m0 *1 9.88,46.2
X$3161 23 38 FILLCELL_X2
* cell instance $3162 r0 *1 6.27,46.2
X$3162 23 38 FILLCELL_X4
* cell instance $3163 r0 *1 7.03,46.2
X$3163 23 38 FILLCELL_X1
* cell instance $3164 r0 *1 7.22,46.2
X$3164 1132 994 1150 23 38 1155 MUX2_X1
* cell instance $3165 r0 *1 8.55,46.2
X$3165 693 23 38 1094 CLKBUF_X3
* cell instance $3166 r0 *1 9.5,46.2
X$3166 1094 23 38 3151 INV_X1
* cell instance $3167 r0 *1 9.88,46.2
X$3167 23 38 FILLCELL_X1
* cell instance $3168 r0 *1 10.07,46.2
X$3168 23 3082 1133 1151 1094 38 DFF_X1
* cell instance $3169 m0 *1 10.45,46.2
X$3169 23 2696 1095 1115 1094 38 DFF_X1
* cell instance $3170 m0 *1 10.26,46.2
X$3170 23 38 FILLCELL_X1
* cell instance $3171 m0 *1 13.68,46.2
X$3171 1095 858 502 23 38 1115 MUX2_X1
* cell instance $3172 m0 *1 15.01,46.2
X$3172 1095 1184 1057 23 38 1117 MUX2_X1
* cell instance $3173 m0 *1 16.34,46.2
X$3173 23 38 FILLCELL_X1
* cell instance $3174 m0 *1 16.53,46.2
X$3174 1117 893 23 38 1096 NOR2_X1
* cell instance $3175 m0 *1 17.1,46.2
X$3175 23 38 FILLCELL_X8
* cell instance $3176 m0 *1 18.62,46.2
X$3176 23 38 FILLCELL_X4
* cell instance $3177 m0 *1 19.38,46.2
X$3177 1058 531 1138 1157 1139 38 23 1119 OAI221_X1
* cell instance $3178 m0 *1 20.52,46.2
X$3178 1158 1097 23 38 1141 NAND2_X1
* cell instance $3179 m0 *1 21.09,46.2
X$3179 23 38 FILLCELL_X2
* cell instance $3180 r0 *1 13.3,46.2
X$3180 1133 858 591 23 38 1151 MUX2_X1
* cell instance $3181 r0 *1 14.63,46.2
X$3181 23 38 FILLCELL_X8
* cell instance $3182 r0 *1 16.15,46.2
X$3182 1155 937 23 38 1134 NOR2_X1
* cell instance $3183 r0 *1 16.72,46.2
X$3183 932 1134 1187 1142 931 877 23 38 1135 OAI33_X1
* cell instance $3184 r0 *1 18.05,46.2
X$3184 23 38 FILLCELL_X2
* cell instance $3185 r0 *1 18.43,46.2
X$3185 1058 531 1136 1137 38 23 1237 OAI22_X2
* cell instance $3186 r0 *1 20.14,46.2
X$3186 1097 1140 23 38 1195 NAND2_X1
* cell instance $3187 r0 *1 20.71,46.2
X$3187 23 3071 1097 1192 991 38 DFF_X1
* cell instance $3188 m0 *1 21.66,46.2
X$3188 1205 1122 23 38 1121 NAND2_X1
* cell instance $3189 m0 *1 21.47,46.2
X$3189 23 38 FILLCELL_X1
* cell instance $3190 m0 *1 22.23,46.2
X$3190 23 38 FILLCELL_X8
* cell instance $3191 m0 *1 23.75,46.2
X$3191 23 38 FILLCELL_X4
* cell instance $3192 m0 *1 24.51,46.2
X$3192 23 38 FILLCELL_X1
* cell instance $3193 m0 *1 24.7,46.2
X$3193 634 38 813 23 BUF_X4
* cell instance $3194 m0 *1 26.03,46.2
X$3194 23 38 FILLCELL_X16
* cell instance $3195 m0 *1 29.07,46.2
X$3195 23 38 FILLCELL_X8
* cell instance $3196 m0 *1 30.59,46.2
X$3196 23 38 FILLCELL_X4
* cell instance $3197 m0 *1 31.35,46.2
X$3197 23 38 FILLCELL_X2
* cell instance $3198 r0 *1 23.94,46.2
X$3198 23 38 FILLCELL_X8
* cell instance $3199 r0 *1 25.46,46.2
X$3199 23 38 FILLCELL_X2
* cell instance $3200 r0 *1 25.84,46.2
X$3200 897 397 1136 1137 38 23 1199 OAI22_X2
* cell instance $3201 r0 *1 27.55,46.2
X$3201 23 38 FILLCELL_X32
* cell instance $3202 m0 *1 33.06,46.2
X$3202 23 38 FILLCELL_X4
* cell instance $3203 m0 *1 31.73,46.2
X$3203 634 38 70 23 BUF_X4
* cell instance $3204 m0 *1 33.82,46.2
X$3204 23 38 FILLCELL_X2
* cell instance $3205 r0 *1 33.63,46.2
X$3205 23 38 FILLCELL_X4
* cell instance $3206 m0 *1 34.39,46.2
X$3206 23 2849 1124 1125 942 38 DFF_X1
* cell instance $3207 m0 *1 34.2,46.2
X$3207 23 38 FILLCELL_X1
* cell instance $3208 m0 *1 37.62,46.2
X$3208 1083 858 319 23 38 1060 MUX2_X1
* cell instance $3209 m0 *1 38.95,46.2
X$3209 23 38 FILLCELL_X2
* cell instance $3210 r0 *1 34.39,46.2
X$3210 23 38 FILLCELL_X2
* cell instance $3211 r0 *1 34.77,46.2
X$3211 23 38 FILLCELL_X1
* cell instance $3212 r0 *1 34.96,46.2
X$3212 1143 1122 23 38 1173 NAND2_X1
* cell instance $3213 r0 *1 35.53,46.2
X$3213 23 38 FILLCELL_X1
* cell instance $3214 r0 *1 35.72,46.2
X$3214 1124 929 319 23 38 1125 MUX2_X1
* cell instance $3215 r0 *1 37.05,46.2
X$3215 23 2972 1087 1160 1174 38 DFF_X1
* cell instance $3216 m0 *1 40.66,46.2
X$3216 23 38 FILLCELL_X1
* cell instance $3217 m0 *1 39.33,46.2
X$3217 1087 941 319 23 38 1160 MUX2_X1
* cell instance $3218 m0 *1 40.85,46.2
X$3218 1098 992 319 23 38 1126 MUX2_X1
* cell instance $3219 m0 *1 42.18,46.2
X$3219 23 2719 1098 1126 1174 38 DFF_X1
* cell instance $3220 m0 *1 45.41,46.2
X$3220 23 38 FILLCELL_X2
* cell instance $3221 r0 *1 40.28,46.2
X$3221 23 38 FILLCELL_X2
* cell instance $3222 r0 *1 40.66,46.2
X$3222 23 38 FILLCELL_X1
* cell instance $3223 r0 *1 40.85,46.2
X$3223 634 38 1099 23 BUF_X4
* cell instance $3224 r0 *1 42.18,46.2
X$3224 23 38 FILLCELL_X16
* cell instance $3225 r0 *1 45.22,46.2
X$3225 23 38 FILLCELL_X4
* cell instance $3226 m0 *1 47.12,46.2
X$3226 23 38 FILLCELL_X2
* cell instance $3227 m0 *1 45.79,46.2
X$3227 1065 38 929 23 BUF_X4
* cell instance $3228 r0 *1 45.98,46.2
X$3228 23 38 FILLCELL_X2
* cell instance $3229 r0 *1 46.36,46.2
X$3229 1175 38 941 23 BUF_X4
* cell instance $3230 m0 *1 47.5,46.2
X$3230 1130 38 858 23 BUF_X4
* cell instance $3231 m0 *1 48.83,46.2
X$3231 1035 23 38 3136 INV_X2
* cell instance $3232 m0 *1 49.4,46.2
X$3232 23 38 FILLCELL_X8
* cell instance $3233 m0 *1 50.92,46.2
X$3233 23 38 FILLCELL_X2
* cell instance $3234 r0 *1 47.69,46.2
X$3234 23 3094 1144 1164 1035 38 DFF_X1
* cell instance $3235 r0 *1 50.92,46.2
X$3235 23 38 FILLCELL_X2
* cell instance $3236 m0 *1 26.79,74.2
X$3236 23 38 FILLCELL_X8
* cell instance $3237 m0 *1 26.22,74.2
X$3237 1926 937 23 38 1941 NOR2_X1
* cell instance $3238 m0 *1 28.31,74.2
X$3238 23 38 FILLCELL_X2
* cell instance $3239 r0 *1 26.22,74.2
X$3239 1940 1177 23 38 2037 NOR2_X1
* cell instance $3240 r0 *1 26.79,74.2
X$3240 23 38 FILLCELL_X8
* cell instance $3241 r0 *1 28.31,74.2
X$3241 23 38 FILLCELL_X2
* cell instance $3242 m0 *1 1.33,15.4
X$3242 23 38 FILLCELL_X8
* cell instance $3243 m0 *1 1.14,15.4
X$3243 23 38 23 38 TAPCELL_X1
* cell instance $3244 m0 *1 2.85,15.4
X$3244 23 2753 293 312 447 38 DFF_X1
* cell instance $3245 m0 *1 6.08,15.4
X$3245 294 257 295 23 38 268 MUX2_X1
* cell instance $3246 m0 *1 7.41,15.4
X$3246 23 38 FILLCELL_X16
* cell instance $3247 m0 *1 10.45,15.4
X$3247 23 38 FILLCELL_X8
* cell instance $3248 m0 *1 11.97,15.4
X$3248 23 38 FILLCELL_X4
* cell instance $3249 m0 *1 12.73,15.4
X$3249 23 38 FILLCELL_X2
* cell instance $3250 r0 *1 1.14,15.4
X$3250 23 38 23 38 TAPCELL_X1
* cell instance $3251 r0 *1 1.33,15.4
X$3251 23 38 FILLCELL_X8
* cell instance $3252 r0 *1 2.85,15.4
X$3252 23 38 FILLCELL_X4
* cell instance $3253 r0 *1 3.14,15.4
X$3253 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $3254 r0 *1 3.14,15.4
X$3254 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $3255 r0 *1 3.14,15.4
X$3255 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $3256 r0 *1 3.61,15.4
X$3256 23 38 FILLCELL_X2
* cell instance $3257 r0 *1 3.99,15.4
X$3257 293 318 295 23 38 312 MUX2_X1
* cell instance $3258 r0 *1 5.32,15.4
X$3258 293 412 294 23 38 337 MUX2_X1
* cell instance $3259 r0 *1 6.65,15.4
X$3259 23 38 FILLCELL_X16
* cell instance $3260 r0 *1 9.69,15.4
X$3260 23 38 FILLCELL_X4
* cell instance $3261 r0 *1 10.45,15.4
X$3261 337 354 23 38 339 NOR2_X1
* cell instance $3262 r0 *1 11.02,15.4
X$3262 23 38 FILLCELL_X4
* cell instance $3263 r0 *1 11.78,15.4
X$3263 23 38 FILLCELL_X1
* cell instance $3264 r0 *1 11.97,15.4
X$3264 27 23 38 295 BUF_X2
* cell instance $3265 r0 *1 12.73,15.4
X$3265 245 254 23 38 431 NOR2_X1
* cell instance $3266 m0 *1 13.3,15.4
X$3266 296 248 23 38 297 NOR2_X1
* cell instance $3267 m0 *1 13.11,15.4
X$3267 23 38 FILLCELL_X1
* cell instance $3268 m0 *1 13.87,15.4
X$3268 23 38 FILLCELL_X8
* cell instance $3269 m0 *1 15.39,15.4
X$3269 247 248 23 38 338 NOR2_X1
* cell instance $3270 m0 *1 15.96,15.4
X$3270 23 38 FILLCELL_X8
* cell instance $3271 m0 *1 17.48,15.4
X$3271 23 38 FILLCELL_X2
* cell instance $3272 r0 *1 13.3,15.4
X$3272 23 38 FILLCELL_X8
* cell instance $3273 r0 *1 14.82,15.4
X$3273 23 38 FILLCELL_X4
* cell instance $3274 r0 *1 15.58,15.4
X$3274 321 254 23 38 322 NOR2_X1
* cell instance $3275 r0 *1 16.15,15.4
X$3275 355 381 23 38 357 NOR2_X1
* cell instance $3276 r0 *1 16.72,15.4
X$3276 356 357 339 360 249 323 23 38 340 OAI33_X1
* cell instance $3277 m0 *1 18.43,15.4
X$3277 23 38 FILLCELL_X8
* cell instance $3278 m0 *1 17.86,15.4
X$3278 203 254 23 38 249 NOR2_X1
* cell instance $3279 m0 *1 19.95,15.4
X$3279 23 38 FILLCELL_X4
* cell instance $3280 m0 *1 20.71,15.4
X$3280 23 38 FILLCELL_X2
* cell instance $3281 r0 *1 18.05,15.4
X$3281 23 38 FILLCELL_X8
* cell instance $3282 r0 *1 19.57,15.4
X$3282 23 38 FILLCELL_X1
* cell instance $3283 r0 *1 19.76,15.4
X$3283 325 257 358 23 38 341 MUX2_X1
* cell instance $3284 m0 *1 21.28,15.4
X$3284 251 254 23 38 417 NOR2_X1
* cell instance $3285 m0 *1 21.09,15.4
X$3285 23 38 FILLCELL_X1
* cell instance $3286 m0 *1 21.85,15.4
X$3286 94 248 23 38 396 NOR2_X1
* cell instance $3287 m0 *1 22.42,15.4
X$3287 23 2805 298 326 324 38 DFF_X1
* cell instance $3288 m0 *1 25.65,15.4
X$3288 23 38 FILLCELL_X2
* cell instance $3289 r0 *1 21.09,15.4
X$3289 23 3041 325 341 324 38 DFF_X1
* cell instance $3290 r0 *1 24.32,15.4
X$3290 298 318 358 23 38 326 MUX2_X1
* cell instance $3291 r0 *1 25.65,15.4
X$3291 23 38 FILLCELL_X1
* cell instance $3292 r0 *1 25.84,15.4
X$3292 298 305 325 23 38 362 MUX2_X1
* cell instance $3293 m0 *1 26.6,15.4
X$3293 23 2768 344 343 73 38 DFF_X1
* cell instance $3294 m0 *1 26.03,15.4
X$3294 276 254 23 38 361 NOR2_X1
* cell instance $3295 m0 *1 29.83,15.4
X$3295 23 38 FILLCELL_X16
* cell instance $3296 m0 *1 32.87,15.4
X$3296 23 38 FILLCELL_X8
* cell instance $3297 m0 *1 34.39,15.4
X$3297 23 38 FILLCELL_X2
* cell instance $3298 r0 *1 27.17,15.4
X$3298 23 38 FILLCELL_X4
* cell instance $3299 r0 *1 27.93,15.4
X$3299 23 38 FILLCELL_X1
* cell instance $3300 r0 *1 28.12,15.4
X$3300 344 318 421 23 38 343 MUX2_X1
* cell instance $3301 r0 *1 29.45,15.4
X$3301 344 305 328 23 38 346 MUX2_X1
* cell instance $3302 r0 *1 30.78,15.4
X$3302 23 38 FILLCELL_X1
* cell instance $3303 r0 *1 30.97,15.4
X$3303 346 354 23 38 363 NOR2_X1
* cell instance $3304 r0 *1 31.54,15.4
X$3304 23 2928 328 387 73 38 DFF_X1
* cell instance $3305 m0 *1 34.96,15.4
X$3305 23 2756 330 317 73 38 DFF_X1
* cell instance $3306 m0 *1 34.77,15.4
X$3306 23 38 FILLCELL_X1
* cell instance $3307 m0 *1 38.19,15.4
X$3307 23 38 FILLCELL_X2
* cell instance $3308 r0 *1 34.77,15.4
X$3308 211 248 23 38 388 NOR2_X1
* cell instance $3309 r0 *1 35.34,15.4
X$3309 23 38 FILLCELL_X1
* cell instance $3310 r0 *1 35.53,15.4
X$3310 23 2869 366 389 329 38 DFF_X1
* cell instance $3311 m0 *1 39.9,15.4
X$3311 23 38 FILLCELL_X4
* cell instance $3312 m0 *1 38.57,15.4
X$3312 330 257 319 23 38 317 MUX2_X1
* cell instance $3313 m0 *1 40.66,15.4
X$3313 23 38 FILLCELL_X2
* cell instance $3314 r0 *1 38.76,15.4
X$3314 23 38 FILLCELL_X1
* cell instance $3315 r0 *1 38.95,15.4
X$3315 366 305 330 23 38 348 MUX2_X1
* cell instance $3316 r0 *1 40.28,15.4
X$3316 348 367 23 38 425 NOR2_X1
* cell instance $3317 r0 *1 40.85,15.4
X$3317 23 2872 368 350 299 38 DFF_X1
* cell instance $3318 m0 *1 41.61,15.4
X$3318 23 2744 300 320 299 38 DFF_X1
* cell instance $3319 m0 *1 41.04,15.4
X$3319 256 248 23 38 429 NOR2_X1
* cell instance $3320 m0 *1 44.84,15.4
X$3320 300 257 398 23 38 320 MUX2_X1
* cell instance $3321 m0 *1 46.17,15.4
X$3321 23 38 FILLCELL_X2
* cell instance $3322 r0 *1 44.08,15.4
X$3322 368 305 300 23 38 369 MUX2_X1
* cell instance $3323 r0 *1 45.41,15.4
X$3323 23 38 FILLCELL_X2
* cell instance $3324 r0 *1 45.79,15.4
X$3324 351 248 23 38 400 NOR2_X1
* cell instance $3325 r0 *1 46.36,15.4
X$3325 23 38 FILLCELL_X4
* cell instance $3326 m0 *1 46.74,15.4
X$3326 302 257 301 23 38 282 MUX2_X1
* cell instance $3327 m0 *1 46.55,15.4
X$3327 23 38 FILLCELL_X1
* cell instance $3328 m0 *1 48.07,15.4
X$3328 259 318 301 23 38 258 MUX2_X1
* cell instance $3329 m0 *1 49.4,15.4
X$3329 66 23 38 301 BUF_X2
* cell instance $3330 m0 *1 50.16,15.4
X$3330 23 38 FILLCELL_X2
* cell instance $3331 r0 *1 47.12,15.4
X$3331 23 3119 463 352 299 38 DFF_X1
* cell instance $3332 r0 *1 50.35,15.4
X$3332 23 38 FILLCELL_X4
* cell instance $3333 m0 *1 51.87,15.4
X$3333 23 38 FILLCELL_X8
* cell instance $3334 m0 *1 50.54,15.4
X$3334 259 305 302 23 38 353 MUX2_X1
* cell instance $3335 m0 *1 53.39,15.4
X$3335 23 38 FILLCELL_X2
* cell instance $3336 r0 *1 51.11,15.4
X$3336 23 38 FILLCELL_X2
* cell instance $3337 r0 *1 51.49,15.4
X$3337 23 38 FILLCELL_X1
* cell instance $3338 r0 *1 51.68,15.4
X$3338 353 367 23 38 371 NOR2_X1
* cell instance $3339 r0 *1 52.25,15.4
X$3339 23 38 FILLCELL_X8
* cell instance $3340 r0 *1 53.77,15.4
X$3340 23 38 FILLCELL_X4
* cell instance $3341 m0 *1 53.96,15.4
X$3341 23 2608 303 332 158 38 DFF_X1
* cell instance $3342 m0 *1 53.77,15.4
X$3342 23 38 FILLCELL_X1
* cell instance $3343 m0 *1 57.19,15.4
X$3343 23 38 FILLCELL_X1
* cell instance $3344 m0 *1 57.38,15.4
X$3344 23 2682 333 349 158 38 DFF_X1
* cell instance $3345 m0 *1 60.61,15.4
X$3345 23 38 FILLCELL_X2
* cell instance $3346 r0 *1 54.53,15.4
X$3346 112 286 303 23 38 332 MUX2_X1
* cell instance $3347 r0 *1 55.86,15.4
X$3347 112 243 333 23 38 349 MUX2_X1
* cell instance $3348 r0 *1 57.19,15.4
X$3348 303 126 333 23 38 424 MUX2_X1
* cell instance $3349 r0 *1 58.52,15.4
X$3349 23 38 FILLCELL_X16
* cell instance $3350 r0 *1 59.14,15.4
X$3350 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $3351 r0 *1 59.14,15.4
X$3351 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $3352 r0 *1 59.14,15.4
X$3352 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $3353 m0 *1 61.18,15.4
X$3353 23 2845 316 304 153 38 DFF_X1
* cell instance $3354 m0 *1 60.99,15.4
X$3354 23 38 FILLCELL_X1
* cell instance $3355 m0 *1 64.41,15.4
X$3355 23 38 FILLCELL_X2
* cell instance $3356 r0 *1 61.56,15.4
X$3356 23 38 FILLCELL_X2
* cell instance $3357 r0 *1 61.94,15.4
X$3357 23 38 FILLCELL_X1
* cell instance $3358 r0 *1 62.13,15.4
X$3358 23 2985 386 347 153 38 DFF_X1
* cell instance $3359 m0 *1 66.12,15.4
X$3359 23 38 FILLCELL_X4
* cell instance $3360 m0 *1 64.79,15.4
X$3360 316 305 290 23 38 306 MUX2_X1
* cell instance $3361 m0 *1 66.88,15.4
X$3361 78 260 315 23 38 288 MUX2_X1
* cell instance $3362 m0 *1 68.21,15.4
X$3362 153 23 38 3140 INV_X1
* cell instance $3363 m0 *1 68.59,15.4
X$3363 23 38 FILLCELL_X1
* cell instance $3364 m0 *1 68.78,15.4
X$3364 23 2590 345 292 334 38 DFF_X1
* cell instance $3365 m0 *1 72.01,15.4
X$3365 23 38 FILLCELL_X32
* cell instance $3366 m0 *1 78.09,15.4
X$3366 23 38 FILLCELL_X4
* cell instance $3367 m0 *1 78.85,15.4
X$3367 23 2586 307 314 334 38 DFF_X1
* cell instance $3368 m0 *1 82.08,15.4
X$3368 23 38 FILLCELL_X16
* cell instance $3369 m0 *1 85.12,15.4
X$3369 23 38 FILLCELL_X4
* cell instance $3370 m0 *1 85.88,15.4
X$3370 49 191 308 23 38 342 MUX2_X1
* cell instance $3371 m0 *1 87.21,15.4
X$3371 23 38 FILLCELL_X2
* cell instance $3372 r0 *1 65.36,15.4
X$3372 23 38 FILLCELL_X4
* cell instance $3373 r0 *1 66.12,15.4
X$3373 23 38 FILLCELL_X1
* cell instance $3374 r0 *1 66.31,15.4
X$3374 139 23 38 153 CLKBUF_X3
* cell instance $3375 r0 *1 67.26,15.4
X$3375 384 373 78 23 38 385 MUX2_X1
* cell instance $3376 r0 *1 68.59,15.4
X$3376 315 305 345 23 38 420 MUX2_X1
* cell instance $3377 r0 *1 69.92,15.4
X$3377 23 38 FILLCELL_X16
* cell instance $3378 r0 *1 72.96,15.4
X$3378 23 38 FILLCELL_X1
* cell instance $3379 r0 *1 73.15,15.4
X$3379 23 2865 375 383 334 38 DFF_X1
* cell instance $3380 r0 *1 76.38,15.4
X$3380 23 2935 376 382 334 38 DFF_X1
* cell instance $3381 r0 *1 79.61,15.4
X$3381 23 38 FILLCELL_X8
* cell instance $3382 r0 *1 81.13,15.4
X$3382 23 38 FILLCELL_X4
* cell instance $3383 r0 *1 81.89,15.4
X$3383 23 38 FILLCELL_X2
* cell instance $3384 r0 *1 83.6,15.4
X$3384 23 38 FILLCELL_X8
* cell instance $3385 r0 *1 85.12,15.4
X$3385 23 2893 308 342 310 38 DFF_X1
* cell instance $3386 m0 *1 88.92,15.4
X$3386 23 38 FILLCELL_X8
* cell instance $3387 m0 *1 87.59,15.4
X$3387 308 263 309 23 38 264 MUX2_X1
* cell instance $3388 m0 *1 90.44,15.4
X$3388 23 38 FILLCELL_X4
* cell instance $3389 m0 *1 91.2,15.4
X$3389 23 38 FILLCELL_X2
* cell instance $3390 r0 *1 88.35,15.4
X$3390 49 187 309 23 38 379 MUX2_X1
* cell instance $3391 r0 *1 89.68,15.4
X$3391 23 38 FILLCELL_X8
* cell instance $3392 r0 *1 91.2,15.4
X$3392 23 38 FILLCELL_X2
* cell instance $3393 m0 *1 1.33,49
X$3393 23 38 FILLCELL_X8
* cell instance $3394 m0 *1 1.14,49
X$3394 23 38 23 38 TAPCELL_X1
* cell instance $3395 m0 *1 2.85,49
X$3395 23 38 FILLCELL_X4
* cell instance $3396 m0 *1 3.61,49
X$3396 23 38 FILLCELL_X2
* cell instance $3397 r0 *1 1.14,49
X$3397 23 38 23 38 TAPCELL_X1
* cell instance $3398 r0 *1 1.33,49
X$3398 23 38 FILLCELL_X8
* cell instance $3399 r0 *1 2.85,49
X$3399 23 38 FILLCELL_X2
* cell instance $3400 r0 *1 3.14,49
X$3400 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $3401 r0 *1 3.14,49
X$3401 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $3402 r0 *1 3.14,49
X$3402 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $3403 r0 *1 3.23,49
X$3403 1232 23 38 1258 BUF_X1
* cell instance $3404 r0 *1 3.8,49
X$3404 1233 23 38 1260 BUF_X2
* cell instance $3405 m0 *1 4.18,49
X$3405 1196 23 38 1201 BUF_X1
* cell instance $3406 m0 *1 3.99,49
X$3406 23 38 FILLCELL_X1
* cell instance $3407 m0 *1 4.75,49
X$3407 23 2739 1150 1168 1094 38 DFF_X1
* cell instance $3408 m0 *1 7.98,49
X$3408 1197 23 38 1200 BUF_X2
* cell instance $3409 m0 *1 8.74,49
X$3409 23 38 FILLCELL_X16
* cell instance $3410 m0 *1 11.78,49
X$3410 23 38 FILLCELL_X4
* cell instance $3411 m0 *1 12.54,49
X$3411 1204 929 591 23 38 1203 MUX2_X1
* cell instance $3412 m0 *1 13.87,49
X$3412 23 38 FILLCELL_X2
* cell instance $3413 r0 *1 4.56,49
X$3413 1202 23 38 1167 BUF_X1
* cell instance $3414 r0 *1 5.13,49
X$3414 1209 23 38 1259 BUF_X2
* cell instance $3415 r0 *1 5.89,49
X$3415 23 38 FILLCELL_X32
* cell instance $3416 r0 *1 11.97,49
X$3416 23 38 FILLCELL_X2
* cell instance $3417 r0 *1 12.35,49
X$3417 23 3095 1204 1203 1326 38 DFF_X1
* cell instance $3418 m0 *1 15.58,49
X$3418 23 38 FILLCELL_X2
* cell instance $3419 m0 *1 14.25,49
X$3419 1133 1184 1204 23 38 1236 MUX2_X1
* cell instance $3420 r0 *1 15.58,49
X$3420 23 38 FILLCELL_X4
* cell instance $3421 m0 *1 16.15,49
X$3421 1236 893 23 38 1187 NOR2_X1
* cell instance $3422 m0 *1 15.96,49
X$3422 23 38 FILLCELL_X1
* cell instance $3423 m0 *1 16.72,49
X$3423 23 38 FILLCELL_X4
* cell instance $3424 m0 *1 17.48,49
X$3424 23 38 FILLCELL_X2
* cell instance $3425 r0 *1 16.34,49
X$3425 23 38 FILLCELL_X1
* cell instance $3426 r0 *1 16.53,49
X$3426 1097 1122 23 38 1238 NAND2_X1
* cell instance $3427 r0 *1 17.1,49
X$3427 1188 1213 1121 38 23 1202 OAI21_X2
* cell instance $3428 m0 *1 19.57,49
X$3428 23 38 FILLCELL_X1
* cell instance $3429 m0 *1 17.86,49
X$3429 1135 614 1136 1137 38 23 1188 OAI22_X2
* cell instance $3430 m0 *1 19.76,49
X$3430 1135 614 1138 1157 1139 38 23 1193 OAI221_X1
* cell instance $3431 m0 *1 20.9,49
X$3431 1206 1141 1119 1208 1195 38 23 1192 OAI221_X1
* cell instance $3432 m0 *1 22.04,49
X$3432 23 38 FILLCELL_X1
* cell instance $3433 m0 *1 22.23,49
X$3433 23 2758 1205 1169 991 38 DFF_X1
* cell instance $3434 m0 *1 25.46,49
X$3434 1199 1210 1244 38 23 1197 OAI21_X4
* cell instance $3435 m0 *1 27.93,49
X$3435 1170 1122 23 38 1244 NAND2_X1
* cell instance $3436 m0 *1 28.5,49
X$3436 23 38 FILLCELL_X2
* cell instance $3437 r0 *1 18.43,49
X$3437 1237 1210 1238 38 23 1232 OAI21_X4
* cell instance $3438 r0 *1 20.9,49
X$3438 23 38 FILLCELL_X1
* cell instance $3439 r0 *1 21.09,49
X$3439 1158 1205 23 38 1207 NAND2_X1
* cell instance $3440 r0 *1 21.66,49
X$3440 1206 1207 1193 1208 1242 38 23 1169 OAI221_X1
* cell instance $3441 r0 *1 22.8,49
X$3441 23 38 FILLCELL_X1
* cell instance $3442 r0 *1 22.99,49
X$3442 1205 1140 23 38 1242 NAND2_X1
* cell instance $3443 r0 *1 23.56,49
X$3443 23 38 FILLCELL_X2
* cell instance $3444 r0 *1 23.94,49
X$3444 1206 1281 1280 1208 1243 38 23 1315 OAI221_X1
* cell instance $3445 r0 *1 25.08,49
X$3445 23 38 FILLCELL_X2
* cell instance $3446 r0 *1 25.46,49
X$3446 897 397 1138 1157 1139 38 23 1280 OAI221_X1
* cell instance $3447 r0 *1 26.6,49
X$3447 23 38 FILLCELL_X2
* cell instance $3448 r0 *1 26.98,49
X$3448 1282 1210 1211 38 23 1209 OAI21_X4
* cell instance $3449 m0 *1 29.45,49
X$3449 23 38 FILLCELL_X4
* cell instance $3450 m0 *1 28.88,49
X$3450 1171 1122 23 38 1211 NAND2_X1
* cell instance $3451 m0 *1 30.21,49
X$3451 1158 1171 23 38 1212 NAND2_X1
* cell instance $3452 m0 *1 30.78,49
X$3452 1206 1212 1172 1208 1263 38 23 1246 OAI221_X1
* cell instance $3453 m0 *1 31.92,49
X$3453 1021 422 1138 1198 1139 38 23 1172 OAI221_X1
* cell instance $3454 m0 *1 33.06,49
X$3454 1194 1213 1173 38 23 1196 OAI21_X4
* cell instance $3455 m0 *1 35.53,49
X$3455 23 997 423 1136 1194 1137 38 OAI22_X4
* cell instance $3456 m0 *1 38.76,49
X$3456 23 38 FILLCELL_X4
* cell instance $3457 m0 *1 39.52,49
X$3457 23 38 FILLCELL_X1
* cell instance $3458 m0 *1 39.71,49
X$3458 620 38 1184 23 BUF_X4
* cell instance $3459 m0 *1 41.04,49
X$3459 23 38 FILLCELL_X4
* cell instance $3460 m0 *1 41.8,49
X$3460 862 38 212 23 BUF_X4
* cell instance $3461 m0 *1 43.13,49
X$3461 988 38 254 23 BUF_X4
* cell instance $3462 m0 *1 44.46,49
X$3462 901 460 1138 1198 1139 38 23 1191 OAI221_X1
* cell instance $3463 m0 *1 45.6,49
X$3463 23 38 FILLCELL_X8
* cell instance $3464 m0 *1 47.12,49
X$3464 23 38 FILLCELL_X4
* cell instance $3465 m0 *1 47.88,49
X$3465 1214 38 992 23 BUF_X4
* cell instance $3466 m0 *1 49.21,49
X$3466 23 38 FILLCELL_X2
* cell instance $3467 r0 *1 29.45,49
X$3467 23 3086 1171 1246 1262 38 DFF_X1
* cell instance $3468 r0 *1 32.68,49
X$3468 1021 422 1136 1137 38 23 1282 OAI22_X2
* cell instance $3469 r0 *1 34.39,49
X$3469 1206 1249 1248 1208 1251 38 23 1264 OAI221_X1
* cell instance $3470 r0 *1 35.53,49
X$3470 997 423 1138 1198 1139 38 23 1248 OAI221_X1
* cell instance $3471 r0 *1 36.67,49
X$3471 23 38 FILLCELL_X2
* cell instance $3472 r0 *1 37.05,49
X$3472 1286 1265 1213 38 23 1285 OAI21_X4
* cell instance $3473 r0 *1 39.52,49
X$3473 23 38 FILLCELL_X2
* cell instance $3474 r0 *1 39.9,49
X$3474 23 38 FILLCELL_X1
* cell instance $3475 r0 *1 40.09,49
X$3475 1174 23 38 CLKBUF_X1
* cell instance $3476 r0 *1 40.66,49
X$3476 1253 1287 1213 38 23 1233 OAI21_X4
* cell instance $3477 r0 *1 43.13,49
X$3477 23 901 460 1136 1253 1137 38 OAI22_X4
* cell instance $3478 r0 *1 46.36,49
X$3478 23 38 FILLCELL_X4
* cell instance $3479 r0 *1 47.12,49
X$3479 23 38 FILLCELL_X2
* cell instance $3480 r0 *1 47.5,49
X$3480 634 38 414 23 BUF_X4
* cell instance $3481 r0 *1 48.83,49
X$3481 23 38 FILLCELL_X4
* cell instance $3482 m0 *1 50.92,49
X$3482 1144 1175 556 23 38 1164 MUX2_X1
* cell instance $3483 m0 *1 49.59,49
X$3483 1254 1214 556 23 38 1215 MUX2_X1
* cell instance $3484 m0 *1 52.25,49
X$3484 23 38 FILLCELL_X1
* cell instance $3485 m0 *1 52.44,49
X$3485 1144 862 1254 23 38 1255 MUX2_X1
* cell instance $3486 m0 *1 53.77,49
X$3486 23 38 FILLCELL_X4
* cell instance $3487 m0 *1 54.53,49
X$3487 23 38 FILLCELL_X1
* cell instance $3488 m0 *1 54.72,49
X$3488 1255 881 23 38 1190 NOR2_X1
* cell instance $3489 m0 *1 55.29,49
X$3489 864 38 1142 23 BUF_X4
* cell instance $3490 m0 *1 56.62,49
X$3490 23 38 FILLCELL_X4
* cell instance $3491 m0 *1 57.38,49
X$3491 23 38 FILLCELL_X2
* cell instance $3492 r0 *1 49.59,49
X$3492 37 23 38 434 CLKBUF_X3
* cell instance $3493 r0 *1 50.54,49
X$3493 23 38 FILLCELL_X1
* cell instance $3494 r0 *1 50.73,49
X$3494 23 3093 1254 1215 1038 38 DFF_X1
* cell instance $3495 r0 *1 53.96,49
X$3495 23 38 FILLCELL_X8
* cell instance $3496 r0 *1 55.48,49
X$3496 23 38 FILLCELL_X4
* cell instance $3497 r0 *1 56.24,49
X$3497 23 38 FILLCELL_X2
* cell instance $3498 r0 *1 56.62,49
X$3498 23 38 FILLCELL_X1
* cell instance $3499 r0 *1 56.81,49
X$3499 23 3092 1216 1256 1038 38 DFF_X1
* cell instance $3500 m0 *1 57.95,49
X$3500 1216 1175 640 23 38 1256 MUX2_X1
* cell instance $3501 m0 *1 57.76,49
X$3501 23 38 FILLCELL_X1
* cell instance $3502 m0 *1 59.28,49
X$3502 1217 1214 640 23 38 1288 MUX2_X1
* cell instance $3503 m0 *1 60.61,49
X$3503 23 38 FILLCELL_X2
* cell instance $3504 r0 *1 59.14,49
X$3504 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $3505 r0 *1 59.14,49
X$3505 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $3506 r0 *1 59.14,49
X$3506 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $3507 r0 *1 60.04,49
X$3507 1216 862 1217 23 38 1257 MUX2_X1
* cell instance $3508 m0 *1 61.18,49
X$3508 1257 881 23 38 1176 NOR2_X1
* cell instance $3509 m0 *1 60.99,49
X$3509 23 38 FILLCELL_X1
* cell instance $3510 m0 *1 61.75,49
X$3510 23 38 FILLCELL_X4
* cell instance $3511 m0 *1 62.51,49
X$3511 23 38 FILLCELL_X1
* cell instance $3512 m0 *1 62.7,49
X$3512 796 38 260 23 BUF_X4
* cell instance $3513 m0 *1 64.03,49
X$3513 23 38 FILLCELL_X8
* cell instance $3514 m0 *1 65.55,49
X$3514 23 38 FILLCELL_X1
* cell instance $3515 m0 *1 65.74,49
X$3515 243 38 187 23 BUF_X4
* cell instance $3516 m0 *1 67.07,49
X$3516 23 38 FILLCELL_X16
* cell instance $3517 m0 *1 70.11,49
X$3517 23 38 FILLCELL_X2
* cell instance $3518 r0 *1 61.37,49
X$3518 23 38 FILLCELL_X1
* cell instance $3519 r0 *1 61.56,49
X$3519 863 38 51 23 BUF_X4
* cell instance $3520 r0 *1 62.89,49
X$3520 23 38 FILLCELL_X2
* cell instance $3521 r0 *1 63.27,49
X$3521 286 38 191 23 BUF_X4
* cell instance $3522 r0 *1 64.6,49
X$3522 23 3090 1302 1284 1301 38 DFF_X1
* cell instance $3523 r0 *1 67.83,49
X$3523 23 38 FILLCELL_X1
* cell instance $3524 r0 *1 68.02,49
X$3524 515 38 227 23 BUF_X4
* cell instance $3525 r0 *1 69.35,49
X$3525 1219 1220 23 600 38 NAND2_X4
* cell instance $3526 m0 *1 73.72,49
X$3526 1221 541 1222 23 38 1252 MUX2_X1
* cell instance $3527 m0 *1 70.49,49
X$3527 23 2779 1221 1186 954 38 DFF_X1
* cell instance $3528 m0 *1 75.05,49
X$3528 1222 520 907 23 38 1185 MUX2_X1
* cell instance $3529 m0 *1 76.38,49
X$3529 1252 1177 23 38 1183 NOR2_X1
* cell instance $3530 m0 *1 76.95,49
X$3530 23 38 FILLCELL_X16
* cell instance $3531 m0 *1 79.99,49
X$3531 23 38 FILLCELL_X4
* cell instance $3532 m0 *1 80.75,49
X$3532 1111 79 1283 23 38 1250 MUX2_X1
* cell instance $3533 m0 *1 82.08,49
X$3533 23 38 FILLCELL_X16
* cell instance $3534 m0 *1 85.12,49
X$3534 474 285 1241 1240 1224 38 23 1182 OAI221_X1
* cell instance $3535 m0 *1 86.26,49
X$3535 1225 1181 1182 1226 1245 38 23 1247 OAI221_X1
* cell instance $3536 m0 *1 87.4,49
X$3536 1228 1178 23 38 1181 NAND2_X1
* cell instance $3537 m0 *1 87.97,49
X$3537 1178 1239 23 38 1245 NAND2_X1
* cell instance $3538 m0 *1 88.54,49
X$3538 23 38 FILLCELL_X8
* cell instance $3539 m0 *1 90.06,49
X$3539 23 38 FILLCELL_X4
* cell instance $3540 m0 *1 90.82,49
X$3540 23 38 FILLCELL_X2
* cell instance $3541 r0 *1 71.06,49
X$3541 1219 1355 23 38 864 NAND2_X2
* cell instance $3542 r0 *1 72.01,49
X$3542 23 38 FILLCELL_X8
* cell instance $3543 r0 *1 73.53,49
X$3543 23 38 FILLCELL_X4
* cell instance $3544 r0 *1 74.29,49
X$3544 23 3112 1222 1185 1223 38 DFF_X1
* cell instance $3545 r0 *1 77.52,49
X$3545 23 38 FILLCELL_X8
* cell instance $3546 r0 *1 79.04,49
X$3546 23 38 FILLCELL_X4
* cell instance $3547 r0 *1 79.8,49
X$3547 23 38 FILLCELL_X2
* cell instance $3548 r0 *1 80.18,49
X$3548 23 3111 1283 1250 1223 38 DFF_X1
* cell instance $3549 r0 *1 83.41,49
X$3549 23 38 FILLCELL_X8
* cell instance $3550 r0 *1 84.93,49
X$3550 23 38 FILLCELL_X2
* cell instance $3551 r0 *1 85.31,49
X$3551 23 38 FILLCELL_X1
* cell instance $3552 r0 *1 85.5,49
X$3552 23 3113 1178 1247 1223 38 DFF_X1
* cell instance $3553 r0 *1 88.73,49
X$3553 1178 1230 23 38 1270 NAND2_X1
* cell instance $3554 r0 *1 89.3,49
X$3554 23 38 FILLCELL_X2
* cell instance $3555 r0 *1 89.68,49
X$3555 483 265 1241 1240 1224 38 23 1279 OAI221_X1
* cell instance $3556 r0 *1 90.82,49
X$3556 23 3117 1272 1271 1227 38 DFF_X1
* cell instance $3557 m0 *1 91.39,49
X$3557 649 608 1241 1240 1224 38 23 1180 OAI221_X1
* cell instance $3558 m0 *1 91.2,49
X$3558 23 38 FILLCELL_X1
* cell instance $3559 m0 *1 92.53,49
X$3559 23 38 FILLCELL_X1
* cell instance $3560 m0 *1 92.72,49
X$3560 1225 1229 1180 1226 1235 38 23 1179 OAI221_X1
* cell instance $3561 m0 *1 93.86,49
X$3561 23 2775 1234 1179 876 38 DFF_X1
* cell instance $3562 r180 *1 97.28,49
X$3562 23 38 23 38 TAPCELL_X1
* cell instance $3563 r0 *1 94.05,49
X$3563 1228 1234 23 38 1229 NAND2_X1
* cell instance $3564 r0 *1 94.62,49
X$3564 1234 1239 23 38 1235 NAND2_X1
* cell instance $3565 r0 *1 95.19,49
X$3565 23 38 FILLCELL_X2
* cell instance $3566 r0 *1 95.57,49
X$3566 23 38 FILLCELL_X1
* cell instance $3567 r0 *1 95.76,49
X$3567 1234 1230 23 38 1231 NAND2_X1
* cell instance $3568 r0 *1 96.33,49
X$3568 1278 23 38 1274 BUF_X1
* cell instance $3569 r0 *1 96.9,49
X$3569 23 38 FILLCELL_X1
* cell instance $3570 m90 *1 97.28,49
X$3570 23 38 23 38 TAPCELL_X1
* cell instance $3571 m0 *1 59.28,96.6
X$3571 23 38 FILLCELL_X2
* cell instance $3572 m0 *1 58.71,96.6
X$3572 2532 23 38 2182 BUF_X1
* cell instance $3573 r0 *1 59.14,96.6
X$3573 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $3574 r0 *1 59.14,96.6
X$3574 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $3575 r0 *1 59.14,96.6
X$3575 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $3576 m0 *1 1.33,57.4
X$3576 23 38 FILLCELL_X2
* cell instance $3577 m0 *1 1.14,57.4
X$3577 23 38 23 38 TAPCELL_X1
* cell instance $3578 r0 *1 1.14,57.4
X$3578 23 38 23 38 TAPCELL_X1
* cell instance $3579 r0 *1 1.33,57.4
X$3579 23 38 FILLCELL_X8
* cell instance $3580 m0 *1 4.94,57.4
X$3580 23 38 FILLCELL_X2
* cell instance $3581 m0 *1 1.71,57.4
X$3581 23 2809 1479 1501 1292 38 DFF_X1
* cell instance $3582 r0 *1 2.85,57.4
X$3582 23 38 FILLCELL_X4
* cell instance $3583 r0 *1 3.14,57.4
X$3583 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $3584 r0 *1 3.14,57.4
X$3584 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $3585 r0 *1 3.14,57.4
X$3585 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $3586 r0 *1 3.61,57.4
X$3586 23 38 FILLCELL_X1
* cell instance $3587 r0 *1 3.8,57.4
X$3587 1325 1493 1479 23 38 1501 MUX2_X1
* cell instance $3588 r0 *1 5.13,57.4
X$3588 23 38 FILLCELL_X2
* cell instance $3589 m0 *1 5.51,57.4
X$3589 1479 70 1481 23 38 1468 MUX2_X1
* cell instance $3590 m0 *1 5.32,57.4
X$3590 23 38 FILLCELL_X1
* cell instance $3591 m0 *1 6.84,57.4
X$3591 23 38 FILLCELL_X2
* cell instance $3592 r0 *1 5.51,57.4
X$3592 23 38 FILLCELL_X1
* cell instance $3593 r0 *1 5.7,57.4
X$3593 1325 1480 1481 23 38 1571 MUX2_X1
* cell instance $3594 r0 *1 7.03,57.4
X$3594 23 38 FILLCELL_X2
* cell instance $3595 m0 *1 7.41,57.4
X$3595 23 2612 1505 1504 1292 38 DFF_X1
* cell instance $3596 m0 *1 7.22,57.4
X$3596 23 38 FILLCELL_X1
* cell instance $3597 m0 *1 10.64,57.4
X$3597 1468 1483 23 38 1467 NOR2_X1
* cell instance $3598 m0 *1 11.21,57.4
X$3598 23 38 FILLCELL_X32
* cell instance $3599 m0 *1 17.29,57.4
X$3599 23 38 FILLCELL_X16
* cell instance $3600 m0 *1 20.33,57.4
X$3600 23 38 FILLCELL_X8
* cell instance $3601 m0 *1 21.85,57.4
X$3601 23 38 FILLCELL_X4
* cell instance $3602 m0 *1 22.61,57.4
X$3602 23 38 FILLCELL_X1
* cell instance $3603 m0 *1 22.8,57.4
X$3603 23 2616 1484 1445 1399 38 DFF_X1
* cell instance $3604 m0 *1 26.03,57.4
X$3604 23 38 FILLCELL_X4
* cell instance $3605 m0 *1 26.79,57.4
X$3605 23 38 FILLCELL_X2
* cell instance $3606 r0 *1 7.41,57.4
X$3606 1361 1544 1505 23 38 1504 MUX2_X1
* cell instance $3607 r0 *1 8.74,57.4
X$3607 1292 23 38 CLKBUF_X1
* cell instance $3608 r0 *1 9.31,57.4
X$3608 23 38 FILLCELL_X1
* cell instance $3609 r0 *1 9.5,57.4
X$3609 1325 1482 1507 23 38 1545 MUX2_X1
* cell instance $3610 r0 *1 10.83,57.4
X$3610 23 38 FILLCELL_X4
* cell instance $3611 r0 *1 11.59,57.4
X$3611 1505 813 1507 23 38 1508 MUX2_X1
* cell instance $3612 r0 *1 12.92,57.4
X$3612 23 38 FILLCELL_X16
* cell instance $3613 r0 *1 15.96,57.4
X$3613 23 38 FILLCELL_X2
* cell instance $3614 r0 *1 16.34,57.4
X$3614 23 2977 1533 1546 1399 38 DFF_X1
* cell instance $3615 r0 *1 19.57,57.4
X$3615 23 38 FILLCELL_X8
* cell instance $3616 r0 *1 21.09,57.4
X$3616 23 38 FILLCELL_X4
* cell instance $3617 r0 *1 21.85,57.4
X$3617 23 38 FILLCELL_X2
* cell instance $3618 r0 *1 22.23,57.4
X$3618 1325 1530 1484 23 38 1445 MUX2_X1
* cell instance $3619 r0 *1 23.56,57.4
X$3619 23 38 FILLCELL_X2
* cell instance $3620 r0 *1 23.94,57.4
X$3620 1508 831 23 38 1514 NOR2_X1
* cell instance $3621 r0 *1 24.51,57.4
X$3621 1361 1492 1534 23 38 1547 MUX2_X1
* cell instance $3622 r0 *1 25.84,57.4
X$3622 23 38 FILLCELL_X1
* cell instance $3623 r0 *1 26.03,57.4
X$3623 1534 792 1484 23 38 1509 MUX2_X1
* cell instance $3624 m0 *1 27.36,57.4
X$3624 1447 893 23 38 1448 NOR2_X1
* cell instance $3625 m0 *1 27.17,57.4
X$3625 23 38 FILLCELL_X1
* cell instance $3626 m0 *1 27.93,57.4
X$3626 1449 937 23 38 1510 NOR2_X1
* cell instance $3627 m0 *1 28.5,57.4
X$3627 1262 23 38 CLKBUF_X1
* cell instance $3628 m0 *1 29.07,57.4
X$3628 1513 1426 1511 1137 38 23 1402 OAI22_X2
* cell instance $3629 m0 *1 30.78,57.4
X$3629 1486 23 38 1262 CLKBUF_X3
* cell instance $3630 m0 *1 31.73,57.4
X$3630 1452 994 1451 23 38 1449 MUX2_X1
* cell instance $3631 m0 *1 33.06,57.4
X$3631 1452 1487 1361 23 38 1453 MUX2_X1
* cell instance $3632 m0 *1 34.39,57.4
X$3632 881 38 1483 23 BUF_X4
* cell instance $3633 m0 *1 35.72,57.4
X$3633 403 23 38 829 CLKBUF_X3
* cell instance $3634 m0 *1 36.67,57.4
X$3634 23 38 FILLCELL_X4
* cell instance $3635 m0 *1 37.43,57.4
X$3635 23 38 FILLCELL_X2
* cell instance $3636 r0 *1 27.36,57.4
X$3636 23 38 FILLCELL_X1
* cell instance $3637 r0 *1 27.55,57.4
X$3637 1509 829 23 38 1512 NOR2_X1
* cell instance $3638 r0 *1 28.12,57.4
X$3638 23 38 FILLCELL_X2
* cell instance $3639 r0 *1 28.5,57.4
X$3639 1485 1510 1448 1142 1514 1512 23 38 1513 OAI33_X1
* cell instance $3640 r0 *1 29.83,57.4
X$3640 23 3008 1451 1517 1262 38 DFF_X1
* cell instance $3641 r0 *1 33.06,57.4
X$3641 1451 1488 1361 23 38 1517 MUX2_X1
* cell instance $3642 r0 *1 34.39,57.4
X$3642 23 38 FILLCELL_X16
* cell instance $3643 r0 *1 37.43,57.4
X$3643 23 38 FILLCELL_X4
* cell instance $3644 m0 *1 38,57.4
X$3644 1158 1368 23 38 1437 NAND2_X1
* cell instance $3645 m0 *1 37.81,57.4
X$3645 23 38 FILLCELL_X1
* cell instance $3646 m0 *1 38.57,57.4
X$3646 23 2808 1489 1522 1174 38 DFF_X1
* cell instance $3647 m0 *1 41.8,57.4
X$3647 1299 38 994 23 BUF_X4
* cell instance $3648 m0 *1 43.13,57.4
X$3648 23 38 FILLCELL_X2
* cell instance $3649 r0 *1 38.19,57.4
X$3649 23 38 FILLCELL_X2
* cell instance $3650 r0 *1 38.57,57.4
X$3650 23 38 FILLCELL_X1
* cell instance $3651 r0 *1 38.76,57.4
X$3651 23 3000 1583 1549 1174 38 DFF_X1
* cell instance $3652 r0 *1 41.99,57.4
X$3652 1489 1488 1490 23 38 1522 MUX2_X1
* cell instance $3653 r0 *1 43.32,57.4
X$3653 403 38 1105 23 BUF_X4
* cell instance $3654 m0 *1 46.74,57.4
X$3654 23 38 FILLCELL_X1
* cell instance $3655 m0 *1 43.51,57.4
X$3655 23 2795 1491 1523 1404 38 DFF_X1
* cell instance $3656 m0 *1 46.93,57.4
X$3656 1405 1403 1490 23 38 1439 MUX2_X1
* cell instance $3657 m0 *1 48.26,57.4
X$3657 1455 1289 1490 23 38 1477 MUX2_X1
* cell instance $3658 m0 *1 49.59,57.4
X$3658 1214 38 1488 23 BUF_X4
* cell instance $3659 m0 *1 50.92,57.4
X$3659 23 38 FILLCELL_X4
* cell instance $3660 m0 *1 51.68,57.4
X$3660 23 38 FILLCELL_X2
* cell instance $3661 r0 *1 44.65,57.4
X$3661 23 38 FILLCELL_X1
* cell instance $3662 r0 *1 44.84,57.4
X$3662 1536 1434 1490 23 38 1554 MUX2_X1
* cell instance $3663 r0 *1 46.17,57.4
X$3663 1491 1446 1490 23 38 1523 MUX2_X1
* cell instance $3664 r0 *1 47.5,57.4
X$3664 1130 38 1446 23 BUF_X4
* cell instance $3665 r0 *1 48.83,57.4
X$3665 23 38 FILLCELL_X4
* cell instance $3666 r0 *1 49.59,57.4
X$3666 1490 1492 1525 23 38 1553 MUX2_X1
* cell instance $3667 r0 *1 50.92,57.4
X$3667 23 38 FILLCELL_X2
* cell instance $3668 r0 *1 51.3,57.4
X$3668 23 38 FILLCELL_X1
* cell instance $3669 r0 *1 51.49,57.4
X$3669 863 38 1544 23 BUF_X4
* cell instance $3670 m0 *1 53.39,57.4
X$3670 23 38 FILLCELL_X4
* cell instance $3671 m0 *1 52.06,57.4
X$3671 796 38 1492 23 BUF_X4
* cell instance $3672 m0 *1 54.15,57.4
X$3672 23 38 FILLCELL_X2
* cell instance $3673 r0 *1 52.82,57.4
X$3673 23 38 FILLCELL_X4
* cell instance $3674 r0 *1 53.58,57.4
X$3674 23 38 FILLCELL_X1
* cell instance $3675 r0 *1 53.77,57.4
X$3675 821 38 1482 23 BUF_X4
* cell instance $3676 m0 *1 57,57.4
X$3676 138 38 1493 23 BUF_X4
* cell instance $3677 m0 *1 54.53,57.4
X$3677 23 1511 38 1300 BUF_X8
* cell instance $3678 m0 *1 58.33,57.4
X$3678 1494 23 38 1407 INV_X1
* cell instance $3679 m0 *1 58.71,57.4
X$3679 1457 1456 23 138 38 NAND2_X4
* cell instance $3680 m0 *1 60.42,57.4
X$3680 23 38 FILLCELL_X1
* cell instance $3681 m0 *1 60.61,57.4
X$3681 1528 23 38 1214 BUF_X2
* cell instance $3682 m0 *1 61.37,57.4
X$3682 1496 1444 38 23 1528 AND2_X1
* cell instance $3683 m0 *1 62.13,57.4
X$3683 23 38 FILLCELL_X1
* cell instance $3684 m0 *1 62.32,57.4
X$3684 1457 1496 23 38 796 NAND2_X2
* cell instance $3685 m0 *1 63.27,57.4
X$3685 1458 1411 23 243 38 NAND2_X4
* cell instance $3686 m0 *1 64.98,57.4
X$3686 23 38 FILLCELL_X2
* cell instance $3687 r0 *1 55.1,57.4
X$3687 23 38 FILLCELL_X2
* cell instance $3688 r0 *1 55.48,57.4
X$3688 68 38 1480 23 BUF_X4
* cell instance $3689 r0 *1 56.81,57.4
X$3689 243 38 1346 23 BUF_X4
* cell instance $3690 r0 *1 58.14,57.4
X$3690 1407 38 403 23 BUF_X4
* cell instance $3691 r0 *1 59.14,57.4
X$3691 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $3692 r0 *1 59.14,57.4
X$3692 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $3693 r0 *1 59.14,57.4
X$3693 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $3694 r0 *1 59.47,57.4
X$3694 23 38 FILLCELL_X1
* cell instance $3695 r0 *1 59.66,57.4
X$3695 1457 1495 23 38 863 NAND2_X2
* cell instance $3696 r0 *1 60.61,57.4
X$3696 1495 1444 38 23 1410 AND2_X1
* cell instance $3697 r0 *1 61.37,57.4
X$3697 1496 1442 38 23 1529 AND2_X1
* cell instance $3698 r0 *1 62.13,57.4
X$3698 1529 23 38 1175 BUF_X2
* cell instance $3699 r0 *1 62.89,57.4
X$3699 1456 1444 38 23 1412 AND2_X1
* cell instance $3700 r0 *1 63.65,57.4
X$3700 1458 1495 23 38 821 NAND2_X2
* cell instance $3701 r0 *1 64.6,57.4
X$3701 1458 1456 23 68 38 NAND2_X4
* cell instance $3702 m0 *1 65.55,57.4
X$3702 23 2568 1413 1476 1301 38 DFF_X1
* cell instance $3703 m0 *1 65.36,57.4
X$3703 23 38 FILLCELL_X1
* cell instance $3704 m0 *1 68.78,57.4
X$3704 1413 1373 1372 23 38 1527 MUX2_X1
* cell instance $3705 m0 *1 70.11,57.4
X$3705 1527 177 23 38 1562 NOR2_X1
* cell instance $3706 m0 *1 70.68,57.4
X$3706 23 38 FILLCELL_X4
* cell instance $3707 m0 *1 71.44,57.4
X$3707 23 38 FILLCELL_X2
* cell instance $3708 r0 *1 66.31,57.4
X$3708 23 38 FILLCELL_X32
* cell instance $3709 m0 *1 72.01,57.4
X$3709 23 2831 1459 1526 1336 38 DFF_X1
* cell instance $3710 m0 *1 71.82,57.4
X$3710 23 38 FILLCELL_X1
* cell instance $3711 m0 *1 75.24,57.4
X$3711 1478 23 38 1460 CLKBUF_X3
* cell instance $3712 m0 *1 76.19,57.4
X$3712 23 38 FILLCELL_X8
* cell instance $3713 m0 *1 77.71,57.4
X$3713 23 38 FILLCELL_X2
* cell instance $3714 r0 *1 72.39,57.4
X$3714 23 38 FILLCELL_X2
* cell instance $3715 r0 *1 72.77,57.4
X$3715 1497 51 1459 23 38 1526 MUX2_X1
* cell instance $3716 r0 *1 74.1,57.4
X$3716 23 38 FILLCELL_X4
* cell instance $3717 r0 *1 74.86,57.4
X$3717 23 38 FILLCELL_X2
* cell instance $3718 r0 *1 75.24,57.4
X$3718 1459 1099 1498 23 38 1499 MUX2_X1
* cell instance $3719 r0 *1 77.9,57.4
X$3719 1499 372 23 38 1539 NOR2_X1
* cell instance $3720 m0 *1 78.66,57.4
X$3720 23 38 FILLCELL_X4
* cell instance $3721 m0 *1 78.09,57.4
X$3721 1524 177 23 38 1471 NOR2_X1
* cell instance $3722 m0 *1 79.42,57.4
X$3722 23 38 FILLCELL_X2
* cell instance $3723 r0 *1 78.47,57.4
X$3723 23 38 FILLCELL_X16
* cell instance $3724 m0 *1 79.99,57.4
X$3724 1332 1520 1375 1319 1521 38 23 1473 OAI221_X1
* cell instance $3725 m0 *1 79.8,57.4
X$3725 23 38 FILLCELL_X1
* cell instance $3726 m0 *1 81.13,57.4
X$3726 1460 1377 23 38 1520 NAND2_X1
* cell instance $3727 m0 *1 81.7,57.4
X$3727 1377 1519 23 38 1521 NAND2_X1
* cell instance $3728 m0 *1 82.27,57.4
X$3728 23 38 FILLCELL_X16
* cell instance $3729 m0 *1 85.31,57.4
X$3729 23 38 FILLCELL_X2
* cell instance $3730 r0 *1 81.51,57.4
X$3730 23 38 FILLCELL_X4
* cell instance $3731 r0 *1 82.27,57.4
X$3731 23 38 FILLCELL_X2
* cell instance $3732 r0 *1 82.65,57.4
X$3732 23 38 FILLCELL_X1
* cell instance $3733 r0 *1 82.84,57.4
X$3733 1073 23 38 1497 CLKBUF_X2
* cell instance $3734 r0 *1 83.6,57.4
X$3734 23 38 FILLCELL_X32
* cell instance $3735 m0 *1 85.88,57.4
X$3735 1225 1518 1418 1226 1516 38 23 1472 OAI221_X1
* cell instance $3736 m0 *1 85.69,57.4
X$3736 23 38 FILLCELL_X1
* cell instance $3737 m0 *1 87.02,57.4
X$3737 1228 1419 23 38 1518 NAND2_X1
* cell instance $3738 m0 *1 87.59,57.4
X$3738 1419 1239 23 38 1516 NAND2_X1
* cell instance $3739 m0 *1 88.16,57.4
X$3739 23 38 FILLCELL_X4
* cell instance $3740 m0 *1 88.92,57.4
X$3740 23 38 FILLCELL_X2
* cell instance $3741 m0 *1 89.49,57.4
X$3741 1146 748 1304 1305 38 23 1500 OAI22_X1
* cell instance $3742 m0 *1 89.3,57.4
X$3742 23 38 FILLCELL_X1
* cell instance $3743 m0 *1 90.44,57.4
X$3743 1146 748 1241 1506 1224 38 23 1461 OAI221_X1
* cell instance $3744 m0 *1 91.58,57.4
X$3744 23 38 FILLCELL_X1
* cell instance $3745 m0 *1 91.77,57.4
X$3745 1154 914 1241 1506 1224 38 23 1462 OAI221_X1
* cell instance $3746 m0 *1 92.91,57.4
X$3746 23 38 FILLCELL_X1
* cell instance $3747 m0 *1 93.1,57.4
X$3747 1306 1503 1463 38 1469 23 OAI21_X1
* cell instance $3748 m0 *1 93.86,57.4
X$3748 23 38 FILLCELL_X1
* cell instance $3749 m0 *1 94.05,57.4
X$3749 1502 1230 23 38 1503 NAND2_X1
* cell instance $3750 m0 *1 94.62,57.4
X$3750 23 38 FILLCELL_X1
* cell instance $3751 m0 *1 94.81,57.4
X$3751 1306 1542 1500 38 1470 23 OAI21_X1
* cell instance $3752 m0 *1 95.57,57.4
X$3752 1469 23 38 1466 BUF_X1
* cell instance $3753 m0 *1 96.14,57.4
X$3753 23 38 FILLCELL_X2
* cell instance $3754 r0 *1 89.68,57.4
X$3754 23 38 FILLCELL_X4
* cell instance $3755 r0 *1 90.44,57.4
X$3755 23 38 FILLCELL_X1
* cell instance $3756 r0 *1 90.63,57.4
X$3756 1227 23 38 3150 INV_X1
* cell instance $3757 r0 *1 91.01,57.4
X$3757 1392 23 38 1227 CLKBUF_X3
* cell instance $3758 r0 *1 91.96,57.4
X$3758 23 3037 1502 1541 1227 38 DFF_X1
* cell instance $3759 r0 *1 95.19,57.4
X$3759 23 38 FILLCELL_X8
* cell instance $3760 r180 *1 97.28,57.4
X$3760 23 38 23 38 TAPCELL_X1
* cell instance $3761 m0 *1 96.52,57.4
X$3761 1306 23 38 1465 BUF_X1
* cell instance $3762 r0 *1 96.71,57.4
X$3762 23 38 FILLCELL_X2
* cell instance $3763 m90 *1 97.28,57.4
X$3763 23 38 23 38 TAPCELL_X1
* cell instance $3764 r0 *1 10.26,1.4
X$3764 23 38 FILLCELL_X8
* cell instance $3765 r0 *1 11.78,1.4
X$3765 23 38 FILLCELL_X2
* cell instance $3766 r0 *1 37.81,1.4
X$3766 23 38 FILLCELL_X1
* cell instance $3767 r0 *1 38.76,1.4
X$3767 23 38 FILLCELL_X32
* cell instance $3768 r0 *1 44.84,1.4
X$3768 23 38 FILLCELL_X2
* cell instance $3769 r0 *1 53.77,1.4
X$3769 23 38 FILLCELL_X1
* cell instance $3770 r0 *1 54.72,1.4
X$3770 23 38 FILLCELL_X16
* cell instance $3771 r0 *1 57.76,1.4
X$3771 23 38 FILLCELL_X8
* cell instance $3772 r0 *1 59.28,1.4
X$3772 23 38 FILLCELL_X1
* cell instance $3773 r0 *1 60.23,1.4
X$3773 23 38 FILLCELL_X32
* cell instance $3774 r0 *1 66.31,1.4
X$3774 23 38 FILLCELL_X4
* cell instance $3775 r0 *1 67.07,1.4
X$3775 23 38 FILLCELL_X2
* cell instance $3776 r0 *1 59.14,1.4
X$3776 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $3777 r0 *1 59.14,1.4
X$3777 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $3778 r0 *1 59.14,1.4
X$3778 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $3779 r0 *1 51.68,1.4
X$3779 23 38 FILLCELL_X1
* cell instance $3780 r0 *1 52.63,1.4
X$3780 23 38 FILLCELL_X4
* cell instance $3781 r0 *1 53.39,1.4
X$3781 23 38 FILLCELL_X2
* cell instance $3782 r0 *1 32.68,1.4
X$3782 23 38 FILLCELL_X1
* cell instance $3783 r0 *1 33.63,1.4
X$3783 23 38 FILLCELL_X16
* cell instance $3784 r0 *1 36.67,1.4
X$3784 23 38 FILLCELL_X4
* cell instance $3785 r0 *1 37.43,1.4
X$3785 23 38 FILLCELL_X2
* cell instance $3786 m0 *1 1.33,26.6
X$3786 23 38 FILLCELL_X1
* cell instance $3787 m0 *1 1.14,26.6
X$3787 23 38 23 38 TAPCELL_X1
* cell instance $3788 m0 *1 1.52,26.6
X$3788 625 23 38 107 BUF_X2
* cell instance $3789 m0 *1 2.28,26.6
X$3789 626 23 38 154 CLKBUF_X2
* cell instance $3790 m0 *1 3.04,26.6
X$3790 23 38 FILLCELL_X2
* cell instance $3791 r0 *1 1.14,26.6
X$3791 23 38 23 38 TAPCELL_X1
* cell instance $3792 r0 *1 1.33,26.6
X$3792 23 38 FILLCELL_X8
* cell instance $3793 r0 *1 2.85,26.6
X$3793 23 38 FILLCELL_X4
* cell instance $3794 r0 *1 3.14,26.6
X$3794 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $3795 r0 *1 3.14,26.6
X$3795 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $3796 r0 *1 3.14,26.6
X$3796 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $3797 m0 *1 6.65,26.6
X$3797 23 38 FILLCELL_X16
* cell instance $3798 m0 *1 3.42,26.6
X$3798 23 2763 590 589 660 38 DFF_X1
* cell instance $3799 m0 *1 9.69,26.6
X$3799 23 38 FILLCELL_X8
* cell instance $3800 m0 *1 11.21,26.6
X$3800 23 38 FILLCELL_X2
* cell instance $3801 r0 *1 3.61,26.6
X$3801 23 38 FILLCELL_X2
* cell instance $3802 r0 *1 3.99,26.6
X$3802 154 659 691 23 38 677 MUX2_X1
* cell instance $3803 r0 *1 5.32,26.6
X$3803 107 23 38 502 BUF_X2
* cell instance $3804 r0 *1 6.08,26.6
X$3804 23 38 FILLCELL_X4
* cell instance $3805 r0 *1 6.84,26.6
X$3805 23 38 FILLCELL_X2
* cell instance $3806 r0 *1 7.22,26.6
X$3806 23 38 FILLCELL_X1
* cell instance $3807 r0 *1 7.41,26.6
X$3807 154 23 38 591 BUF_X2
* cell instance $3808 r0 *1 8.17,26.6
X$3808 23 38 FILLCELL_X1
* cell instance $3809 r0 *1 8.36,26.6
X$3809 27 659 692 23 38 679 MUX2_X1
* cell instance $3810 r0 *1 9.69,26.6
X$3810 24 659 661 23 38 681 MUX2_X1
* cell instance $3811 r0 *1 11.02,26.6
X$3811 23 38 FILLCELL_X8
* cell instance $3812 m0 *1 11.78,26.6
X$3812 593 627 592 23 38 595 MUX2_X1
* cell instance $3813 m0 *1 11.59,26.6
X$3813 23 38 FILLCELL_X1
* cell instance $3814 m0 *1 13.11,26.6
X$3814 23 38 FILLCELL_X16
* cell instance $3815 m0 *1 16.15,26.6
X$3815 23 38 FILLCELL_X8
* cell instance $3816 m0 *1 17.67,26.6
X$3816 24 23 38 453 BUF_X2
* cell instance $3817 m0 *1 18.43,26.6
X$3817 453 628 629 23 38 652 MUX2_X1
* cell instance $3818 m0 *1 19.76,26.6
X$3818 23 38 FILLCELL_X8
* cell instance $3819 m0 *1 21.28,26.6
X$3819 23 38 FILLCELL_X2
* cell instance $3820 r0 *1 12.54,26.6
X$3820 23 38 FILLCELL_X4
* cell instance $3821 r0 *1 13.3,26.6
X$3821 23 38 FILLCELL_X2
* cell instance $3822 r0 *1 13.68,26.6
X$3822 23 38 FILLCELL_X1
* cell instance $3823 r0 *1 13.87,26.6
X$3823 154 632 695 23 38 719 MUX2_X1
* cell instance $3824 r0 *1 15.2,26.6
X$3824 23 38 FILLCELL_X8
* cell instance $3825 r0 *1 16.72,26.6
X$3825 23 38 FILLCELL_X4
* cell instance $3826 r0 *1 17.48,26.6
X$3826 23 38 FILLCELL_X1
* cell instance $3827 r0 *1 17.67,26.6
X$3827 23 3013 629 652 653 38 DFF_X1
* cell instance $3828 r0 *1 20.9,26.6
X$3828 23 38 FILLCELL_X2
* cell instance $3829 r0 *1 21.28,26.6
X$3829 23 3010 631 630 653 38 DFF_X1
* cell instance $3830 m0 *1 21.85,26.6
X$3830 358 628 631 23 38 630 MUX2_X1
* cell instance $3831 m0 *1 21.66,26.6
X$3831 23 38 FILLCELL_X1
* cell instance $3832 m0 *1 23.18,26.6
X$3832 23 2806 685 684 653 38 DFF_X1
* cell instance $3833 m0 *1 26.41,26.6
X$3833 23 38 FILLCELL_X8
* cell instance $3834 m0 *1 27.93,26.6
X$3834 23 38 FILLCELL_X4
* cell instance $3835 m0 *1 28.69,26.6
X$3835 23 38 FILLCELL_X1
* cell instance $3836 m0 *1 28.88,26.6
X$3836 29 23 38 421 BUF_X2
* cell instance $3837 m0 *1 29.64,26.6
X$3837 23 38 FILLCELL_X16
* cell instance $3838 m0 *1 32.68,26.6
X$3838 634 38 305 23 BUF_X4
* cell instance $3839 m0 *1 34.01,26.6
X$3839 23 2843 688 633 655 38 DFF_X1
* cell instance $3840 m0 *1 37.24,26.6
X$3840 23 38 FILLCELL_X16
* cell instance $3841 m0 *1 40.28,26.6
X$3841 23 38 FILLCELL_X8
* cell instance $3842 m0 *1 41.8,26.6
X$3842 23 38 FILLCELL_X4
* cell instance $3843 m0 *1 42.56,26.6
X$3843 23 38 FILLCELL_X1
* cell instance $3844 m0 *1 42.75,26.6
X$3844 23 2735 637 635 636 38 DFF_X1
* cell instance $3845 m0 *1 45.98,26.6
X$3845 23 38 FILLCELL_X4
* cell instance $3846 m0 *1 46.74,26.6
X$3846 23 38 FILLCELL_X2
* cell instance $3847 r0 *1 24.51,26.6
X$3847 26 632 685 23 38 684 MUX2_X1
* cell instance $3848 r0 *1 25.84,26.6
X$3848 634 38 412 23 BUF_X4
* cell instance $3849 r0 *1 27.17,26.6
X$3849 23 38 FILLCELL_X2
* cell instance $3850 r0 *1 27.55,26.6
X$3850 23 38 FILLCELL_X1
* cell instance $3851 r0 *1 27.74,26.6
X$3851 23 3058 686 662 329 38 DFF_X1
* cell instance $3852 r0 *1 30.97,26.6
X$3852 23 3053 725 663 655 38 DFF_X1
* cell instance $3853 r0 *1 34.2,26.6
X$3853 25 632 688 23 38 633 MUX2_X1
* cell instance $3854 r0 *1 35.53,26.6
X$3854 23 38 FILLCELL_X16
* cell instance $3855 r0 *1 38.57,26.6
X$3855 23 38 FILLCELL_X8
* cell instance $3856 r0 *1 40.09,26.6
X$3856 23 38 FILLCELL_X2
* cell instance $3857 r0 *1 40.47,26.6
X$3857 23 38 FILLCELL_X1
* cell instance $3858 r0 *1 40.66,26.6
X$3858 634 38 144 23 BUF_X4
* cell instance $3859 r0 *1 41.99,26.6
X$3859 23 38 FILLCELL_X2
* cell instance $3860 r0 *1 42.37,26.6
X$3860 23 38 FILLCELL_X1
* cell instance $3861 r0 *1 42.56,26.6
X$3861 75 632 637 23 38 635 MUX2_X1
* cell instance $3862 r0 *1 43.89,26.6
X$3862 23 3047 665 664 636 38 DFF_X1
* cell instance $3863 m0 *1 47.31,26.6
X$3863 620 38 627 23 BUF_X4
* cell instance $3864 m0 *1 47.12,26.6
X$3864 23 38 FILLCELL_X1
* cell instance $3865 m0 *1 48.64,26.6
X$3865 23 38 FILLCELL_X32
* cell instance $3866 m0 *1 54.72,26.6
X$3866 23 38 FILLCELL_X1
* cell instance $3867 m0 *1 54.91,26.6
X$3867 23 2752 638 658 666 38 DFF_X1
* cell instance $3868 m0 *1 58.14,26.6
X$3868 638 597 640 23 38 658 MUX2_X1
* cell instance $3869 m0 *1 59.47,26.6
X$3869 23 38 FILLCELL_X8
* cell instance $3870 m0 *1 60.99,26.6
X$3870 23 38 FILLCELL_X4
* cell instance $3871 m0 *1 61.75,26.6
X$3871 23 38 FILLCELL_X1
* cell instance $3872 m0 *1 61.94,26.6
X$3872 641 599 640 23 38 657 MUX2_X1
* cell instance $3873 m0 *1 63.27,26.6
X$3873 23 2732 641 657 543 38 DFF_X1
* cell instance $3874 m0 *1 66.5,26.6
X$3874 139 23 38 543 CLKBUF_X3
* cell instance $3875 m0 *1 67.45,26.6
X$3875 23 38 FILLCELL_X16
* cell instance $3876 m0 *1 70.49,26.6
X$3876 23 38 FILLCELL_X4
* cell instance $3877 m0 *1 71.25,26.6
X$3877 23 2723 606 605 445 38 DFF_X1
* cell instance $3878 m0 *1 74.48,26.6
X$3878 642 520 524 23 38 654 MUX2_X1
* cell instance $3879 m0 *1 75.81,26.6
X$3879 23 38 FILLCELL_X32
* cell instance $3880 m0 *1 81.89,26.6
X$3880 23 38 FILLCELL_X8
* cell instance $3881 m0 *1 83.41,26.6
X$3881 651 88 524 23 38 643 MUX2_X1
* cell instance $3882 m0 *1 84.74,26.6
X$3882 23 38 FILLCELL_X2
* cell instance $3883 r0 *1 47.12,26.6
X$3883 23 38 FILLCELL_X2
* cell instance $3884 r0 *1 47.5,26.6
X$3884 634 38 80 23 BUF_X4
* cell instance $3885 r0 *1 48.83,26.6
X$3885 23 38 FILLCELL_X1
* cell instance $3886 r0 *1 49.02,26.6
X$3886 23 3120 667 689 666 38 DFF_X1
* cell instance $3887 r0 *1 52.25,26.6
X$3887 23 38 FILLCELL_X8
* cell instance $3888 r0 *1 53.77,26.6
X$3888 23 38 FILLCELL_X4
* cell instance $3889 r0 *1 54.53,26.6
X$3889 23 3033 669 687 666 38 DFF_X1
* cell instance $3890 r0 *1 57.76,26.6
X$3890 638 305 669 23 38 639 MUX2_X1
* cell instance $3891 r0 *1 59.14,26.6
X$3891 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $3892 r0 *1 59.14,26.6
X$3892 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $3893 r0 *1 59.14,26.6
X$3893 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $3894 r0 *1 59.09,26.6
X$3894 669 557 640 23 38 687 MUX2_X1
* cell instance $3895 r0 *1 60.42,26.6
X$3895 671 598 640 23 38 670 MUX2_X1
* cell instance $3896 r0 *1 61.75,26.6
X$3896 671 438 641 23 38 656 MUX2_X1
* cell instance $3897 r0 *1 63.08,26.6
X$3897 23 38 FILLCELL_X32
* cell instance $3898 r0 *1 69.16,26.6
X$3898 23 38 FILLCELL_X16
* cell instance $3899 r0 *1 72.2,26.6
X$3899 23 2924 642 654 705 38 DFF_X1
* cell instance $3900 r0 *1 75.43,26.6
X$3900 23 38 FILLCELL_X8
* cell instance $3901 r0 *1 76.95,26.6
X$3901 23 38 FILLCELL_X2
* cell instance $3902 r0 *1 77.33,26.6
X$3902 23 38 FILLCELL_X1
* cell instance $3903 r0 *1 77.52,26.6
X$3903 23 2936 682 683 673 38 DFF_X1
* cell instance $3904 r0 *1 80.75,26.6
X$3904 23 38 FILLCELL_X8
* cell instance $3905 r0 *1 82.27,26.6
X$3905 23 38 FILLCELL_X4
* cell instance $3906 r0 *1 83.03,26.6
X$3906 23 38 FILLCELL_X2
* cell instance $3907 r0 *1 83.41,26.6
X$3907 23 38 FILLCELL_X1
* cell instance $3908 r0 *1 83.6,26.6
X$3908 23 2871 651 643 673 38 DFF_X1
* cell instance $3909 m0 *1 85.31,26.6
X$3909 651 724 644 23 38 650 MUX2_X1
* cell instance $3910 m0 *1 85.12,26.6
X$3910 23 38 FILLCELL_X1
* cell instance $3911 m0 *1 86.64,26.6
X$3911 644 130 524 23 38 645 MUX2_X1
* cell instance $3912 m0 *1 87.97,26.6
X$3912 23 38 FILLCELL_X8
* cell instance $3913 m0 *1 89.49,26.6
X$3913 23 38 FILLCELL_X1
* cell instance $3914 m0 *1 89.68,26.6
X$3914 23 2790 680 648 647 38 DFF_X1
* cell instance $3915 m0 *1 92.91,26.6
X$3915 23 38 FILLCELL_X2
* cell instance $3916 r0 *1 86.83,26.6
X$3916 23 38 FILLCELL_X2
* cell instance $3917 r0 *1 87.21,26.6
X$3917 23 2859 644 645 673 38 DFF_X1
* cell instance $3918 r0 *1 90.44,26.6
X$3918 23 38 FILLCELL_X4
* cell instance $3919 r0 *1 91.2,26.6
X$3919 675 191 680 23 38 648 MUX2_X1
* cell instance $3920 r0 *1 92.53,26.6
X$3920 23 38 FILLCELL_X4
* cell instance $3921 m0 *1 93.48,26.6
X$3921 23 2825 646 676 647 38 DFF_X1
* cell instance $3922 m0 *1 93.29,26.6
X$3922 23 38 FILLCELL_X1
* cell instance $3923 m0 *1 96.71,26.6
X$3923 23 38 FILLCELL_X2
* cell instance $3924 r0 *1 93.29,26.6
X$3924 680 263 646 23 38 678 MUX2_X1
* cell instance $3925 r0 *1 94.62,26.6
X$3925 23 38 FILLCELL_X4
* cell instance $3926 r0 *1 95.38,26.6
X$3926 675 187 646 23 38 676 MUX2_X1
* cell instance $3927 r0 *1 96.71,26.6
X$3927 23 38 FILLCELL_X2
* cell instance $3928 m0 *1 1.33,35
X$3928 23 38 FILLCELL_X1
* cell instance $3929 m0 *1 1.14,35
X$3929 23 38 23 38 TAPCELL_X1
* cell instance $3930 m0 *1 1.52,35
X$3930 23 2769 790 807 789 38 DFF_X1
* cell instance $3931 m0 *1 4.75,35
X$3931 23 38 FILLCELL_X1
* cell instance $3932 m0 *1 4.94,35
X$3932 23 2764 825 808 789 38 DFF_X1
* cell instance $3933 m0 *1 8.17,35
X$3933 23 38 FILLCELL_X1
* cell instance $3934 m0 *1 8.36,35
X$3934 23 2767 810 809 789 38 DFF_X1
* cell instance $3935 m0 *1 11.59,35
X$3935 23 38 FILLCELL_X1
* cell instance $3936 m0 *1 11.78,35
X$3936 23 2693 826 874 660 38 DFF_X1
* cell instance $3937 m0 *1 15.01,35
X$3937 812 792 694 23 38 849 MUX2_X1
* cell instance $3938 m0 *1 16.34,35
X$3938 502 628 791 23 38 781 MUX2_X1
* cell instance $3939 m0 *1 17.67,35
X$3939 791 792 733 23 38 827 MUX2_X1
* cell instance $3940 m0 *1 19,35
X$3940 23 38 FILLCELL_X16
* cell instance $3941 m0 *1 22.04,35
X$3941 23 38 FILLCELL_X4
* cell instance $3942 m0 *1 22.8,35
X$3942 23 38 FILLCELL_X2
* cell instance $3943 r0 *1 1.14,35
X$3943 23 38 23 38 TAPCELL_X1
* cell instance $3944 r0 *1 1.33,35
X$3944 23 38 FILLCELL_X8
* cell instance $3945 r0 *1 2.85,35
X$3945 23 38 FILLCELL_X4
* cell instance $3946 r0 *1 3.14,35
X$3946 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $3947 r0 *1 3.14,35
X$3947 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $3948 r0 *1 3.14,35
X$3948 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $3949 r0 *1 3.61,35
X$3949 23 38 FILLCELL_X2
* cell instance $3950 r0 *1 3.99,35
X$3950 591 762 845 23 38 870 MUX2_X1
* cell instance $3951 r0 *1 5.32,35
X$3951 23 38 FILLCELL_X8
* cell instance $3952 r0 *1 6.84,35
X$3952 790 813 732 23 38 871 MUX2_X1
* cell instance $3953 r0 *1 8.17,35
X$3953 23 38 FILLCELL_X1
* cell instance $3954 r0 *1 8.36,35
X$3954 825 813 692 23 38 873 MUX2_X1
* cell instance $3955 r0 *1 9.69,35
X$3955 23 38 FILLCELL_X4
* cell instance $3956 r0 *1 10.45,35
X$3956 23 38 FILLCELL_X1
* cell instance $3957 r0 *1 10.64,35
X$3957 810 813 661 23 38 875 MUX2_X1
* cell instance $3958 r0 *1 11.97,35
X$3958 23 38 FILLCELL_X4
* cell instance $3959 r0 *1 12.73,35
X$3959 295 628 812 23 38 847 MUX2_X1
* cell instance $3960 r0 *1 14.06,35
X$3960 591 628 826 23 38 874 MUX2_X1
* cell instance $3961 r0 *1 15.39,35
X$3961 23 38 FILLCELL_X2
* cell instance $3962 r0 *1 15.77,35
X$3962 826 792 695 23 38 857 MUX2_X1
* cell instance $3963 r0 *1 17.1,35
X$3963 23 38 FILLCELL_X2
* cell instance $3964 r0 *1 17.48,35
X$3964 849 829 23 38 889 NOR2_X1
* cell instance $3965 r0 *1 18.05,35
X$3965 23 38 FILLCELL_X8
* cell instance $3966 r0 *1 19.57,35
X$3966 851 858 358 23 38 879 MUX2_X1
* cell instance $3967 r0 *1 20.9,35
X$3967 23 3012 851 879 763 38 DFF_X1
* cell instance $3968 m0 *1 23.37,35
X$3968 358 762 764 23 38 782 MUX2_X1
* cell instance $3969 m0 *1 23.18,35
X$3969 23 38 FILLCELL_X1
* cell instance $3970 m0 *1 24.7,35
X$3970 764 813 697 23 38 852 MUX2_X1
* cell instance $3971 m0 *1 26.03,35
X$3971 23 38 FILLCELL_X1
* cell instance $3972 m0 *1 26.22,35
X$3972 421 762 793 23 38 815 MUX2_X1
* cell instance $3973 m0 *1 27.55,35
X$3973 23 2731 793 815 763 38 DFF_X1
* cell instance $3974 m0 *1 30.78,35
X$3974 793 144 735 23 38 830 MUX2_X1
* cell instance $3975 m0 *1 32.11,35
X$3975 23 38 FILLCELL_X1
* cell instance $3976 m0 *1 32.3,35
X$3976 510 762 767 23 38 766 MUX2_X1
* cell instance $3977 m0 *1 33.63,35
X$3977 23 38 FILLCELL_X1
* cell instance $3978 m0 *1 33.82,35
X$3978 767 144 699 23 38 832 MUX2_X1
* cell instance $3979 m0 *1 35.15,35
X$3979 23 38 FILLCELL_X2
* cell instance $3980 r0 *1 24.13,35
X$3980 23 38 FILLCELL_X8
* cell instance $3981 r0 *1 25.65,35
X$3981 23 38 FILLCELL_X4
* cell instance $3982 r0 *1 26.41,35
X$3982 693 23 38 763 CLKBUF_X3
* cell instance $3983 r0 *1 27.36,35
X$3983 763 23 38 CLKBUF_X1
* cell instance $3984 r0 *1 27.93,35
X$3984 23 38 FILLCELL_X16
* cell instance $3985 r0 *1 30.97,35
X$3985 23 38 FILLCELL_X1
* cell instance $3986 r0 *1 31.16,35
X$3986 828 829 23 38 993 NOR2_X1
* cell instance $3987 r0 *1 31.73,35
X$3987 830 831 23 38 1023 NOR2_X1
* cell instance $3988 r0 *1 32.3,35
X$3988 23 38 FILLCELL_X8
* cell instance $3989 r0 *1 33.82,35
X$3989 23 38 FILLCELL_X4
* cell instance $3990 r0 *1 34.58,35
X$3990 23 38 FILLCELL_X1
* cell instance $3991 r0 *1 34.77,35
X$3991 832 831 23 38 946 NOR2_X1
* cell instance $3992 r0 *1 35.34,35
X$3992 700 829 23 38 859 NOR2_X1
* cell instance $3993 m0 *1 38.76,35
X$3993 23 38 FILLCELL_X16
* cell instance $3994 m0 *1 35.53,35
X$3994 23 2846 833 817 655 38 DFF_X1
* cell instance $3995 m0 *1 41.8,35
X$3995 23 38 FILLCELL_X8
* cell instance $3996 m0 *1 43.32,35
X$3996 23 38 FILLCELL_X2
* cell instance $3997 r0 *1 35.91,35
X$3997 23 38 FILLCELL_X2
* cell instance $3998 r0 *1 36.29,35
X$3998 319 762 833 23 38 817 MUX2_X1
* cell instance $3999 r0 *1 37.62,35
X$3999 833 144 768 23 38 1053 MUX2_X1
* cell instance $4000 r0 *1 38.95,35
X$4000 23 38 FILLCELL_X4
* cell instance $4001 r0 *1 39.71,35
X$4001 23 38 FILLCELL_X2
* cell instance $4002 r0 *1 40.09,35
X$4002 834 858 398 23 38 860 MUX2_X1
* cell instance $4003 r0 *1 41.42,35
X$4003 23 38 FILLCELL_X8
* cell instance $4004 r0 *1 42.94,35
X$4004 23 38 FILLCELL_X2
* cell instance $4005 r0 *1 43.32,35
X$4005 23 3049 836 835 636 38 DFF_X1
* cell instance $4006 m0 *1 43.89,35
X$4006 693 23 38 636 CLKBUF_X3
* cell instance $4007 m0 *1 43.7,35
X$4007 23 38 FILLCELL_X1
* cell instance $4008 m0 *1 44.84,35
X$4008 23 38 FILLCELL_X16
* cell instance $4009 m0 *1 47.88,35
X$4009 23 38 FILLCELL_X1
* cell instance $4010 m0 *1 48.07,35
X$4010 301 762 820 23 38 838 MUX2_X1
* cell instance $4011 m0 *1 49.4,35
X$4011 23 38 FILLCELL_X4
* cell instance $4012 m0 *1 50.16,35
X$4012 23 38 FILLCELL_X1
* cell instance $4013 m0 *1 50.35,35
X$4013 796 23 38 628 CLKBUF_X3
* cell instance $4014 m0 *1 51.3,35
X$4014 820 144 738 23 38 795 MUX2_X1
* cell instance $4015 m0 *1 52.63,35
X$4015 23 38 FILLCELL_X4
* cell instance $4016 m0 *1 53.39,35
X$4016 23 38 FILLCELL_X2
* cell instance $4017 r0 *1 46.55,35
X$4017 23 38 FILLCELL_X8
* cell instance $4018 r0 *1 48.07,35
X$4018 23 38 FILLCELL_X1
* cell instance $4019 r0 *1 48.26,35
X$4019 23 3097 820 838 839 38 DFF_X1
* cell instance $4020 r0 *1 51.49,35
X$4020 23 38 FILLCELL_X4
* cell instance $4021 r0 *1 52.25,35
X$4021 23 38 FILLCELL_X1
* cell instance $4022 r0 *1 52.44,35
X$4022 702 261 23 38 861 NOR2_X1
* cell instance $4023 r0 *1 53.01,35
X$4023 23 38 FILLCELL_X4
* cell instance $4024 r0 *1 53.77,35
X$4024 23 38 FILLCELL_X1
* cell instance $4025 m0 *1 53.96,35
X$4025 556 796 797 23 38 822 MUX2_X1
* cell instance $4026 m0 *1 53.77,35
X$4026 23 38 FILLCELL_X1
* cell instance $4027 m0 *1 55.29,35
X$4027 797 602 772 23 38 823 MUX2_X1
* cell instance $4028 m0 *1 56.62,35
X$4028 823 261 23 38 798 NOR2_X1
* cell instance $4029 m0 *1 57.19,35
X$4029 23 38 FILLCELL_X4
* cell instance $4030 m0 *1 57.95,35
X$4030 23 2813 773 824 666 38 DFF_X1
* cell instance $4031 m0 *1 61.18,35
X$4031 774 602 773 23 38 855 MUX2_X1
* cell instance $4032 m0 *1 62.51,35
X$4032 23 38 FILLCELL_X8
* cell instance $4033 m0 *1 64.03,35
X$4033 23 38 FILLCELL_X1
* cell instance $4034 m0 *1 64.22,35
X$4034 23 2703 739 819 705 38 DFF_X1
* cell instance $4035 m0 *1 67.45,35
X$4035 739 88 799 23 38 819 MUX2_X1
* cell instance $4036 m0 *1 68.78,35
X$4036 771 38 240 23 BUF_X4
* cell instance $4037 m0 *1 70.11,35
X$4037 23 38 FILLCELL_X1
* cell instance $4038 m0 *1 70.3,35
X$4038 672 51 800 23 38 854 MUX2_X1
* cell instance $4039 m0 *1 71.63,35
X$4039 23 38 FILLCELL_X16
* cell instance $4040 m0 *1 74.67,35
X$4040 23 2796 784 816 801 38 DFF_X1
* cell instance $4041 m0 *1 77.9,35
X$4041 751 840 23 38 850 NOR2_X1
* cell instance $4042 m0 *1 78.47,35
X$4042 23 38 FILLCELL_X1
* cell instance $4043 m0 *1 78.66,35
X$4043 802 274 23 38 814 NOR2_X1
* cell instance $4044 m0 *1 79.23,35
X$4044 23 38 FILLCELL_X16
* cell instance $4045 m0 *1 82.27,35
X$4045 23 38 FILLCELL_X8
* cell instance $4046 m0 *1 83.79,35
X$4046 23 38 FILLCELL_X4
* cell instance $4047 m0 *1 84.55,35
X$4047 23 38 FILLCELL_X2
* cell instance $4048 r0 *1 53.96,35
X$4048 862 38 126 23 BUF_X4
* cell instance $4049 r0 *1 55.29,35
X$4049 839 23 38 CLKBUF_X1
* cell instance $4050 r0 *1 55.86,35
X$4050 23 38 FILLCELL_X4
* cell instance $4051 r0 *1 56.62,35
X$4051 112 821 905 23 38 886 MUX2_X1
* cell instance $4052 r0 *1 57.95,35
X$4052 23 38 FILLCELL_X4
* cell instance $4053 r0 *1 58.71,35
X$4053 23 38 FILLCELL_X2
* cell instance $4054 r0 *1 59.14,35
X$4054 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $4055 r0 *1 59.14,35
X$4055 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $4056 r0 *1 59.14,35
X$4056 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $4057 r0 *1 59.09,35
X$4057 121 821 856 23 38 884 MUX2_X1
* cell instance $4058 r0 *1 60.42,35
X$4058 23 38 FILLCELL_X8
* cell instance $4059 r0 *1 61.94,35
X$4059 23 38 FILLCELL_X2
* cell instance $4060 r0 *1 62.32,35
X$4060 855 261 23 38 1163 NOR2_X1
* cell instance $4061 r0 *1 62.89,35
X$4061 23 38 FILLCELL_X16
* cell instance $4062 r0 *1 65.93,35
X$4062 23 38 FILLCELL_X8
* cell instance $4063 r0 *1 67.45,35
X$4063 23 38 FILLCELL_X4
* cell instance $4064 r0 *1 68.21,35
X$4064 23 38 FILLCELL_X1
* cell instance $4065 r0 *1 68.4,35
X$4065 23 3068 800 854 705 38 DFF_X1
* cell instance $4066 r0 *1 71.63,35
X$4066 23 38 FILLCELL_X2
* cell instance $4067 r0 *1 72.01,35
X$4067 23 38 FILLCELL_X1
* cell instance $4068 r0 *1 72.2,35
X$4068 883 840 23 38 865 NOR2_X1
* cell instance $4069 r0 *1 72.77,35
X$4069 706 865 864 853 818 475 23 38 841 OAI33_X1
* cell instance $4070 r0 *1 74.1,35
X$4070 23 38 FILLCELL_X8
* cell instance $4071 r0 *1 75.62,35
X$4071 23 38 FILLCELL_X1
* cell instance $4072 r0 *1 75.81,35
X$4072 840 23 38 274 CLKBUF_X3
* cell instance $4073 r0 *1 76.76,35
X$4073 23 38 FILLCELL_X4
* cell instance $4074 r0 *1 77.52,35
X$4074 23 38 FILLCELL_X2
* cell instance $4075 r0 *1 77.9,35
X$4075 882 850 600 814 803 227 23 38 1088 OAI33_X1
* cell instance $4076 r0 *1 79.23,35
X$4076 23 38 FILLCELL_X32
* cell instance $4077 m0 *1 85.12,35
X$4077 804 223 799 23 38 848 MUX2_X1
* cell instance $4078 m0 *1 84.93,35
X$4078 23 38 FILLCELL_X1
* cell instance $4079 m0 *1 86.45,35
X$4079 23 2818 804 848 647 38 DFF_X1
* cell instance $4080 m0 *1 89.68,35
X$4080 804 188 776 23 38 805 MUX2_X1
* cell instance $4081 m0 *1 91.01,35
X$4081 23 2789 846 811 647 38 DFF_X1
* cell instance $4082 m0 *1 94.24,35
X$4082 806 133 843 23 38 844 MUX2_X1
* cell instance $4083 m0 *1 95.57,35
X$4083 23 38 FILLCELL_X8
* cell instance $4084 r180 *1 97.28,35
X$4084 23 38 23 38 TAPCELL_X1
* cell instance $4085 r0 *1 85.31,35
X$4085 23 38 FILLCELL_X16
* cell instance $4086 r0 *1 88.35,35
X$4086 23 38 FILLCELL_X8
* cell instance $4087 r0 *1 89.87,35
X$4087 23 38 FILLCELL_X2
* cell instance $4088 r0 *1 90.25,35
X$4088 806 79 846 23 38 811 MUX2_X1
* cell instance $4089 r0 *1 91.58,35
X$4089 843 126 846 23 38 872 MUX2_X1
* cell instance $4090 r0 *1 92.91,35
X$4090 23 2864 843 844 647 38 DFF_X1
* cell instance $4091 r0 *1 96.14,35
X$4091 842 23 38 675 CLKBUF_X2
* cell instance $4092 r0 *1 96.9,35
X$4092 23 38 FILLCELL_X1
* cell instance $4093 m90 *1 97.28,35
X$4093 23 38 23 38 TAPCELL_X1
* cell instance $4094 r0 *1 27.74,1.4
X$4094 23 38 FILLCELL_X1
* cell instance $4095 r0 *1 28.5,1.4
X$4095 23 38 FILLCELL_X16
* cell instance $4096 r0 *1 31.54,1.4
X$4096 23 38 FILLCELL_X4
* cell instance $4097 r0 *1 32.3,1.4
X$4097 23 38 FILLCELL_X2
* cell instance $4098 m0 *1 1.33,29.4
X$4098 23 38 FILLCELL_X4
* cell instance $4099 m0 *1 1.14,29.4
X$4099 23 38 23 38 TAPCELL_X1
* cell instance $4100 m0 *1 2.09,29.4
X$4100 23 2770 691 677 660 38 DFF_X1
* cell instance $4101 m0 *1 5.32,29.4
X$4101 23 38 FILLCELL_X1
* cell instance $4102 m0 *1 5.51,29.4
X$4102 23 2766 692 679 660 38 DFF_X1
* cell instance $4103 m0 *1 8.74,29.4
X$4103 23 38 FILLCELL_X2
* cell instance $4104 r0 *1 1.14,29.4
X$4104 23 38 23 38 TAPCELL_X1
* cell instance $4105 r0 *1 1.33,29.4
X$4105 23 38 FILLCELL_X8
* cell instance $4106 r0 *1 2.85,29.4
X$4106 23 38 FILLCELL_X4
* cell instance $4107 r0 *1 3.14,29.4
X$4107 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $4108 r0 *1 3.14,29.4
X$4108 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $4109 r0 *1 3.14,29.4
X$4109 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $4110 r0 *1 3.61,29.4
X$4110 23 38 FILLCELL_X1
* cell instance $4111 r0 *1 3.8,29.4
X$4111 107 659 732 23 38 715 MUX2_X1
* cell instance $4112 r0 *1 5.13,29.4
X$4112 23 3022 732 715 660 38 DFF_X1
* cell instance $4113 r0 *1 8.36,29.4
X$4113 660 23 38 CLKBUF_X1
* cell instance $4114 r0 *1 8.93,29.4
X$4114 693 23 38 660 CLKBUF_X3
* cell instance $4115 m0 *1 12.35,29.4
X$4115 23 38 FILLCELL_X8
* cell instance $4116 m0 *1 9.12,29.4
X$4116 23 2771 661 681 660 38 DFF_X1
* cell instance $4117 m0 *1 13.87,29.4
X$4117 23 38 FILLCELL_X2
* cell instance $4118 r0 *1 9.88,29.4
X$4118 23 38 FILLCELL_X1
* cell instance $4119 r0 *1 10.07,29.4
X$4119 23 3081 694 718 660 38 DFF_X1
* cell instance $4120 r0 *1 13.3,29.4
X$4120 23 38 FILLCELL_X4
* cell instance $4121 r0 *1 14.06,29.4
X$4121 27 632 694 23 38 718 MUX2_X1
* cell instance $4122 m0 *1 17.48,29.4
X$4122 23 2787 696 720 653 38 DFF_X1
* cell instance $4123 m0 *1 14.25,29.4
X$4123 23 2778 695 719 653 38 DFF_X1
* cell instance $4124 m0 *1 20.71,29.4
X$4124 24 632 696 23 38 720 MUX2_X1
* cell instance $4125 m0 *1 22.04,29.4
X$4125 693 23 38 653 CLKBUF_X3
* cell instance $4126 m0 *1 22.99,29.4
X$4126 26 23 38 358 BUF_X2
* cell instance $4127 m0 *1 23.75,29.4
X$4127 23 38 FILLCELL_X4
* cell instance $4128 m0 *1 24.51,29.4
X$4128 23 38 FILLCELL_X1
* cell instance $4129 m0 *1 24.7,29.4
X$4129 631 602 685 23 38 698 MUX2_X1
* cell instance $4130 m0 *1 26.03,29.4
X$4130 23 38 FILLCELL_X4
* cell instance $4131 m0 *1 26.79,29.4
X$4131 23 38 FILLCELL_X1
* cell instance $4132 m0 *1 26.98,29.4
X$4132 29 632 686 23 38 662 MUX2_X1
* cell instance $4133 m0 *1 28.31,29.4
X$4133 23 38 FILLCELL_X2
* cell instance $4134 r0 *1 15.39,29.4
X$4134 23 38 FILLCELL_X1
* cell instance $4135 r0 *1 15.58,29.4
X$4135 107 632 733 23 38 749 MUX2_X1
* cell instance $4136 r0 *1 16.91,29.4
X$4136 23 38 FILLCELL_X8
* cell instance $4137 r0 *1 18.43,29.4
X$4137 23 38 FILLCELL_X4
* cell instance $4138 r0 *1 19.19,29.4
X$4138 23 38 FILLCELL_X2
* cell instance $4139 r0 *1 19.57,29.4
X$4139 653 23 38 CLKBUF_X1
* cell instance $4140 r0 *1 20.14,29.4
X$4140 629 602 696 23 38 878 MUX2_X1
* cell instance $4141 r0 *1 21.47,29.4
X$4141 23 38 FILLCELL_X2
* cell instance $4142 r0 *1 21.85,29.4
X$4142 26 659 697 23 38 734 MUX2_X1
* cell instance $4143 r0 *1 23.18,29.4
X$4143 23 38 FILLCELL_X16
* cell instance $4144 r0 *1 26.22,29.4
X$4144 23 38 FILLCELL_X8
* cell instance $4145 r0 *1 27.74,29.4
X$4145 23 38 FILLCELL_X4
* cell instance $4146 r0 *1 28.5,29.4
X$4146 23 38 FILLCELL_X2
* cell instance $4147 m0 *1 30.02,29.4
X$4147 23 38 FILLCELL_X4
* cell instance $4148 m0 *1 28.69,29.4
X$4148 29 659 735 23 38 723 MUX2_X1
* cell instance $4149 m0 *1 30.78,29.4
X$4149 23 38 FILLCELL_X1
* cell instance $4150 m0 *1 30.97,29.4
X$4150 510 628 725 23 38 663 MUX2_X1
* cell instance $4151 m0 *1 32.3,29.4
X$4151 23 38 FILLCELL_X8
* cell instance $4152 m0 *1 33.82,29.4
X$4152 23 38 FILLCELL_X2
* cell instance $4153 r0 *1 28.88,29.4
X$4153 23 38 FILLCELL_X1
* cell instance $4154 r0 *1 29.07,29.4
X$4154 23 3060 735 723 655 38 DFF_X1
* cell instance $4155 r0 *1 32.3,29.4
X$4155 23 38 FILLCELL_X2
* cell instance $4156 r0 *1 32.68,29.4
X$4156 23 38 FILLCELL_X1
* cell instance $4157 r0 *1 32.87,29.4
X$4157 25 23 38 510 BUF_X2
* cell instance $4158 r0 *1 33.63,29.4
X$4158 25 659 699 23 38 752 MUX2_X1
* cell instance $4159 m0 *1 34.39,29.4
X$4159 725 602 688 23 38 700 MUX2_X1
* cell instance $4160 m0 *1 34.2,29.4
X$4160 23 38 FILLCELL_X1
* cell instance $4161 m0 *1 35.72,29.4
X$4161 23 38 FILLCELL_X4
* cell instance $4162 m0 *1 36.48,29.4
X$4162 319 628 690 23 38 726 MUX2_X1
* cell instance $4163 m0 *1 37.81,29.4
X$4163 23 38 FILLCELL_X1
* cell instance $4164 m0 *1 38,29.4
X$4164 23 2690 690 726 655 38 DFF_X1
* cell instance $4165 m0 *1 41.23,29.4
X$4165 23 38 FILLCELL_X8
* cell instance $4166 m0 *1 42.75,29.4
X$4166 23 38 FILLCELL_X2
* cell instance $4167 r0 *1 34.96,29.4
X$4167 23 38 FILLCELL_X8
* cell instance $4168 r0 *1 36.48,29.4
X$4168 23 38 FILLCELL_X2
* cell instance $4169 r0 *1 36.86,29.4
X$4169 23 38 FILLCELL_X1
* cell instance $4170 r0 *1 37.05,29.4
X$4170 23 3051 736 727 655 38 DFF_X1
* cell instance $4171 r0 *1 40.28,29.4
X$4171 98 632 736 23 38 727 MUX2_X1
* cell instance $4172 r0 *1 41.61,29.4
X$4172 23 38 FILLCELL_X4
* cell instance $4173 r0 *1 42.37,29.4
X$4173 23 38 FILLCELL_X2
* cell instance $4174 r0 *1 42.75,29.4
X$4174 23 38 FILLCELL_X1
* cell instance $4175 r0 *1 42.94,29.4
X$4175 634 38 724 23 BUF_X4
* cell instance $4176 m0 *1 43.32,29.4
X$4176 398 628 665 23 38 664 MUX2_X1
* cell instance $4177 m0 *1 43.13,29.4
X$4177 23 38 FILLCELL_X1
* cell instance $4178 m0 *1 44.65,29.4
X$4178 23 38 FILLCELL_X2
* cell instance $4179 r0 *1 44.27,29.4
X$4179 23 38 FILLCELL_X2
* cell instance $4180 r0 *1 44.65,29.4
X$4180 75 659 737 23 38 756 MUX2_X1
* cell instance $4181 m0 *1 45.22,29.4
X$4181 665 602 637 23 38 701 MUX2_X1
* cell instance $4182 m0 *1 45.03,29.4
X$4182 23 38 FILLCELL_X1
* cell instance $4183 m0 *1 46.55,29.4
X$4183 23 38 FILLCELL_X16
* cell instance $4184 m0 *1 49.59,29.4
X$4184 23 38 FILLCELL_X1
* cell instance $4185 m0 *1 49.78,29.4
X$4185 301 628 667 23 38 689 MUX2_X1
* cell instance $4186 m0 *1 51.11,29.4
X$4186 667 602 668 23 38 702 MUX2_X1
* cell instance $4187 m0 *1 52.44,29.4
X$4187 66 632 668 23 38 729 MUX2_X1
* cell instance $4188 m0 *1 53.77,29.4
X$4188 23 38 FILLCELL_X32
* cell instance $4189 m0 *1 59.85,29.4
X$4189 23 38 FILLCELL_X2
* cell instance $4190 r0 *1 45.98,29.4
X$4190 23 38 FILLCELL_X1
* cell instance $4191 r0 *1 46.17,29.4
X$4191 701 261 23 38 837 NOR2_X1
* cell instance $4192 r0 *1 46.74,29.4
X$4192 23 38 FILLCELL_X16
* cell instance $4193 r0 *1 49.78,29.4
X$4193 66 659 738 23 38 757 MUX2_X1
* cell instance $4194 r0 *1 51.11,29.4
X$4194 23 38 FILLCELL_X2
* cell instance $4195 r0 *1 51.49,29.4
X$4195 23 38 FILLCELL_X1
* cell instance $4196 r0 *1 51.68,29.4
X$4196 23 3046 668 729 666 38 DFF_X1
* cell instance $4197 r0 *1 54.91,29.4
X$4197 23 38 FILLCELL_X2
* cell instance $4198 r0 *1 55.29,29.4
X$4198 23 38 FILLCELL_X1
* cell instance $4199 r0 *1 55.48,29.4
X$4199 744 23 38 666 CLKBUF_X3
* cell instance $4200 r0 *1 56.43,29.4
X$4200 23 38 FILLCELL_X32
* cell instance $4201 r0 *1 59.14,29.4
X$4201 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $4202 r0 *1 59.14,29.4
X$4202 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $4203 r0 *1 59.14,29.4
X$4203 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $4204 m0 *1 60.42,29.4
X$4204 23 2815 671 670 543 38 DFF_X1
* cell instance $4205 m0 *1 60.23,29.4
X$4205 23 38 FILLCELL_X1
* cell instance $4206 m0 *1 63.65,29.4
X$4206 23 38 FILLCELL_X8
* cell instance $4207 m0 *1 65.17,29.4
X$4207 23 2702 703 731 543 38 DFF_X1
* cell instance $4208 m0 *1 68.4,29.4
X$4208 704 441 672 23 38 730 MUX2_X1
* cell instance $4209 m0 *1 69.73,29.4
X$4209 23 2718 704 730 705 38 DFF_X1
* cell instance $4210 m0 *1 72.96,29.4
X$4210 23 38 FILLCELL_X16
* cell instance $4211 m0 *1 76,29.4
X$4211 23 38 FILLCELL_X1
* cell instance $4212 m0 *1 76.19,29.4
X$4212 682 223 672 23 38 683 MUX2_X1
* cell instance $4213 m0 *1 77.52,29.4
X$4213 23 2799 709 708 673 38 DFF_X1
* cell instance $4214 m0 *1 80.75,29.4
X$4214 23 38 FILLCELL_X8
* cell instance $4215 m0 *1 82.27,29.4
X$4215 23 38 FILLCELL_X4
* cell instance $4216 m0 *1 83.03,29.4
X$4216 744 23 38 673 CLKBUF_X3
* cell instance $4217 m0 *1 83.98,29.4
X$4217 23 2841 711 722 673 38 DFF_X1
* cell instance $4218 m0 *1 87.21,29.4
X$4218 23 38 FILLCELL_X16
* cell instance $4219 m0 *1 90.25,29.4
X$4219 23 38 FILLCELL_X4
* cell instance $4220 m0 *1 91.01,29.4
X$4220 23 38 FILLCELL_X2
* cell instance $4221 r0 *1 62.51,29.4
X$4221 23 38 FILLCELL_X16
* cell instance $4222 r0 *1 65.55,29.4
X$4222 23 38 FILLCELL_X4
* cell instance $4223 r0 *1 66.31,29.4
X$4223 23 38 FILLCELL_X2
* cell instance $4224 r0 *1 66.69,29.4
X$4224 23 38 FILLCELL_X1
* cell instance $4225 r0 *1 66.88,29.4
X$4225 703 373 672 23 38 731 MUX2_X1
* cell instance $4226 r0 *1 68.21,29.4
X$4226 704 126 703 23 38 741 MUX2_X1
* cell instance $4227 r0 *1 69.54,29.4
X$4227 23 38 FILLCELL_X4
* cell instance $4228 r0 *1 70.3,29.4
X$4228 23 2897 743 728 705 38 DFF_X1
* cell instance $4229 r0 *1 73.53,29.4
X$4229 743 520 672 23 38 728 MUX2_X1
* cell instance $4230 r0 *1 74.86,29.4
X$4230 707 370 23 38 706 NOR2_X1
* cell instance $4231 r0 *1 75.43,29.4
X$4231 23 38 FILLCELL_X8
* cell instance $4232 r0 *1 76.95,29.4
X$4232 754 88 672 23 38 755 MUX2_X1
* cell instance $4233 r0 *1 78.28,29.4
X$4233 709 174 672 23 38 708 MUX2_X1
* cell instance $4234 r0 *1 79.61,29.4
X$4234 682 80 709 23 38 783 MUX2_X1
* cell instance $4235 r0 *1 80.94,29.4
X$4235 23 38 FILLCELL_X8
* cell instance $4236 r0 *1 82.46,29.4
X$4236 711 438 712 23 38 751 MUX2_X1
* cell instance $4237 r0 *1 83.79,29.4
X$4237 23 38 FILLCELL_X1
* cell instance $4238 r0 *1 83.98,29.4
X$4238 710 191 711 23 38 722 MUX2_X1
* cell instance $4239 r0 *1 85.31,29.4
X$4239 710 187 712 23 38 721 MUX2_X1
* cell instance $4240 r0 *1 86.64,29.4
X$4240 23 2915 712 721 673 38 DFF_X1
* cell instance $4241 r0 *1 89.87,29.4
X$4241 23 2916 713 717 647 38 DFF_X1
* cell instance $4242 m0 *1 91.96,29.4
X$4242 23 38 FILLCELL_X8
* cell instance $4243 m0 *1 91.39,29.4
X$4243 678 274 23 38 674 NOR2_X1
* cell instance $4244 m0 *1 93.48,29.4
X$4244 23 2827 714 716 647 38 DFF_X1
* cell instance $4245 m0 *1 96.71,29.4
X$4245 23 38 FILLCELL_X2
* cell instance $4246 r0 *1 93.1,29.4
X$4246 675 133 713 23 38 717 MUX2_X1
* cell instance $4247 r0 *1 94.43,29.4
X$4247 23 38 FILLCELL_X1
* cell instance $4248 r0 *1 94.62,29.4
X$4248 675 79 714 23 38 716 MUX2_X1
* cell instance $4249 r0 *1 95.95,29.4
X$4249 23 38 FILLCELL_X4
* cell instance $4250 r0 *1 96.71,29.4
X$4250 23 38 FILLCELL_X2
* cell instance $4251 m0 *1 1.33,88.2
X$4251 23 38 FILLCELL_X4
* cell instance $4252 m0 *1 1.14,88.2
X$4252 23 38 23 38 TAPCELL_X1
* cell instance $4253 m0 *1 2.09,88.2
X$4253 23 38 FILLCELL_X1
* cell instance $4254 m0 *1 2.28,88.2
X$4254 23 2652 2272 2271 2045 38 DFF_X1
* cell instance $4255 m0 *1 5.51,88.2
X$4255 23 2683 2325 2273 2045 38 DFF_X1
* cell instance $4256 m0 *1 8.74,88.2
X$4256 23 38 FILLCELL_X2
* cell instance $4257 r0 *1 1.14,88.2
X$4257 23 38 23 38 TAPCELL_X1
* cell instance $4258 r0 *1 1.33,88.2
X$4258 23 38 FILLCELL_X16
* cell instance $4259 r0 *1 3.14,88.2
X$4259 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $4260 r0 *1 3.14,88.2
X$4260 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $4261 r0 *1 3.14,88.2
X$4261 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $4262 r0 *1 4.37,88.2
X$4262 2272 412 2325 23 38 2375 MUX2_X1
* cell instance $4263 r0 *1 5.7,88.2
X$4263 2272 1383 1820 23 38 2271 MUX2_X1
* cell instance $4264 r0 *1 7.03,88.2
X$4264 23 38 FILLCELL_X1
* cell instance $4265 r0 *1 7.22,88.2
X$4265 23 2969 2327 2326 2045 38 DFF_X1
* cell instance $4266 m0 *1 9.31,88.2
X$4266 2297 1403 1820 23 38 2296 MUX2_X1
* cell instance $4267 m0 *1 9.12,88.2
X$4267 23 38 FILLCELL_X1
* cell instance $4268 m0 *1 10.64,88.2
X$4268 23 38 FILLCELL_X2
* cell instance $4269 r0 *1 10.45,88.2
X$4269 2327 1289 1820 23 38 2326 MUX2_X1
* cell instance $4270 m0 *1 11.21,88.2
X$4270 2297 627 2327 23 38 2328 MUX2_X1
* cell instance $4271 m0 *1 11.02,88.2
X$4271 23 38 FILLCELL_X1
* cell instance $4272 m0 *1 12.54,88.2
X$4272 23 38 FILLCELL_X1
* cell instance $4273 m0 *1 12.73,88.2
X$4273 23 2680 2329 2341 2434 38 DFF_X1
* cell instance $4274 m0 *1 15.96,88.2
X$4274 2274 1369 1822 23 38 2299 MUX2_X1
* cell instance $4275 m0 *1 17.29,88.2
X$4275 23 38 FILLCELL_X2
* cell instance $4276 r0 *1 11.78,88.2
X$4276 2375 1650 23 38 2349 NOR2_X1
* cell instance $4277 r0 *1 12.35,88.2
X$4277 23 38 FILLCELL_X1
* cell instance $4278 r0 *1 12.54,88.2
X$4278 2328 1579 23 38 2350 NOR2_X1
* cell instance $4279 r0 *1 13.11,88.2
X$4279 23 38 FILLCELL_X2
* cell instance $4280 r0 *1 13.49,88.2
X$4280 23 38 FILLCELL_X1
* cell instance $4281 r0 *1 13.68,88.2
X$4281 2329 1383 1822 23 38 2341 MUX2_X1
* cell instance $4282 r0 *1 15.01,88.2
X$4282 23 38 FILLCELL_X2
* cell instance $4283 r0 *1 15.39,88.2
X$4283 2329 412 2274 23 38 2380 MUX2_X1
* cell instance $4284 r0 *1 16.72,88.2
X$4284 2380 1650 23 38 2420 NOR2_X1
* cell instance $4285 r0 *1 17.29,88.2
X$4285 23 38 FILLCELL_X8
* cell instance $4286 m0 *1 17.86,88.2
X$4286 23 2685 2330 2344 2144 38 DFF_X1
* cell instance $4287 m0 *1 17.67,88.2
X$4287 23 38 FILLCELL_X1
* cell instance $4288 m0 *1 21.09,88.2
X$4288 2275 1289 1822 23 38 2239 MUX2_X1
* cell instance $4289 m0 *1 22.42,88.2
X$4289 1909 23 38 2144 CLKBUF_X3
* cell instance $4290 m0 *1 23.37,88.2
X$4290 23 2640 2276 2302 2144 38 DFF_X1
* cell instance $4291 m0 *1 26.6,88.2
X$4291 2276 412 2277 23 38 2305 MUX2_X1
* cell instance $4292 m0 *1 27.93,88.2
X$4292 23 2642 2240 2303 2145 38 DFF_X1
* cell instance $4293 m0 *1 31.16,88.2
X$4293 23 38 FILLCELL_X2
* cell instance $4294 r0 *1 18.81,88.2
X$4294 2330 1403 1822 23 38 2344 MUX2_X1
* cell instance $4295 r0 *1 20.14,88.2
X$4295 2382 1579 23 38 2381 NOR2_X1
* cell instance $4296 r0 *1 20.71,88.2
X$4296 2330 627 2275 23 38 2382 MUX2_X1
* cell instance $4297 r0 *1 22.04,88.2
X$4297 23 38 FILLCELL_X8
* cell instance $4298 r0 *1 23.56,88.2
X$4298 23 3027 2277 2383 2144 38 DFF_X1
* cell instance $4299 r0 *1 26.79,88.2
X$4299 2277 1369 1725 23 38 2383 MUX2_X1
* cell instance $4300 r0 *1 28.12,88.2
X$4300 2356 1289 1725 23 38 2354 MUX2_X1
* cell instance $4301 r0 *1 29.45,88.2
X$4301 23 38 FILLCELL_X4
* cell instance $4302 r0 *1 30.21,88.2
X$4302 2240 627 2356 23 38 2384 MUX2_X1
* cell instance $4303 m0 *1 31.73,88.2
X$4303 2305 1650 23 38 2278 NOR2_X1
* cell instance $4304 m0 *1 31.54,88.2
X$4304 23 38 FILLCELL_X1
* cell instance $4305 m0 *1 32.3,88.2
X$4305 23 38 FILLCELL_X8
* cell instance $4306 m0 *1 33.82,88.2
X$4306 23 38 FILLCELL_X4
* cell instance $4307 m0 *1 34.58,88.2
X$4307 23 38 FILLCELL_X2
* cell instance $4308 r0 *1 31.54,88.2
X$4308 2384 1579 23 38 2385 NOR2_X1
* cell instance $4309 r0 *1 32.11,88.2
X$4309 23 38 FILLCELL_X1
* cell instance $4310 r0 *1 32.3,88.2
X$4310 1425 2385 2278 548 2357 2468 23 38 2008 OAI33_X1
* cell instance $4311 r0 *1 33.63,88.2
X$4311 23 38 FILLCELL_X2
* cell instance $4312 r0 *1 34.01,88.2
X$4312 23 38 FILLCELL_X1
* cell instance $4313 r0 *1 34.2,88.2
X$4313 23 3024 2358 2386 2333 38 DFF_X1
* cell instance $4314 m0 *1 38.19,88.2
X$4314 23 38 FILLCELL_X8
* cell instance $4315 m0 *1 34.96,88.2
X$4315 23 2635 2331 2347 2333 38 DFF_X1
* cell instance $4316 m0 *1 39.71,88.2
X$4316 2308 1383 1730 23 38 2307 MUX2_X1
* cell instance $4317 m0 *1 41.04,88.2
X$4317 23 38 FILLCELL_X2
* cell instance $4318 r0 *1 37.43,88.2
X$4318 2331 1289 1730 23 38 2347 MUX2_X1
* cell instance $4319 r0 *1 38.76,88.2
X$4319 23 38 FILLCELL_X2
* cell instance $4320 r0 *1 39.14,88.2
X$4320 23 3083 2332 2348 2333 38 DFF_X1
* cell instance $4321 m0 *1 42.75,88.2
X$4321 23 38 FILLCELL_X16
* cell instance $4322 m0 *1 41.42,88.2
X$4322 2332 1369 1730 23 38 2348 MUX2_X1
* cell instance $4323 m0 *1 45.79,88.2
X$4323 23 38 FILLCELL_X8
* cell instance $4324 m0 *1 47.31,88.2
X$4324 23 38 FILLCELL_X4
* cell instance $4325 m0 *1 48.07,88.2
X$4325 2241 627 2279 23 38 2346 MUX2_X1
* cell instance $4326 m0 *1 49.4,88.2
X$4326 23 38 FILLCELL_X2
* cell instance $4327 r0 *1 42.37,88.2
X$4327 2308 724 2332 23 38 2361 MUX2_X1
* cell instance $4328 r0 *1 43.7,88.2
X$4328 23 38 FILLCELL_X2
* cell instance $4329 r0 *1 44.08,88.2
X$4329 23 3074 2334 2392 2333 38 DFF_X1
* cell instance $4330 r0 *1 47.31,88.2
X$4330 2334 1403 1813 23 38 2392 MUX2_X1
* cell instance $4331 r0 *1 48.64,88.2
X$4331 23 38 FILLCELL_X4
* cell instance $4332 r0 *1 49.4,88.2
X$4332 2397 1383 1813 23 38 2395 MUX2_X1
* cell instance $4333 m0 *1 49.97,88.2
X$4333 2346 1579 23 38 2310 NOR2_X1
* cell instance $4334 m0 *1 49.78,88.2
X$4334 23 38 FILLCELL_X1
* cell instance $4335 m0 *1 50.54,88.2
X$4335 23 38 FILLCELL_X16
* cell instance $4336 m0 *1 53.58,88.2
X$4336 23 38 FILLCELL_X8
* cell instance $4337 m0 *1 55.1,88.2
X$4337 23 38 FILLCELL_X4
* cell instance $4338 m0 *1 55.86,88.2
X$4338 2151 1406 2280 23 38 2314 MUX2_X1
* cell instance $4339 m0 *1 57.19,88.2
X$4339 23 2592 2280 2314 2316 38 DFF_X1
* cell instance $4340 m0 *1 60.42,88.2
X$4340 23 38 FILLCELL_X8
* cell instance $4341 m0 *1 61.94,88.2
X$4341 23 38 FILLCELL_X2
* cell instance $4342 r0 *1 50.73,88.2
X$4342 23 3114 2397 2395 2316 38 DFF_X1
* cell instance $4343 r0 *1 53.96,88.2
X$4343 23 38 FILLCELL_X8
* cell instance $4344 r0 *1 55.48,88.2
X$4344 23 38 FILLCELL_X2
* cell instance $4345 r0 *1 55.86,88.2
X$4345 2398 1483 23 38 2244 NOR2_X1
* cell instance $4346 r0 *1 56.43,88.2
X$4346 23 38 FILLCELL_X32
* cell instance $4347 r0 *1 59.14,88.2
X$4347 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $4348 r0 *1 59.14,88.2
X$4348 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $4349 r0 *1 59.14,88.2
X$4349 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $4350 m0 *1 62.51,88.2
X$4350 2223 23 38 2213 INV_X1
* cell instance $4351 m0 *1 62.32,88.2
X$4351 23 38 FILLCELL_X1
* cell instance $4352 m0 *1 62.89,88.2
X$4352 23 38 FILLCELL_X4
* cell instance $4353 m0 *1 63.65,88.2
X$4353 1949 2213 23 38 2335 NOR2_X1
* cell instance $4354 m0 *1 64.22,88.2
X$4354 1496 2236 23 38 2345 NAND2_X1
* cell instance $4355 m0 *1 64.79,88.2
X$4355 2116 2223 23 38 2281 NOR2_X1
* cell instance $4356 m0 *1 65.36,88.2
X$4356 23 38 FILLCELL_X2
* cell instance $4357 r0 *1 62.51,88.2
X$4357 23 38 FILLCELL_X4
* cell instance $4358 r0 *1 63.27,88.2
X$4358 23 38 FILLCELL_X1
* cell instance $4359 r0 *1 63.46,88.2
X$4359 2335 2394 2281 23 38 2396 MUX2_X1
* cell instance $4360 r0 *1 64.79,88.2
X$4360 2058 23 38 2246 CLKBUF_X3
* cell instance $4361 r0 *1 65.74,88.2
X$4361 2345 2065 2232 23 2394 38 AOI21_X1
* cell instance $4362 m0 *1 68.97,88.2
X$4362 23 38 FILLCELL_X2
* cell instance $4363 m0 *1 65.74,88.2
X$4363 23 2577 2320 2319 2246 38 DFF_X1
* cell instance $4364 r0 *1 66.5,88.2
X$4364 2364 23 38 2223 CLKBUF_X2
* cell instance $4365 r0 *1 67.26,88.2
X$4365 23 38 FILLCELL_X8
* cell instance $4366 r0 *1 68.78,88.2
X$4366 23 2472 2283 1980 2246 38 DFF_X1
* cell instance $4367 m0 *1 69.54,88.2
X$4367 2322 2057 38 23 2282 AND2_X1
* cell instance $4368 m0 *1 69.35,88.2
X$4368 23 38 FILLCELL_X1
* cell instance $4369 m0 *1 70.3,88.2
X$4369 2283 1460 38 23 2321 AND2_X1
* cell instance $4370 m0 *1 71.06,88.2
X$4370 2324 2283 2322 38 23 2285 HA_X1
* cell instance $4371 m0 *1 72.96,88.2
X$4371 2283 2284 2187 2160 23 38 2286 NAND4_X1
* cell instance $4372 m0 *1 73.91,88.2
X$4372 2286 2190 2232 23 2323 38 AOI21_X1
* cell instance $4373 m0 *1 74.67,88.2
X$4373 23 38 FILLCELL_X8
* cell instance $4374 m0 *1 76.19,88.2
X$4374 23 38 FILLCELL_X4
* cell instance $4375 m0 *1 76.95,88.2
X$4375 2190 23 38 2249 INV_X1
* cell instance $4376 m0 *1 77.33,88.2
X$4376 23 1300 38 2287 BUF_X8
* cell instance $4377 m0 *1 79.8,88.2
X$4377 2287 38 1686 23 BUF_X4
* cell instance $4378 m0 *1 81.13,88.2
X$4378 23 38 FILLCELL_X16
* cell instance $4379 m0 *1 84.17,88.2
X$4379 23 38 FILLCELL_X1
* cell instance $4380 m0 *1 84.36,88.2
X$4380 2288 23 38 2342 INV_X1
* cell instance $4381 m0 *1 84.74,88.2
X$4381 23 38 FILLCELL_X4
* cell instance $4382 m0 *1 85.5,88.2
X$4382 23 38 FILLCELL_X1
* cell instance $4383 m0 *1 85.69,88.2
X$4383 2289 2290 23 38 2337 NOR2_X1
* cell instance $4384 m0 *1 86.26,88.2
X$4384 23 38 FILLCELL_X2
* cell instance $4385 r0 *1 72.01,88.2
X$4385 2187 23 38 2324 BUF_X1
* cell instance $4386 r0 *1 72.58,88.2
X$4386 23 38 FILLCELL_X4
* cell instance $4387 r0 *1 73.34,88.2
X$4387 2285 2160 23 38 2366 NAND2_X1
* cell instance $4388 r0 *1 73.91,88.2
X$4388 2248 2320 2336 38 23 2367 HA_X1
* cell instance $4389 r0 *1 75.81,88.2
X$4389 23 38 FILLCELL_X16
* cell instance $4390 r0 *1 78.85,88.2
X$4390 23 38 FILLCELL_X8
* cell instance $4391 r0 *1 80.37,88.2
X$4391 23 38 FILLCELL_X4
* cell instance $4392 r0 *1 81.13,88.2
X$4392 23 38 FILLCELL_X1
* cell instance $4393 r0 *1 81.32,88.2
X$4393 2369 1460 38 23 2368 AND2_X1
* cell instance $4394 r0 *1 82.08,88.2
X$4394 2388 2343 2368 23 38 2389 MUX2_X1
* cell instance $4395 r0 *1 83.41,88.2
X$4395 1949 2369 23 38 2388 NOR2_X1
* cell instance $4396 r0 *1 83.98,88.2
X$4396 23 38 FILLCELL_X2
* cell instance $4397 r0 *1 84.36,88.2
X$4397 2370 2342 2232 2190 23 38 2343 NAND4_X1
* cell instance $4398 r0 *1 85.31,88.2
X$4398 23 38 FILLCELL_X2
* cell instance $4399 r0 *1 85.69,88.2
X$4399 2370 2193 2369 23 38 2378 NAND3_X1
* cell instance $4400 r0 *1 86.45,88.2
X$4400 2161 2063 2337 2338 23 38 2339 NAND4_X1
* cell instance $4401 m0 *1 86.83,88.2
X$4401 2288 1300 2065 23 38 2300 NOR3_X1
* cell instance $4402 m0 *1 86.64,88.2
X$4402 23 38 FILLCELL_X1
* cell instance $4403 m0 *1 87.59,88.2
X$4403 23 38 FILLCELL_X4
* cell instance $4404 m0 *1 88.35,88.2
X$4404 23 2591 2251 2306 2026 38 DFF_X1
* cell instance $4405 m0 *1 91.58,88.2
X$4405 2225 2113 38 23 2291 AND2_X1
* cell instance $4406 m0 *1 92.34,88.2
X$4406 2291 2300 2292 23 38 2340 MUX2_X1
* cell instance $4407 m0 *1 93.67,88.2
X$4407 23 38 FILLCELL_X8
* cell instance $4408 m0 *1 95.19,88.2
X$4408 2293 23 38 2225 CLKBUF_X2
* cell instance $4409 m0 *1 95.95,88.2
X$4409 23 38 FILLCELL_X4
* cell instance $4410 m0 *1 96.71,88.2
X$4410 23 38 FILLCELL_X2
* cell instance $4411 r0 *1 87.4,88.2
X$4411 2339 1300 2065 23 38 2379 NOR3_X1
* cell instance $4412 r0 *1 88.16,88.2
X$4412 1949 2338 23 38 2377 NOR2_X1
* cell instance $4413 r0 *1 88.73,88.2
X$4413 23 38 FILLCELL_X2
* cell instance $4414 r0 *1 89.11,88.2
X$4414 2338 1460 38 23 2371 AND2_X1
* cell instance $4415 r0 *1 89.87,88.2
X$4415 23 38 FILLCELL_X8
* cell instance $4416 r0 *1 91.39,88.2
X$4416 23 38 FILLCELL_X4
* cell instance $4417 r0 *1 92.15,88.2
X$4417 23 38 FILLCELL_X1
* cell instance $4418 r0 *1 92.34,88.2
X$4418 23 3099 2293 2340 2373 38 DFF_X1
* cell instance $4419 r0 *1 95.57,88.2
X$4419 23 38 FILLCELL_X8
* cell instance $4420 m90 *1 97.28,88.2
X$4420 23 38 23 38 TAPCELL_X1
* cell instance $4421 r180 *1 97.28,88.2
X$4421 23 38 23 38 TAPCELL_X1
* cell instance $4422 m0 *1 1.33,82.6
X$4422 23 38 FILLCELL_X4
* cell instance $4423 m0 *1 1.14,82.6
X$4423 23 38 23 38 TAPCELL_X1
* cell instance $4424 m0 *1 2.09,82.6
X$4424 23 2660 2175 2174 1902 38 DFF_X1
* cell instance $4425 m0 *1 5.32,82.6
X$4425 2175 1358 2165 23 38 2202 MUX2_X1
* cell instance $4426 m0 *1 6.65,82.6
X$4426 23 38 FILLCELL_X4
* cell instance $4427 m0 *1 7.41,82.6
X$4427 1820 1544 2140 23 38 2198 MUX2_X1
* cell instance $4428 m0 *1 8.74,82.6
X$4428 23 38 FILLCELL_X4
* cell instance $4429 m0 *1 9.5,82.6
X$4429 23 38 FILLCELL_X1
* cell instance $4430 m0 *1 9.69,82.6
X$4430 2140 813 2141 23 38 2126 MUX2_X1
* cell instance $4431 m0 *1 11.02,82.6
X$4431 23 38 FILLCELL_X4
* cell instance $4432 m0 *1 11.78,82.6
X$4432 23 38 FILLCELL_X2
* cell instance $4433 r0 *1 1.14,82.6
X$4433 23 38 23 38 TAPCELL_X1
* cell instance $4434 r0 *1 1.33,82.6
X$4434 23 38 FILLCELL_X4
* cell instance $4435 r0 *1 2.09,82.6
X$4435 23 38 FILLCELL_X1
* cell instance $4436 r0 *1 2.28,82.6
X$4436 1935 1406 2175 23 38 2174 MUX2_X1
* cell instance $4437 r0 *1 3.14,82.6
X$4437 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $4438 r0 *1 3.14,82.6
X$4438 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $4439 r0 *1 3.14,82.6
X$4439 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $4440 r0 *1 3.61,82.6
X$4440 1935 1346 2165 23 38 2197 MUX2_X1
* cell instance $4441 r0 *1 4.94,82.6
X$4441 23 38 FILLCELL_X4
* cell instance $4442 r0 *1 5.7,82.6
X$4442 23 38 FILLCELL_X2
* cell instance $4443 r0 *1 6.08,82.6
X$4443 23 3122 2140 2198 2045 38 DFF_X1
* cell instance $4444 r0 *1 9.31,82.6
X$4444 2199 1482 2141 23 38 2216 MUX2_X1
* cell instance $4445 r0 *1 10.64,82.6
X$4445 23 38 FILLCELL_X8
* cell instance $4446 m0 *1 12.35,82.6
X$4446 2202 1535 23 38 2166 NOR2_X1
* cell instance $4447 m0 *1 12.16,82.6
X$4447 23 38 FILLCELL_X1
* cell instance $4448 m0 *1 12.92,82.6
X$4448 2199 1530 2176 23 38 2203 MUX2_X1
* cell instance $4449 m0 *1 14.25,82.6
X$4449 23 38 FILLCELL_X2
* cell instance $4450 r0 *1 12.16,82.6
X$4450 23 38 FILLCELL_X2
* cell instance $4451 r0 *1 12.54,82.6
X$4451 23 2959 2176 2203 1902 38 DFF_X1
* cell instance $4452 m0 *1 17.86,82.6
X$4452 23 38 FILLCELL_X2
* cell instance $4453 m0 *1 14.63,82.6
X$4453 23 2664 2105 2142 1848 38 DFF_X1
* cell instance $4454 r0 *1 15.77,82.6
X$4454 23 38 FILLCELL_X8
* cell instance $4455 r0 *1 17.29,82.6
X$4455 23 38 FILLCELL_X4
* cell instance $4456 r0 *1 18.05,82.6
X$4456 23 38 FILLCELL_X2
* cell instance $4457 m0 *1 18.43,82.6
X$4457 23 2663 2127 2143 2144 38 DFF_X1
* cell instance $4458 m0 *1 18.24,82.6
X$4458 23 38 FILLCELL_X1
* cell instance $4459 m0 *1 21.66,82.6
X$4459 23 38 FILLCELL_X2
* cell instance $4460 r0 *1 18.43,82.6
X$4460 23 38 FILLCELL_X1
* cell instance $4461 r0 *1 18.62,82.6
X$4461 23 2938 2177 2229 2144 38 DFF_X1
* cell instance $4462 r0 *1 21.85,82.6
X$4462 23 38 FILLCELL_X4
* cell instance $4463 m0 *1 22.23,82.6
X$4463 23 2631 2128 2167 2145 38 DFF_X1
* cell instance $4464 m0 *1 22.04,82.6
X$4464 23 38 FILLCELL_X1
* cell instance $4465 m0 *1 25.46,82.6
X$4465 23 38 FILLCELL_X2
* cell instance $4466 r0 *1 22.61,82.6
X$4466 23 3017 2178 2231 2145 38 DFF_X1
* cell instance $4467 r0 *1 25.84,82.6
X$4467 23 38 FILLCELL_X8
* cell instance $4468 m0 *1 26.03,82.6
X$4468 23 2632 2106 2205 2145 38 DFF_X1
* cell instance $4469 m0 *1 25.84,82.6
X$4469 23 38 FILLCELL_X1
* cell instance $4470 m0 *1 29.26,82.6
X$4470 23 38 FILLCELL_X8
* cell instance $4471 m0 *1 30.78,82.6
X$4471 23 38 FILLCELL_X4
* cell instance $4472 m0 *1 31.54,82.6
X$4472 23 2622 2180 2208 2145 38 DFF_X1
* cell instance $4473 m0 *1 34.77,82.6
X$4473 23 38 FILLCELL_X8
* cell instance $4474 m0 *1 36.29,82.6
X$4474 23 38 FILLCELL_X2
* cell instance $4475 r0 *1 27.36,82.6
X$4475 23 38 FILLCELL_X2
* cell instance $4476 r0 *1 27.74,82.6
X$4476 2218 1530 2206 23 38 2179 MUX2_X1
* cell instance $4477 r0 *1 29.07,82.6
X$4477 1909 23 38 2145 CLKBUF_X3
* cell instance $4478 r0 *1 30.02,82.6
X$4478 23 38 FILLCELL_X8
* cell instance $4479 r0 *1 31.54,82.6
X$4479 23 38 FILLCELL_X4
* cell instance $4480 r0 *1 32.3,82.6
X$4480 23 38 FILLCELL_X1
* cell instance $4481 r0 *1 32.49,82.6
X$4481 2218 1482 2180 23 38 2208 MUX2_X1
* cell instance $4482 r0 *1 33.82,82.6
X$4482 23 38 FILLCELL_X1
* cell instance $4483 r0 *1 34.01,82.6
X$4483 1725 1544 2107 23 38 2233 MUX2_X1
* cell instance $4484 r0 *1 35.34,82.6
X$4484 23 38 FILLCELL_X4
* cell instance $4485 r0 *1 36.1,82.6
X$4485 23 3023 2219 2234 1933 38 DFF_X1
* cell instance $4486 m0 *1 36.86,82.6
X$4486 1730 1492 2146 23 38 2173 MUX2_X1
* cell instance $4487 m0 *1 36.67,82.6
X$4487 23 38 FILLCELL_X1
* cell instance $4488 m0 *1 38.19,82.6
X$4488 2146 792 2219 23 38 2091 MUX2_X1
* cell instance $4489 m0 *1 39.52,82.6
X$4489 23 38 FILLCELL_X4
* cell instance $4490 m0 *1 40.28,82.6
X$4490 23 38 FILLCELL_X2
* cell instance $4491 r0 *1 39.33,82.6
X$4491 23 38 FILLCELL_X8
* cell instance $4492 m0 *1 43.89,82.6
X$4492 23 38 FILLCELL_X16
* cell instance $4493 m0 *1 40.66,82.6
X$4493 23 2627 2108 2148 2149 38 DFF_X1
* cell instance $4494 m0 *1 46.93,82.6
X$4494 23 38 FILLCELL_X2
* cell instance $4495 r0 *1 40.85,82.6
X$4495 23 3059 2221 2235 2149 38 DFF_X1
* cell instance $4496 r0 *1 44.08,82.6
X$4496 23 38 FILLCELL_X2
* cell instance $4497 r0 *1 44.46,82.6
X$4497 23 38 FILLCELL_X1
* cell instance $4498 r0 *1 44.65,82.6
X$4498 2149 23 38 CLKBUF_X1
* cell instance $4499 r0 *1 45.22,82.6
X$4499 23 38 FILLCELL_X8
* cell instance $4500 r0 *1 46.74,82.6
X$4500 23 38 FILLCELL_X4
* cell instance $4501 m0 *1 50.54,82.6
X$4501 23 38 FILLCELL_X4
* cell instance $4502 m0 *1 47.31,82.6
X$4502 23 2724 2181 2209 2149 38 DFF_X1
* cell instance $4503 m0 *1 51.3,82.6
X$4503 23 38 FILLCELL_X2
* cell instance $4504 r0 *1 47.5,82.6
X$4504 23 38 FILLCELL_X2
* cell instance $4505 r0 *1 47.88,82.6
X$4505 23 38 FILLCELL_X1
* cell instance $4506 r0 *1 48.07,82.6
X$4506 2182 1482 2181 23 38 2209 MUX2_X1
* cell instance $4507 r0 *1 49.4,82.6
X$4507 2182 23 38 1813 BUF_X2
* cell instance $4508 r0 *1 50.16,82.6
X$4508 23 38 FILLCELL_X8
* cell instance $4509 r0 *1 51.68,82.6
X$4509 2238 1369 1767 23 38 2184 MUX2_X1
* cell instance $4510 m0 *1 51.87,82.6
X$4510 23 2595 2138 2150 1960 38 DFF_X1
* cell instance $4511 m0 *1 51.68,82.6
X$4511 23 38 FILLCELL_X1
* cell instance $4512 m0 *1 55.1,82.6
X$4512 2151 1482 2211 23 38 2210 MUX2_X1
* cell instance $4513 m0 *1 56.43,82.6
X$4513 23 38 FILLCELL_X4
* cell instance $4514 m0 *1 57.19,82.6
X$4514 23 38 FILLCELL_X2
* cell instance $4515 r0 *1 53.01,82.6
X$4515 1960 23 38 CLKBUF_X1
* cell instance $4516 r0 *1 53.58,82.6
X$4516 23 38 FILLCELL_X1
* cell instance $4517 r0 *1 53.77,82.6
X$4517 23 2974 2211 2210 1960 38 DFF_X1
* cell instance $4518 r0 *1 57,82.6
X$4518 23 38 FILLCELL_X16
* cell instance $4519 m0 *1 58.9,82.6
X$4519 23 38 FILLCELL_X16
* cell instance $4520 m0 *1 57.57,82.6
X$4520 2151 1530 2020 23 38 2152 MUX2_X1
* cell instance $4521 m0 *1 61.94,82.6
X$4521 23 38 FILLCELL_X4
* cell instance $4522 m0 *1 62.7,82.6
X$4522 1458 1496 23 771 38 NAND2_X4
* cell instance $4523 m0 *1 64.41,82.6
X$4523 23 38 FILLCELL_X1
* cell instance $4524 m0 *1 64.6,82.6
X$4524 2186 2154 3134 38 23 1597 HA_X1
* cell instance $4525 m0 *1 66.5,82.6
X$4525 23 38 FILLCELL_X2
* cell instance $4526 r0 *1 59.14,82.6
X$4526 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $4527 r0 *1 59.14,82.6
X$4527 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $4528 r0 *1 59.14,82.6
X$4528 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $4529 r0 *1 60.04,82.6
X$4529 23 38 FILLCELL_X8
* cell instance $4530 r0 *1 61.56,82.6
X$4530 23 38 FILLCELL_X2
* cell instance $4531 r0 *1 61.94,82.6
X$4531 23 38 FILLCELL_X1
* cell instance $4532 r0 *1 62.13,82.6
X$4532 2237 23 38 1457 CLKBUF_X3
* cell instance $4533 r0 *1 63.08,82.6
X$4533 2213 2185 2155 38 1444 23 NOR3_X2
* cell instance $4534 r0 *1 64.41,82.6
X$4534 2223 2185 2155 38 1442 23 NOR3_X2
* cell instance $4535 r0 *1 65.74,82.6
X$4535 23 38 FILLCELL_X8
* cell instance $4536 m0 *1 67.07,82.6
X$4536 2155 2156 1951 23 2157 38 AOI21_X1
* cell instance $4537 m0 *1 66.88,82.6
X$4537 23 38 FILLCELL_X1
* cell instance $4538 m0 *1 67.83,82.6
X$4538 2171 2157 2215 23 38 2214 MUX2_X1
* cell instance $4539 m0 *1 69.16,82.6
X$4539 2186 1460 38 23 2215 AND2_X1
* cell instance $4540 m0 *1 69.92,82.6
X$4540 23 38 FILLCELL_X2
* cell instance $4541 r0 *1 67.26,82.6
X$4541 23 38 FILLCELL_X1
* cell instance $4542 r0 *1 67.45,82.6
X$4542 23 2214 1981 2186 2102 38 DFF_X2
* cell instance $4543 m0 *1 73.91,82.6
X$4543 2058 23 38 1981 CLKBUF_X3
* cell instance $4544 m0 *1 70.3,82.6
X$4544 23 2158 1981 2056 2187 38 DFF_X2
* cell instance $4545 m0 *1 74.86,82.6
X$4545 23 38 FILLCELL_X1
* cell instance $4546 m0 *1 75.05,82.6
X$4546 23 2649 2115 2212 1981 38 DFF_X1
* cell instance $4547 m0 *1 78.28,82.6
X$4547 23 38 FILLCELL_X16
* cell instance $4548 m0 *1 81.32,82.6
X$4548 23 38 FILLCELL_X2
* cell instance $4549 r0 *1 71.06,82.6
X$4549 23 38 FILLCELL_X2
* cell instance $4550 r0 *1 71.44,82.6
X$4550 1949 2187 23 38 2137 NOR2_X1
* cell instance $4551 r0 *1 72.01,82.6
X$4551 2187 1478 38 23 2170 AND2_X1
* cell instance $4552 r0 *1 72.77,82.6
X$4552 23 38 FILLCELL_X4
* cell instance $4553 r0 *1 73.53,82.6
X$4553 23 38 FILLCELL_X2
* cell instance $4554 r0 *1 73.91,82.6
X$4554 23 38 FILLCELL_X1
* cell instance $4555 r0 *1 74.1,82.6
X$4555 771 1951 2232 23 2114 38 AOI21_X1
* cell instance $4556 r0 *1 74.86,82.6
X$4556 23 38 FILLCELL_X8
* cell instance $4557 r0 *1 76.38,82.6
X$4557 23 38 FILLCELL_X4
* cell instance $4558 r0 *1 77.14,82.6
X$4558 23 38 FILLCELL_X1
* cell instance $4559 r0 *1 77.33,82.6
X$4559 2188 2115 38 2189 23 XOR2_X2
* cell instance $4560 r0 *1 79.04,82.6
X$4560 2116 2188 23 38 2262 NOR2_X1
* cell instance $4561 r0 *1 79.61,82.6
X$4561 2188 2113 38 23 2230 AND2_X1
* cell instance $4562 r0 *1 80.37,82.6
X$4562 23 38 FILLCELL_X8
* cell instance $4563 m0 *1 81.7,82.6
X$4563 23 38 FILLCELL_X1
* cell instance $4564 m0 *1 81.89,82.6
X$4564 2156 2190 2062 2160 23 38 2159 NAND4_X1
* cell instance $4565 m0 *1 82.84,82.6
X$4565 2156 2190 2160 23 38 2025 NAND3_X2
* cell instance $4566 m0 *1 84.17,82.6
X$4566 23 38 FILLCELL_X16
* cell instance $4567 m0 *1 87.21,82.6
X$4567 23 38 FILLCELL_X4
* cell instance $4568 m0 *1 87.97,82.6
X$4568 23 38 FILLCELL_X2
* cell instance $4569 r0 *1 81.89,82.6
X$4569 23 38 FILLCELL_X4
* cell instance $4570 r0 *1 82.65,82.6
X$4570 23 3130 2192 2191 1917 38 DFF_X1
* cell instance $4571 r0 *1 85.88,82.6
X$4571 23 38 FILLCELL_X4
* cell instance $4572 r0 *1 86.64,82.6
X$4572 2063 2207 38 23 2193 AND2_X1
* cell instance $4573 r0 *1 87.4,82.6
X$4573 23 38 FILLCELL_X4
* cell instance $4574 r0 *1 88.16,82.6
X$4574 23 38 FILLCELL_X1
* cell instance $4575 m0 *1 88.35,82.6
X$4575 23 38 FILLCELL_X1
* cell instance $4576 m0 *1 88.54,82.6
X$4576 2062 2064 2069 38 23 2207 AND3_X1
* cell instance $4577 m0 *1 89.49,82.6
X$4577 23 38 FILLCELL_X8
* cell instance $4578 m0 *1 91.01,82.6
X$4578 23 38 FILLCELL_X2
* cell instance $4579 r0 *1 88.35,82.6
X$4579 2251 1460 38 23 2194 AND2_X1
* cell instance $4580 r0 *1 89.11,82.6
X$4580 23 38 FILLCELL_X1
* cell instance $4581 r0 *1 89.3,82.6
X$4581 2207 2063 2225 23 38 2204 NAND3_X1
* cell instance $4582 r0 *1 90.06,82.6
X$4582 23 38 FILLCELL_X1
* cell instance $4583 r0 *1 90.25,82.6
X$4583 2204 1686 2065 23 38 2195 NOR3_X1
* cell instance $4584 r0 *1 91.01,82.6
X$4584 2227 2195 2201 23 38 2200 MUX2_X1
* cell instance $4585 m0 *1 92.15,82.6
X$4585 2116 2226 23 38 2201 NOR2_X1
* cell instance $4586 m0 *1 91.39,82.6
X$4586 2069 2113 38 23 2120 AND2_X1
* cell instance $4587 m0 *1 92.72,82.6
X$4587 2116 2069 23 38 2066 NOR2_X1
* cell instance $4588 m0 *1 93.29,82.6
X$4588 23 38 FILLCELL_X1
* cell instance $4589 m0 *1 93.48,82.6
X$4589 2058 23 38 2026 CLKBUF_X3
* cell instance $4590 m0 *1 94.43,82.6
X$4590 2026 23 38 CLKBUF_X1
* cell instance $4591 m0 *1 95,82.6
X$4591 23 38 FILLCELL_X8
* cell instance $4592 m0 *1 96.52,82.6
X$4592 2069 23 38 2162 BUF_X1
* cell instance $4593 r180 *1 97.28,82.6
X$4593 23 38 23 38 TAPCELL_X1
* cell instance $4594 r0 *1 92.34,82.6
X$4594 23 38 FILLCELL_X4
* cell instance $4595 r0 *1 93.1,82.6
X$4595 23 38 FILLCELL_X1
* cell instance $4596 r0 *1 93.29,82.6
X$4596 23 3108 2196 2200 2026 38 DFF_X1
* cell instance $4597 r0 *1 96.52,82.6
X$4597 23 38 FILLCELL_X2
* cell instance $4598 r0 *1 96.9,82.6
X$4598 23 38 FILLCELL_X1
* cell instance $4599 m90 *1 97.28,82.6
X$4599 23 38 23 38 TAPCELL_X1
* cell instance $4600 m0 *1 1.33,77
X$4600 23 38 FILLCELL_X4
* cell instance $4601 m0 *1 1.14,77
X$4601 23 38 23 38 TAPCELL_X1
* cell instance $4602 m0 *1 2.09,77
X$4602 23 38 FILLCELL_X1
* cell instance $4603 m0 *1 2.28,77
X$4603 23 2661 1950 1967 1902 38 DFF_X1
* cell instance $4604 m0 *1 5.51,77
X$4604 1935 1480 1968 23 38 2029 MUX2_X1
* cell instance $4605 m0 *1 6.84,77
X$4605 23 38 FILLCELL_X4
* cell instance $4606 m0 *1 7.6,77
X$4606 1791 1544 2000 23 38 2031 MUX2_X1
* cell instance $4607 m0 *1 8.93,77
X$4607 23 38 FILLCELL_X8
* cell instance $4608 m0 *1 10.45,77
X$4608 23 38 FILLCELL_X4
* cell instance $4609 m0 *1 11.21,77
X$4609 1935 23 38 1791 BUF_X2
* cell instance $4610 m0 *1 11.97,77
X$4610 23 38 FILLCELL_X8
* cell instance $4611 m0 *1 13.49,77
X$4611 23 38 FILLCELL_X2
* cell instance $4612 r0 *1 1.14,77
X$4612 23 38 23 38 TAPCELL_X1
* cell instance $4613 r0 *1 1.33,77
X$4613 23 38 FILLCELL_X8
* cell instance $4614 r0 *1 2.85,77
X$4614 23 38 FILLCELL_X2
* cell instance $4615 r0 *1 3.14,77
X$4615 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $4616 r0 *1 3.14,77
X$4616 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $4617 r0 *1 3.14,77
X$4617 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $4618 r0 *1 3.23,77
X$4618 23 38 FILLCELL_X1
* cell instance $4619 r0 *1 3.42,77
X$4619 23 2970 1968 2029 1902 38 DFF_X1
* cell instance $4620 r0 *1 6.65,77
X$4620 23 2937 2000 2031 1902 38 DFF_X1
* cell instance $4621 r0 *1 9.88,77
X$4621 2000 813 2046 23 38 2078 MUX2_X1
* cell instance $4622 r0 *1 11.21,77
X$4622 23 38 FILLCELL_X2
* cell instance $4623 r0 *1 11.59,77
X$4623 23 38 FILLCELL_X1
* cell instance $4624 r0 *1 11.78,77
X$4624 1935 1530 2047 23 38 2072 MUX2_X1
* cell instance $4625 r0 *1 13.11,77
X$4625 23 38 FILLCELL_X1
* cell instance $4626 r0 *1 13.3,77
X$4626 23 2939 2033 2075 1848 38 DFF_X1
* cell instance $4627 m0 *1 14.06,77
X$4627 23 2578 1936 1988 1848 38 DFF_X1
* cell instance $4628 m0 *1 13.87,77
X$4628 23 38 FILLCELL_X1
* cell instance $4629 m0 *1 17.29,77
X$4629 23 2662 1937 1969 1848 38 DFF_X1
* cell instance $4630 m0 *1 20.52,77
X$4630 1485 1992 1991 1142 2001 2035 23 38 2005 OAI33_X1
* cell instance $4631 m0 *1 21.85,77
X$4631 23 38 FILLCELL_X4
* cell instance $4632 m0 *1 22.61,77
X$4632 2002 1446 1822 23 38 2036 MUX2_X1
* cell instance $4633 m0 *1 23.94,77
X$4633 23 38 FILLCELL_X1
* cell instance $4634 m0 *1 24.13,77
X$4634 2002 1184 1939 23 38 1940 MUX2_X1
* cell instance $4635 m0 *1 25.46,77
X$4635 23 38 FILLCELL_X2
* cell instance $4636 r0 *1 16.53,77
X$4636 1791 1492 2033 23 38 2075 MUX2_X1
* cell instance $4637 r0 *1 17.86,77
X$4637 1937 1434 1820 23 38 1969 MUX2_X1
* cell instance $4638 r0 *1 19.19,77
X$4638 1848 23 38 CLKBUF_X1
* cell instance $4639 r0 *1 19.76,77
X$4639 2048 1537 23 38 1925 NOR2_X1
* cell instance $4640 r0 *1 20.33,77
X$4640 2078 1605 23 38 1970 NOR2_X1
* cell instance $4641 r0 *1 20.9,77
X$4641 23 38 FILLCELL_X1
* cell instance $4642 r0 *1 21.09,77
X$4642 2126 1605 23 38 2001 NOR2_X1
* cell instance $4643 r0 *1 21.66,77
X$4643 23 3014 2002 2036 2145 38 DFF_X1
* cell instance $4644 r0 *1 24.89,77
X$4644 434 23 38 1909 CLKBUF_X3
* cell instance $4645 m0 *1 26.03,77
X$4645 1485 1941 2037 1142 2003 2004 23 38 1971 OAI33_X1
* cell instance $4646 m0 *1 25.84,77
X$4646 23 38 FILLCELL_X1
* cell instance $4647 m0 *1 27.36,77
X$4647 23 38 FILLCELL_X2
* cell instance $4648 r0 *1 25.84,77
X$4648 2080 1605 23 38 2003 NOR2_X1
* cell instance $4649 r0 *1 26.41,77
X$4649 23 38 FILLCELL_X2
* cell instance $4650 r0 *1 26.79,77
X$4650 2049 1537 23 38 2004 NOR2_X1
* cell instance $4651 r0 *1 27.36,77
X$4651 23 38 FILLCELL_X8
* cell instance $4652 m0 *1 28.88,77
X$4652 1971 1972 1511 1787 38 23 2084 OAI22_X2
* cell instance $4653 m0 *1 27.74,77
X$4653 2005 2081 1629 1157 1727 38 23 2039 OAI221_X1
* cell instance $4654 m0 *1 30.59,77
X$4654 23 38 FILLCELL_X1
* cell instance $4655 m0 *1 30.78,77
X$4655 23 2646 1963 2038 1795 38 DFF_X1
* cell instance $4656 m0 *1 34.01,77
X$4656 1485 1910 1911 1142 2040 2006 23 38 2007 OAI33_X1
* cell instance $4657 m0 *1 35.34,77
X$4657 23 38 FILLCELL_X2
* cell instance $4658 r0 *1 28.88,77
X$4658 23 38 FILLCELL_X1
* cell instance $4659 r0 *1 29.07,77
X$4659 2005 2081 1511 1787 38 23 2082 OAI22_X2
* cell instance $4660 r0 *1 30.78,77
X$4660 23 3080 2050 2086 1795 38 DFF_X1
* cell instance $4661 r0 *1 34.01,77
X$4661 1963 1728 23 38 2085 NAND2_X1
* cell instance $4662 r0 *1 34.58,77
X$4662 2088 1537 23 38 2006 NOR2_X1
* cell instance $4663 r0 *1 35.15,77
X$4663 23 38 FILLCELL_X1
* cell instance $4664 r0 *1 35.34,77
X$4664 2051 1605 23 38 2040 NOR2_X1
* cell instance $4665 m0 *1 36.86,77
X$4665 1743 1999 1997 1804 2041 38 23 1966 OAI221_X1
* cell instance $4666 m0 *1 35.72,77
X$4666 2007 2008 1629 1506 1727 38 23 1997 OAI221_X1
* cell instance $4667 m0 *1 38,77
X$4667 1944 1638 23 38 2041 NAND2_X1
* cell instance $4668 m0 *1 38.57,77
X$4668 1944 1728 23 38 2011 NAND2_X1
* cell instance $4669 m0 *1 39.14,77
X$4669 23 38 FILLCELL_X2
* cell instance $4670 r0 *1 35.91,77
X$4670 2007 2008 1511 1787 38 23 2090 OAI22_X2
* cell instance $4671 r0 *1 37.62,77
X$4671 23 38 FILLCELL_X1
* cell instance $4672 r0 *1 37.81,77
X$4672 2091 1537 23 38 2009 NOR2_X1
* cell instance $4673 r0 *1 38.38,77
X$4673 2090 2010 2011 38 23 2147 OAI21_X2
* cell instance $4674 m0 *1 39.71,77
X$4674 1485 1998 1796 1142 1974 2009 23 38 2012 OAI33_X1
* cell instance $4675 m0 *1 39.52,77
X$4675 23 38 FILLCELL_X1
* cell instance $4676 m0 *1 41.04,77
X$4676 2012 2013 1629 1506 1727 38 23 2043 OAI221_X1
* cell instance $4677 m0 *1 42.18,77
X$4677 1743 1975 2043 1804 2042 38 23 2014 OAI221_X1
* cell instance $4678 m0 *1 43.32,77
X$4678 1945 1728 23 38 2094 NAND2_X1
* cell instance $4679 m0 *1 43.89,77
X$4679 23 38 FILLCELL_X16
* cell instance $4680 m0 *1 46.93,77
X$4680 23 38 FILLCELL_X4
* cell instance $4681 m0 *1 47.69,77
X$4681 23 38 FILLCELL_X1
* cell instance $4682 m0 *1 47.88,77
X$4682 1485 1875 1996 1142 2015 1995 23 38 1976 OAI33_X1
* cell instance $4683 m0 *1 49.21,77
X$4683 1994 1537 23 38 1995 NOR2_X1
* cell instance $4684 m0 *1 49.78,77
X$4684 2044 1605 23 38 2015 NOR2_X1
* cell instance $4685 m0 *1 50.35,77
X$4685 23 38 FILLCELL_X2
* cell instance $4686 r0 *1 39.71,77
X$4686 23 38 FILLCELL_X2
* cell instance $4687 r0 *1 40.09,77
X$4687 1909 23 38 1933 CLKBUF_X3
* cell instance $4688 r0 *1 41.04,77
X$4688 2012 2013 1511 1787 38 23 2093 OAI22_X2
* cell instance $4689 r0 *1 42.75,77
X$4689 2093 2010 2094 38 23 2052 OAI21_X2
* cell instance $4690 r0 *1 44.08,77
X$4690 1933 23 38 CLKBUF_X1
* cell instance $4691 r0 *1 44.65,77
X$4691 23 38 FILLCELL_X2
* cell instance $4692 r0 *1 45.03,77
X$4692 23 38 FILLCELL_X1
* cell instance $4693 r0 *1 45.22,77
X$4693 23 1331 2010 38 BUF_X16
* cell instance $4694 r0 *1 49.97,77
X$4694 23 38 FILLCELL_X2
* cell instance $4695 r0 *1 50.35,77
X$4695 1976 2016 1511 1787 38 23 2097 OAI22_X2
* cell instance $4696 m0 *1 50.92,77
X$4696 1976 2016 1629 1506 1727 38 23 2098 OAI221_X1
* cell instance $4697 m0 *1 50.73,77
X$4697 23 38 FILLCELL_X1
* cell instance $4698 m0 *1 52.06,77
X$4698 23 38 FILLCELL_X2
* cell instance $4699 r0 *1 52.06,77
X$4699 2097 2010 2100 38 23 2183 OAI21_X2
* cell instance $4700 m0 *1 53.01,77
X$4700 1636 1977 23 38 2017 NAND2_X1
* cell instance $4701 m0 *1 52.44,77
X$4701 1977 1728 23 38 2100 NAND2_X1
* cell instance $4702 m0 *1 53.58,77
X$4702 1977 1638 23 38 2018 NAND2_X1
* cell instance $4703 m0 *1 54.15,77
X$4703 23 38 FILLCELL_X1
* cell instance $4704 m0 *1 54.34,77
X$4704 1987 1537 23 38 1978 NOR2_X1
* cell instance $4705 m0 *1 54.91,77
X$4705 1947 2019 1629 1506 1727 38 23 1990 OAI221_X1
* cell instance $4706 m0 *1 56.05,77
X$4706 1636 1948 23 38 1989 NAND2_X1
* cell instance $4707 m0 *1 56.62,77
X$4707 23 38 FILLCELL_X1
* cell instance $4708 m0 *1 56.81,77
X$4708 1767 1492 1979 23 38 2034 MUX2_X1
* cell instance $4709 m0 *1 58.14,77
X$4709 23 2654 1979 2034 1915 38 DFF_X1
* cell instance $4710 m0 *1 61.37,77
X$4710 23 38 FILLCELL_X16
* cell instance $4711 m0 *1 64.41,77
X$4711 23 38 FILLCELL_X1
* cell instance $4712 m0 *1 64.6,77
X$4712 2058 23 38 1915 CLKBUF_X3
* cell instance $4713 m0 *1 65.55,77
X$4713 1915 23 38 3139 INV_X1
* cell instance $4714 m0 *1 65.93,77
X$4714 23 38 FILLCELL_X8
* cell instance $4715 m0 *1 67.45,77
X$4715 23 38 FILLCELL_X4
* cell instance $4716 m0 *1 68.21,77
X$4716 23 38 FILLCELL_X2
* cell instance $4717 r0 *1 53.39,77
X$4717 1743 2017 2098 1804 2018 38 23 1993 OAI221_X1
* cell instance $4718 r0 *1 54.53,77
X$4718 23 38 FILLCELL_X2
* cell instance $4719 r0 *1 54.91,77
X$4719 1947 2019 1511 1787 38 23 2053 OAI22_X2
* cell instance $4720 r0 *1 56.62,77
X$4720 23 38 FILLCELL_X1
* cell instance $4721 r0 *1 56.81,77
X$4721 1519 23 38 1638 CLKBUF_X3
* cell instance $4722 r0 *1 57.76,77
X$4722 2054 1605 23 38 1956 NOR2_X1
* cell instance $4723 r0 *1 58.33,77
X$4723 1948 1728 23 38 2103 NAND2_X1
* cell instance $4724 r0 *1 58.9,77
X$4724 23 38 FILLCELL_X32
* cell instance $4725 r0 *1 59.14,77
X$4725 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $4726 r0 *1 59.14,77
X$4726 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $4727 r0 *1 59.14,77
X$4727 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $4728 r0 *1 64.98,77
X$4728 2104 23 38 1456 BUF_X2
* cell instance $4729 r0 *1 65.74,77
X$4729 23 38 FILLCELL_X4
* cell instance $4730 r0 *1 66.5,77
X$4730 23 38 FILLCELL_X1
* cell instance $4731 r0 *1 66.69,77
X$4731 2021 23 38 1494 CLKBUF_X2
* cell instance $4732 r0 *1 67.45,77
X$4732 23 38 FILLCELL_X8
* cell instance $4733 m0 *1 71.82,77
X$4733 1982 23 38 1219 BUF_X2
* cell instance $4734 m0 *1 68.59,77
X$4734 23 2587 1355 1980 1981 38 DFF_X1
* cell instance $4735 m0 *1 72.58,77
X$4735 23 38 FILLCELL_X16
* cell instance $4736 m0 *1 75.62,77
X$4736 23 38 FILLCELL_X8
* cell instance $4737 m0 *1 77.14,77
X$4737 23 38 FILLCELL_X4
* cell instance $4738 m0 *1 77.9,77
X$4738 23 38 FILLCELL_X2
* cell instance $4739 r0 *1 68.97,77
X$4739 23 38 FILLCELL_X4
* cell instance $4740 r0 *1 69.73,77
X$4740 23 2922 2021 2099 1981 38 DFF_X1
* cell instance $4741 r0 *1 72.96,77
X$4741 23 38 FILLCELL_X32
* cell instance $4742 m0 *1 78.47,77
X$4742 1478 23 38 1983 INV_X2
* cell instance $4743 m0 *1 78.28,77
X$4743 23 38 FILLCELL_X1
* cell instance $4744 m0 *1 79.04,77
X$4744 1983 23 38 1949 CLKBUF_X3
* cell instance $4745 m0 *1 79.99,77
X$4745 1983 1519 1318 23 38 NOR2_X4
* cell instance $4746 m0 *1 81.7,77
X$4746 1951 38 1198 23 BUF_X4
* cell instance $4747 m0 *1 83.03,77
X$4747 23 38 FILLCELL_X16
* cell instance $4748 m0 *1 86.07,77
X$4748 23 38 FILLCELL_X8
* cell instance $4749 m0 *1 87.59,77
X$4749 23 38 FILLCELL_X4
* cell instance $4750 m0 *1 88.35,77
X$4750 2023 1460 38 23 2024 AND2_X1
* cell instance $4751 m0 *1 89.11,77
X$4751 23 38 FILLCELL_X16
* cell instance $4752 m0 *1 92.15,77
X$4752 23 38 FILLCELL_X8
* cell instance $4753 m0 *1 93.67,77
X$4753 23 38 FILLCELL_X2
* cell instance $4754 r0 *1 79.04,77
X$4754 23 38 FILLCELL_X4
* cell instance $4755 r0 *1 79.8,77
X$4755 1983 38 1319 23 BUF_X4
* cell instance $4756 r0 *1 81.13,77
X$4756 1951 38 1240 23 BUF_X4
* cell instance $4757 r0 *1 82.46,77
X$4757 23 38 FILLCELL_X4
* cell instance $4758 r0 *1 83.22,77
X$4758 23 38 FILLCELL_X2
* cell instance $4759 r0 *1 83.6,77
X$4759 23 38 FILLCELL_X1
* cell instance $4760 r0 *1 83.79,77
X$4760 2058 23 38 1917 CLKBUF_X3
* cell instance $4761 r0 *1 84.74,77
X$4761 1917 23 38 3152 INV_X1
* cell instance $4762 r0 *1 85.12,77
X$4762 23 38 FILLCELL_X1
* cell instance $4763 r0 *1 85.31,77
X$4763 2089 2025 2032 23 38 2092 MUX2_X1
* cell instance $4764 r0 *1 86.64,77
X$4764 2022 1460 38 23 2032 AND2_X1
* cell instance $4765 r0 *1 87.4,77
X$4765 23 38 FILLCELL_X2
* cell instance $4766 r0 *1 87.78,77
X$4766 23 38 FILLCELL_X1
* cell instance $4767 r0 *1 87.97,77
X$4767 2118 2025 2024 23 38 2079 MUX2_X1
* cell instance $4768 r0 *1 89.3,77
X$4768 23 2079 2026 3132 2023 38 DFF_X2
* cell instance $4769 r0 *1 92.91,77
X$4769 23 3105 2064 2067 2026 38 DFF_X1
* cell instance $4770 m0 *1 94.81,77
X$4770 23 38 FILLCELL_X4
* cell instance $4771 m0 *1 94.05,77
X$4771 1226 2030 2025 23 1986 38 AOI21_X1
* cell instance $4772 m0 *1 95.57,77
X$4772 23 38 FILLCELL_X1
* cell instance $4773 m0 *1 95.76,77
X$4773 2027 1985 23 38 2030 NAND2_X1
* cell instance $4774 m0 *1 96.33,77
X$4774 23 38 FILLCELL_X1
* cell instance $4775 m0 *1 96.52,77
X$4775 1985 23 38 2028 BUF_X1
* cell instance $4776 r180 *1 97.28,77
X$4776 23 38 23 38 TAPCELL_X1
* cell instance $4777 r0 *1 96.14,77
X$4777 23 38 FILLCELL_X2
* cell instance $4778 r0 *1 96.52,77
X$4778 2068 23 38 2027 INV_X1
* cell instance $4779 r0 *1 96.9,77
X$4779 23 38 FILLCELL_X1
* cell instance $4780 m90 *1 97.28,77
X$4780 23 38 23 38 TAPCELL_X1
* cell instance $4781 m0 *1 1.33,23.8
X$4781 23 38 FILLCELL_X4
* cell instance $4782 m0 *1 1.14,23.8
X$4782 23 38 23 38 TAPCELL_X1
* cell instance $4783 m0 *1 2.09,23.8
X$4783 23 38 FILLCELL_X1
* cell instance $4784 m0 *1 2.28,23.8
X$4784 23 2750 610 569 447 38 DFF_X1
* cell instance $4785 m0 *1 5.51,23.8
X$4785 23 38 FILLCELL_X2
* cell instance $4786 r0 *1 1.14,23.8
X$4786 23 38 23 38 TAPCELL_X1
* cell instance $4787 r0 *1 1.33,23.8
X$4787 23 38 FILLCELL_X8
* cell instance $4788 r0 *1 2.85,23.8
X$4788 23 38 FILLCELL_X4
* cell instance $4789 r0 *1 3.14,23.8
X$4789 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $4790 r0 *1 3.14,23.8
X$4790 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $4791 r0 *1 3.14,23.8
X$4791 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $4792 r0 *1 3.61,23.8
X$4792 23 38 FILLCELL_X2
* cell instance $4793 r0 *1 3.99,23.8
X$4793 590 318 591 23 38 589 MUX2_X1
* cell instance $4794 r0 *1 5.32,23.8
X$4794 23 38 FILLCELL_X2
* cell instance $4795 r0 *1 5.7,23.8
X$4795 23 38 FILLCELL_X1
* cell instance $4796 r0 *1 5.89,23.8
X$4796 610 257 591 23 38 569 MUX2_X1
* cell instance $4797 m0 *1 7.22,23.8
X$4797 23 38 FILLCELL_X4
* cell instance $4798 m0 *1 5.89,23.8
X$4798 590 412 610 23 38 528 MUX2_X1
* cell instance $4799 m0 *1 7.98,23.8
X$4799 23 2746 592 571 447 38 DFF_X1
* cell instance $4800 m0 *1 11.21,23.8
X$4800 592 437 591 23 38 571 MUX2_X1
* cell instance $4801 m0 *1 12.54,23.8
X$4801 356 594 547 548 431 297 23 38 614 OAI33_X1
* cell instance $4802 m0 *1 13.87,23.8
X$4802 23 38 FILLCELL_X8
* cell instance $4803 m0 *1 15.39,23.8
X$4803 23 38 FILLCELL_X2
* cell instance $4804 r0 *1 7.22,23.8
X$4804 23 38 FILLCELL_X8
* cell instance $4805 r0 *1 8.74,23.8
X$4805 23 38 FILLCELL_X2
* cell instance $4806 r0 *1 9.12,23.8
X$4806 23 2981 593 611 503 38 DFF_X1
* cell instance $4807 r0 *1 12.35,23.8
X$4807 593 393 591 23 38 611 MUX2_X1
* cell instance $4808 r0 *1 13.68,23.8
X$4808 595 381 23 38 594 NOR2_X1
* cell instance $4809 r0 *1 14.25,23.8
X$4809 23 38 FILLCELL_X4
* cell instance $4810 r0 *1 15.01,23.8
X$4810 23 38 FILLCELL_X2
* cell instance $4811 r0 *1 15.39,23.8
X$4811 23 2992 549 574 503 38 DFF_X1
* cell instance $4812 m0 *1 17.1,23.8
X$4812 23 38 FILLCELL_X4
* cell instance $4813 m0 *1 15.77,23.8
X$4813 549 393 502 23 38 574 MUX2_X1
* cell instance $4814 m0 *1 17.86,23.8
X$4814 23 2740 504 550 503 38 DFF_X1
* cell instance $4815 m0 *1 21.09,23.8
X$4815 23 38 FILLCELL_X8
* cell instance $4816 m0 *1 22.61,23.8
X$4816 23 38 FILLCELL_X4
* cell instance $4817 m0 *1 23.37,23.8
X$4817 23 38 FILLCELL_X1
* cell instance $4818 m0 *1 23.56,23.8
X$4818 576 437 358 23 38 615 MUX2_X1
* cell instance $4819 m0 *1 24.89,23.8
X$4819 23 38 FILLCELL_X2
* cell instance $4820 r0 *1 18.62,23.8
X$4820 23 38 FILLCELL_X16
* cell instance $4821 r0 *1 21.66,23.8
X$4821 23 38 FILLCELL_X2
* cell instance $4822 r0 *1 22.04,23.8
X$4822 23 38 FILLCELL_X1
* cell instance $4823 r0 *1 22.23,23.8
X$4823 23 2993 576 615 653 38 DFF_X1
* cell instance $4824 m0 *1 25.46,23.8
X$4824 507 393 421 23 38 506 MUX2_X1
* cell instance $4825 m0 *1 25.27,23.8
X$4825 23 38 FILLCELL_X1
* cell instance $4826 m0 *1 26.79,23.8
X$4826 23 38 FILLCELL_X4
* cell instance $4827 m0 *1 27.55,23.8
X$4827 23 38 FILLCELL_X2
* cell instance $4828 r0 *1 25.46,23.8
X$4828 23 38 FILLCELL_X32
* cell instance $4829 m0 *1 31.16,23.8
X$4829 23 38 FILLCELL_X2
* cell instance $4830 m0 *1 27.93,23.8
X$4830 23 2783 551 508 329 38 DFF_X1
* cell instance $4831 m0 *1 31.73,23.8
X$4831 509 257 510 23 38 596 MUX2_X1
* cell instance $4832 m0 *1 31.54,23.8
X$4832 23 38 FILLCELL_X1
* cell instance $4833 m0 *1 33.06,23.8
X$4833 23 38 FILLCELL_X1
* cell instance $4834 m0 *1 33.25,23.8
X$4834 149 23 38 329 CLKBUF_X3
* cell instance $4835 m0 *1 34.2,23.8
X$4835 23 2749 540 552 329 38 DFF_X1
* cell instance $4836 m0 *1 37.43,23.8
X$4836 554 393 319 23 38 553 MUX2_X1
* cell instance $4837 m0 *1 38.76,23.8
X$4837 578 437 319 23 38 542 MUX2_X1
* cell instance $4838 m0 *1 40.09,23.8
X$4838 554 472 578 23 38 579 MUX2_X1
* cell instance $4839 m0 *1 41.42,23.8
X$4839 23 38 FILLCELL_X4
* cell instance $4840 m0 *1 42.18,23.8
X$4840 23 38 FILLCELL_X2
* cell instance $4841 r0 *1 31.54,23.8
X$4841 23 38 FILLCELL_X1
* cell instance $4842 r0 *1 31.73,23.8
X$4842 23 2950 509 596 329 38 DFF_X1
* cell instance $4843 r0 *1 34.96,23.8
X$4843 23 38 FILLCELL_X32
* cell instance $4844 r0 *1 41.04,23.8
X$4844 23 38 FILLCELL_X2
* cell instance $4845 r0 *1 41.42,23.8
X$4845 23 38 FILLCELL_X1
* cell instance $4846 r0 *1 41.61,23.8
X$4846 620 38 602 23 BUF_X4
* cell instance $4847 m0 *1 42.75,23.8
X$4847 23 2743 512 581 299 38 DFF_X1
* cell instance $4848 m0 *1 42.56,23.8
X$4848 23 38 FILLCELL_X1
* cell instance $4849 m0 *1 45.98,23.8
X$4849 23 38 FILLCELL_X4
* cell instance $4850 m0 *1 46.74,23.8
X$4850 23 38 FILLCELL_X1
* cell instance $4851 m0 *1 46.93,23.8
X$4851 620 23 38 472 CLKBUF_X3
* cell instance $4852 m0 *1 47.88,23.8
X$4852 599 23 38 437 CLKBUF_X3
* cell instance $4853 m0 *1 48.83,23.8
X$4853 557 38 257 23 BUF_X4
* cell instance $4854 m0 *1 50.16,23.8
X$4854 513 598 556 23 38 545 MUX2_X1
* cell instance $4855 m0 *1 51.49,23.8
X$4855 555 599 556 23 38 621 MUX2_X1
* cell instance $4856 m0 *1 52.82,23.8
X$4856 23 38 FILLCELL_X1
* cell instance $4857 m0 *1 53.01,23.8
X$4857 558 597 556 23 38 586 MUX2_X1
* cell instance $4858 m0 *1 54.34,23.8
X$4858 514 557 556 23 38 499 MUX2_X1
* cell instance $4859 m0 *1 55.67,23.8
X$4859 23 38 FILLCELL_X1
* cell instance $4860 m0 *1 55.86,23.8
X$4860 558 305 514 23 38 588 MUX2_X1
* cell instance $4861 m0 *1 57.19,23.8
X$4861 23 38 FILLCELL_X2
* cell instance $4862 r0 *1 42.94,23.8
X$4862 75 23 38 398 BUF_X2
* cell instance $4863 r0 *1 43.7,23.8
X$4863 23 38 FILLCELL_X8
* cell instance $4864 r0 *1 45.22,23.8
X$4864 23 38 FILLCELL_X4
* cell instance $4865 r0 *1 45.98,23.8
X$4865 23 38 FILLCELL_X2
* cell instance $4866 r0 *1 46.36,23.8
X$4866 598 23 38 393 CLKBUF_X3
* cell instance $4867 r0 *1 47.31,23.8
X$4867 23 38 FILLCELL_X4
* cell instance $4868 r0 *1 48.07,23.8
X$4868 23 38 FILLCELL_X1
* cell instance $4869 r0 *1 48.26,23.8
X$4869 597 38 318 23 BUF_X4
* cell instance $4870 r0 *1 49.59,23.8
X$4870 23 38 FILLCELL_X2
* cell instance $4871 r0 *1 49.97,23.8
X$4871 23 38 FILLCELL_X1
* cell instance $4872 r0 *1 50.16,23.8
X$4872 23 2913 555 621 158 38 DFF_X1
* cell instance $4873 r0 *1 53.39,23.8
X$4873 23 38 FILLCELL_X4
* cell instance $4874 r0 *1 54.15,23.8
X$4874 23 38 FILLCELL_X2
* cell instance $4875 r0 *1 54.53,23.8
X$4875 112 23 38 556 BUF_X2
* cell instance $4876 r0 *1 55.29,23.8
X$4876 23 38 FILLCELL_X2
* cell instance $4877 r0 *1 55.67,23.8
X$4877 23 38 FILLCELL_X1
* cell instance $4878 r0 *1 55.86,23.8
X$4878 600 38 548 23 BUF_X4
* cell instance $4879 r0 *1 57.19,23.8
X$4879 23 38 FILLCELL_X8
* cell instance $4880 m0 *1 58.52,23.8
X$4880 23 38 FILLCELL_X8
* cell instance $4881 m0 *1 57.57,23.8
X$4881 600 23 38 360 CLKBUF_X3
* cell instance $4882 m0 *1 60.04,23.8
X$4882 23 38 FILLCELL_X2
* cell instance $4883 r0 *1 58.71,23.8
X$4883 23 38 FILLCELL_X4
* cell instance $4884 r0 *1 59.14,23.8
X$4884 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $4885 r0 *1 59.14,23.8
X$4885 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $4886 r0 *1 59.14,23.8
X$4886 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $4887 r0 *1 59.47,23.8
X$4887 639 367 23 38 622 NOR2_X1
* cell instance $4888 r0 *1 60.04,23.8
X$4888 23 38 FILLCELL_X8
* cell instance $4889 m0 *1 60.99,23.8
X$4889 585 559 48 23 38 584 MUX2_X1
* cell instance $4890 m0 *1 60.42,23.8
X$4890 473 372 23 38 623 NOR2_X1
* cell instance $4891 m0 *1 62.32,23.8
X$4891 585 602 519 23 38 583 MUX2_X1
* cell instance $4892 m0 *1 63.65,23.8
X$4892 23 38 FILLCELL_X4
* cell instance $4893 m0 *1 64.41,23.8
X$4893 23 38 FILLCELL_X1
* cell instance $4894 m0 *1 64.6,23.8
X$4894 583 367 23 38 560 NOR2_X1
* cell instance $4895 m0 *1 65.17,23.8
X$4895 23 38 FILLCELL_X2
* cell instance $4896 r0 *1 61.56,23.8
X$4896 656 370 23 38 601 NOR2_X1
* cell instance $4897 r0 *1 62.13,23.8
X$4897 515 601 622 600 623 603 23 38 624 OAI33_X1
* cell instance $4898 r0 *1 63.46,23.8
X$4898 23 38 FILLCELL_X4
* cell instance $4899 r0 *1 64.22,23.8
X$4899 23 38 FILLCELL_X2
* cell instance $4900 r0 *1 64.6,23.8
X$4900 23 38 FILLCELL_X1
* cell instance $4901 r0 *1 64.79,23.8
X$4901 543 23 38 CLKBUF_X1
* cell instance $4902 r0 *1 65.36,23.8
X$4902 23 38 FILLCELL_X16
* cell instance $4903 m0 *1 65.74,23.8
X$4903 23 2797 538 582 543 38 DFF_X1
* cell instance $4904 m0 *1 65.55,23.8
X$4904 23 38 FILLCELL_X1
* cell instance $4905 m0 *1 68.97,23.8
X$4905 561 559 78 23 38 604 MUX2_X1
* cell instance $4906 m0 *1 70.3,23.8
X$4906 23 38 FILLCELL_X8
* cell instance $4907 m0 *1 71.82,23.8
X$4907 23 38 FILLCELL_X2
* cell instance $4908 r0 *1 68.4,23.8
X$4908 23 38 FILLCELL_X1
* cell instance $4909 r0 *1 68.59,23.8
X$4909 23 2919 561 604 543 38 DFF_X1
* cell instance $4910 r0 *1 71.82,23.8
X$4910 23 38 FILLCELL_X2
* cell instance $4911 r0 *1 1.33,1.4
X$4911 23 38 FILLCELL_X32
* cell instance $4912 r0 *1 1.14,1.4
X$4912 23 38 23 38 TAPCELL_X1
* cell instance $4913 r0 *1 7.41,1.4
X$4913 23 38 FILLCELL_X4
* cell instance $4914 r0 *1 8.17,1.4
X$4914 23 38 FILLCELL_X1
* cell instance $4915 r0 *1 9.12,1.4
X$4915 23 38 FILLCELL_X2
* cell instance $4916 r0 *1 3.14,1.4
X$4916 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $4917 r0 *1 3.14,1.4
X$4917 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $4918 r0 *1 3.14,1.4
X$4918 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $4919 m90 *1 97.28,26.6
X$4919 23 38 23 38 TAPCELL_X1
* cell instance $4920 r180 *1 97.28,26.6
X$4920 23 38 23 38 TAPCELL_X1
* cell instance $4921 r180 *1 97.28,96.6
X$4921 23 38 23 38 TAPCELL_X1
* cell instance $4922 m0 *1 96.9,96.6
X$4922 23 38 FILLCELL_X1
* cell instance $4923 r180 *1 97.28,29.4
X$4923 23 38 23 38 TAPCELL_X1
* cell instance $4924 m90 *1 97.28,29.4
X$4924 23 38 23 38 TAPCELL_X1
* cell instance $4925 m0 *1 1.33,4.2
X$4925 23 38 FILLCELL_X32
* cell instance $4926 m0 *1 1.14,4.2
X$4926 23 38 23 38 TAPCELL_X1
* cell instance $4927 m0 *1 7.41,4.2
X$4927 23 38 FILLCELL_X8
* cell instance $4928 m0 *1 8.93,4.2
X$4928 23 38 FILLCELL_X4
* cell instance $4929 m0 *1 9.69,4.2
X$4929 23 38 FILLCELL_X1
* cell instance $4930 m0 *1 13.11,4.2
X$4930 23 38 FILLCELL_X2
* cell instance $4931 r0 *1 1.14,4.2
X$4931 23 38 23 38 TAPCELL_X1
* cell instance $4932 r0 *1 1.33,4.2
X$4932 23 38 FILLCELL_X32
* cell instance $4933 r0 *1 3.14,4.2
X$4933 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $4934 r0 *1 3.14,4.2
X$4934 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $4935 r0 *1 3.14,4.2
X$4935 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $4936 r0 *1 7.41,4.2
X$4936 23 38 FILLCELL_X16
* cell instance $4937 r0 *1 10.45,4.2
X$4937 23 38 FILLCELL_X1
* cell instance $4938 r0 *1 10.64,4.2
X$4938 107 42 69 23 38 55 MUX2_X1
* cell instance $4939 r0 *1 11.97,4.2
X$4939 23 38 FILLCELL_X2
* cell instance $4940 r0 *1 12.35,4.2
X$4940 23 38 FILLCELL_X1
* cell instance $4941 r0 *1 12.54,4.2
X$4941 107 40 87 23 38 114 MUX2_X1
* cell instance $4942 m0 *1 14.82,4.2
X$4942 23 38 FILLCELL_X4
* cell instance $4943 m0 *1 15.58,4.2
X$4943 23 2757 71 41 28 38 DFF_X1
* cell instance $4944 m0 *1 18.81,4.2
X$4944 23 38 FILLCELL_X4
* cell instance $4945 m0 *1 19.57,4.2
X$4945 23 38 FILLCELL_X1
* cell instance $4946 m0 *1 19.76,4.2
X$4946 23 2760 43 57 28 38 DFF_X1
* cell instance $4947 m0 *1 22.99,4.2
X$4947 23 38 FILLCELL_X8
* cell instance $4948 m0 *1 24.51,4.2
X$4948 23 38 FILLCELL_X2
* cell instance $4949 r0 *1 13.87,4.2
X$4949 69 70 87 23 38 247 MUX2_X1
* cell instance $4950 r0 *1 15.2,4.2
X$4950 23 38 FILLCELL_X1
* cell instance $4951 r0 *1 15.39,4.2
X$4951 27 42 71 23 38 41 MUX2_X1
* cell instance $4952 r0 *1 16.72,4.2
X$4952 23 38 FILLCELL_X2
* cell instance $4953 r0 *1 17.1,4.2
X$4953 71 70 56 23 38 204 MUX2_X1
* cell instance $4954 r0 *1 18.43,4.2
X$4954 23 3030 131 93 28 38 DFF_X1
* cell instance $4955 r0 *1 21.66,4.2
X$4955 24 40 43 23 38 57 MUX2_X1
* cell instance $4956 r0 *1 22.99,4.2
X$4956 23 38 FILLCELL_X4
* cell instance $4957 r0 *1 23.75,4.2
X$4957 23 38 FILLCELL_X2
* cell instance $4958 r0 *1 24.13,4.2
X$4958 23 38 FILLCELL_X1
* cell instance $4959 m0 *1 26.22,4.2
X$4959 23 38 FILLCELL_X4
* cell instance $4960 m0 *1 26.98,4.2
X$4960 23 38 FILLCELL_X1
* cell instance $4961 m0 *1 27.17,4.2
X$4961 29 40 59 23 38 58 MUX2_X1
* cell instance $4962 m0 *1 28.5,4.2
X$4962 23 2765 59 58 73 38 DFF_X1
* cell instance $4963 m0 *1 31.73,4.2
X$4963 23 38 FILLCELL_X32
* cell instance $4964 m0 *1 37.81,4.2
X$4964 23 38 FILLCELL_X4
* cell instance $4965 m0 *1 38.57,4.2
X$4965 23 2700 44 61 74 38 DFF_X1
* cell instance $4966 m0 *1 41.8,4.2
X$4966 23 38 FILLCELL_X4
* cell instance $4967 m0 *1 42.56,4.2
X$4967 23 38 FILLCELL_X2
* cell instance $4968 r0 *1 27.55,4.2
X$4968 23 38 FILLCELL_X4
* cell instance $4969 r0 *1 28.31,4.2
X$4969 23 38 FILLCELL_X2
* cell instance $4970 r0 *1 28.69,4.2
X$4970 23 38 FILLCELL_X1
* cell instance $4971 r0 *1 28.88,4.2
X$4971 23 2932 116 96 73 38 DFF_X1
* cell instance $4972 r0 *1 32.11,4.2
X$4972 23 2894 117 111 74 38 DFF_X1
* cell instance $4973 r0 *1 35.34,4.2
X$4973 25 40 118 23 38 97 MUX2_X1
* cell instance $4974 r0 *1 36.67,4.2
X$4974 23 2885 119 89 74 38 DFF_X1
* cell instance $4975 r0 *1 39.9,4.2
X$4975 98 40 44 23 38 61 MUX2_X1
* cell instance $4976 r0 *1 41.23,4.2
X$4976 23 38 FILLCELL_X4
* cell instance $4977 r0 *1 41.99,4.2
X$4977 23 38 FILLCELL_X1
* cell instance $4978 r0 *1 42.18,4.2
X$4978 23 2905 120 91 30 38 DFF_X1
* cell instance $4979 m0 *1 46.17,4.2
X$4979 23 38 FILLCELL_X8
* cell instance $4980 m0 *1 42.94,4.2
X$4980 23 2707 31 62 30 38 DFF_X1
* cell instance $4981 m0 *1 47.69,4.2
X$4981 23 2722 45 64 30 38 DFF_X1
* cell instance $4982 m0 *1 50.92,4.2
X$4982 23 38 FILLCELL_X8
* cell instance $4983 m0 *1 52.44,4.2
X$4983 23 38 FILLCELL_X4
* cell instance $4984 m0 *1 53.2,4.2
X$4984 23 38 FILLCELL_X2
* cell instance $4985 r0 *1 45.41,4.2
X$4985 75 40 31 23 38 62 MUX2_X1
* cell instance $4986 r0 *1 46.74,4.2
X$4986 23 38 FILLCELL_X4
* cell instance $4987 r0 *1 47.5,4.2
X$4987 23 38 FILLCELL_X2
* cell instance $4988 r0 *1 47.88,4.2
X$4988 23 3091 99 92 76 38 DFF_X1
* cell instance $4989 r0 *1 51.11,4.2
X$4989 66 40 45 23 38 64 MUX2_X1
* cell instance $4990 r0 *1 52.44,4.2
X$4990 23 38 FILLCELL_X4
* cell instance $4991 r0 *1 53.2,4.2
X$4991 23 2957 135 113 76 38 DFF_X1
* cell instance $4992 m0 *1 54.53,4.2
X$4992 23 2671 46 67 76 38 DFF_X1
* cell instance $4993 m0 *1 53.58,4.2
X$4993 68 23 38 40 CLKBUF_X3
* cell instance $4994 m0 *1 57.76,4.2
X$4994 23 38 FILLCELL_X8
* cell instance $4995 m0 *1 59.28,4.2
X$4995 23 38 FILLCELL_X1
* cell instance $4996 m0 *1 59.47,4.2
X$4996 23 2715 122 102 32 38 DFF_X1
* cell instance $4997 m0 *1 62.7,4.2
X$4997 23 38 FILLCELL_X4
* cell instance $4998 m0 *1 63.46,4.2
X$4998 23 38 FILLCELL_X1
* cell instance $4999 m0 *1 63.65,4.2
X$4999 23 2684 47 65 32 38 DFF_X1
* cell instance $5000 m0 *1 69.54,4.2
X$5000 23 38 FILLCELL_X2
* cell instance $5001 r0 *1 56.43,4.2
X$5001 112 68 46 23 38 67 MUX2_X1
* cell instance $5002 r0 *1 57.76,4.2
X$5002 23 38 FILLCELL_X1
* cell instance $5003 r0 *1 57.95,4.2
X$5003 23 2967 103 101 76 38 DFF_X1
* cell instance $5004 r0 *1 59.14,4.2
X$5004 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $5005 r0 *1 59.14,4.2
X$5005 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $5006 r0 *1 59.14,4.2
X$5006 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $5007 r0 *1 61.18,4.2
X$5007 23 38 FILLCELL_X8
* cell instance $5008 r0 *1 62.7,4.2
X$5008 48 51 90 23 38 104 MUX2_X1
* cell instance $5009 r0 *1 64.03,4.2
X$5009 32 23 38 CLKBUF_X1
* cell instance $5010 r0 *1 64.6,4.2
X$5010 90 80 47 23 38 105 MUX2_X1
* cell instance $5011 r0 *1 65.93,4.2
X$5011 68 38 79 23 BUF_X4
* cell instance $5012 r0 *1 67.26,4.2
X$5012 77 23 38 48 CLKBUF_X2
* cell instance $5013 r0 *1 68.02,4.2
X$5013 23 38 FILLCELL_X8
* cell instance $5014 r0 *1 69.54,4.2
X$5014 23 38 FILLCELL_X2
* cell instance $5015 m0 *1 1.33,7
X$5015 23 38 FILLCELL_X32
* cell instance $5016 m0 *1 1.14,7
X$5016 23 38 23 38 TAPCELL_X1
* cell instance $5017 m0 *1 7.41,7
X$5017 23 38 FILLCELL_X1
* cell instance $5018 m0 *1 10.83,7
X$5018 154 42 106 23 38 129 MUX2_X1
* cell instance $5019 m0 *1 12.16,7
X$5019 23 38 FILLCELL_X2
* cell instance $5020 r0 *1 1.14,7
X$5020 23 38 23 38 TAPCELL_X1
* cell instance $5021 r0 *1 1.33,7
X$5021 23 38 FILLCELL_X32
* cell instance $5022 r0 *1 3.14,7
X$5022 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $5023 r0 *1 3.14,7
X$5023 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $5024 r0 *1 3.14,7
X$5024 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $5025 r0 *1 7.41,7
X$5025 23 38 FILLCELL_X4
* cell instance $5026 r0 *1 8.17,7
X$5026 23 38 FILLCELL_X2
* cell instance $5027 r0 *1 8.55,7
X$5027 23 38 FILLCELL_X1
* cell instance $5028 r0 *1 8.74,7
X$5028 23 3032 148 147 28 38 DFF_X1
* cell instance $5029 r0 *1 11.97,7
X$5029 154 40 148 23 38 147 MUX2_X1
* cell instance $5030 m0 *1 15.77,7
X$5030 23 38 FILLCELL_X1
* cell instance $5031 m0 *1 12.54,7
X$5031 23 2781 87 114 28 38 DFF_X1
* cell instance $5032 m0 *1 15.96,7
X$5032 149 23 38 28 CLKBUF_X3
* cell instance $5033 m0 *1 16.91,7
X$5033 23 38 FILLCELL_X8
* cell instance $5034 m0 *1 18.43,7
X$5034 23 38 FILLCELL_X1
* cell instance $5035 m0 *1 18.62,7
X$5035 24 42 131 23 38 93 MUX2_X1
* cell instance $5036 m0 *1 19.95,7
X$5036 23 38 FILLCELL_X4
* cell instance $5037 m0 *1 20.71,7
X$5037 23 38 FILLCELL_X2
* cell instance $5038 r0 *1 13.3,7
X$5038 23 38 FILLCELL_X8
* cell instance $5039 r0 *1 14.82,7
X$5039 23 3029 136 156 28 38 DFF_X1
* cell instance $5040 r0 *1 18.05,7
X$5040 23 38 FILLCELL_X16
* cell instance $5041 m0 *1 21.28,7
X$5041 131 70 43 23 38 94 MUX2_X1
* cell instance $5042 m0 *1 21.09,7
X$5042 23 38 FILLCELL_X1
* cell instance $5043 m0 *1 22.61,7
X$5043 23 38 FILLCELL_X8
* cell instance $5044 m0 *1 24.13,7
X$5044 23 38 FILLCELL_X1
* cell instance $5045 m0 *1 24.32,7
X$5045 26 40 115 23 38 72 MUX2_X1
* cell instance $5046 m0 *1 26.98,7
X$5046 23 38 FILLCELL_X8
* cell instance $5047 m0 *1 28.5,7
X$5047 23 38 FILLCELL_X2
* cell instance $5048 r0 *1 21.09,7
X$5048 23 38 FILLCELL_X8
* cell instance $5049 r0 *1 22.61,7
X$5049 23 38 FILLCELL_X2
* cell instance $5050 r0 *1 22.99,7
X$5050 23 38 FILLCELL_X1
* cell instance $5051 r0 *1 24.13,7
X$5051 23 38 FILLCELL_X32
* cell instance $5052 m0 *1 29.07,7
X$5052 29 42 116 23 38 96 MUX2_X1
* cell instance $5053 m0 *1 28.88,7
X$5053 23 38 FILLCELL_X1
* cell instance $5054 m0 *1 30.4,7
X$5054 23 38 FILLCELL_X1
* cell instance $5055 m0 *1 30.59,7
X$5055 116 70 59 23 38 278 MUX2_X1
* cell instance $5056 m0 *1 31.92,7
X$5056 23 38 FILLCELL_X2
* cell instance $5057 r0 *1 30.21,7
X$5057 23 38 FILLCELL_X32
* cell instance $5058 m0 *1 32.49,7
X$5058 25 42 117 23 38 111 MUX2_X1
* cell instance $5059 m0 *1 32.3,7
X$5059 23 38 FILLCELL_X1
* cell instance $5060 m0 *1 33.82,7
X$5060 117 70 118 23 38 211 MUX2_X1
* cell instance $5061 m0 *1 35.15,7
X$5061 23 38 FILLCELL_X4
* cell instance $5062 m0 *1 35.91,7
X$5062 23 2759 118 97 74 38 DFF_X1
* cell instance $5063 m0 *1 39.14,7
X$5063 98 42 119 23 38 89 MUX2_X1
* cell instance $5064 m0 *1 40.47,7
X$5064 23 38 FILLCELL_X1
* cell instance $5065 m0 *1 40.66,7
X$5065 119 80 44 23 38 256 MUX2_X1
* cell instance $5066 m0 *1 41.99,7
X$5066 23 38 FILLCELL_X4
* cell instance $5067 m0 *1 42.75,7
X$5067 23 38 FILLCELL_X2
* cell instance $5068 r0 *1 36.29,7
X$5068 23 38 FILLCELL_X4
* cell instance $5069 r0 *1 37.05,7
X$5069 23 38 FILLCELL_X1
* cell instance $5070 r0 *1 37.24,7
X$5070 149 23 38 74 CLKBUF_X3
* cell instance $5071 r0 *1 38.19,7
X$5071 23 38 FILLCELL_X32
* cell instance $5072 m0 *1 43.32,7
X$5072 75 42 120 23 38 91 MUX2_X1
* cell instance $5073 m0 *1 43.13,7
X$5073 23 38 FILLCELL_X1
* cell instance $5074 m0 *1 44.65,7
X$5074 120 80 31 23 38 351 MUX2_X1
* cell instance $5075 m0 *1 45.98,7
X$5075 23 38 FILLCELL_X16
* cell instance $5076 m0 *1 49.02,7
X$5076 66 42 99 23 38 92 MUX2_X1
* cell instance $5077 m0 *1 50.35,7
X$5077 99 80 45 23 38 100 MUX2_X1
* cell instance $5078 m0 *1 51.68,7
X$5078 23 38 FILLCELL_X8
* cell instance $5079 m0 *1 53.2,7
X$5079 138 23 38 42 CLKBUF_X3
* cell instance $5080 m0 *1 54.15,7
X$5080 112 138 135 23 38 113 MUX2_X1
* cell instance $5081 m0 *1 55.48,7
X$5081 23 38 FILLCELL_X4
* cell instance $5082 m0 *1 56.24,7
X$5082 23 38 FILLCELL_X1
* cell instance $5083 m0 *1 56.43,7
X$5083 135 80 46 23 38 134 MUX2_X1
* cell instance $5084 m0 *1 57.76,7
X$5084 23 38 FILLCELL_X1
* cell instance $5085 m0 *1 57.95,7
X$5085 121 138 103 23 38 101 MUX2_X1
* cell instance $5086 m0 *1 59.28,7
X$5086 23 38 FILLCELL_X1
* cell instance $5087 m0 *1 59.47,7
X$5087 121 68 122 23 38 102 MUX2_X1
* cell instance $5088 m0 *1 60.8,7
X$5088 23 38 FILLCELL_X1
* cell instance $5089 m0 *1 60.99,7
X$5089 103 80 122 23 38 123 MUX2_X1
* cell instance $5090 m0 *1 62.32,7
X$5090 23 38 FILLCELL_X1
* cell instance $5091 m0 *1 62.51,7
X$5091 23 2641 90 104 32 38 DFF_X1
* cell instance $5092 m0 *1 65.74,7
X$5092 23 38 FILLCELL_X1
* cell instance $5093 m0 *1 65.93,7
X$5093 23 2645 124 152 32 38 DFF_X1
* cell instance $5094 m0 *1 69.16,7
X$5094 23 38 FILLCELL_X4
* cell instance $5095 m0 *1 69.92,7
X$5095 23 38 FILLCELL_X1
* cell instance $5096 m0 *1 70.11,7
X$5096 77 133 141 23 38 151 MUX2_X1
* cell instance $5097 m0 *1 71.44,7
X$5097 23 38 FILLCELL_X8
* cell instance $5098 m0 *1 72.96,7
X$5098 23 38 FILLCELL_X1
* cell instance $5099 m0 *1 73.15,7
X$5099 23 2698 81 125 34 38 DFF_X1
* cell instance $5100 m0 *1 76.38,7
X$5100 23 38 FILLCELL_X8
* cell instance $5101 m0 *1 77.9,7
X$5101 23 38 FILLCELL_X1
* cell instance $5102 m0 *1 78.09,7
X$5102 23 2636 82 132 36 38 DFF_X1
* cell instance $5103 m0 *1 81.32,7
X$5103 23 38 FILLCELL_X4
* cell instance $5104 m0 *1 82.08,7
X$5104 23 38 FILLCELL_X1
* cell instance $5105 m0 *1 82.27,7
X$5105 145 130 78 23 38 109 MUX2_X1
* cell instance $5106 m0 *1 83.6,7
X$5106 23 38 FILLCELL_X16
* cell instance $5107 m0 *1 86.64,7
X$5107 23 38 FILLCELL_X2
* cell instance $5108 r0 *1 44.27,7
X$5108 23 38 FILLCELL_X16
* cell instance $5109 r0 *1 47.31,7
X$5109 23 38 FILLCELL_X8
* cell instance $5110 r0 *1 48.83,7
X$5110 23 38 FILLCELL_X4
* cell instance $5111 r0 *1 49.59,7
X$5111 23 38 FILLCELL_X1
* cell instance $5112 r0 *1 49.78,7
X$5112 23 3052 137 164 76 38 DFF_X1
* cell instance $5113 r0 *1 53.01,7
X$5113 23 38 FILLCELL_X8
* cell instance $5114 r0 *1 54.53,7
X$5114 23 38 FILLCELL_X4
* cell instance $5115 r0 *1 55.29,7
X$5115 23 38 FILLCELL_X2
* cell instance $5116 r0 *1 55.67,7
X$5116 23 38 FILLCELL_X1
* cell instance $5117 r0 *1 55.86,7
X$5117 139 23 38 76 CLKBUF_X3
* cell instance $5118 r0 *1 56.81,7
X$5118 23 38 FILLCELL_X16
* cell instance $5119 r0 *1 59.14,7
X$5119 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $5120 r0 *1 59.14,7
X$5120 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $5121 r0 *1 59.14,7
X$5121 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $5122 r0 *1 59.85,7
X$5122 23 38 FILLCELL_X4
* cell instance $5123 r0 *1 60.61,7
X$5123 23 38 FILLCELL_X2
* cell instance $5124 r0 *1 60.99,7
X$5124 23 38 FILLCELL_X1
* cell instance $5125 r0 *1 61.18,7
X$5125 138 38 133 23 BUF_X4
* cell instance $5126 r0 *1 62.51,7
X$5126 23 38 FILLCELL_X8
* cell instance $5127 r0 *1 64.03,7
X$5127 139 23 38 32 CLKBUF_X3
* cell instance $5128 r0 *1 64.98,7
X$5128 23 3015 140 163 32 38 DFF_X1
* cell instance $5129 r0 *1 68.21,7
X$5129 124 88 48 23 38 152 MUX2_X1
* cell instance $5130 r0 *1 69.54,7
X$5130 23 38 FILLCELL_X2
* cell instance $5131 r0 *1 69.92,7
X$5131 23 3044 141 151 153 38 DFF_X1
* cell instance $5132 r0 *1 73.15,7
X$5132 141 126 81 23 38 142 MUX2_X1
* cell instance $5133 r0 *1 74.48,7
X$5133 23 38 FILLCELL_X4
* cell instance $5134 r0 *1 75.24,7
X$5134 23 38 FILLCELL_X1
* cell instance $5135 r0 *1 75.43,7
X$5135 34 23 38 CLKBUF_X1
* cell instance $5136 r0 *1 76,7
X$5136 139 23 38 34 CLKBUF_X3
* cell instance $5137 r0 *1 76.95,7
X$5137 23 38 FILLCELL_X2
* cell instance $5138 r0 *1 77.33,7
X$5138 150 130 52 23 38 143 MUX2_X1
* cell instance $5139 r0 *1 78.66,7
X$5139 23 38 FILLCELL_X4
* cell instance $5140 r0 *1 79.42,7
X$5140 23 38 FILLCELL_X2
* cell instance $5141 r0 *1 79.8,7
X$5141 23 38 FILLCELL_X1
* cell instance $5142 r0 *1 79.99,7
X$5142 82 144 150 23 38 233 MUX2_X1
* cell instance $5143 r0 *1 81.32,7
X$5143 23 38 FILLCELL_X8
* cell instance $5144 r0 *1 82.84,7
X$5144 36 23 38 3145 INV_X1
* cell instance $5145 r0 *1 83.22,7
X$5145 86 144 145 23 38 162 MUX2_X1
* cell instance $5146 r0 *1 84.55,7
X$5146 139 23 38 36 CLKBUF_X3
* cell instance $5147 r0 *1 85.5,7
X$5147 23 38 FILLCELL_X16
* cell instance $5148 m0 *1 87.21,7
X$5148 49 133 54 23 38 108 MUX2_X1
* cell instance $5149 m0 *1 87.02,7
X$5149 23 38 FILLCELL_X1
* cell instance $5150 m0 *1 88.54,7
X$5150 54 126 85 23 38 146 MUX2_X1
* cell instance $5151 m0 *1 89.87,7
X$5151 23 38 FILLCELL_X8
* cell instance $5152 m0 *1 91.39,7
X$5152 53 79 127 23 38 128 MUX2_X1
* cell instance $5153 m0 *1 92.72,7
X$5153 23 2712 127 128 83 38 DFF_X1
* cell instance $5154 m0 *1 95.95,7
X$5154 23 38 FILLCELL_X4
* cell instance $5155 m0 *1 96.71,7
X$5155 23 38 FILLCELL_X2
* cell instance $5156 r0 *1 88.54,7
X$5156 23 38 FILLCELL_X8
* cell instance $5157 r0 *1 90.06,7
X$5157 83 23 38 CLKBUF_X1
* cell instance $5158 r0 *1 90.63,7
X$5158 139 23 38 83 CLKBUF_X3
* cell instance $5159 r0 *1 91.58,7
X$5159 23 3128 159 161 83 38 DFF_X1
* cell instance $5160 r0 *1 94.81,7
X$5160 23 38 FILLCELL_X8
* cell instance $5161 r0 *1 96.33,7
X$5161 23 38 FILLCELL_X4
* cell instance $5162 r180 *1 97.28,7
X$5162 23 38 23 38 TAPCELL_X1
* cell instance $5163 m90 *1 97.28,7
X$5163 23 38 23 38 TAPCELL_X1
* cell instance $5164 m0 *1 1.33,9.8
X$5164 23 38 FILLCELL_X32
* cell instance $5165 m0 *1 1.14,9.8
X$5165 23 38 23 38 TAPCELL_X1
* cell instance $5166 m0 *1 7.41,9.8
X$5166 23 38 FILLCELL_X8
* cell instance $5167 m0 *1 8.93,9.8
X$5167 23 38 FILLCELL_X4
* cell instance $5168 m0 *1 9.69,9.8
X$5168 23 38 FILLCELL_X2
* cell instance $5169 r0 *1 1.14,9.8
X$5169 23 38 23 38 TAPCELL_X1
* cell instance $5170 r0 *1 1.33,9.8
X$5170 23 38 FILLCELL_X32
* cell instance $5171 r0 *1 3.14,9.8
X$5171 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $5172 r0 *1 3.14,9.8
X$5172 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $5173 r0 *1 3.14,9.8
X$5173 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $5174 r0 *1 7.41,9.8
X$5174 23 38 FILLCELL_X4
* cell instance $5175 r0 *1 8.17,9.8
X$5175 23 38 FILLCELL_X2
* cell instance $5176 r0 *1 8.55,9.8
X$5176 23 38 FILLCELL_X1
* cell instance $5177 r0 *1 8.74,9.8
X$5177 154 171 201 23 38 200 MUX2_X1
* cell instance $5178 m0 *1 10.07,9.8
X$5178 23 38 FILLCELL_X1
* cell instance $5179 m0 *1 11.59,9.8
X$5179 23 38 FILLCELL_X1
* cell instance $5180 m0 *1 11.78,9.8
X$5180 106 70 148 23 38 296 MUX2_X1
* cell instance $5181 m0 *1 13.11,9.8
X$5181 23 38 FILLCELL_X4
* cell instance $5182 m0 *1 13.87,9.8
X$5182 23 38 FILLCELL_X1
* cell instance $5183 m0 *1 14.06,9.8
X$5183 27 155 136 23 38 156 MUX2_X1
* cell instance $5184 m0 *1 15.39,9.8
X$5184 23 2755 189 166 28 38 DFF_X1
* cell instance $5185 m0 *1 18.62,9.8
X$5185 23 38 FILLCELL_X16
* cell instance $5186 m0 *1 21.66,9.8
X$5186 23 38 FILLCELL_X2
* cell instance $5187 r0 *1 10.07,9.8
X$5187 23 3036 202 230 28 38 DFF_X1
* cell instance $5188 r0 *1 13.3,9.8
X$5188 154 155 202 23 38 230 MUX2_X1
* cell instance $5189 r0 *1 14.63,9.8
X$5189 23 38 FILLCELL_X4
* cell instance $5190 r0 *1 15.39,9.8
X$5190 27 171 189 23 38 166 MUX2_X1
* cell instance $5191 r0 *1 16.72,9.8
X$5191 189 212 136 23 38 203 MUX2_X1
* cell instance $5192 r0 *1 21.28,9.8
X$5192 24 155 273 23 38 167 MUX2_X1
* cell instance $5193 m0 *1 22.61,9.8
X$5193 26 155 165 23 38 193 MUX2_X1
* cell instance $5194 m0 *1 27.17,9.8
X$5194 23 38 FILLCELL_X8
* cell instance $5195 m0 *1 28.69,9.8
X$5195 23 38 FILLCELL_X1
* cell instance $5196 m0 *1 28.88,9.8
X$5196 23 2762 169 207 73 38 DFF_X1
* cell instance $5197 m0 *1 32.11,9.8
X$5197 23 2748 170 194 74 38 DFF_X1
* cell instance $5198 m0 *1 35.34,9.8
X$5198 25 171 170 23 38 194 MUX2_X1
* cell instance $5199 m0 *1 36.67,9.8
X$5199 23 38 FILLCELL_X1
* cell instance $5200 m0 *1 36.86,9.8
X$5200 23 2751 157 196 74 38 DFF_X1
* cell instance $5201 m0 *1 40.09,9.8
X$5201 98 155 157 23 38 196 MUX2_X1
* cell instance $5202 m0 *1 41.42,9.8
X$5202 23 38 FILLCELL_X1
* cell instance $5203 m0 *1 41.61,9.8
X$5203 23 2704 172 197 30 38 DFF_X1
* cell instance $5204 m0 *1 44.84,9.8
X$5204 23 38 FILLCELL_X8
* cell instance $5205 m0 *1 46.36,9.8
X$5205 149 23 38 30 CLKBUF_X3
* cell instance $5206 m0 *1 47.31,9.8
X$5206 30 23 38 CLKBUF_X1
* cell instance $5207 m0 *1 47.88,9.8
X$5207 23 38 FILLCELL_X8
* cell instance $5208 m0 *1 49.4,9.8
X$5208 66 171 137 23 38 164 MUX2_X1
* cell instance $5209 m0 *1 50.73,9.8
X$5209 23 2617 242 199 158 38 DFF_X1
* cell instance $5210 m0 *1 53.96,9.8
X$5210 23 38 FILLCELL_X8
* cell instance $5211 m0 *1 55.48,9.8
X$5211 23 38 FILLCELL_X1
* cell instance $5212 m0 *1 55.67,9.8
X$5212 23 2624 173 198 76 38 DFF_X1
* cell instance $5213 m0 *1 58.9,9.8
X$5213 23 38 FILLCELL_X8
* cell instance $5214 m0 *1 60.42,9.8
X$5214 23 2844 220 244 32 38 DFF_X1
* cell instance $5215 m0 *1 63.65,9.8
X$5215 23 38 FILLCELL_X8
* cell instance $5216 m0 *1 65.17,9.8
X$5216 23 38 FILLCELL_X4
* cell instance $5217 m0 *1 65.93,9.8
X$5217 23 38 FILLCELL_X1
* cell instance $5218 m0 *1 66.12,9.8
X$5218 140 130 48 23 38 163 MUX2_X1
* cell instance $5219 m0 *1 67.45,9.8
X$5219 23 38 FILLCELL_X2
* cell instance $5220 r0 *1 22.61,9.8
X$5220 23 38 FILLCELL_X8
* cell instance $5221 r0 *1 24.13,9.8
X$5221 23 38 FILLCELL_X1
* cell instance $5222 r0 *1 27.55,9.8
X$5222 23 38 FILLCELL_X2
* cell instance $5223 r0 *1 27.93,9.8
X$5223 23 38 FILLCELL_X1
* cell instance $5224 r0 *1 28.12,9.8
X$5224 29 155 169 23 38 207 MUX2_X1
* cell instance $5225 r0 *1 29.45,9.8
X$5225 23 2934 209 208 73 38 DFF_X1
* cell instance $5226 r0 *1 32.68,9.8
X$5226 23 38 FILLCELL_X4
* cell instance $5227 r0 *1 33.44,9.8
X$5227 23 38 FILLCELL_X2
* cell instance $5228 r0 *1 33.82,9.8
X$5228 23 3028 235 210 74 38 DFF_X1
* cell instance $5229 r0 *1 37.05,9.8
X$5229 23 38 FILLCELL_X8
* cell instance $5230 r0 *1 38.57,9.8
X$5230 23 2909 214 213 74 38 DFF_X1
* cell instance $5231 r0 *1 41.8,9.8
X$5231 23 38 FILLCELL_X4
* cell instance $5232 r0 *1 42.56,9.8
X$5232 75 171 172 23 38 197 MUX2_X1
* cell instance $5233 r0 *1 43.89,9.8
X$5233 23 2907 216 215 30 38 DFF_X1
* cell instance $5234 r0 *1 47.12,9.8
X$5234 23 38 FILLCELL_X16
* cell instance $5235 r0 *1 50.16,9.8
X$5235 23 38 FILLCELL_X4
* cell instance $5236 r0 *1 50.92,9.8
X$5236 23 38 FILLCELL_X1
* cell instance $5237 r0 *1 51.11,9.8
X$5237 66 155 242 23 38 199 MUX2_X1
* cell instance $5238 r0 *1 52.44,9.8
X$5238 23 38 FILLCELL_X2
* cell instance $5239 r0 *1 52.82,9.8
X$5239 23 38 FILLCELL_X1
* cell instance $5240 r0 *1 53.01,9.8
X$5240 137 126 242 23 38 405 MUX2_X1
* cell instance $5241 r0 *1 54.34,9.8
X$5241 243 23 38 155 CLKBUF_X3
* cell instance $5242 r0 *1 55.29,9.8
X$5242 121 243 173 23 38 198 MUX2_X1
* cell instance $5243 r0 *1 56.62,9.8
X$5243 23 38 FILLCELL_X2
* cell instance $5244 r0 *1 57,9.8
X$5244 23 3061 218 217 76 38 DFF_X1
* cell instance $5245 r0 *1 59.14,9.8
X$5245 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $5246 r0 *1 59.14,9.8
X$5246 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $5247 r0 *1 59.14,9.8
X$5247 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $5248 r0 *1 60.23,9.8
X$5248 218 126 173 23 38 473 MUX2_X1
* cell instance $5249 r0 *1 61.56,9.8
X$5249 23 38 FILLCELL_X4
* cell instance $5250 r0 *1 62.32,9.8
X$5250 23 38 FILLCELL_X2
* cell instance $5251 r0 *1 62.7,9.8
X$5251 23 38 FILLCELL_X1
* cell instance $5252 r0 *1 62.89,9.8
X$5252 220 174 48 23 38 244 MUX2_X1
* cell instance $5253 r0 *1 64.22,9.8
X$5253 23 38 FILLCELL_X16
* cell instance $5254 r0 *1 67.26,9.8
X$5254 23 38 FILLCELL_X4
* cell instance $5255 m0 *1 68.02,9.8
X$5255 124 144 140 23 38 195 MUX2_X1
* cell instance $5256 m0 *1 67.83,9.8
X$5256 23 38 FILLCELL_X1
* cell instance $5257 m0 *1 69.35,9.8
X$5257 23 38 FILLCELL_X16
* cell instance $5258 m0 *1 72.39,9.8
X$5258 23 38 FILLCELL_X8
* cell instance $5259 m0 *1 73.91,9.8
X$5259 142 177 23 38 175 NOR2_X1
* cell instance $5260 m0 *1 74.48,9.8
X$5260 23 38 FILLCELL_X16
* cell instance $5261 m0 *1 77.52,9.8
X$5261 23 2637 150 143 34 38 DFF_X1
* cell instance $5262 m0 *1 80.75,9.8
X$5262 23 38 FILLCELL_X2
* cell instance $5263 r0 *1 68.02,9.8
X$5263 77 240 290 23 38 241 MUX2_X1
* cell instance $5264 r0 *1 69.35,9.8
X$5264 23 38 FILLCELL_X4
* cell instance $5265 r0 *1 70.11,9.8
X$5265 23 38 FILLCELL_X2
* cell instance $5266 r0 *1 70.49,9.8
X$5266 195 190 23 38 289 NOR2_X1
* cell instance $5267 r0 *1 71.06,9.8
X$5267 23 38 FILLCELL_X8
* cell instance $5268 r0 *1 72.58,9.8
X$5268 23 38 FILLCELL_X1
* cell instance $5269 r0 *1 72.77,9.8
X$5269 77 191 237 23 38 238 MUX2_X1
* cell instance $5270 r0 *1 74.1,9.8
X$5270 77 187 176 23 38 236 MUX2_X1
* cell instance $5271 r0 *1 75.43,9.8
X$5271 23 3106 176 236 34 38 DFF_X1
* cell instance $5272 r0 *1 78.66,9.8
X$5272 23 38 FILLCELL_X2
* cell instance $5273 r0 *1 79.04,9.8
X$5273 23 3100 284 234 36 38 DFF_X1
* cell instance $5274 m0 *1 84.36,9.8
X$5274 23 2589 180 179 36 38 DFF_X1
* cell instance $5275 m0 *1 81.13,9.8
X$5275 23 2655 178 192 36 38 DFF_X1
* cell instance $5276 m0 *1 87.59,9.8
X$5276 162 190 23 38 181 NOR2_X1
* cell instance $5277 m0 *1 88.16,9.8
X$5277 23 38 FILLCELL_X2
* cell instance $5278 r0 *1 82.27,9.8
X$5278 178 174 78 23 38 192 MUX2_X1
* cell instance $5279 r0 *1 83.6,9.8
X$5279 233 190 23 38 231 NOR2_X1
* cell instance $5280 r0 *1 84.17,9.8
X$5280 180 174 52 23 38 179 MUX2_X1
* cell instance $5281 r0 *1 85.5,9.8
X$5281 23 2901 183 224 36 38 DFF_X1
* cell instance $5282 m0 *1 89.11,9.8
X$5282 23 38 FILLCELL_X8
* cell instance $5283 m0 *1 88.54,9.8
X$5283 146 177 23 38 182 NOR2_X1
* cell instance $5284 m0 *1 90.63,9.8
X$5284 159 126 127 23 38 184 MUX2_X1
* cell instance $5285 m0 *1 91.96,9.8
X$5285 53 133 159 23 38 161 MUX2_X1
* cell instance $5286 m0 *1 93.29,9.8
X$5286 23 38 FILLCELL_X16
* cell instance $5287 m0 *1 96.33,9.8
X$5287 23 38 FILLCELL_X4
* cell instance $5288 r180 *1 97.28,9.8
X$5288 23 38 23 38 TAPCELL_X1
* cell instance $5289 r0 *1 88.73,9.8
X$5289 183 188 180 23 38 226 MUX2_X1
* cell instance $5290 r0 *1 90.06,9.8
X$5290 23 38 FILLCELL_X4
* cell instance $5291 r0 *1 90.82,9.8
X$5291 23 38 FILLCELL_X2
* cell instance $5292 r0 *1 91.2,9.8
X$5292 23 38 FILLCELL_X1
* cell instance $5293 r0 *1 91.39,9.8
X$5293 184 177 23 38 229 NOR2_X1
* cell instance $5294 r0 *1 91.96,9.8
X$5294 23 38 FILLCELL_X1
* cell instance $5295 r0 *1 92.15,9.8
X$5295 53 187 185 23 38 186 MUX2_X1
* cell instance $5296 r0 *1 93.48,9.8
X$5296 23 3103 185 186 83 38 DFF_X1
* cell instance $5297 r0 *1 96.71,9.8
X$5297 23 38 FILLCELL_X2
* cell instance $5298 m90 *1 97.28,9.8
X$5298 23 38 23 38 TAPCELL_X1
* cell instance $5299 m0 *1 1.33,85.4
X$5299 23 38 FILLCELL_X32
* cell instance $5300 m0 *1 1.14,85.4
X$5300 23 38 23 38 TAPCELL_X1
* cell instance $5301 m0 *1 7.41,85.4
X$5301 23 38 FILLCELL_X2
* cell instance $5302 r0 *1 1.14,85.4
X$5302 23 38 23 38 TAPCELL_X1
* cell instance $5303 r0 *1 1.33,85.4
X$5303 23 38 FILLCELL_X16
* cell instance $5304 r0 *1 3.14,85.4
X$5304 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $5305 r0 *1 3.14,85.4
X$5305 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $5306 r0 *1 3.14,85.4
X$5306 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $5307 r0 *1 4.37,85.4
X$5307 23 38 FILLCELL_X2
* cell instance $5308 r0 *1 4.75,85.4
X$5308 23 38 FILLCELL_X1
* cell instance $5309 r0 *1 4.94,85.4
X$5309 2325 1369 1820 23 38 2273 MUX2_X1
* cell instance $5310 r0 *1 6.27,85.4
X$5310 23 38 FILLCELL_X8
* cell instance $5311 m0 *1 7.98,85.4
X$5311 23 2659 2141 2216 2045 38 DFF_X1
* cell instance $5312 m0 *1 7.79,85.4
X$5312 23 38 FILLCELL_X1
* cell instance $5313 m0 *1 11.21,85.4
X$5313 23 38 FILLCELL_X32
* cell instance $5314 m0 *1 17.29,85.4
X$5314 23 38 FILLCELL_X8
* cell instance $5315 m0 *1 18.81,85.4
X$5315 2217 23 38 1822 CLKBUF_X2
* cell instance $5316 m0 *1 19.57,85.4
X$5316 23 38 FILLCELL_X4
* cell instance $5317 m0 *1 20.33,85.4
X$5317 23 38 FILLCELL_X2
* cell instance $5318 r0 *1 7.79,85.4
X$5318 23 38 FILLCELL_X1
* cell instance $5319 r0 *1 7.98,85.4
X$5319 1909 23 38 2045 CLKBUF_X3
* cell instance $5320 r0 *1 8.93,85.4
X$5320 23 2960 2297 2296 2045 38 DFF_X1
* cell instance $5321 r0 *1 12.16,85.4
X$5321 23 38 FILLCELL_X4
* cell instance $5322 r0 *1 12.92,85.4
X$5322 23 38 FILLCELL_X2
* cell instance $5323 r0 *1 13.3,85.4
X$5323 23 38 FILLCELL_X1
* cell instance $5324 r0 *1 13.49,85.4
X$5324 2199 23 38 1820 BUF_X2
* cell instance $5325 r0 *1 14.25,85.4
X$5325 23 38 FILLCELL_X8
* cell instance $5326 r0 *1 15.77,85.4
X$5326 23 2955 2274 2299 2144 38 DFF_X1
* cell instance $5327 r0 *1 19,85.4
X$5327 23 38 FILLCELL_X8
* cell instance $5328 r0 *1 20.52,85.4
X$5328 23 38 FILLCELL_X4
* cell instance $5329 m0 *1 22.04,85.4
X$5329 23 38 FILLCELL_X1
* cell instance $5330 m0 *1 20.71,85.4
X$5330 2217 1482 2177 23 38 2229 MUX2_X1
* cell instance $5331 m0 *1 22.23,85.4
X$5331 2217 1530 2178 23 38 2231 MUX2_X1
* cell instance $5332 m0 *1 23.56,85.4
X$5332 23 38 FILLCELL_X16
* cell instance $5333 m0 *1 26.6,85.4
X$5333 23 38 FILLCELL_X4
* cell instance $5334 m0 *1 27.36,85.4
X$5334 23 38 FILLCELL_X2
* cell instance $5335 r0 *1 21.28,85.4
X$5335 23 3018 2275 2239 2144 38 DFF_X1
* cell instance $5336 r0 *1 24.51,85.4
X$5336 23 38 FILLCELL_X8
* cell instance $5337 r0 *1 26.03,85.4
X$5337 2276 1383 1725 23 38 2302 MUX2_X1
* cell instance $5338 r0 *1 27.36,85.4
X$5338 23 38 FILLCELL_X8
* cell instance $5339 m0 *1 27.93,85.4
X$5339 23 2648 2206 2179 2145 38 DFF_X1
* cell instance $5340 m0 *1 27.74,85.4
X$5340 23 38 FILLCELL_X1
* cell instance $5341 m0 *1 31.16,85.4
X$5341 2218 23 38 1725 BUF_X2
* cell instance $5342 m0 *1 31.92,85.4
X$5342 23 38 FILLCELL_X4
* cell instance $5343 m0 *1 32.68,85.4
X$5343 23 38 FILLCELL_X1
* cell instance $5344 m0 *1 32.87,85.4
X$5344 23 2621 2107 2233 2145 38 DFF_X1
* cell instance $5345 m0 *1 36.1,85.4
X$5345 23 38 FILLCELL_X4
* cell instance $5346 m0 *1 36.86,85.4
X$5346 23 38 FILLCELL_X2
* cell instance $5347 r0 *1 28.88,85.4
X$5347 23 38 FILLCELL_X2
* cell instance $5348 r0 *1 29.26,85.4
X$5348 23 38 FILLCELL_X1
* cell instance $5349 r0 *1 29.45,85.4
X$5349 2240 1403 1725 23 38 2303 MUX2_X1
* cell instance $5350 r0 *1 30.78,85.4
X$5350 23 38 FILLCELL_X32
* cell instance $5351 r0 *1 36.86,85.4
X$5351 23 38 FILLCELL_X4
* cell instance $5352 m0 *1 37.43,85.4
X$5352 2220 1530 2219 23 38 2234 MUX2_X1
* cell instance $5353 m0 *1 37.24,85.4
X$5353 23 38 FILLCELL_X1
* cell instance $5354 m0 *1 38.76,85.4
X$5354 23 38 FILLCELL_X8
* cell instance $5355 m0 *1 40.28,85.4
X$5355 23 38 FILLCELL_X4
* cell instance $5356 m0 *1 41.04,85.4
X$5356 2220 1482 2221 23 38 2235 MUX2_X1
* cell instance $5357 m0 *1 42.37,85.4
X$5357 23 38 FILLCELL_X4
* cell instance $5358 m0 *1 43.13,85.4
X$5358 23 38 FILLCELL_X1
* cell instance $5359 m0 *1 43.32,85.4
X$5359 1909 23 38 2149 CLKBUF_X3
* cell instance $5360 m0 *1 44.27,85.4
X$5360 23 2658 2241 2263 2149 38 DFF_X1
* cell instance $5361 m0 *1 47.5,85.4
X$5361 2241 1403 1767 23 38 2263 MUX2_X1
* cell instance $5362 m0 *1 48.83,85.4
X$5362 23 38 FILLCELL_X4
* cell instance $5363 m0 *1 49.59,85.4
X$5363 23 38 FILLCELL_X2
* cell instance $5364 r0 *1 37.62,85.4
X$5364 23 38 FILLCELL_X2
* cell instance $5365 r0 *1 38,85.4
X$5365 23 38 FILLCELL_X1
* cell instance $5366 r0 *1 38.19,85.4
X$5366 2220 23 38 1730 BUF_X2
* cell instance $5367 r0 *1 38.95,85.4
X$5367 23 3066 2308 2307 2149 38 DFF_X1
* cell instance $5368 r0 *1 42.18,85.4
X$5368 23 38 FILLCELL_X16
* cell instance $5369 r0 *1 45.22,85.4
X$5369 23 38 FILLCELL_X1
* cell instance $5370 r0 *1 45.41,85.4
X$5370 23 3019 2279 2309 2149 38 DFF_X1
* cell instance $5371 r0 *1 48.64,85.4
X$5371 2279 1289 1767 23 38 2309 MUX2_X1
* cell instance $5372 m0 *1 51.3,85.4
X$5372 23 2593 2238 2184 1960 38 DFF_X1
* cell instance $5373 m0 *1 49.97,85.4
X$5373 2242 1383 1767 23 38 2311 MUX2_X1
* cell instance $5374 m0 *1 54.53,85.4
X$5374 23 38 FILLCELL_X2
* cell instance $5375 r0 *1 49.97,85.4
X$5375 23 38 FILLCELL_X2
* cell instance $5376 r0 *1 50.35,85.4
X$5376 23 3087 2242 2311 1960 38 DFF_X1
* cell instance $5377 r0 *1 53.58,85.4
X$5377 2242 724 2238 23 38 2243 MUX2_X1
* cell instance $5378 m0 *1 55.1,85.4
X$5378 2243 1650 23 38 2312 NOR2_X1
* cell instance $5379 m0 *1 54.91,85.4
X$5379 23 38 FILLCELL_X1
* cell instance $5380 m0 *1 55.67,85.4
X$5380 23 38 FILLCELL_X2
* cell instance $5381 r0 *1 54.91,85.4
X$5381 1425 2310 2312 548 2269 2244 23 38 2019 OAI33_X1
* cell instance $5382 m0 *1 56.81,85.4
X$5382 2245 1535 23 38 2269 NOR2_X1
* cell instance $5383 m0 *1 56.05,85.4
X$5383 2151 23 38 1767 BUF_X2
* cell instance $5384 m0 *1 57.38,85.4
X$5384 2151 1346 2270 23 38 2313 MUX2_X1
* cell instance $5385 m0 *1 58.71,85.4
X$5385 23 38 FILLCELL_X8
* cell instance $5386 m0 *1 60.23,85.4
X$5386 23 38 FILLCELL_X4
* cell instance $5387 m0 *1 60.99,85.4
X$5387 23 38 FILLCELL_X2
* cell instance $5388 r0 *1 56.24,85.4
X$5388 23 38 FILLCELL_X1
* cell instance $5389 r0 *1 56.43,85.4
X$5389 2280 1358 2270 23 38 2245 MUX2_X1
* cell instance $5390 r0 *1 57.76,85.4
X$5390 23 3085 2270 2313 2246 38 DFF_X1
* cell instance $5391 r0 *1 59.14,85.4
X$5391 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $5392 r0 *1 59.14,85.4
X$5392 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $5393 r0 *1 59.14,85.4
X$5393 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $5394 r0 *1 60.99,85.4
X$5394 23 38 FILLCELL_X4
* cell instance $5395 m0 *1 62.32,85.4
X$5395 2222 23 38 1458 CLKBUF_X3
* cell instance $5396 m0 *1 61.37,85.4
X$5396 2236 2185 2213 38 23 2237 AND3_X1
* cell instance $5397 m0 *1 63.27,85.4
X$5397 2102 2154 3135 38 23 2268 HA_X1
* cell instance $5398 m0 *1 65.17,85.4
X$5398 2102 2154 2223 2236 23 38 2317 NAND4_X1
* cell instance $5399 m0 *1 66.12,85.4
X$5399 23 38 FILLCELL_X1
* cell instance $5400 m0 *1 66.31,85.4
X$5400 2185 2113 38 23 2247 AND2_X1
* cell instance $5401 m0 *1 67.07,85.4
X$5401 2116 2185 23 38 2318 NOR2_X1
* cell instance $5402 m0 *1 67.64,85.4
X$5402 23 38 FILLCELL_X16
* cell instance $5403 m0 *1 70.68,85.4
X$5403 23 38 FILLCELL_X8
* cell instance $5404 m0 *1 72.2,85.4
X$5404 23 38 FILLCELL_X2
* cell instance $5405 r0 *1 61.75,85.4
X$5405 23 38 FILLCELL_X2
* cell instance $5406 r0 *1 62.13,85.4
X$5406 23 38 FILLCELL_X1
* cell instance $5407 r0 *1 62.32,85.4
X$5407 2236 2185 2223 38 23 2222 AND3_X1
* cell instance $5408 r0 *1 63.27,85.4
X$5408 23 38 FILLCELL_X4
* cell instance $5409 r0 *1 64.03,85.4
X$5409 23 38 FILLCELL_X2
* cell instance $5410 r0 *1 64.41,85.4
X$5410 23 38 FILLCELL_X1
* cell instance $5411 r0 *1 64.6,85.4
X$5411 2268 23 38 1496 BUF_X2
* cell instance $5412 r0 *1 65.36,85.4
X$5412 2317 1951 2232 23 2267 38 AOI21_X1
* cell instance $5413 r0 *1 66.12,85.4
X$5413 23 38 FILLCELL_X2
* cell instance $5414 r0 *1 66.5,85.4
X$5414 2247 2267 2318 23 38 2319 MUX2_X1
* cell instance $5415 r0 *1 67.83,85.4
X$5415 2320 23 38 2185 BUF_X2
* cell instance $5416 r0 *1 68.59,85.4
X$5416 23 38 FILLCELL_X8
* cell instance $5417 r0 *1 70.11,85.4
X$5417 2282 1984 2321 23 38 1980 MUX2_X1
* cell instance $5418 r0 *1 71.44,85.4
X$5418 23 2248 2224 2101 1981 38 DFF_X1
* cell instance $5419 m0 *1 73.91,85.4
X$5419 1319 2224 23 38 2266 NOR2_X1
* cell instance $5420 m0 *1 72.58,85.4
X$5420 2265 2323 2266 23 38 2101 MUX2_X1
* cell instance $5421 m0 *1 74.48,85.4
X$5421 2224 2057 38 23 2265 AND2_X1
* cell instance $5422 m0 *1 75.24,85.4
X$5422 23 2647 2188 2261 1981 38 DFF_X1
* cell instance $5423 m0 *1 78.47,85.4
X$5423 2230 2264 2262 23 38 2261 MUX2_X1
* cell instance $5424 m0 *1 79.8,85.4
X$5424 23 38 FILLCELL_X8
* cell instance $5425 m0 *1 81.32,85.4
X$5425 23 38 FILLCELL_X4
* cell instance $5426 m0 *1 82.08,85.4
X$5426 2259 2250 2260 23 38 2191 MUX2_X1
* cell instance $5427 m0 *1 83.41,85.4
X$5427 23 38 FILLCELL_X2
* cell instance $5428 r0 *1 74.67,85.4
X$5428 2224 2284 2285 2160 23 38 2315 NAND4_X1
* cell instance $5429 r0 *1 75.62,85.4
X$5429 2315 2190 2232 23 2264 38 AOI21_X1
* cell instance $5430 r0 *1 76.38,85.4
X$5430 2287 2249 1953 23 38 NOR2_X4
* cell instance $5431 r0 *1 78.09,85.4
X$5431 2249 38 1951 23 BUF_X4
* cell instance $5432 r0 *1 79.42,85.4
X$5432 2160 2287 1951 38 23 1984 OAI21_X2
* cell instance $5433 r0 *1 80.75,85.4
X$5433 23 38 FILLCELL_X8
* cell instance $5434 r0 *1 82.27,85.4
X$5434 2288 2289 1686 1951 23 38 2250 NOR4_X1
* cell instance $5435 r0 *1 83.22,85.4
X$5435 23 38 FILLCELL_X8
* cell instance $5436 m0 *1 84.36,85.4
X$5436 1949 2290 23 38 2259 NOR2_X1
* cell instance $5437 m0 *1 83.79,85.4
X$5437 2116 2192 23 38 2260 NOR2_X1
* cell instance $5438 m0 *1 84.93,85.4
X$5438 23 38 FILLCELL_X8
* cell instance $5439 m0 *1 86.45,85.4
X$5439 23 38 FILLCELL_X1
* cell instance $5440 m0 *1 86.64,85.4
X$5440 2193 2257 2232 2190 23 38 2228 NAND4_X1
* cell instance $5441 m0 *1 87.59,85.4
X$5441 23 38 FILLCELL_X2
* cell instance $5442 r0 *1 84.74,85.4
X$5442 23 38 FILLCELL_X4
* cell instance $5443 r0 *1 85.5,85.4
X$5443 2192 23 38 2290 INV_X1
* cell instance $5444 r0 *1 85.88,85.4
X$5444 23 38 FILLCELL_X4
* cell instance $5445 r0 *1 86.64,85.4
X$5445 2161 2063 23 38 2288 NAND2_X1
* cell instance $5446 r0 *1 87.21,85.4
X$5446 23 38 FILLCELL_X4
* cell instance $5447 r0 *1 87.97,85.4
X$5447 1949 2251 23 38 2258 NOR2_X1
* cell instance $5448 m0 *1 89.3,85.4
X$5448 2225 2226 2252 38 23 2257 AND3_X1
* cell instance $5449 m0 *1 87.97,85.4
X$5449 2258 2228 2194 23 38 2306 MUX2_X1
* cell instance $5450 m0 *1 90.25,85.4
X$5450 2161 2063 2226 2225 23 38 2301 NAND4_X1
* cell instance $5451 m0 *1 91.2,85.4
X$5451 2226 2113 38 23 2227 AND2_X1
* cell instance $5452 m0 *1 91.96,85.4
X$5452 2116 2252 23 38 2254 NOR2_X1
* cell instance $5453 m0 *1 92.53,85.4
X$5453 23 2255 2026 3131 2252 38 DFF_X2
* cell instance $5454 m0 *1 96.14,85.4
X$5454 23 38 FILLCELL_X2
* cell instance $5455 r0 *1 88.54,85.4
X$5455 2252 2226 2225 2251 23 2289 38 NAND4_X2
* cell instance $5456 r0 *1 90.25,85.4
X$5456 2252 2113 38 23 2298 AND2_X1
* cell instance $5457 r0 *1 91.01,85.4
X$5457 2301 1686 2065 23 38 2253 NOR3_X1
* cell instance $5458 r0 *1 91.77,85.4
X$5458 2298 2253 2254 23 38 2255 MUX2_X1
* cell instance $5459 r0 *1 93.1,85.4
X$5459 2116 2225 23 38 2292 NOR2_X1
* cell instance $5460 r0 *1 93.67,85.4
X$5460 23 38 FILLCELL_X4
* cell instance $5461 r0 *1 94.43,85.4
X$5461 23 38 FILLCELL_X2
* cell instance $5462 r0 *1 94.81,85.4
X$5462 2251 23 38 2294 BUF_X1
* cell instance $5463 r0 *1 95.38,85.4
X$5463 23 38 FILLCELL_X2
* cell instance $5464 r0 *1 95.76,85.4
X$5464 23 38 FILLCELL_X1
* cell instance $5465 r0 *1 95.95,85.4
X$5465 2252 23 38 2295 BUF_X1
* cell instance $5466 r0 *1 96.52,85.4
X$5466 2196 23 38 2256 BUF_X1
* cell instance $5467 r180 *1 97.28,85.4
X$5467 23 38 23 38 TAPCELL_X1
* cell instance $5468 m0 *1 96.52,85.4
X$5468 2196 23 38 2226 BUF_X1
* cell instance $5469 m90 *1 97.28,85.4
X$5469 23 38 23 38 TAPCELL_X1
* cell instance $5470 m0 *1 1.33,32.2
X$5470 23 38 FILLCELL_X32
* cell instance $5471 m0 *1 1.14,32.2
X$5471 23 38 23 38 TAPCELL_X1
* cell instance $5472 m0 *1 7.41,32.2
X$5472 23 38 FILLCELL_X32
* cell instance $5473 m0 *1 13.49,32.2
X$5473 23 38 FILLCELL_X8
* cell instance $5474 m0 *1 15.01,32.2
X$5474 23 38 FILLCELL_X2
* cell instance $5475 r0 *1 1.14,32.2
X$5475 23 38 23 38 TAPCELL_X1
* cell instance $5476 r0 *1 1.33,32.2
X$5476 23 38 FILLCELL_X8
* cell instance $5477 r0 *1 2.85,32.2
X$5477 23 38 FILLCELL_X4
* cell instance $5478 r0 *1 3.14,32.2
X$5478 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $5479 r0 *1 3.14,32.2
X$5479 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $5480 r0 *1 3.14,32.2
X$5480 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $5481 r0 *1 3.61,32.2
X$5481 502 762 790 23 38 807 MUX2_X1
* cell instance $5482 r0 *1 4.94,32.2
X$5482 23 38 FILLCELL_X4
* cell instance $5483 r0 *1 5.7,32.2
X$5483 23 38 FILLCELL_X1
* cell instance $5484 r0 *1 5.89,32.2
X$5484 295 762 825 23 38 808 MUX2_X1
* cell instance $5485 r0 *1 7.22,32.2
X$5485 23 38 FILLCELL_X8
* cell instance $5486 r0 *1 8.74,32.2
X$5486 453 762 810 23 38 809 MUX2_X1
* cell instance $5487 r0 *1 10.07,32.2
X$5487 23 38 FILLCELL_X4
* cell instance $5488 r0 *1 10.83,32.2
X$5488 23 38 FILLCELL_X2
* cell instance $5489 r0 *1 11.21,32.2
X$5489 23 38 FILLCELL_X1
* cell instance $5490 r0 *1 11.4,32.2
X$5490 23 3076 812 847 660 38 DFF_X1
* cell instance $5491 r0 *1 14.63,32.2
X$5491 23 3011 791 781 653 38 DFF_X1
* cell instance $5492 m0 *1 15.58,32.2
X$5492 23 2772 733 749 653 38 DFF_X1
* cell instance $5493 m0 *1 15.39,32.2
X$5493 23 38 FILLCELL_X1
* cell instance $5494 m0 *1 18.81,32.2
X$5494 23 38 FILLCELL_X16
* cell instance $5495 m0 *1 21.85,32.2
X$5495 23 2803 697 734 763 38 DFF_X1
* cell instance $5496 m0 *1 25.08,32.2
X$5496 23 38 FILLCELL_X8
* cell instance $5497 m0 *1 26.6,32.2
X$5497 23 38 FILLCELL_X4
* cell instance $5498 m0 *1 27.36,32.2
X$5498 23 38 FILLCELL_X2
* cell instance $5499 r0 *1 17.86,32.2
X$5499 23 38 FILLCELL_X16
* cell instance $5500 r0 *1 20.9,32.2
X$5500 23 38 FILLCELL_X2
* cell instance $5501 r0 *1 21.28,32.2
X$5501 23 38 FILLCELL_X1
* cell instance $5502 r0 *1 21.47,32.2
X$5502 23 2997 764 782 763 38 DFF_X1
* cell instance $5503 r0 *1 24.7,32.2
X$5503 23 38 FILLCELL_X1
* cell instance $5504 r0 *1 24.89,32.2
X$5504 434 23 38 693 CLKBUF_X3
* cell instance $5505 r0 *1 25.84,32.2
X$5505 693 23 38 3155 CLKBUF_X3
* cell instance $5506 r0 *1 26.79,32.2
X$5506 23 3064 750 765 763 38 DFF_X1
* cell instance $5507 m0 *1 29.07,32.2
X$5507 23 38 FILLCELL_X1
* cell instance $5508 m0 *1 27.74,32.2
X$5508 421 628 750 23 38 765 MUX2_X1
* cell instance $5509 m0 *1 29.26,32.2
X$5509 750 602 686 23 38 828 MUX2_X1
* cell instance $5510 m0 *1 30.59,32.2
X$5510 23 38 FILLCELL_X8
* cell instance $5511 m0 *1 32.11,32.2
X$5511 23 38 FILLCELL_X4
* cell instance $5512 m0 *1 32.87,32.2
X$5512 23 2733 699 752 655 38 DFF_X1
* cell instance $5513 m0 *1 36.1,32.2
X$5513 693 23 38 655 CLKBUF_X3
* cell instance $5514 m0 *1 37.05,32.2
X$5514 655 23 38 CLKBUF_X1
* cell instance $5515 m0 *1 37.62,32.2
X$5515 690 602 736 23 38 794 MUX2_X1
* cell instance $5516 m0 *1 38.95,32.2
X$5516 98 659 768 23 38 785 MUX2_X1
* cell instance $5517 m0 *1 40.28,32.2
X$5517 23 38 FILLCELL_X16
* cell instance $5518 m0 *1 43.32,32.2
X$5518 23 38 FILLCELL_X2
* cell instance $5519 r0 *1 30.02,32.2
X$5519 23 38 FILLCELL_X1
* cell instance $5520 r0 *1 30.21,32.2
X$5520 23 3057 767 766 763 38 DFF_X1
* cell instance $5521 r0 *1 33.44,32.2
X$5521 23 38 FILLCELL_X16
* cell instance $5522 r0 *1 36.48,32.2
X$5522 23 38 FILLCELL_X8
* cell instance $5523 r0 *1 38,32.2
X$5523 23 38 FILLCELL_X2
* cell instance $5524 r0 *1 38.38,32.2
X$5524 23 3048 768 785 655 38 DFF_X1
* cell instance $5525 r0 *1 41.61,32.2
X$5525 23 38 FILLCELL_X2
* cell instance $5526 r0 *1 41.99,32.2
X$5526 636 23 38 3147 INV_X1
* cell instance $5527 r0 *1 42.37,32.2
X$5527 398 762 769 23 38 786 MUX2_X1
* cell instance $5528 m0 *1 43.89,32.2
X$5528 23 2689 737 756 636 38 DFF_X1
* cell instance $5529 m0 *1 43.7,32.2
X$5529 23 38 FILLCELL_X1
* cell instance $5530 m0 *1 47.12,32.2
X$5530 23 38 FILLCELL_X8
* cell instance $5531 m0 *1 48.64,32.2
X$5531 23 38 FILLCELL_X2
* cell instance $5532 r0 *1 43.7,32.2
X$5532 23 3050 769 786 636 38 DFF_X1
* cell instance $5533 r0 *1 46.93,32.2
X$5533 769 144 737 23 38 770 MUX2_X1
* cell instance $5534 r0 *1 48.26,32.2
X$5534 23 38 FILLCELL_X8
* cell instance $5535 m0 *1 49.21,32.2
X$5535 23 2777 738 757 666 38 DFF_X1
* cell instance $5536 m0 *1 49.02,32.2
X$5536 23 38 FILLCELL_X1
* cell instance $5537 m0 *1 52.44,32.2
X$5537 771 23 38 632 CLKBUF_X3
* cell instance $5538 m0 *1 53.39,32.2
X$5538 23 38 FILLCELL_X4
* cell instance $5539 m0 *1 54.15,32.2
X$5539 23 38 FILLCELL_X1
* cell instance $5540 m0 *1 54.34,32.2
X$5540 23 2761 772 759 666 38 DFF_X1
* cell instance $5541 m0 *1 57.57,32.2
X$5541 23 38 FILLCELL_X4
* cell instance $5542 m0 *1 58.33,32.2
X$5542 23 38 FILLCELL_X1
* cell instance $5543 m0 *1 58.52,32.2
X$5543 121 23 38 640 BUF_X2
* cell instance $5544 m0 *1 59.28,32.2
X$5544 23 38 FILLCELL_X1
* cell instance $5545 m0 *1 59.47,32.2
X$5545 23 2822 774 761 666 38 DFF_X1
* cell instance $5546 m0 *1 62.7,32.2
X$5546 23 38 FILLCELL_X16
* cell instance $5547 m0 *1 65.74,32.2
X$5547 23 38 FILLCELL_X4
* cell instance $5548 m0 *1 66.5,32.2
X$5548 23 38 FILLCELL_X1
* cell instance $5549 m0 *1 66.69,32.2
X$5549 739 724 740 23 38 760 MUX2_X1
* cell instance $5550 m0 *1 68.02,32.2
X$5550 23 38 FILLCELL_X4
* cell instance $5551 m0 *1 68.78,32.2
X$5551 23 38 FILLCELL_X2
* cell instance $5552 r0 *1 49.78,32.2
X$5552 23 38 FILLCELL_X4
* cell instance $5553 r0 *1 50.54,32.2
X$5553 23 38 FILLCELL_X2
* cell instance $5554 r0 *1 50.92,32.2
X$5554 821 23 38 659 CLKBUF_X3
* cell instance $5555 r0 *1 51.87,32.2
X$5555 23 38 FILLCELL_X8
* cell instance $5556 r0 *1 53.39,32.2
X$5556 23 3034 797 822 839 38 DFF_X1
* cell instance $5557 r0 *1 56.62,32.2
X$5557 112 771 772 23 38 759 MUX2_X1
* cell instance $5558 r0 *1 57.95,32.2
X$5558 23 38 FILLCELL_X4
* cell instance $5559 r0 *1 58.71,32.2
X$5559 121 771 773 23 38 824 MUX2_X1
* cell instance $5560 r0 *1 59.14,32.2
X$5560 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $5561 r0 *1 59.14,32.2
X$5561 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $5562 r0 *1 59.14,32.2
X$5562 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $5563 r0 *1 60.04,32.2
X$5563 23 38 FILLCELL_X4
* cell instance $5564 r0 *1 60.8,32.2
X$5564 23 38 FILLCELL_X2
* cell instance $5565 r0 *1 61.18,32.2
X$5565 640 796 774 23 38 761 MUX2_X1
* cell instance $5566 r0 *1 62.51,32.2
X$5566 23 38 FILLCELL_X4
* cell instance $5567 r0 *1 63.27,32.2
X$5567 23 38 FILLCELL_X2
* cell instance $5568 r0 *1 63.65,32.2
X$5568 23 38 FILLCELL_X1
* cell instance $5569 r0 *1 63.84,32.2
X$5569 23 3054 740 788 705 38 DFF_X1
* cell instance $5570 r0 *1 67.07,32.2
X$5570 23 38 FILLCELL_X2
* cell instance $5571 r0 *1 67.45,32.2
X$5571 740 130 799 23 38 788 MUX2_X1
* cell instance $5572 r0 *1 68.78,32.2
X$5572 23 38 FILLCELL_X1
* cell instance $5573 r0 *1 68.97,32.2
X$5573 705 23 38 CLKBUF_X1
* cell instance $5574 m0 *1 69.35,32.2
X$5574 760 190 23 38 747 NOR2_X1
* cell instance $5575 m0 *1 69.16,32.2
X$5575 23 38 FILLCELL_X1
* cell instance $5576 m0 *1 69.92,32.2
X$5576 744 23 38 705 CLKBUF_X3
* cell instance $5577 m0 *1 70.87,32.2
X$5577 742 559 672 23 38 758 MUX2_X1
* cell instance $5578 m0 *1 72.2,32.2
X$5578 742 263 743 23 38 787 MUX2_X1
* cell instance $5579 m0 *1 73.53,32.2
X$5579 23 38 FILLCELL_X2
* cell instance $5580 r0 *1 69.54,32.2
X$5580 23 3069 742 758 705 38 DFF_X1
* cell instance $5581 r0 *1 72.77,32.2
X$5581 741 177 23 38 818 NOR2_X1
* cell instance $5582 r0 *1 73.34,32.2
X$5582 787 274 23 38 853 NOR2_X1
* cell instance $5583 r0 *1 73.91,32.2
X$5583 744 23 38 3154 CLKBUF_X3
* cell instance $5584 m0 *1 74.86,32.2
X$5584 23 38 FILLCELL_X2
* cell instance $5585 m0 *1 73.91,32.2
X$5585 434 23 38 744 CLKBUF_X3
* cell instance $5586 r0 *1 74.86,32.2
X$5586 23 38 FILLCELL_X1
* cell instance $5587 r0 *1 75.05,32.2
X$5587 784 130 672 23 38 816 MUX2_X1
* cell instance $5588 m0 *1 78.47,32.2
X$5588 23 38 FILLCELL_X8
* cell instance $5589 m0 *1 75.24,32.2
X$5589 23 2794 754 755 801 38 DFF_X1
* cell instance $5590 m0 *1 79.99,32.2
X$5590 23 38 FILLCELL_X2
* cell instance $5591 r0 *1 76.38,32.2
X$5591 23 38 FILLCELL_X2
* cell instance $5592 r0 *1 76.76,32.2
X$5592 23 38 FILLCELL_X1
* cell instance $5593 r0 *1 76.95,32.2
X$5593 754 263 784 23 38 802 MUX2_X1
* cell instance $5594 r0 *1 78.28,32.2
X$5594 23 38 FILLCELL_X2
* cell instance $5595 r0 *1 78.66,32.2
X$5595 23 38 FILLCELL_X1
* cell instance $5596 r0 *1 78.85,32.2
X$5596 710 23 38 672 BUF_X2
* cell instance $5597 r0 *1 79.61,32.2
X$5597 783 374 23 38 803 NOR2_X1
* cell instance $5598 r0 *1 80.18,32.2
X$5598 23 2921 753 775 673 38 DFF_X1
* cell instance $5599 m0 *1 81.7,32.2
X$5599 23 38 FILLCELL_X2
* cell instance $5600 m0 *1 80.37,32.2
X$5600 672 260 753 23 38 775 MUX2_X1
* cell instance $5601 m0 *1 83.41,32.2
X$5601 23 38 FILLCELL_X1
* cell instance $5602 m0 *1 82.08,32.2
X$5602 753 438 745 23 38 707 MUX2_X1
* cell instance $5603 m0 *1 83.6,32.2
X$5603 23 2713 745 746 673 38 DFF_X1
* cell instance $5604 m0 *1 86.83,32.2
X$5604 23 38 FILLCELL_X16
* cell instance $5605 m0 *1 89.87,32.2
X$5605 23 38 FILLCELL_X2
* cell instance $5606 r0 *1 83.41,32.2
X$5606 710 240 745 23 38 746 MUX2_X1
* cell instance $5607 r0 *1 84.74,32.2
X$5607 23 38 FILLCELL_X4
* cell instance $5608 r0 *1 85.5,32.2
X$5608 776 174 799 23 38 780 MUX2_X1
* cell instance $5609 r0 *1 86.83,32.2
X$5609 23 2862 776 780 647 38 DFF_X1
* cell instance $5610 r0 *1 90.06,32.2
X$5610 23 38 FILLCELL_X2
* cell instance $5611 m0 *1 90.44,32.2
X$5611 227 777 747 225 674 779 23 38 748 OAI33_X1
* cell instance $5612 m0 *1 90.25,32.2
X$5612 23 38 FILLCELL_X1
* cell instance $5613 m0 *1 91.77,32.2
X$5613 23 38 FILLCELL_X2
* cell instance $5614 r0 *1 90.44,32.2
X$5614 23 38 FILLCELL_X1
* cell instance $5615 r0 *1 90.63,32.2
X$5615 805 261 23 38 777 NOR2_X1
* cell instance $5616 r0 *1 91.2,32.2
X$5616 23 38 FILLCELL_X4
* cell instance $5617 r0 *1 91.96,32.2
X$5617 23 38 FILLCELL_X2
* cell instance $5618 m0 *1 93.1,32.2
X$5618 23 38 FILLCELL_X2
* cell instance $5619 m0 *1 92.15,32.2
X$5619 744 23 38 647 CLKBUF_X3
* cell instance $5620 r0 *1 92.34,32.2
X$5620 778 177 23 38 779 NOR2_X1
* cell instance $5621 r0 *1 92.91,32.2
X$5621 23 38 FILLCELL_X16
* cell instance $5622 m0 *1 94.81,32.2
X$5622 23 38 FILLCELL_X8
* cell instance $5623 m0 *1 93.48,32.2
X$5623 713 126 714 23 38 778 MUX2_X1
* cell instance $5624 m0 *1 96.33,32.2
X$5624 23 38 FILLCELL_X4
* cell instance $5625 r180 *1 97.28,32.2
X$5625 23 38 23 38 TAPCELL_X1
* cell instance $5626 r0 *1 95.95,32.2
X$5626 23 38 FILLCELL_X4
* cell instance $5627 r0 *1 96.71,32.2
X$5627 23 38 FILLCELL_X2
* cell instance $5628 m90 *1 97.28,32.2
X$5628 23 38 23 38 TAPCELL_X1
* cell instance $5629 m0 *1 1.33,74.2
X$5629 23 38 FILLCELL_X32
* cell instance $5630 m0 *1 1.14,74.2
X$5630 23 38 23 38 TAPCELL_X1
* cell instance $5631 m0 *1 7.41,74.2
X$5631 23 38 FILLCELL_X4
* cell instance $5632 m0 *1 8.17,74.2
X$5632 23 38 FILLCELL_X1
* cell instance $5633 m0 *1 8.36,74.2
X$5633 23 2619 1903 1952 1902 38 DFF_X1
* cell instance $5634 m0 *1 11.59,74.2
X$5634 1903 627 1868 23 38 1924 MUX2_X1
* cell instance $5635 m0 *1 12.92,74.2
X$5635 1924 381 23 38 1922 NOR2_X1
* cell instance $5636 m0 *1 13.49,74.2
X$5636 23 38 FILLCELL_X8
* cell instance $5637 m0 *1 15.01,74.2
X$5637 23 38 FILLCELL_X4
* cell instance $5638 m0 *1 15.77,74.2
X$5638 23 38 FILLCELL_X1
* cell instance $5639 m0 *1 15.96,74.2
X$5639 1870 1446 1791 23 38 1923 MUX2_X1
* cell instance $5640 m0 *1 17.29,74.2
X$5640 23 38 FILLCELL_X8
* cell instance $5641 m0 *1 18.81,74.2
X$5641 23 38 FILLCELL_X4
* cell instance $5642 m0 *1 19.57,74.2
X$5642 23 38 FILLCELL_X1
* cell instance $5643 m0 *1 19.76,74.2
X$5643 1485 1793 1904 1142 1970 1925 23 38 1905 OAI33_X1
* cell instance $5644 m0 *1 21.09,74.2
X$5644 23 38 FILLCELL_X2
* cell instance $5645 r0 *1 1.14,74.2
X$5645 23 38 23 38 TAPCELL_X1
* cell instance $5646 r0 *1 1.33,74.2
X$5646 23 38 FILLCELL_X8
* cell instance $5647 r0 *1 2.85,74.2
X$5647 1935 1493 1950 23 38 1967 MUX2_X1
* cell instance $5648 r0 *1 3.14,74.2
X$5648 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $5649 r0 *1 3.14,74.2
X$5649 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $5650 r0 *1 3.14,74.2
X$5650 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $5651 r0 *1 4.18,74.2
X$5651 23 38 FILLCELL_X4
* cell instance $5652 r0 *1 4.94,74.2
X$5652 23 38 FILLCELL_X1
* cell instance $5653 r0 *1 5.13,74.2
X$5653 1950 70 1968 23 38 1954 MUX2_X1
* cell instance $5654 r0 *1 6.46,74.2
X$5654 23 38 FILLCELL_X16
* cell instance $5655 r0 *1 9.5,74.2
X$5655 23 38 FILLCELL_X2
* cell instance $5656 r0 *1 9.88,74.2
X$5656 1903 1403 1791 23 38 1952 MUX2_X1
* cell instance $5657 r0 *1 11.21,74.2
X$5657 1954 1483 23 38 1955 NOR2_X1
* cell instance $5658 r0 *1 11.78,74.2
X$5658 1425 1922 1869 548 2166 1955 23 38 1927 OAI33_X1
* cell instance $5659 r0 *1 13.11,74.2
X$5659 23 38 FILLCELL_X8
* cell instance $5660 r0 *1 14.63,74.2
X$5660 23 38 FILLCELL_X2
* cell instance $5661 r0 *1 15.01,74.2
X$5661 23 38 FILLCELL_X1
* cell instance $5662 r0 *1 15.2,74.2
X$5662 1936 1446 1820 23 38 1988 MUX2_X1
* cell instance $5663 r0 *1 16.53,74.2
X$5663 23 38 FILLCELL_X4
* cell instance $5664 r0 *1 17.29,74.2
X$5664 23 38 FILLCELL_X1
* cell instance $5665 r0 *1 17.48,74.2
X$5665 1936 1184 1937 23 38 1938 MUX2_X1
* cell instance $5666 r0 *1 18.81,74.2
X$5666 23 38 FILLCELL_X1
* cell instance $5667 r0 *1 19,74.2
X$5667 1909 23 38 1848 CLKBUF_X3
* cell instance $5668 r0 *1 19.95,74.2
X$5668 1938 893 23 38 1991 NOR2_X1
* cell instance $5669 r0 *1 20.52,74.2
X$5669 23 2940 1939 1959 1848 38 DFF_X1
* cell instance $5670 m0 *1 22.04,74.2
X$5670 23 38 FILLCELL_X16
* cell instance $5671 m0 *1 21.47,74.2
X$5671 1872 937 23 38 1992 NOR2_X1
* cell instance $5672 m0 *1 25.08,74.2
X$5672 23 38 FILLCELL_X4
* cell instance $5673 m0 *1 25.84,74.2
X$5673 23 38 FILLCELL_X2
* cell instance $5674 r0 *1 23.75,74.2
X$5674 1939 1434 1822 23 38 1959 MUX2_X1
* cell instance $5675 r0 *1 25.08,74.2
X$5675 23 38 FILLCELL_X4
* cell instance $5676 r0 *1 25.84,74.2
X$5676 23 38 FILLCELL_X2
* cell instance $5677 m0 *1 1.33,12.6
X$5677 23 38 FILLCELL_X32
* cell instance $5678 m0 *1 1.14,12.6
X$5678 23 38 23 38 TAPCELL_X1
* cell instance $5679 m0 *1 7.41,12.6
X$5679 23 38 FILLCELL_X4
* cell instance $5680 m0 *1 11.4,12.6
X$5680 201 212 202 23 38 245 MUX2_X1
* cell instance $5681 m0 *1 12.73,12.6
X$5681 23 38 FILLCELL_X4
* cell instance $5682 m0 *1 13.49,12.6
X$5682 23 38 FILLCELL_X1
* cell instance $5683 m0 *1 13.68,12.6
X$5683 107 155 270 23 38 271 MUX2_X1
* cell instance $5684 m0 *1 18.24,12.6
X$5684 23 38 FILLCELL_X1
* cell instance $5685 m0 *1 18.43,12.6
X$5685 24 171 250 23 38 205 MUX2_X1
* cell instance $5686 m0 *1 19.76,12.6
X$5686 23 38 FILLCELL_X2
* cell instance $5687 r0 *1 1.14,12.6
X$5687 23 38 23 38 TAPCELL_X1
* cell instance $5688 r0 *1 1.33,12.6
X$5688 23 38 FILLCELL_X8
* cell instance $5689 r0 *1 2.85,12.6
X$5689 23 38 FILLCELL_X2
* cell instance $5690 r0 *1 3.14,12.6
X$5690 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $5691 r0 *1 3.14,12.6
X$5691 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $5692 r0 *1 3.14,12.6
X$5692 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $5693 r0 *1 3.23,12.6
X$5693 23 38 FILLCELL_X1
* cell instance $5694 r0 *1 6.65,12.6
X$5694 23 38 FILLCELL_X8
* cell instance $5695 r0 *1 8.17,12.6
X$5695 23 38 FILLCELL_X4
* cell instance $5696 r0 *1 8.93,12.6
X$5696 23 38 FILLCELL_X2
* cell instance $5697 r0 *1 9.31,12.6
X$5697 107 171 246 23 38 269 MUX2_X1
* cell instance $5698 r0 *1 13.87,12.6
X$5698 246 212 270 23 38 321 MUX2_X1
* cell instance $5699 r0 *1 15.2,12.6
X$5699 23 38 FILLCELL_X8
* cell instance $5700 r0 *1 16.72,12.6
X$5700 23 38 FILLCELL_X4
* cell instance $5701 r0 *1 17.48,12.6
X$5701 23 38 FILLCELL_X2
* cell instance $5702 r0 *1 17.86,12.6
X$5702 204 248 23 38 323 NOR2_X1
* cell instance $5703 r0 *1 18.43,12.6
X$5703 23 38 FILLCELL_X8
* cell instance $5704 r0 *1 19.95,12.6
X$5704 23 38 FILLCELL_X4
* cell instance $5705 m0 *1 23.37,12.6
X$5705 23 38 FILLCELL_X4
* cell instance $5706 m0 *1 24.13,12.6
X$5706 23 38 FILLCELL_X1
* cell instance $5707 m0 *1 24.32,12.6
X$5707 26 171 206 23 38 168 MUX2_X1
* cell instance $5708 m0 *1 25.65,12.6
X$5708 206 212 165 23 38 276 MUX2_X1
* cell instance $5709 m0 *1 26.98,12.6
X$5709 23 38 FILLCELL_X8
* cell instance $5710 m0 *1 28.5,12.6
X$5710 23 38 FILLCELL_X4
* cell instance $5711 m0 *1 29.26,12.6
X$5711 23 38 FILLCELL_X1
* cell instance $5712 m0 *1 29.45,12.6
X$5712 29 171 209 23 38 208 MUX2_X1
* cell instance $5713 m0 *1 30.78,12.6
X$5713 209 212 169 23 38 252 MUX2_X1
* cell instance $5714 m0 *1 32.11,12.6
X$5714 149 23 38 73 CLKBUF_X3
* cell instance $5715 m0 *1 33.06,12.6
X$5715 73 23 38 CLKBUF_X1
* cell instance $5716 m0 *1 33.63,12.6
X$5716 25 155 235 23 38 210 MUX2_X1
* cell instance $5717 m0 *1 34.96,12.6
X$5717 170 212 235 23 38 279 MUX2_X1
* cell instance $5718 m0 *1 36.29,12.6
X$5718 23 38 FILLCELL_X8
* cell instance $5719 m0 *1 37.81,12.6
X$5719 23 38 FILLCELL_X4
* cell instance $5720 m0 *1 38.57,12.6
X$5720 98 171 214 23 38 213 MUX2_X1
* cell instance $5721 m0 *1 39.9,12.6
X$5721 214 212 157 23 38 255 MUX2_X1
* cell instance $5722 m0 *1 41.23,12.6
X$5722 23 38 FILLCELL_X8
* cell instance $5723 m0 *1 42.75,12.6
X$5723 23 38 FILLCELL_X1
* cell instance $5724 m0 *1 42.94,12.6
X$5724 172 212 216 23 38 280 MUX2_X1
* cell instance $5725 m0 *1 44.27,12.6
X$5725 75 155 216 23 38 215 MUX2_X1
* cell instance $5726 m0 *1 45.6,12.6
X$5726 23 38 FILLCELL_X8
* cell instance $5727 m0 *1 47.12,12.6
X$5727 23 38 FILLCELL_X2
* cell instance $5728 r0 *1 20.71,12.6
X$5728 250 212 273 23 38 251 MUX2_X1
* cell instance $5729 r0 *1 22.04,12.6
X$5729 23 38 FILLCELL_X16
* cell instance $5730 r0 *1 25.08,12.6
X$5730 23 38 FILLCELL_X4
* cell instance $5731 r0 *1 25.84,12.6
X$5731 23 38 FILLCELL_X2
* cell instance $5732 r0 *1 26.22,12.6
X$5732 23 38 FILLCELL_X1
* cell instance $5733 r0 *1 26.41,12.6
X$5733 95 248 23 38 327 NOR2_X1
* cell instance $5734 r0 *1 26.98,12.6
X$5734 23 38 FILLCELL_X16
* cell instance $5735 r0 *1 30.02,12.6
X$5735 23 38 FILLCELL_X8
* cell instance $5736 r0 *1 31.54,12.6
X$5736 23 38 FILLCELL_X1
* cell instance $5737 r0 *1 31.73,12.6
X$5737 278 248 23 38 365 NOR2_X1
* cell instance $5738 r0 *1 32.3,12.6
X$5738 252 254 23 38 364 NOR2_X1
* cell instance $5739 r0 *1 32.87,12.6
X$5739 23 38 FILLCELL_X8
* cell instance $5740 r0 *1 34.39,12.6
X$5740 23 38 FILLCELL_X2
* cell instance $5741 r0 *1 34.77,12.6
X$5741 23 38 FILLCELL_X1
* cell instance $5742 r0 *1 34.96,12.6
X$5742 279 254 23 38 253 NOR2_X1
* cell instance $5743 r0 *1 35.53,12.6
X$5743 23 38 FILLCELL_X16
* cell instance $5744 r0 *1 38.57,12.6
X$5744 23 38 FILLCELL_X8
* cell instance $5745 r0 *1 40.09,12.6
X$5745 23 38 FILLCELL_X2
* cell instance $5746 r0 *1 40.47,12.6
X$5746 23 38 FILLCELL_X1
* cell instance $5747 r0 *1 40.66,12.6
X$5747 255 254 23 38 331 NOR2_X1
* cell instance $5748 r0 *1 41.23,12.6
X$5748 23 38 FILLCELL_X8
* cell instance $5749 r0 *1 42.75,12.6
X$5749 23 38 FILLCELL_X4
* cell instance $5750 r0 *1 43.51,12.6
X$5750 23 38 FILLCELL_X2
* cell instance $5751 r0 *1 43.89,12.6
X$5751 23 38 FILLCELL_X1
* cell instance $5752 r0 *1 44.08,12.6
X$5752 280 254 23 38 430 NOR2_X1
* cell instance $5753 r0 *1 44.65,12.6
X$5753 23 38 FILLCELL_X8
* cell instance $5754 r0 *1 46.17,12.6
X$5754 23 38 FILLCELL_X4
* cell instance $5755 r0 *1 46.93,12.6
X$5755 23 38 FILLCELL_X1
* cell instance $5756 r0 *1 47.12,12.6
X$5756 23 3098 302 282 30 38 DFF_X1
* cell instance $5757 m0 *1 50.73,12.6
X$5757 23 38 FILLCELL_X2
* cell instance $5758 m0 *1 47.5,12.6
X$5758 23 2725 259 258 30 38 DFF_X1
* cell instance $5759 r0 *1 50.35,12.6
X$5759 23 38 FILLCELL_X4
* cell instance $5760 m0 *1 52.06,12.6
X$5760 23 38 FILLCELL_X16
* cell instance $5761 m0 *1 51.11,12.6
X$5761 286 23 38 171 CLKBUF_X3
* cell instance $5762 m0 *1 55.1,12.6
X$5762 23 38 FILLCELL_X8
* cell instance $5763 m0 *1 56.62,12.6
X$5763 23 38 FILLCELL_X1
* cell instance $5764 m0 *1 56.81,12.6
X$5764 121 286 218 23 38 217 MUX2_X1
* cell instance $5765 m0 *1 58.14,12.6
X$5765 23 2839 219 287 76 38 DFF_X1
* cell instance $5766 m0 *1 61.37,12.6
X$5766 23 38 FILLCELL_X2
* cell instance $5767 r0 *1 51.11,12.6
X$5767 23 38 FILLCELL_X2
* cell instance $5768 r0 *1 51.49,12.6
X$5768 100 248 23 38 390 NOR2_X1
* cell instance $5769 r0 *1 52.06,12.6
X$5769 23 38 FILLCELL_X32
* cell instance $5770 r0 *1 58.14,12.6
X$5770 23 38 FILLCELL_X16
* cell instance $5771 r0 *1 59.14,12.6
X$5771 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $5772 r0 *1 59.14,12.6
X$5772 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $5773 r0 *1 59.14,12.6
X$5773 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $5774 r0 *1 61.18,12.6
X$5774 23 38 FILLCELL_X8
* cell instance $5775 m0 *1 61.94,12.6
X$5775 219 223 48 23 38 287 MUX2_X1
* cell instance $5776 m0 *1 61.75,12.6
X$5776 23 38 FILLCELL_X1
* cell instance $5777 m0 *1 63.27,12.6
X$5777 219 188 220 23 38 291 MUX2_X1
* cell instance $5778 m0 *1 64.6,12.6
X$5778 23 38 FILLCELL_X4
* cell instance $5779 m0 *1 65.36,12.6
X$5779 23 38 FILLCELL_X2
* cell instance $5780 r0 *1 62.7,12.6
X$5780 23 38 FILLCELL_X4
* cell instance $5781 r0 *1 63.46,12.6
X$5781 23 38 FILLCELL_X2
* cell instance $5782 r0 *1 63.84,12.6
X$5782 48 260 316 23 38 304 MUX2_X1
* cell instance $5783 r0 *1 65.17,12.6
X$5783 23 38 FILLCELL_X4
* cell instance $5784 m0 *1 68.97,12.6
X$5784 23 38 FILLCELL_X4
* cell instance $5785 m0 *1 65.74,12.6
X$5785 23 2716 290 241 153 38 DFF_X1
* cell instance $5786 m0 *1 69.73,12.6
X$5786 291 261 23 38 239 NOR2_X1
* cell instance $5787 m0 *1 70.3,12.6
X$5787 23 38 FILLCELL_X8
* cell instance $5788 m0 *1 71.82,12.6
X$5788 23 38 FILLCELL_X1
* cell instance $5789 m0 *1 72.01,12.6
X$5789 23 2691 237 238 34 38 DFF_X1
* cell instance $5790 m0 *1 75.24,12.6
X$5790 221 274 23 38 222 NOR2_X1
* cell instance $5791 m0 *1 75.81,12.6
X$5791 23 38 FILLCELL_X16
* cell instance $5792 m0 *1 78.85,12.6
X$5792 23 38 FILLCELL_X4
* cell instance $5793 m0 *1 79.61,12.6
X$5793 23 38 FILLCELL_X2
* cell instance $5794 r0 *1 65.93,12.6
X$5794 23 38 FILLCELL_X1
* cell instance $5795 r0 *1 66.12,12.6
X$5795 23 2941 315 288 153 38 DFF_X1
* cell instance $5796 r0 *1 69.35,12.6
X$5796 23 38 FILLCELL_X2
* cell instance $5797 r0 *1 69.73,12.6
X$5797 49 240 345 23 38 292 MUX2_X1
* cell instance $5798 r0 *1 71.06,12.6
X$5798 23 38 FILLCELL_X8
* cell instance $5799 r0 *1 72.58,12.6
X$5799 23 38 FILLCELL_X2
* cell instance $5800 r0 *1 72.96,12.6
X$5800 227 239 289 225 222 175 23 38 285 OAI33_X1
* cell instance $5801 r0 *1 74.29,12.6
X$5801 237 263 176 23 38 221 MUX2_X1
* cell instance $5802 r0 *1 75.62,12.6
X$5802 23 38 FILLCELL_X16
* cell instance $5803 r0 *1 78.66,12.6
X$5803 23 38 FILLCELL_X4
* cell instance $5804 r0 *1 79.42,12.6
X$5804 23 38 FILLCELL_X2
* cell instance $5805 r0 *1 79.8,12.6
X$5805 53 240 307 23 38 314 MUX2_X1
* cell instance $5806 m0 *1 81.32,12.6
X$5806 23 38 FILLCELL_X2
* cell instance $5807 m0 *1 79.99,12.6
X$5807 284 223 78 23 38 234 MUX2_X1
* cell instance $5808 r0 *1 81.13,12.6
X$5808 23 38 FILLCELL_X32
* cell instance $5809 m0 *1 81.89,12.6
X$5809 284 188 178 23 38 283 MUX2_X1
* cell instance $5810 m0 *1 81.7,12.6
X$5810 23 38 FILLCELL_X1
* cell instance $5811 m0 *1 83.22,12.6
X$5811 23 38 FILLCELL_X8
* cell instance $5812 m0 *1 84.74,12.6
X$5812 283 261 23 38 232 NOR2_X1
* cell instance $5813 m0 *1 85.31,12.6
X$5813 23 38 FILLCELL_X2
* cell instance $5814 m0 *1 87.02,12.6
X$5814 23 38 FILLCELL_X2
* cell instance $5815 m0 *1 85.69,12.6
X$5815 183 223 52 23 38 224 MUX2_X1
* cell instance $5816 r0 *1 87.21,12.6
X$5816 23 38 FILLCELL_X4
* cell instance $5817 m0 *1 87.4,12.6
X$5817 23 38 FILLCELL_X1
* cell instance $5818 m0 *1 87.59,12.6
X$5818 227 232 181 225 281 182 23 38 265 OAI33_X1
* cell instance $5819 m0 *1 88.92,12.6
X$5819 23 38 FILLCELL_X2
* cell instance $5820 r0 *1 87.97,12.6
X$5820 23 38 FILLCELL_X2
* cell instance $5821 r0 *1 88.35,12.6
X$5821 264 274 23 38 281 NOR2_X1
* cell instance $5822 r0 *1 88.92,12.6
X$5822 23 38 FILLCELL_X8
* cell instance $5823 m0 *1 89.49,12.6
X$5823 226 261 23 38 228 NOR2_X1
* cell instance $5824 m0 *1 89.3,12.6
X$5824 23 38 FILLCELL_X1
* cell instance $5825 m0 *1 90.06,12.6
X$5825 227 228 231 225 266 229 23 38 277 OAI33_X1
* cell instance $5826 m0 *1 91.39,12.6
X$5826 23 2665 267 275 83 38 DFF_X1
* cell instance $5827 m0 *1 94.62,12.6
X$5827 23 38 FILLCELL_X4
* cell instance $5828 m0 *1 95.38,12.6
X$5828 23 38 FILLCELL_X2
* cell instance $5829 r0 *1 90.44,12.6
X$5829 23 38 FILLCELL_X4
* cell instance $5830 r0 *1 91.2,12.6
X$5830 272 274 23 38 266 NOR2_X1
* cell instance $5831 r0 *1 91.77,12.6
X$5831 53 191 267 23 38 275 MUX2_X1
* cell instance $5832 r0 *1 93.1,12.6
X$5832 267 263 185 23 38 272 MUX2_X1
* cell instance $5833 r0 *1 94.43,12.6
X$5833 23 38 FILLCELL_X8
* cell instance $5834 m0 *1 95.95,12.6
X$5834 160 23 38 377 BUF_X1
* cell instance $5835 m0 *1 95.76,12.6
X$5835 23 38 FILLCELL_X1
* cell instance $5836 m0 *1 96.52,12.6
X$5836 23 38 FILLCELL_X2
* cell instance $5837 r0 *1 95.95,12.6
X$5837 23 38 FILLCELL_X4
* cell instance $5838 r0 *1 96.71,12.6
X$5838 23 38 FILLCELL_X2
* cell instance $5839 r180 *1 97.28,12.6
X$5839 23 38 23 38 TAPCELL_X1
* cell instance $5840 m0 *1 96.9,12.6
X$5840 23 38 FILLCELL_X1
* cell instance $5841 m90 *1 97.28,12.6
X$5841 23 38 23 38 TAPCELL_X1
* cell instance $5842 m0 *1 1.33,96.6
X$5842 23 38 FILLCELL_X32
* cell instance $5843 m0 *1 1.14,96.6
X$5843 23 38 23 38 TAPCELL_X1
* cell instance $5844 m0 *1 7.41,96.6
X$5844 23 38 FILLCELL_X16
* cell instance $5845 m0 *1 10.45,96.6
X$5845 23 38 FILLCELL_X8
* cell instance $5846 m0 *1 11.97,96.6
X$5846 23 38 FILLCELL_X4
* cell instance $5847 m0 *1 12.73,96.6
X$5847 23 38 FILLCELL_X2
* cell instance $5848 r0 *1 3.14,96.6
X$5848 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $5849 r0 *1 3.14,96.6
X$5849 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $5850 r0 *1 3.14,96.6
X$5850 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $5851 m0 *1 1.33,91
X$5851 23 38 FILLCELL_X32
* cell instance $5852 m0 *1 1.14,91
X$5852 23 38 23 38 TAPCELL_X1
* cell instance $5853 m0 *1 7.41,91
X$5853 23 38 FILLCELL_X16
* cell instance $5854 m0 *1 10.45,91
X$5854 23 38 FILLCELL_X1
* cell instance $5855 m0 *1 10.64,91
X$5855 2418 1535 23 38 2419 NOR2_X1
* cell instance $5856 m0 *1 11.21,91
X$5856 23 38 FILLCELL_X4
* cell instance $5857 m0 *1 11.97,91
X$5857 1425 2350 2349 548 2419 2351 23 38 2081 OAI33_X1
* cell instance $5858 m0 *1 13.3,91
X$5858 23 38 FILLCELL_X16
* cell instance $5859 m0 *1 16.34,91
X$5859 23 38 FILLCELL_X8
* cell instance $5860 m0 *1 17.86,91
X$5860 23 38 FILLCELL_X2
* cell instance $5861 r0 *1 1.14,91
X$5861 23 38 23 38 TAPCELL_X1
* cell instance $5862 r0 *1 1.33,91
X$5862 23 38 FILLCELL_X16
* cell instance $5863 r0 *1 3.14,91
X$5863 23 VIA_via1_2_960_340_1_3_300_300
* cell instance $5864 r0 *1 3.14,91
X$5864 23 VIA_via2_3_960_340_1_3_320_320
* cell instance $5865 r0 *1 3.14,91
X$5865 23 VIA_via3_4_960_340_1_3_320_320
* cell instance $5866 r0 *1 4.37,91
X$5866 23 38 FILLCELL_X4
* cell instance $5867 r0 *1 5.13,91
X$5867 23 2968 2432 2460 2045 38 DFF_X1
* cell instance $5868 r0 *1 8.36,91
X$5868 2199 1406 2432 23 38 2460 MUX2_X1
* cell instance $5869 r0 *1 9.69,91
X$5869 23 38 FILLCELL_X2
* cell instance $5870 r0 *1 10.07,91
X$5870 23 38 FILLCELL_X1
* cell instance $5871 r0 *1 10.26,91
X$5871 2199 1493 2433 23 38 2461 MUX2_X1
* cell instance $5872 r0 *1 11.59,91
X$5872 23 38 FILLCELL_X1
* cell instance $5873 r0 *1 11.78,91
X$5873 2433 1373 2463 23 38 2464 MUX2_X1
* cell instance $5874 r0 *1 13.11,91
X$5874 2464 1483 23 38 2351 NOR2_X1
* cell instance $5875 r0 *1 13.68,91
X$5875 23 38 FILLCELL_X1
* cell instance $5876 r0 *1 13.87,91
X$5876 1909 23 38 2434 CLKBUF_X3
* cell instance $5877 r0 *1 14.82,91
X$5877 23 38 FILLCELL_X1
* cell instance $5878 r0 *1 15.01,91
X$5878 23 2964 2475 2465 2434 38 DFF_X1
* cell instance $5879 m0 *1 18.43,91
X$5879 2466 1535 23 38 2421 NOR2_X1
* cell instance $5880 m0 *1 18.24,91
X$5880 23 38 FILLCELL_X1
* cell instance $5881 m0 *1 19,91
X$5881 23 38 FILLCELL_X2
* cell instance $5882 r0 *1 18.24,91
X$5882 23 38 FILLCELL_X4
* cell instance $5883 r0 *1 19,91
X$5883 23 38 FILLCELL_X1
* cell instance $5884 r0 *1 19.19,91
X$5884 2217 1480 2437 23 38 2436 MUX2_X1
* cell instance $5885 m0 *1 20.71,91
X$5885 23 38 FILLCELL_X1
* cell instance $5886 m0 *1 19.38,91
X$5886 1425 2381 2420 548 2421 2352 23 38 1972 OAI33_X1
* cell instance $5887 m0 *1 20.9,91
X$5887 2353 1483 23 38 2352 NOR2_X1
* cell instance $5888 m0 *1 21.47,91
X$5888 23 38 FILLCELL_X32
* cell instance $5889 m0 *1 27.55,91
X$5889 23 38 FILLCELL_X2
* cell instance $5890 r0 *1 20.52,91
X$5890 2438 1373 2437 23 38 2353 MUX2_X1
* cell instance $5891 r0 *1 21.85,91
X$5891 23 3016 2438 2439 2144 38 DFF_X1
* cell instance $5892 r0 *1 25.08,91
X$5892 23 38 FILLCELL_X4
* cell instance $5893 r0 *1 25.84,91
X$5893 23 38 FILLCELL_X2
* cell instance $5894 r0 *1 26.22,91
X$5894 2218 1480 2440 23 38 2490 MUX2_X1
* cell instance $5895 r0 *1 27.55,91
X$5895 23 38 FILLCELL_X2
* cell instance $5896 r0 *1 80.94,1.4
X$5896 23 38 FILLCELL_X32
* cell instance $5897 r0 *1 87.02,1.4
X$5897 23 38 FILLCELL_X16
* cell instance $5898 r0 *1 90.06,1.4
X$5898 23 38 FILLCELL_X8
* cell instance $5899 r0 *1 91.58,1.4
X$5899 23 38 FILLCELL_X4
* cell instance $5900 r0 *1 93.1,1.4
X$5900 23 38 FILLCELL_X16
* cell instance $5901 r0 *1 96.14,1.4
X$5901 23 38 FILLCELL_X4
* cell instance $5902 r0 *1 96.9,1.4
X$5902 23 38 FILLCELL_X1
* cell instance $5903 m90 *1 97.28,1.4
X$5903 23 38 23 38 TAPCELL_X1
* cell instance $5904 r0 *1 19.095,4.83
X$5904 24 VIA_via2_5
* cell instance $5905 r0 *1 19.095,2.59
X$5905 24 VIA_via2_5
* cell instance $5906 r0 *1 19.095,10.29
X$5906 24 VIA_via2_5
* cell instance $5907 r0 *1 18.715,11.13
X$5907 24 VIA_via2_5
* cell instance $5908 r0 *1 19.095,11.13
X$5908 24 VIA_via2_5
* cell instance $5909 r0 *1 17.765,27.09
X$5909 24 VIA_via2_5
* cell instance $5910 r0 *1 21.185,25.97
X$5910 24 VIA_via2_5
* cell instance $5911 r0 *1 21.945,4.83
X$5911 24 VIA_via1_4
* cell instance $5912 r0 *1 21.945,4.83
X$5912 24 VIA_via2_5
* cell instance $5913 r0 *1 9.975,2.45
X$5913 24 VIA_via1_4
* cell instance $5914 r0 *1 9.975,2.45
X$5914 24 VIA_via2_5
* cell instance $5915 r0 *1 21.565,10.43
X$5915 24 VIA_via1_4
* cell instance $5916 r0 *1 21.565,10.29
X$5916 24 VIA_via2_5
* cell instance $5917 r0 *1 18.905,6.37
X$5917 24 VIA_via1_4
* cell instance $5918 r0 *1 18.715,11.97
X$5918 24 VIA_via1_4
* cell instance $5919 r0 *1 18.715,11.97
X$5919 24 VIA_via2_5
* cell instance $5920 r0 *1 18.855,11.97
X$5920 24 VIA_via3_2
* cell instance $5921 r0 *1 9.975,27.23
X$5921 24 VIA_via1_4
* cell instance $5922 r0 *1 9.975,27.09
X$5922 24 VIA_via2_5
* cell instance $5923 r0 *1 17.765,25.97
X$5923 24 VIA_via1_4
* cell instance $5924 r0 *1 17.765,25.97
X$5924 24 VIA_via2_5
* cell instance $5925 r0 *1 20.995,28.77
X$5925 24 VIA_via1_4
* cell instance $5926 r0 *1 18.855,25.97
X$5926 24 VIA_via3_2
* cell instance $5927 r0 *1 34.105,29.61
X$5927 25 VIA_via2_5
* cell instance $5928 r0 *1 32.775,6.65
X$5928 25 VIA_via2_5
* cell instance $5929 r0 *1 33.915,6.65
X$5929 25 VIA_via2_5
* cell instance $5930 r0 *1 35.625,6.65
X$5930 25 VIA_via2_5
* cell instance $5931 r0 *1 32.775,6.37
X$5931 25 VIA_via1_4
* cell instance $5932 r0 *1 35.625,9.17
X$5932 25 VIA_via1_4
* cell instance $5933 r0 *1 33.915,11.97
X$5933 25 VIA_via1_4
* cell instance $5934 r0 *1 33.345,2.45
X$5934 25 VIA_via1_4
* cell instance $5935 r0 *1 35.625,4.83
X$5935 25 VIA_via1_4
* cell instance $5936 r0 *1 32.965,30.03
X$5936 25 VIA_via1_4
* cell instance $5937 r0 *1 32.965,29.89
X$5937 25 VIA_via2_5
* cell instance $5938 r0 *1 33.915,30.03
X$5938 25 VIA_via1_4
* cell instance $5939 r0 *1 34.485,27.23
X$5939 25 VIA_via1_4
* cell instance $5940 r0 *1 24.605,2.45
X$5940 26 VIA_via2_5
* cell instance $5941 r0 *1 24.795,27.65
X$5941 26 VIA_via2_5
* cell instance $5942 r0 *1 24.985,16.31
X$5942 26 VIA_via2_5
* cell instance $5943 r0 *1 25.175,2.45
X$5943 26 VIA_via2_5
* cell instance $5944 r0 *1 24.605,16.31
X$5944 26 VIA_via2_5
* cell instance $5945 r0 *1 24.605,8.89
X$5945 26 VIA_via2_5
* cell instance $5946 r0 *1 22.895,8.89
X$5946 26 VIA_via2_5
* cell instance $5947 r0 *1 23.085,27.65
X$5947 26 VIA_via2_5
* cell instance $5948 r0 *1 22.325,28.77
X$5948 26 VIA_via2_5
* cell instance $5949 r0 *1 19.285,2.45
X$5949 26 VIA_via1_4
* cell instance $5950 r0 *1 19.285,2.45
X$5950 26 VIA_via2_5
* cell instance $5951 r0 *1 24.605,11.97
X$5951 26 VIA_via1_4
* cell instance $5952 r0 *1 24.605,6.37
X$5952 26 VIA_via1_4
* cell instance $5953 r0 *1 22.895,9.17
X$5953 26 VIA_via1_4
* cell instance $5954 r0 *1 25.175,3.57
X$5954 26 VIA_via1_4
* cell instance $5955 r0 *1 23.085,28.77
X$5955 26 VIA_via1_4
* cell instance $5956 r0 *1 23.085,28.77
X$5956 26 VIA_via2_5
* cell instance $5957 r0 *1 22.135,30.03
X$5957 26 VIA_via1_4
* cell instance $5958 r0 *1 24.795,27.23
X$5958 26 VIA_via1_4
* cell instance $5959 r0 *1 14.345,8.89
X$5959 27 VIA_via2_5
* cell instance $5960 r0 *1 15.675,8.89
X$5960 27 VIA_via2_5
* cell instance $5961 r0 *1 15.865,8.89
X$5961 27 VIA_via2_5
* cell instance $5962 r0 *1 11.685,27.23
X$5962 27 VIA_via2_5
* cell instance $5963 r0 *1 13.775,3.29
X$5963 27 VIA_via2_5
* cell instance $5964 r0 *1 15.675,3.29
X$5964 27 VIA_via2_5
* cell instance $5965 r0 *1 12.445,8.89
X$5965 27 VIA_via2_5
* cell instance $5966 r0 *1 14.345,27.23
X$5966 27 VIA_via2_5
* cell instance $5967 r0 *1 8.835,3.29
X$5967 27 VIA_via2_5
* cell instance $5968 r0 *1 8.835,2.45
X$5968 27 VIA_via1_4
* cell instance $5969 r0 *1 14.345,9.17
X$5969 27 VIA_via1_4
* cell instance $5970 r0 *1 15.675,4.83
X$5970 27 VIA_via1_4
* cell instance $5971 r0 *1 13.775,3.57
X$5971 27 VIA_via1_4
* cell instance $5972 r0 *1 15.675,10.43
X$5972 27 VIA_via1_4
* cell instance $5973 r0 *1 12.065,16.03
X$5973 27 VIA_via1_4
* cell instance $5974 r0 *1 8.645,27.23
X$5974 27 VIA_via1_4
* cell instance $5975 r0 *1 8.645,27.23
X$5975 27 VIA_via2_5
* cell instance $5976 r0 *1 14.345,30.03
X$5976 27 VIA_via1_4
* cell instance $5977 r0 *1 20.045,3.57
X$5977 28 VIA_via2_5
* cell instance $5978 r0 *1 16.435,6.37
X$5978 28 VIA_via2_5
* cell instance $5979 r0 *1 14.155,7.63
X$5979 28 VIA_via2_5
* cell instance $5980 r0 *1 16.435,8.33
X$5980 28 VIA_via2_5
* cell instance $5981 r0 *1 17.005,8.33
X$5981 28 VIA_via2_5
* cell instance $5982 r0 *1 16.815,3.57
X$5982 28 VIA_via2_5
* cell instance $5983 r0 *1 11.685,7.63
X$5983 28 VIA_via2_5
* cell instance $5984 r0 *1 11.685,10.43
X$5984 28 VIA_via1_4
* cell instance $5985 r0 *1 21.375,3.57
X$5985 28 VIA_via1_4
* cell instance $5986 r0 *1 21.375,3.57
X$5986 28 VIA_via2_5
* cell instance $5987 r0 *1 10.355,7.63
X$5987 28 VIA_via1_4
* cell instance $5988 r0 *1 10.355,7.63
X$5988 28 VIA_via2_5
* cell instance $5989 r0 *1 20.045,4.83
X$5989 28 VIA_via1_4
* cell instance $5990 r0 *1 16.435,7.63
X$5990 28 VIA_via1_4
* cell instance $5991 r0 *1 14.155,6.37
X$5991 28 VIA_via1_4
* cell instance $5992 r0 *1 14.155,6.37
X$5992 28 VIA_via2_5
* cell instance $5993 r0 *1 16.815,5.95
X$5993 28 VIA_via1_4
* cell instance $5994 r0 *1 16.435,6.65
X$5994 28 VIA_via1_4
* cell instance $5995 r0 *1 17.195,3.57
X$5995 28 VIA_via1_4
* cell instance $5996 r0 *1 17.195,3.57
X$5996 28 VIA_via2_5
* cell instance $5997 r0 *1 17.005,9.17
X$5997 28 VIA_via1_4
* cell instance $5998 r0 *1 28.405,2.59
X$5998 29 VIA_via1_7
* cell instance $5999 r0 *1 29.165,10.57
X$5999 29 VIA_via2_5
* cell instance $6000 r0 *1 29.165,11.97
X$6000 29 VIA_via2_5
* cell instance $6001 r0 *1 29.355,6.37
X$6001 29 VIA_via1_4
* cell instance $6002 r0 *1 29.735,11.97
X$6002 29 VIA_via1_4
* cell instance $6003 r0 *1 29.735,11.97
X$6003 29 VIA_via2_5
* cell instance $6004 r0 *1 28.405,10.43
X$6004 29 VIA_via1_4
* cell instance $6005 r0 *1 28.405,10.57
X$6005 29 VIA_via2_5
* cell instance $6006 r0 *1 27.455,3.57
X$6006 29 VIA_via1_4
* cell instance $6007 r0 *1 27.265,28.77
X$6007 29 VIA_via1_4
* cell instance $6008 r0 *1 27.265,28.77
X$6008 29 VIA_via2_5
* cell instance $6009 r0 *1 28.975,28.77
X$6009 29 VIA_via1_4
* cell instance $6010 r0 *1 28.975,28.77
X$6010 29 VIA_via2_5
* cell instance $6011 r0 *1 28.975,25.97
X$6011 29 VIA_via1_4
* cell instance $6012 r0 *1 49.115,8.75
X$6012 30 VIA_via2_5
* cell instance $6013 r0 *1 46.075,3.57
X$6013 30 VIA_via2_5
* cell instance $6014 r0 *1 43.225,8.75
X$6014 30 VIA_via2_5
* cell instance $6015 r0 *1 46.075,8.75
X$6015 30 VIA_via2_5
* cell instance $6016 r0 *1 45.505,8.75
X$6016 30 VIA_via2_5
* cell instance $6017 r0 *1 47.405,8.75
X$6017 30 VIA_via2_5
* cell instance $6018 r0 *1 48.735,13.23
X$6018 30 VIA_via1_4
* cell instance $6019 r0 *1 49.115,11.97
X$6019 30 VIA_via1_4
* cell instance $6020 r0 *1 47.405,9.17
X$6020 30 VIA_via1_4
* cell instance $6021 r0 *1 43.225,9.17
X$6021 30 VIA_via1_4
* cell instance $6022 r0 *1 45.505,10.43
X$6022 30 VIA_via1_4
* cell instance $6023 r0 *1 46.835,8.75
X$6023 30 VIA_via1_4
* cell instance $6024 r0 *1 46.835,8.75
X$6024 30 VIA_via2_5
* cell instance $6025 r0 *1 44.555,3.57
X$6025 30 VIA_via1_4
* cell instance $6026 r0 *1 44.555,3.57
X$6026 30 VIA_via2_5
* cell instance $6027 r0 *1 43.795,4.83
X$6027 30 VIA_via1_4
* cell instance $6028 r0 *1 49.305,3.57
X$6028 30 VIA_via1_4
* cell instance $6029 r0 *1 49.305,3.57
X$6029 30 VIA_via2_5
* cell instance $6030 r0 *1 45.505,5.11
X$6030 31 VIA_via2_5
* cell instance $6031 r0 *1 46.265,5.11
X$6031 31 VIA_via2_5
* cell instance $6032 r0 *1 45.885,5.11
X$6032 31 VIA_via2_5
* cell instance $6033 r0 *1 45.505,6.37
X$6033 31 VIA_via1_4
* cell instance $6034 r0 *1 46.075,3.29
X$6034 31 VIA_via1_4
* cell instance $6035 r0 *1 46.265,4.83
X$6035 31 VIA_via1_4
* cell instance $6036 r0 *1 66.595,6.37
X$6036 32 VIA_via2_5
* cell instance $6037 r0 *1 69.255,3.57
X$6037 32 VIA_via2_5
* cell instance $6038 r0 *1 67.545,3.57
X$6038 32 VIA_via2_5
* cell instance $6039 r0 *1 62.035,7.35
X$6039 32 VIA_via2_5
* cell instance $6040 r0 *1 64.125,3.57
X$6040 32 VIA_via2_5
* cell instance $6041 r0 *1 69.255,2.03
X$6041 32 VIA_via1_4
* cell instance $6042 r0 *1 67.545,6.37
X$6042 32 VIA_via1_4
* cell instance $6043 r0 *1 67.545,6.37
X$6043 32 VIA_via2_5
* cell instance $6044 r0 *1 61.085,3.57
X$6044 32 VIA_via1_4
* cell instance $6045 r0 *1 61.085,3.57
X$6045 32 VIA_via2_5
* cell instance $6046 r0 *1 64.125,6.37
X$6046 32 VIA_via1_4
* cell instance $6047 r0 *1 62.035,9.17
X$6047 32 VIA_via1_4
* cell instance $6048 r0 *1 66.595,7.63
X$6048 32 VIA_via1_4
* cell instance $6049 r0 *1 64.505,7.35
X$6049 32 VIA_via1_4
* cell instance $6050 r0 *1 64.505,7.35
X$6050 32 VIA_via2_5
* cell instance $6051 r0 *1 64.125,4.83
X$6051 32 VIA_via1_4
* cell instance $6052 r0 *1 65.265,3.57
X$6052 32 VIA_via1_4
* cell instance $6053 r0 *1 65.265,3.57
X$6053 32 VIA_via2_5
* cell instance $6054 r0 *1 74.575,3.43
X$6054 33 VIA_via1_4
* cell instance $6055 r0 *1 74.575,3.43
X$6055 33 VIA_via2_5
* cell instance $6056 r0 *1 70.775,4.83
X$6056 33 VIA_via1_4
* cell instance $6057 r0 *1 70.965,3.57
X$6057 33 VIA_via1_4
* cell instance $6058 r0 *1 70.965,3.43
X$6058 33 VIA_via2_5
* cell instance $6059 r0 *1 76.475,8.33
X$6059 34 VIA_via2_5
* cell instance $6060 r0 *1 79.135,8.33
X$6060 34 VIA_via2_5
* cell instance $6061 r0 *1 76.475,7.63
X$6061 34 VIA_via2_5
* cell instance $6062 r0 *1 73.055,6.37
X$6062 34 VIA_via2_5
* cell instance $6063 r0 *1 74.765,7.63
X$6063 34 VIA_via2_5
* cell instance $6064 r0 *1 73.815,10.43
X$6064 34 VIA_via2_5
* cell instance $6065 r0 *1 76.475,10.43
X$6065 34 VIA_via2_5
* cell instance $6066 r0 *1 76.475,8.05
X$6066 34 VIA_via1_4
* cell instance $6067 r0 *1 79.135,9.17
X$6067 34 VIA_via1_4
* cell instance $6068 r0 *1 77.045,10.43
X$6068 34 VIA_via1_4
* cell instance $6069 r0 *1 77.045,10.43
X$6069 34 VIA_via2_5
* cell instance $6070 r0 *1 73.625,11.97
X$6070 34 VIA_via1_4
* cell instance $6071 r0 *1 75.525,7.63
X$6071 34 VIA_via1_4
* cell instance $6072 r0 *1 75.525,7.63
X$6072 34 VIA_via2_5
* cell instance $6073 r0 *1 77.615,2.03
X$6073 34 VIA_via1_4
* cell instance $6074 r0 *1 76.285,3.57
X$6074 34 VIA_via1_4
* cell instance $6075 r0 *1 74.765,6.37
X$6075 34 VIA_via1_4
* cell instance $6076 r0 *1 74.765,6.37
X$6076 34 VIA_via2_5
* cell instance $6077 r0 *1 73.055,3.57
X$6077 34 VIA_via1_4
* cell instance $6078 r0 *1 82.555,4.41
X$6078 35 VIA_via1_7
* cell instance $6079 r0 *1 83.125,3.57
X$6079 35 VIA_via1_4
* cell instance $6080 r0 *1 87.115,9.17
X$6080 36 VIA_via2_5
* cell instance $6081 r0 *1 85.405,9.17
X$6081 36 VIA_via2_5
* cell instance $6082 r0 *1 82.935,9.17
X$6082 36 VIA_via2_5
* cell instance $6083 r0 *1 79.705,9.17
X$6083 36 VIA_via2_5
* cell instance $6084 r0 *1 80.655,9.17
X$6084 36 VIA_via2_5
* cell instance $6085 r0 *1 82.935,7.63
X$6085 36 VIA_via1_4
* cell instance $6086 r0 *1 82.745,9.17
X$6086 36 VIA_via1_4
* cell instance $6087 r0 *1 82.745,9.17
X$6087 36 VIA_via2_5
* cell instance $6088 r0 *1 85.405,8.05
X$6088 36 VIA_via1_4
* cell instance $6089 r0 *1 80.655,10.43
X$6089 36 VIA_via1_4
* cell instance $6090 r0 *1 79.705,6.37
X$6090 36 VIA_via1_4
* cell instance $6091 r0 *1 83.885,3.57
X$6091 36 VIA_via1_4
* cell instance $6092 r0 *1 87.115,10.43
X$6092 36 VIA_via1_4
* cell instance $6093 r0 *1 85.975,9.17
X$6093 36 VIA_via1_4
* cell instance $6094 r0 *1 85.975,9.17
X$6094 36 VIA_via2_5
* cell instance $6095 r0 *1 49.685,49.63
X$6095 37 VIA_via1_4
* cell instance $6096 r0 *1 49.685,49.63
X$6096 37 VIA_via2_5
* cell instance $6097 r0 *1 72.335,3.43
X$6097 37 VIA_via4_0
* cell instance $6098 r0 *1 49.935,26.25
X$6098 37 VIA_via3_2
* cell instance $6099 r0 *1 49.935,49.63
X$6099 37 VIA_via3_2
* cell instance $6100 r0 *1 72.335,26.25
X$6100 37 VIA_via3_2
* cell instance $6101 r0 *1 31.14,67.2
X$6101 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6102 r0 *1 31.14,67.2
X$6102 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6103 r0 *1 31.14,67.2
X$6103 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6104 r0 *1 87.14,67.2
X$6104 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6105 r0 *1 87.14,67.2
X$6105 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6106 r0 *1 87.14,67.2
X$6106 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6107 r0 *1 87.14,14
X$6107 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6108 r0 *1 87.14,14
X$6108 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6109 r0 *1 87.14,14
X$6109 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6110 r0 *1 31.14,50.4
X$6110 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6111 r0 *1 31.14,50.4
X$6111 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6112 r0 *1 31.14,50.4
X$6112 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6113 r0 *1 87.14,50.4
X$6113 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6114 r0 *1 87.14,50.4
X$6114 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6115 r0 *1 87.14,50.4
X$6115 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6116 r0 *1 31.14,84
X$6116 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6117 r0 *1 31.14,84
X$6117 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6118 r0 *1 31.14,84
X$6118 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6119 r0 *1 87.14,84
X$6119 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6120 r0 *1 87.14,84
X$6120 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6121 r0 *1 87.14,84
X$6121 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6122 r0 *1 87.14,48.4
X$6122 38 VIA_via5_6_960_2800_5_2_600_600
* cell instance $6123 r0 *1 87.14,48.4
X$6123 38 VIA_via4_5_960_2800_5_2_600_600
* cell instance $6124 r0 *1 87.14,48.4
X$6124 38 VIA_via6_7_960_2800_4_1_600_600
* cell instance $6125 r0 *1 87.14,18.4
X$6125 38 VIA_via5_6_960_2800_5_2_600_600
* cell instance $6126 r0 *1 87.14,18.4
X$6126 38 VIA_via4_5_960_2800_5_2_600_600
* cell instance $6127 r0 *1 87.14,18.4
X$6127 38 VIA_via6_7_960_2800_4_1_600_600
* cell instance $6128 r0 *1 31.14,18.4
X$6128 38 VIA_via5_6_960_2800_5_2_600_600
* cell instance $6129 r0 *1 31.14,18.4
X$6129 38 VIA_via4_5_960_2800_5_2_600_600
* cell instance $6130 r0 *1 31.14,18.4
X$6130 38 VIA_via6_7_960_2800_4_1_600_600
* cell instance $6131 r0 *1 31.14,48.4
X$6131 38 VIA_via5_6_960_2800_5_2_600_600
* cell instance $6132 r0 *1 31.14,48.4
X$6132 38 VIA_via4_5_960_2800_5_2_600_600
* cell instance $6133 r0 *1 31.14,48.4
X$6133 38 VIA_via6_7_960_2800_4_1_600_600
* cell instance $6134 r0 *1 31.14,92.4
X$6134 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6135 r0 *1 31.14,92.4
X$6135 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6136 r0 *1 31.14,92.4
X$6136 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6137 r0 *1 87.14,92.4
X$6137 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6138 r0 *1 87.14,92.4
X$6138 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6139 r0 *1 87.14,92.4
X$6139 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6140 r0 *1 31.14,47.6
X$6140 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6141 r0 *1 31.14,47.6
X$6141 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6142 r0 *1 31.14,47.6
X$6142 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6143 r0 *1 87.14,47.6
X$6143 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6144 r0 *1 87.14,47.6
X$6144 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6145 r0 *1 87.14,47.6
X$6145 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6146 r0 *1 31.14,39.2
X$6146 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6147 r0 *1 31.14,39.2
X$6147 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6148 r0 *1 31.14,39.2
X$6148 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6149 r0 *1 87.14,39.2
X$6149 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6150 r0 *1 87.14,39.2
X$6150 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6151 r0 *1 87.14,39.2
X$6151 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6152 r0 *1 31.14,81.2
X$6152 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6153 r0 *1 31.14,81.2
X$6153 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6154 r0 *1 31.14,81.2
X$6154 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6155 r0 *1 31.14,44.8
X$6155 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6156 r0 *1 31.14,44.8
X$6156 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6157 r0 *1 31.14,44.8
X$6157 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6158 r0 *1 87.14,64.4
X$6158 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6159 r0 *1 87.14,64.4
X$6159 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6160 r0 *1 87.14,64.4
X$6160 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6161 r0 *1 31.14,16.8
X$6161 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6162 r0 *1 31.14,16.8
X$6162 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6163 r0 *1 31.14,16.8
X$6163 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6164 r0 *1 31.14,11.2
X$6164 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6165 r0 *1 31.14,11.2
X$6165 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6166 r0 *1 31.14,11.2
X$6166 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6167 r0 *1 87.14,11.2
X$6167 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6168 r0 *1 87.14,11.2
X$6168 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6169 r0 *1 87.14,11.2
X$6169 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6170 r0 *1 31.14,86.8
X$6170 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6171 r0 *1 31.14,86.8
X$6171 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6172 r0 *1 31.14,86.8
X$6172 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6173 r0 *1 87.14,86.8
X$6173 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6174 r0 *1 87.14,86.8
X$6174 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6175 r0 *1 87.14,86.8
X$6175 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6176 r0 *1 87.14,81.2
X$6176 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6177 r0 *1 87.14,81.2
X$6177 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6178 r0 *1 87.14,81.2
X$6178 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6179 r0 *1 31.14,53.2
X$6179 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6180 r0 *1 31.14,53.2
X$6180 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6181 r0 *1 31.14,53.2
X$6181 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6182 r0 *1 87.14,53.2
X$6182 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6183 r0 *1 87.14,53.2
X$6183 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6184 r0 *1 87.14,53.2
X$6184 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6185 r0 *1 31.14,78.4
X$6185 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6186 r0 *1 31.14,78.4
X$6186 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6187 r0 *1 31.14,78.4
X$6187 38 VIA_via4_5_960_2800_5_2_600_600
* cell instance $6188 r0 *1 31.14,78.4
X$6188 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6189 r0 *1 31.14,78.4
X$6189 38 VIA_via5_6_960_2800_5_2_600_600
* cell instance $6190 r0 *1 31.14,78.4
X$6190 38 VIA_via6_7_960_2800_4_1_600_600
* cell instance $6191 r0 *1 87.14,78.4
X$6191 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6192 r0 *1 87.14,78.4
X$6192 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6193 r0 *1 87.14,78.4
X$6193 38 VIA_via4_5_960_2800_5_2_600_600
* cell instance $6194 r0 *1 87.14,78.4
X$6194 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6195 r0 *1 87.14,78.4
X$6195 38 VIA_via5_6_960_2800_5_2_600_600
* cell instance $6196 r0 *1 87.14,78.4
X$6196 38 VIA_via6_7_960_2800_4_1_600_600
* cell instance $6197 r0 *1 31.14,95.2
X$6197 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6198 r0 *1 31.14,95.2
X$6198 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6199 r0 *1 31.14,95.2
X$6199 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6200 r0 *1 87.14,95.2
X$6200 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6201 r0 *1 87.14,95.2
X$6201 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6202 r0 *1 87.14,95.2
X$6202 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6203 r0 *1 31.14,89.6
X$6203 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6204 r0 *1 31.14,89.6
X$6204 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6205 r0 *1 31.14,89.6
X$6205 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6206 r0 *1 87.14,89.6
X$6206 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6207 r0 *1 87.14,89.6
X$6207 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6208 r0 *1 87.14,89.6
X$6208 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6209 r0 *1 31.14,61.6
X$6209 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6210 r0 *1 31.14,61.6
X$6210 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6211 r0 *1 31.14,61.6
X$6211 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6212 r0 *1 87.14,61.6
X$6212 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6213 r0 *1 87.14,61.6
X$6213 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6214 r0 *1 87.14,61.6
X$6214 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6215 r0 *1 31.14,42
X$6215 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6216 r0 *1 31.14,42
X$6216 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6217 r0 *1 31.14,42
X$6217 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6218 r0 *1 87.14,42
X$6218 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6219 r0 *1 87.14,42
X$6219 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6220 r0 *1 87.14,42
X$6220 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6221 r0 *1 31.14,25.2
X$6221 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6222 r0 *1 31.14,25.2
X$6222 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6223 r0 *1 31.14,25.2
X$6223 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6224 r0 *1 87.14,25.2
X$6224 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6225 r0 *1 87.14,25.2
X$6225 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6226 r0 *1 87.14,25.2
X$6226 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6227 r0 *1 31.14,14
X$6227 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6228 r0 *1 31.14,14
X$6228 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6229 r0 *1 31.14,14
X$6229 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6230 r0 *1 31.14,28
X$6230 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6231 r0 *1 31.14,28
X$6231 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6232 r0 *1 31.14,28
X$6232 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6233 r0 *1 87.14,28
X$6233 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6234 r0 *1 87.14,28
X$6234 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6235 r0 *1 87.14,28
X$6235 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6236 r0 *1 31.14,33.6
X$6236 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6237 r0 *1 31.14,33.6
X$6237 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6238 r0 *1 31.14,33.6
X$6238 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6239 r0 *1 87.14,33.6
X$6239 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6240 r0 *1 87.14,33.6
X$6240 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6241 r0 *1 87.14,33.6
X$6241 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6242 r0 *1 31.14,22.4
X$6242 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6243 r0 *1 31.14,22.4
X$6243 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6244 r0 *1 31.14,22.4
X$6244 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6245 r0 *1 87.14,22.4
X$6245 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6246 r0 *1 87.14,22.4
X$6246 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6247 r0 *1 87.14,22.4
X$6247 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6248 r0 *1 87.14,44.8
X$6248 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6249 r0 *1 87.14,44.8
X$6249 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6250 r0 *1 87.14,44.8
X$6250 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6251 r0 *1 31.14,36.4
X$6251 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6252 r0 *1 31.14,36.4
X$6252 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6253 r0 *1 31.14,36.4
X$6253 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6254 r0 *1 87.14,36.4
X$6254 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6255 r0 *1 87.14,36.4
X$6255 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6256 r0 *1 87.14,36.4
X$6256 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6257 r0 *1 31.14,30.8
X$6257 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6258 r0 *1 31.14,30.8
X$6258 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6259 r0 *1 31.14,30.8
X$6259 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6260 r0 *1 87.14,30.8
X$6260 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6261 r0 *1 87.14,30.8
X$6261 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6262 r0 *1 87.14,30.8
X$6262 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6263 r0 *1 87.14,72.8
X$6263 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6264 r0 *1 87.14,72.8
X$6264 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6265 r0 *1 87.14,72.8
X$6265 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6266 r0 *1 31.14,75.6
X$6266 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6267 r0 *1 31.14,75.6
X$6267 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6268 r0 *1 31.14,75.6
X$6268 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6269 r0 *1 87.14,75.6
X$6269 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6270 r0 *1 87.14,75.6
X$6270 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6271 r0 *1 87.14,75.6
X$6271 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6272 r0 *1 31.14,64.4
X$6272 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6273 r0 *1 31.14,64.4
X$6273 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6274 r0 *1 31.14,64.4
X$6274 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6275 r0 *1 31.14,56
X$6275 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6276 r0 *1 31.14,56
X$6276 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6277 r0 *1 31.14,56
X$6277 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6278 r0 *1 87.14,56
X$6278 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6279 r0 *1 87.14,56
X$6279 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6280 r0 *1 87.14,56
X$6280 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6281 r0 *1 31.14,58.8
X$6281 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6282 r0 *1 31.14,58.8
X$6282 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6283 r0 *1 31.14,58.8
X$6283 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6284 r0 *1 87.14,58.8
X$6284 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6285 r0 *1 87.14,58.8
X$6285 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6286 r0 *1 87.14,58.8
X$6286 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6287 r0 *1 31.14,72.8
X$6287 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6288 r0 *1 31.14,72.8
X$6288 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6289 r0 *1 31.14,72.8
X$6289 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6290 r0 *1 87.14,16.8
X$6290 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6291 r0 *1 87.14,16.8
X$6291 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6292 r0 *1 87.14,16.8
X$6292 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6293 r0 *1 31.14,70
X$6293 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6294 r0 *1 31.14,70
X$6294 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6295 r0 *1 31.14,70
X$6295 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6296 r0 *1 87.14,70
X$6296 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6297 r0 *1 87.14,70
X$6297 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6298 r0 *1 87.14,70
X$6298 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6299 r0 *1 31.14,19.6
X$6299 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6300 r0 *1 31.14,19.6
X$6300 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6301 r0 *1 31.14,19.6
X$6301 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6302 r0 *1 87.14,19.6
X$6302 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6303 r0 *1 87.14,19.6
X$6303 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6304 r0 *1 87.14,19.6
X$6304 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6305 r0 *1 31.14,2.8
X$6305 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6306 r0 *1 31.14,2.8
X$6306 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6307 r0 *1 31.14,2.8
X$6307 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6308 r0 *1 31.14,8.4
X$6308 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6309 r0 *1 31.14,8.4
X$6309 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6310 r0 *1 31.14,8.4
X$6310 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6311 r0 *1 87.14,8.4
X$6311 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6312 r0 *1 87.14,8.4
X$6312 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6313 r0 *1 87.14,8.4
X$6313 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6314 r0 *1 87.14,2.8
X$6314 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6315 r0 *1 87.14,2.8
X$6315 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6316 r0 *1 87.14,2.8
X$6316 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6317 r0 *1 31.14,5.6
X$6317 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6318 r0 *1 31.14,5.6
X$6318 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6319 r0 *1 31.14,5.6
X$6319 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6320 r0 *1 87.14,5.6
X$6320 38 VIA_via1_2_960_340_1_3_300_300
* cell instance $6321 r0 *1 87.14,5.6
X$6321 38 VIA_via2_3_960_340_1_3_320_320
* cell instance $6322 r0 *1 87.14,5.6
X$6322 38 VIA_via3_4_960_340_1_3_320_320
* cell instance $6323 r0 *1 26.125,3.01
X$6323 39 VIA_via1_7
* cell instance $6324 r0 *1 26.125,3.01
X$6324 39 VIA_via2_5
* cell instance $6325 r0 *1 25.365,3.01
X$6325 39 VIA_via2_5
* cell instance $6326 r0 *1 25.365,2.03
X$6326 39 VIA_via1_4
* cell instance $6327 r0 *1 35.435,4.97
X$6327 40 VIA_via1_7
* cell instance $6328 r0 *1 35.435,4.97
X$6328 40 VIA_via2_5
* cell instance $6329 r0 *1 12.635,4.97
X$6329 40 VIA_via1_7
* cell instance $6330 r0 *1 12.065,7.56
X$6330 40 VIA_via1_7
* cell instance $6331 r0 *1 51.205,4.55
X$6331 40 VIA_via2_5
* cell instance $6332 r0 *1 54.055,4.55
X$6332 40 VIA_via2_5
* cell instance $6333 r0 *1 24.415,4.27
X$6333 40 VIA_via2_5
* cell instance $6334 r0 *1 21.755,4.27
X$6334 40 VIA_via2_5
* cell instance $6335 r0 *1 45.505,4.55
X$6335 40 VIA_via2_5
* cell instance $6336 r0 *1 39.995,5.25
X$6336 40 VIA_via2_5
* cell instance $6337 r0 *1 12.635,4.27
X$6337 40 VIA_via2_5
* cell instance $6338 r0 *1 13.585,4.27
X$6338 40 VIA_via2_5
* cell instance $6339 r0 *1 35.435,5.25
X$6339 40 VIA_via2_5
* cell instance $6340 r0 *1 27.455,4.27
X$6340 40 VIA_via2_5
* cell instance $6341 r0 *1 27.455,4.97
X$6341 40 VIA_via2_5
* cell instance $6342 r0 *1 13.585,3.57
X$6342 40 VIA_via1_4
* cell instance $6343 r0 *1 21.755,4.83
X$6343 40 VIA_via1_4
* cell instance $6344 r0 *1 24.415,6.37
X$6344 40 VIA_via1_4
* cell instance $6345 r0 *1 27.265,3.57
X$6345 40 VIA_via1_4
* cell instance $6346 r0 *1 45.505,4.83
X$6346 40 VIA_via1_4
* cell instance $6347 r0 *1 39.995,4.83
X$6347 40 VIA_via1_4
* cell instance $6348 r0 *1 39.995,4.69
X$6348 40 VIA_via2_5
* cell instance $6349 r0 *1 54.055,3.85
X$6349 40 VIA_via1_4
* cell instance $6350 r0 *1 51.205,4.83
X$6350 40 VIA_via1_4
* cell instance $6351 r0 *1 16.625,4.41
X$6351 41 VIA_via1_7
* cell instance $6352 r0 *1 16.435,3.57
X$6352 41 VIA_via1_4
* cell instance $6353 r0 *1 29.165,6.23
X$6353 42 VIA_via1_7
* cell instance $6354 r0 *1 29.165,6.23
X$6354 42 VIA_via2_5
* cell instance $6355 r0 *1 10.925,6.23
X$6355 42 VIA_via1_7
* cell instance $6356 r0 *1 10.925,6.23
X$6356 42 VIA_via2_5
* cell instance $6357 r0 *1 18.715,6.23
X$6357 42 VIA_via1_7
* cell instance $6358 r0 *1 10.735,4.97
X$6358 42 VIA_via1_7
* cell instance $6359 r0 *1 18.905,4.55
X$6359 42 VIA_via2_5
* cell instance $6360 r0 *1 15.485,6.23
X$6360 42 VIA_via2_5
* cell instance $6361 r0 *1 15.485,4.55
X$6361 42 VIA_via2_5
* cell instance $6362 r0 *1 39.235,6.65
X$6362 42 VIA_via2_5
* cell instance $6363 r0 *1 32.585,6.79
X$6363 42 VIA_via2_5
* cell instance $6364 r0 *1 29.545,6.37
X$6364 42 VIA_via2_5
* cell instance $6365 r0 *1 29.165,4.41
X$6365 42 VIA_via2_5
* cell instance $6366 r0 *1 25.365,4.41
X$6366 42 VIA_via2_5
* cell instance $6367 r0 *1 29.545,6.79
X$6367 42 VIA_via2_5
* cell instance $6368 r0 *1 15.485,4.83
X$6368 42 VIA_via1_4
* cell instance $6369 r0 *1 49.115,6.37
X$6369 42 VIA_via1_4
* cell instance $6370 r0 *1 49.115,6.51
X$6370 42 VIA_via2_5
* cell instance $6371 r0 *1 32.585,6.37
X$6371 42 VIA_via1_4
* cell instance $6372 r0 *1 24.985,3.57
X$6372 42 VIA_via1_4
* cell instance $6373 r0 *1 39.235,6.37
X$6373 42 VIA_via1_4
* cell instance $6374 r0 *1 43.415,6.37
X$6374 42 VIA_via1_4
* cell instance $6375 r0 *1 43.415,6.51
X$6375 42 VIA_via2_5
* cell instance $6376 r0 *1 53.675,6.51
X$6376 42 VIA_via1_4
* cell instance $6377 r0 *1 53.675,6.51
X$6377 42 VIA_via2_5
* cell instance $6378 r0 *1 22.515,4.83
X$6378 43 VIA_via1_4
* cell instance $6379 r0 *1 22.895,3.85
X$6379 43 VIA_via1_4
* cell instance $6380 r0 *1 22.135,6.37
X$6380 43 VIA_via1_4
* cell instance $6381 r0 *1 41.515,6.37
X$6381 44 VIA_via1_4
* cell instance $6382 r0 *1 41.705,3.85
X$6382 44 VIA_via1_4
* cell instance $6383 r0 *1 40.755,4.83
X$6383 44 VIA_via1_4
* cell instance $6384 r0 *1 50.825,3.85
X$6384 45 VIA_via1_4
* cell instance $6385 r0 *1 51.965,4.83
X$6385 45 VIA_via1_4
* cell instance $6386 r0 *1 51.205,6.37
X$6386 45 VIA_via1_4
* cell instance $6387 r0 *1 57.285,6.37
X$6387 46 VIA_via1_4
* cell instance $6388 r0 *1 57.285,4.83
X$6388 46 VIA_via1_4
* cell instance $6389 r0 *1 57.665,3.85
X$6389 46 VIA_via1_4
* cell instance $6390 r0 *1 67.735,3.85
X$6390 47 VIA_via2_5
* cell instance $6391 r0 *1 65.455,3.85
X$6391 47 VIA_via2_5
* cell instance $6392 r0 *1 67.735,3.57
X$6392 47 VIA_via1_4
* cell instance $6393 r0 *1 65.455,4.83
X$6393 47 VIA_via1_4
* cell instance $6394 r0 *1 66.785,3.85
X$6394 47 VIA_via1_4
* cell instance $6395 r0 *1 66.785,3.85
X$6395 47 VIA_via2_5
* cell instance $6396 r0 *1 69.065,8.33
X$6396 48 VIA_via2_5
* cell instance $6397 r0 *1 63.745,8.33
X$6397 48 VIA_via2_5
* cell instance $6398 r0 *1 69.065,7.07
X$6398 48 VIA_via2_5
* cell instance $6399 r0 *1 67.925,7.07
X$6399 48 VIA_via2_5
* cell instance $6400 r0 *1 62.795,10.29
X$6400 48 VIA_via2_5
* cell instance $6401 r0 *1 66.975,8.33
X$6401 48 VIA_via2_5
* cell instance $6402 r0 *1 63.175,5.67
X$6402 48 VIA_via2_5
* cell instance $6403 r0 *1 63.745,5.67
X$6403 48 VIA_via2_5
* cell instance $6404 r0 *1 62.795,12.25
X$6404 48 VIA_via2_5
* cell instance $6405 r0 *1 64.125,12.25
X$6405 48 VIA_via2_5
* cell instance $6406 r0 *1 63.175,18.69
X$6406 48 VIA_via2_5
* cell instance $6407 r0 *1 63.745,18.69
X$6407 48 VIA_via2_5
* cell instance $6408 r0 *1 64.125,18.69
X$6408 48 VIA_via2_5
* cell instance $6409 r0 *1 63.555,22.89
X$6409 48 VIA_via2_5
* cell instance $6410 r0 *1 61.275,18.83
X$6410 48 VIA_via1_4
* cell instance $6411 r0 *1 61.275,18.69
X$6411 48 VIA_via2_5
* cell instance $6412 r0 *1 63.175,17.57
X$6412 48 VIA_via1_4
* cell instance $6413 r0 *1 64.125,13.23
X$6413 48 VIA_via1_4
* cell instance $6414 r0 *1 63.555,21.63
X$6414 48 VIA_via1_4
* cell instance $6415 r0 *1 61.845,23.17
X$6415 48 VIA_via1_4
* cell instance $6416 r0 *1 61.845,23.17
X$6416 48 VIA_via2_5
* cell instance $6417 r0 *1 67.735,4.55
X$6417 48 VIA_via1_4
* cell instance $6418 r0 *1 62.985,4.83
X$6418 48 VIA_via1_4
* cell instance $6419 r0 *1 69.065,7.63
X$6419 48 VIA_via1_4
* cell instance $6420 r0 *1 62.795,11.97
X$6420 48 VIA_via1_4
* cell instance $6421 r0 *1 63.745,10.43
X$6421 48 VIA_via1_4
* cell instance $6422 r0 *1 63.745,10.29
X$6422 48 VIA_via2_5
* cell instance $6423 r0 *1 66.975,9.17
X$6423 48 VIA_via1_4
* cell instance $6424 r0 *1 90.345,4.27
X$6424 49 VIA_via2_5
* cell instance $6425 r0 *1 87.495,4.27
X$6425 49 VIA_via2_5
* cell instance $6426 r0 *1 75.905,4.27
X$6426 49 VIA_via2_5
* cell instance $6427 r0 *1 80.275,4.27
X$6427 49 VIA_via2_5
* cell instance $6428 r0 *1 88.635,15.05
X$6428 49 VIA_via2_5
* cell instance $6429 r0 *1 87.495,15.05
X$6429 49 VIA_via2_5
* cell instance $6430 r0 *1 86.165,15.05
X$6430 49 VIA_via2_5
* cell instance $6431 r0 *1 69.825,4.27
X$6431 49 VIA_via2_5
* cell instance $6432 r0 *1 70.395,4.27
X$6432 49 VIA_via2_5
* cell instance $6433 r0 *1 88.635,16.03
X$6433 49 VIA_via1_4
* cell instance $6434 r0 *1 80.275,3.85
X$6434 49 VIA_via1_4
* cell instance $6435 r0 *1 87.495,6.37
X$6435 49 VIA_via1_4
* cell instance $6436 r0 *1 90.345,4.83
X$6436 49 VIA_via1_4
* cell instance $6437 r0 *1 75.905,4.83
X$6437 49 VIA_via1_4
* cell instance $6438 r0 *1 70.015,13.23
X$6438 49 VIA_via1_4
* cell instance $6439 r0 *1 70.395,3.57
X$6439 49 VIA_via1_4
* cell instance $6440 r0 *1 86.165,14.77
X$6440 49 VIA_via1_4
* cell instance $6441 r0 *1 77.805,3.57
X$6441 50 VIA_via2_5
* cell instance $6442 r0 *1 78.755,3.57
X$6442 50 VIA_via1_4
* cell instance $6443 r0 *1 78.755,3.57
X$6443 50 VIA_via2_5
* cell instance $6444 r0 *1 77.615,4.83
X$6444 50 VIA_via1_4
* cell instance $6445 r0 *1 77.805,3.85
X$6445 50 VIA_via1_4
* cell instance $6446 r0 *1 70.395,34.23
X$6446 51 VIA_via1_7
* cell instance $6447 r0 *1 70.395,34.23
X$6447 51 VIA_via2_5
* cell instance $6448 r0 *1 77.805,72.17
X$6448 51 VIA_via1_7
* cell instance $6449 r0 *1 64.125,72.17
X$6449 51 VIA_via1_7
* cell instance $6450 r0 *1 64.125,72.17
X$6450 51 VIA_via2_5
* cell instance $6451 r0 *1 64.215,72.17
X$6451 51 VIA_via3_2
* cell instance $6452 r0 *1 77.995,3.85
X$6452 51 VIA_via2_5
* cell instance $6453 r0 *1 77.995,21.07
X$6453 51 VIA_via2_5
* cell instance $6454 r0 *1 64.125,72.87
X$6454 51 VIA_via2_5
* cell instance $6455 r0 *1 68.305,3.85
X$6455 51 VIA_via2_5
* cell instance $6456 r0 *1 68.305,4.69
X$6456 51 VIA_via2_5
* cell instance $6457 r0 *1 67.545,50.19
X$6457 51 VIA_via2_5
* cell instance $6458 r0 *1 77.805,72.87
X$6458 51 VIA_via2_5
* cell instance $6459 r0 *1 71.345,42.49
X$6459 51 VIA_via2_5
* cell instance $6460 r0 *1 70.395,42.49
X$6460 51 VIA_via2_5
* cell instance $6461 r0 *1 67.925,46.13
X$6461 51 VIA_via2_5
* cell instance $6462 r0 *1 71.345,46.13
X$6462 51 VIA_via2_5
* cell instance $6463 r0 *1 76.095,46.13
X$6463 51 VIA_via2_5
* cell instance $6464 r0 *1 76.095,45.57
X$6464 51 VIA_via1_4
* cell instance $6465 r0 *1 67.735,45.57
X$6465 51 VIA_via1_4
* cell instance $6466 r0 *1 77.995,3.57
X$6466 51 VIA_via1_4
* cell instance $6467 r0 *1 77.995,20.37
X$6467 51 VIA_via1_4
* cell instance $6468 r0 *1 62.605,50.05
X$6468 51 VIA_via1_4
* cell instance $6469 r0 *1 62.605,50.05
X$6469 51 VIA_via2_5
* cell instance $6470 r0 *1 62.795,4.83
X$6470 51 VIA_via1_4
* cell instance $6471 r0 *1 62.795,4.69
X$6471 51 VIA_via2_5
* cell instance $6472 r0 *1 68.305,3.57
X$6472 51 VIA_via1_4
* cell instance $6473 r0 *1 72.865,58.03
X$6473 51 VIA_via1_4
* cell instance $6474 r0 *1 72.865,57.89
X$6474 51 VIA_via2_5
* cell instance $6475 r0 *1 64.215,50.19
X$6475 51 VIA_via3_2
* cell instance $6476 r0 *1 64.215,57.89
X$6476 51 VIA_via3_2
* cell instance $6477 r0 *1 73.455,21.07
X$6477 51 VIA_via3_2
* cell instance $6478 r0 *1 73.455,34.23
X$6478 51 VIA_via3_2
* cell instance $6479 r0 *1 78.215,3.85
X$6479 51 VIA_via3_2
* cell instance $6480 r0 *1 78.215,21.07
X$6480 51 VIA_via3_2
* cell instance $6481 r0 *1 85.975,3.99
X$6481 52 VIA_via1_7
* cell instance $6482 r0 *1 77.615,17.29
X$6482 52 VIA_via2_5
* cell instance $6483 r0 *1 76.665,17.29
X$6483 52 VIA_via2_5
* cell instance $6484 r0 *1 78.185,17.29
X$6484 52 VIA_via2_5
* cell instance $6485 r0 *1 77.995,4.69
X$6485 52 VIA_via2_5
* cell instance $6486 r0 *1 85.975,4.41
X$6486 52 VIA_via2_5
* cell instance $6487 r0 *1 80.655,4.41
X$6487 52 VIA_via2_5
* cell instance $6488 r0 *1 86.545,11.69
X$6488 52 VIA_via2_5
* cell instance $6489 r0 *1 85.025,4.41
X$6489 52 VIA_via2_5
* cell instance $6490 r0 *1 85.025,11.55
X$6490 52 VIA_via2_5
* cell instance $6491 r0 *1 75.145,21.35
X$6491 52 VIA_via2_5
* cell instance $6492 r0 *1 73.435,17.29
X$6492 52 VIA_via2_5
* cell instance $6493 r0 *1 73.435,21.35
X$6493 52 VIA_via2_5
* cell instance $6494 r0 *1 78.185,7.63
X$6494 52 VIA_via1_4
* cell instance $6495 r0 *1 80.655,4.83
X$6495 52 VIA_via1_4
* cell instance $6496 r0 *1 80.655,4.69
X$6496 52 VIA_via2_5
* cell instance $6497 r0 *1 86.545,11.97
X$6497 52 VIA_via1_4
* cell instance $6498 r0 *1 78.185,3.57
X$6498 52 VIA_via1_4
* cell instance $6499 r0 *1 75.145,21.63
X$6499 52 VIA_via1_4
* cell instance $6500 r0 *1 85.025,10.43
X$6500 52 VIA_via1_4
* cell instance $6501 r0 *1 76.665,17.57
X$6501 52 VIA_via1_4
* cell instance $6502 r0 *1 77.615,17.57
X$6502 52 VIA_via1_4
* cell instance $6503 r0 *1 73.055,23.17
X$6503 52 VIA_via1_4
* cell instance $6504 r0 *1 73.435,18.83
X$6504 52 VIA_via1_4
* cell instance $6505 r0 *1 92.815,3.71
X$6505 53 VIA_via2_5
* cell instance $6506 r0 *1 91.675,3.71
X$6506 53 VIA_via2_5
* cell instance $6507 r0 *1 92.055,10.85
X$6507 53 VIA_via2_5
* cell instance $6508 r0 *1 92.245,8.47
X$6508 53 VIA_via2_5
* cell instance $6509 r0 *1 92.435,10.85
X$6509 53 VIA_via2_5
* cell instance $6510 r0 *1 92.625,8.47
X$6510 53 VIA_via2_5
* cell instance $6511 r0 *1 80.085,3.71
X$6511 53 VIA_via2_5
* cell instance $6512 r0 *1 91.675,9.03
X$6512 53 VIA_via2_5
* cell instance $6513 r0 *1 92.055,13.23
X$6513 53 VIA_via1_4
* cell instance $6514 r0 *1 92.435,10.43
X$6514 53 VIA_via1_4
* cell instance $6515 r0 *1 92.245,9.17
X$6515 53 VIA_via1_4
* cell instance $6516 r0 *1 92.245,9.03
X$6516 53 VIA_via2_5
* cell instance $6517 r0 *1 85.595,3.57
X$6517 53 VIA_via1_4
* cell instance $6518 r0 *1 85.595,3.71
X$6518 53 VIA_via2_5
* cell instance $6519 r0 *1 91.675,6.37
X$6519 53 VIA_via1_4
* cell instance $6520 r0 *1 92.815,2.45
X$6520 53 VIA_via1_4
* cell instance $6521 r0 *1 79.895,2.03
X$6521 53 VIA_via1_4
* cell instance $6522 r0 *1 80.085,13.23
X$6522 53 VIA_via1_4
* cell instance $6523 r0 *1 89.585,6.37
X$6523 54 VIA_via2_5
* cell instance $6524 r0 *1 88.825,6.37
X$6524 54 VIA_via1_4
* cell instance $6525 r0 *1 88.825,6.37
X$6525 54 VIA_via2_5
* cell instance $6526 r0 *1 88.065,6.37
X$6526 54 VIA_via1_4
* cell instance $6527 r0 *1 88.065,6.37
X$6527 54 VIA_via2_5
* cell instance $6528 r0 *1 89.965,4.55
X$6528 54 VIA_via1_4
* cell instance $6529 r0 *1 11.875,4.41
X$6529 55 VIA_via1_7
* cell instance $6530 r0 *1 11.875,3.57
X$6530 55 VIA_via2_5
* cell instance $6531 r0 *1 10.735,3.57
X$6531 55 VIA_via1_4
* cell instance $6532 r0 *1 10.735,3.57
X$6532 55 VIA_via2_5
* cell instance $6533 r0 *1 15.295,3.71
X$6533 56 VIA_via2_5
* cell instance $6534 r0 *1 17.955,3.71
X$6534 56 VIA_via2_5
* cell instance $6535 r0 *1 15.295,2.03
X$6535 56 VIA_via1_4
* cell instance $6536 r0 *1 17.955,4.83
X$6536 56 VIA_via1_4
* cell instance $6537 r0 *1 14.345,3.57
X$6537 56 VIA_via1_4
* cell instance $6538 r0 *1 14.345,3.71
X$6538 56 VIA_via2_5
* cell instance $6539 r0 *1 22.895,4.41
X$6539 57 VIA_via1_7
* cell instance $6540 r0 *1 22.895,4.41
X$6540 57 VIA_via2_5
* cell instance $6541 r0 *1 20.615,4.41
X$6541 57 VIA_via2_5
* cell instance $6542 r0 *1 20.615,3.57
X$6542 57 VIA_via1_4
* cell instance $6543 r0 *1 28.405,3.57
X$6543 58 VIA_via1_4
* cell instance $6544 r0 *1 29.355,3.57
X$6544 58 VIA_via1_4
* cell instance $6545 r0 *1 31.445,6.37
X$6545 59 VIA_via1_4
* cell instance $6546 r0 *1 28.025,3.57
X$6546 59 VIA_via1_4
* cell instance $6547 r0 *1 28.025,3.57
X$6547 59 VIA_via2_5
* cell instance $6548 r0 *1 31.635,3.57
X$6548 59 VIA_via1_4
* cell instance $6549 r0 *1 31.635,3.57
X$6549 59 VIA_via2_5
* cell instance $6550 r0 *1 75.525,3.57
X$6550 60 VIA_via1_4
* cell instance $6551 r0 *1 75.525,3.71
X$6551 60 VIA_via2_5
* cell instance $6552 r0 *1 79.135,3.71
X$6552 60 VIA_via1_4
* cell instance $6553 r0 *1 79.135,3.71
X$6553 60 VIA_via2_5
* cell instance $6554 r0 *1 41.135,4.41
X$6554 61 VIA_via1_7
* cell instance $6555 r0 *1 41.135,4.41
X$6555 61 VIA_via2_5
* cell instance $6556 r0 *1 39.425,4.41
X$6556 61 VIA_via2_5
* cell instance $6557 r0 *1 39.425,3.57
X$6557 61 VIA_via1_4
* cell instance $6558 r0 *1 46.645,4.41
X$6558 62 VIA_via1_7
* cell instance $6559 r0 *1 46.645,4.41
X$6559 62 VIA_via2_5
* cell instance $6560 r0 *1 43.795,4.41
X$6560 62 VIA_via2_5
* cell instance $6561 r0 *1 43.795,3.57
X$6561 62 VIA_via1_4
* cell instance $6562 r0 *1 71.345,3.57
X$6562 63 VIA_via1_4
* cell instance $6563 r0 *1 71.345,3.57
X$6563 63 VIA_via2_5
* cell instance $6564 r0 *1 72.295,3.57
X$6564 63 VIA_via1_4
* cell instance $6565 r0 *1 72.295,3.57
X$6565 63 VIA_via2_5
* cell instance $6566 r0 *1 52.345,4.41
X$6566 64 VIA_via1_7
* cell instance $6567 r0 *1 52.345,4.41
X$6567 64 VIA_via2_5
* cell instance $6568 r0 *1 48.545,4.41
X$6568 64 VIA_via2_5
* cell instance $6569 r0 *1 48.545,3.57
X$6569 64 VIA_via1_4
* cell instance $6570 r0 *1 68.115,3.71
X$6570 65 VIA_via1_4
* cell instance $6571 r0 *1 68.115,3.71
X$6571 65 VIA_via2_5
* cell instance $6572 r0 *1 64.505,3.57
X$6572 65 VIA_via1_4
* cell instance $6573 r0 *1 64.505,3.71
X$6573 65 VIA_via2_5
* cell instance $6574 r0 *1 50.065,10.43
X$6574 66 VIA_via2_5
* cell instance $6575 r0 *1 52.155,6.65
X$6575 66 VIA_via2_5
* cell instance $6576 r0 *1 49.305,6.65
X$6576 66 VIA_via2_5
* cell instance $6577 r0 *1 49.685,6.65
X$6577 66 VIA_via2_5
* cell instance $6578 r0 *1 51.395,4.13
X$6578 66 VIA_via2_5
* cell instance $6579 r0 *1 52.155,4.13
X$6579 66 VIA_via2_5
* cell instance $6580 r0 *1 52.345,4.13
X$6580 66 VIA_via2_5
* cell instance $6581 r0 *1 49.685,28.63
X$6581 66 VIA_via2_5
* cell instance $6582 r0 *1 49.305,6.37
X$6582 66 VIA_via1_4
* cell instance $6583 r0 *1 49.685,9.17
X$6583 66 VIA_via1_4
* cell instance $6584 r0 *1 51.395,10.43
X$6584 66 VIA_via1_4
* cell instance $6585 r0 *1 51.395,10.43
X$6585 66 VIA_via2_5
* cell instance $6586 r0 *1 49.495,14.77
X$6586 66 VIA_via1_4
* cell instance $6587 r0 *1 52.725,28.77
X$6587 66 VIA_via1_4
* cell instance $6588 r0 *1 52.725,28.63
X$6588 66 VIA_via2_5
* cell instance $6589 r0 *1 50.065,30.03
X$6589 66 VIA_via1_4
* cell instance $6590 r0 *1 52.345,2.45
X$6590 66 VIA_via1_4
* cell instance $6591 r0 *1 51.395,4.83
X$6591 66 VIA_via1_4
* cell instance $6592 r0 *1 57.665,4.41
X$6592 67 VIA_via1_7
* cell instance $6593 r0 *1 57.665,4.41
X$6593 67 VIA_via2_5
* cell instance $6594 r0 *1 55.385,4.41
X$6594 67 VIA_via2_5
* cell instance $6595 r0 *1 55.385,3.57
X$6595 67 VIA_via1_4
* cell instance $6596 r0 *1 66.025,57.75
X$6596 68 VIA_via1_7
* cell instance $6597 r0 *1 66.025,57.75
X$6597 68 VIA_via2_5
* cell instance $6598 r0 *1 56.525,4.97
X$6598 68 VIA_via1_7
* cell instance $6599 r0 *1 56.525,5.11
X$6599 68 VIA_via2_5
* cell instance $6600 r0 *1 59.565,6.23
X$6600 68 VIA_via1_7
* cell instance $6601 r0 *1 60.135,6.65
X$6601 68 VIA_via2_5
* cell instance $6602 r0 *1 55.575,57.75
X$6602 68 VIA_via2_5
* cell instance $6603 r0 *1 59.565,5.11
X$6603 68 VIA_via2_5
* cell instance $6604 r0 *1 59.565,5.95
X$6604 68 VIA_via2_5
* cell instance $6605 r0 *1 56.905,5.11
X$6605 68 VIA_via2_5
* cell instance $6606 r0 *1 56.905,3.57
X$6606 68 VIA_via2_5
* cell instance $6607 r0 *1 60.135,5.95
X$6607 68 VIA_via2_5
* cell instance $6608 r0 *1 66.025,6.37
X$6608 68 VIA_via2_5
* cell instance $6609 r0 *1 66.025,6.65
X$6609 68 VIA_via2_5
* cell instance $6610 r0 *1 53.675,3.57
X$6610 68 VIA_via1_4
* cell instance $6611 r0 *1 53.675,3.57
X$6611 68 VIA_via2_5
* cell instance $6612 r0 *1 55.575,58.03
X$6612 68 VIA_via1_4
* cell instance $6613 r0 *1 66.025,4.83
X$6613 68 VIA_via1_4
* cell instance $6614 r0 *1 56.655,57.75
X$6614 68 VIA_via4_0
* cell instance $6615 r0 *1 56.655,57.75
X$6615 68 VIA_via3_2
* cell instance $6616 r0 *1 66.175,57.75
X$6616 68 VIA_via3_2
* cell instance $6617 r0 *1 66.175,57.75
X$6617 68 VIA_via4_0
* cell instance $6618 r0 *1 66.175,6.37
X$6618 68 VIA_via3_2
* cell instance $6619 r0 *1 13.015,4.83
X$6619 69 VIA_via2_5
* cell instance $6620 r0 *1 14.155,4.83
X$6620 69 VIA_via1_4
* cell instance $6621 r0 *1 14.155,4.69
X$6621 69 VIA_via2_5
* cell instance $6622 r0 *1 13.015,3.85
X$6622 69 VIA_via1_4
* cell instance $6623 r0 *1 11.495,4.83
X$6623 69 VIA_via1_4
* cell instance $6624 r0 *1 11.495,4.83
X$6624 69 VIA_via2_5
* cell instance $6625 r0 *1 11.875,9.03
X$6625 70 VIA_via1_7
* cell instance $6626 r0 *1 13.965,4.97
X$6626 70 VIA_via1_7
* cell instance $6627 r0 *1 13.965,4.97
X$6627 70 VIA_via2_5
* cell instance $6628 r0 *1 17.195,4.97
X$6628 70 VIA_via1_7
* cell instance $6629 r0 *1 17.195,4.97
X$6629 70 VIA_via2_5
* cell instance $6630 r0 *1 8.075,58.31
X$6630 70 VIA_via2_5
* cell instance $6631 r0 *1 6.745,58.31
X$6631 70 VIA_via2_5
* cell instance $6632 r0 *1 9.025,56.07
X$6632 70 VIA_via2_5
* cell instance $6633 r0 *1 8.075,56.07
X$6633 70 VIA_via2_5
* cell instance $6634 r0 *1 5.225,73.57
X$6634 70 VIA_via2_5
* cell instance $6635 r0 *1 7.505,73.57
X$6635 70 VIA_via2_5
* cell instance $6636 r0 *1 21.375,4.97
X$6636 70 VIA_via2_5
* cell instance $6637 r0 *1 13.965,8.61
X$6637 70 VIA_via2_5
* cell instance $6638 r0 *1 9.215,45.43
X$6638 70 VIA_via2_5
* cell instance $6639 r0 *1 11.875,8.61
X$6639 70 VIA_via2_5
* cell instance $6640 r0 *1 5.605,58.31
X$6640 70 VIA_via2_5
* cell instance $6641 r0 *1 21.375,6.37
X$6641 70 VIA_via1_4
* cell instance $6642 r0 *1 21.375,6.51
X$6642 70 VIA_via2_5
* cell instance $6643 r0 *1 30.685,6.37
X$6643 70 VIA_via1_4
* cell instance $6644 r0 *1 30.685,6.51
X$6644 70 VIA_via2_5
* cell instance $6645 r0 *1 33.915,6.37
X$6645 70 VIA_via1_4
* cell instance $6646 r0 *1 33.915,6.23
X$6646 70 VIA_via2_5
* cell instance $6647 r0 *1 25.745,6.37
X$6647 70 VIA_via1_4
* cell instance $6648 r0 *1 25.745,6.51
X$6648 70 VIA_via2_5
* cell instance $6649 r0 *1 32.395,45.15
X$6649 70 VIA_via1_4
* cell instance $6650 r0 *1 32.395,45.15
X$6650 70 VIA_via2_5
* cell instance $6651 r0 *1 7.125,62.37
X$6651 70 VIA_via1_4
* cell instance $6652 r0 *1 5.605,56.77
X$6652 70 VIA_via1_4
* cell instance $6653 r0 *1 5.225,74.83
X$6653 70 VIA_via1_4
* cell instance $6654 r0 *1 32.575,45.15
X$6654 70 VIA_via3_2
* cell instance $6655 r0 *1 32.575,6.37
X$6655 70 VIA_via3_2
* cell instance $6656 r0 *1 18.715,4.83
X$6656 71 VIA_via2_5
* cell instance $6657 r0 *1 16.245,4.83
X$6657 71 VIA_via1_4
* cell instance $6658 r0 *1 16.245,4.83
X$6658 71 VIA_via2_5
* cell instance $6659 r0 *1 18.715,3.85
X$6659 71 VIA_via1_4
* cell instance $6660 r0 *1 17.385,4.83
X$6660 71 VIA_via1_4
* cell instance $6661 r0 *1 17.385,4.83
X$6661 71 VIA_via2_5
* cell instance $6662 r0 *1 25.555,5.81
X$6662 72 VIA_via1_7
* cell instance $6663 r0 *1 25.175,4.83
X$6663 72 VIA_via1_4
* cell instance $6664 r0 *1 32.965,14.77
X$6664 73 VIA_via2_5
* cell instance $6665 r0 *1 33.155,14.77
X$6665 73 VIA_via2_5
* cell instance $6666 r0 *1 31.065,10.99
X$6666 73 VIA_via2_5
* cell instance $6667 r0 *1 32.585,10.99
X$6667 73 VIA_via2_5
* cell instance $6668 r0 *1 31.065,10.43
X$6668 73 VIA_via1_4
* cell instance $6669 r0 *1 30.495,9.17
X$6669 73 VIA_via1_4
* cell instance $6670 r0 *1 32.585,11.55
X$6670 73 VIA_via1_4
* cell instance $6671 r0 *1 32.965,12.39
X$6671 73 VIA_via1_7
* cell instance $6672 r0 *1 33.155,11.97
X$6672 73 VIA_via1_4
* cell instance $6673 r0 *1 30.495,4.83
X$6673 73 VIA_via1_4
* cell instance $6674 r0 *1 30.115,3.57
X$6674 73 VIA_via1_4
* cell instance $6675 r0 *1 33.155,16.03
X$6675 73 VIA_via1_4
* cell instance $6676 r0 *1 36.575,14.77
X$6676 73 VIA_via1_4
* cell instance $6677 r0 *1 36.575,14.77
X$6677 73 VIA_via2_5
* cell instance $6678 r0 *1 28.215,14.77
X$6678 73 VIA_via1_4
* cell instance $6679 r0 *1 28.215,14.77
X$6679 73 VIA_via2_5
* cell instance $6680 r0 *1 38.285,4.55
X$6680 74 VIA_via2_5
* cell instance $6681 r0 *1 38.475,10.43
X$6681 74 VIA_via2_5
* cell instance $6682 r0 *1 40.185,4.55
X$6682 74 VIA_via2_5
* cell instance $6683 r0 *1 33.725,10.43
X$6683 74 VIA_via2_5
* cell instance $6684 r0 *1 33.725,9.17
X$6684 74 VIA_via1_4
* cell instance $6685 r0 *1 35.435,10.43
X$6685 74 VIA_via1_4
* cell instance $6686 r0 *1 35.435,10.43
X$6686 74 VIA_via2_5
* cell instance $6687 r0 *1 33.725,4.83
X$6687 74 VIA_via1_4
* cell instance $6688 r0 *1 37.525,6.37
X$6688 74 VIA_via1_4
* cell instance $6689 r0 *1 38.475,9.17
X$6689 74 VIA_via1_4
* cell instance $6690 r0 *1 37.715,7.35
X$6690 74 VIA_via1_4
* cell instance $6691 r0 *1 38.095,8.05
X$6691 74 VIA_via1_4
* cell instance $6692 r0 *1 40.185,10.43
X$6692 74 VIA_via1_4
* cell instance $6693 r0 *1 40.185,10.43
X$6693 74 VIA_via2_5
* cell instance $6694 r0 *1 40.185,3.57
X$6694 74 VIA_via1_4
* cell instance $6695 r0 *1 38.285,4.83
X$6695 74 VIA_via1_4
* cell instance $6696 r0 *1 42.94,10.36
X$6696 75 VIA_via1_7
* cell instance $6697 r0 *1 42.845,30.03
X$6697 75 VIA_via2_5
* cell instance $6698 r0 *1 43.605,12.11
X$6698 75 VIA_via2_5
* cell instance $6699 r0 *1 43.605,10.57
X$6699 75 VIA_via2_5
* cell instance $6700 r0 *1 43.035,10.57
X$6700 75 VIA_via2_5
* cell instance $6701 r0 *1 45.695,10.57
X$6701 75 VIA_via2_5
* cell instance $6702 r0 *1 43.035,24.43
X$6702 75 VIA_via1_4
* cell instance $6703 r0 *1 43.605,6.37
X$6703 75 VIA_via1_4
* cell instance $6704 r0 *1 44.555,11.97
X$6704 75 VIA_via1_4
* cell instance $6705 r0 *1 44.555,12.11
X$6705 75 VIA_via2_5
* cell instance $6706 r0 *1 45.695,2.45
X$6706 75 VIA_via1_4
* cell instance $6707 r0 *1 45.695,4.83
X$6707 75 VIA_via1_4
* cell instance $6708 r0 *1 44.935,30.03
X$6708 75 VIA_via1_4
* cell instance $6709 r0 *1 44.935,30.03
X$6709 75 VIA_via2_5
* cell instance $6710 r0 *1 42.845,27.23
X$6710 75 VIA_via1_4
* cell instance $6711 r0 *1 57.285,10.29
X$6711 76 VIA_via2_5
* cell instance $6712 r0 *1 59.565,10.43
X$6712 76 VIA_via2_5
* cell instance $6713 r0 *1 49.495,6.23
X$6713 76 VIA_via2_5
* cell instance $6714 r0 *1 51.395,6.23
X$6714 76 VIA_via2_5
* cell instance $6715 r0 *1 56.335,9.17
X$6715 76 VIA_via2_5
* cell instance $6716 r0 *1 56.145,6.23
X$6716 76 VIA_via2_5
* cell instance $6717 r0 *1 59.755,10.43
X$6717 76 VIA_via2_5
* cell instance $6718 r0 *1 56.145,4.83
X$6718 76 VIA_via2_5
* cell instance $6719 r0 *1 58.615,10.43
X$6719 76 VIA_via1_4
* cell instance $6720 r0 *1 58.615,10.43
X$6720 76 VIA_via2_5
* cell instance $6721 r0 *1 59.755,11.97
X$6721 76 VIA_via1_4
* cell instance $6722 r0 *1 54.815,4.83
X$6722 76 VIA_via1_4
* cell instance $6723 r0 *1 54.815,4.83
X$6723 76 VIA_via2_5
* cell instance $6724 r0 *1 49.495,4.83
X$6724 76 VIA_via1_4
* cell instance $6725 r0 *1 57.285,9.17
X$6725 76 VIA_via1_4
* cell instance $6726 r0 *1 57.285,9.17
X$6726 76 VIA_via2_5
* cell instance $6727 r0 *1 56.335,8.05
X$6727 76 VIA_via1_4
* cell instance $6728 r0 *1 51.395,7.63
X$6728 76 VIA_via1_4
* cell instance $6729 r0 *1 56.145,3.57
X$6729 76 VIA_via1_4
* cell instance $6730 r0 *1 59.565,4.83
X$6730 76 VIA_via1_4
* cell instance $6731 r0 *1 72.105,2.59
X$6731 77 VIA_via1_7
* cell instance $6732 r0 *1 69.635,10.29
X$6732 77 VIA_via2_5
* cell instance $6733 r0 *1 69.635,6.23
X$6733 77 VIA_via2_5
* cell instance $6734 r0 *1 67.355,5.53
X$6734 77 VIA_via2_5
* cell instance $6735 r0 *1 72.105,6.23
X$6735 77 VIA_via2_5
* cell instance $6736 r0 *1 69.635,5.53
X$6736 77 VIA_via2_5
* cell instance $6737 r0 *1 73.435,6.23
X$6737 77 VIA_via2_5
* cell instance $6738 r0 *1 74.385,10.43
X$6738 77 VIA_via1_4
* cell instance $6739 r0 *1 74.385,10.29
X$6739 77 VIA_via2_5
* cell instance $6740 r0 *1 73.435,4.83
X$6740 77 VIA_via1_4
* cell instance $6741 r0 *1 70.395,6.37
X$6741 77 VIA_via1_4
* cell instance $6742 r0 *1 70.395,6.23
X$6742 77 VIA_via2_5
* cell instance $6743 r0 *1 68.305,10.43
X$6743 77 VIA_via1_4
* cell instance $6744 r0 *1 68.305,10.29
X$6744 77 VIA_via2_5
* cell instance $6745 r0 *1 73.055,10.43
X$6745 77 VIA_via1_4
* cell instance $6746 r0 *1 73.055,10.29
X$6746 77 VIA_via2_5
* cell instance $6747 r0 *1 67.165,3.57
X$6747 77 VIA_via1_4
* cell instance $6748 r0 *1 67.355,4.83
X$6748 77 VIA_via1_4
* cell instance $6749 r0 *1 76.285,4.41
X$6749 78 VIA_via1_7
* cell instance $6750 r0 *1 67.925,12.95
X$6750 78 VIA_via2_5
* cell instance $6751 r0 *1 67.545,12.95
X$6751 78 VIA_via2_5
* cell instance $6752 r0 *1 67.545,15.75
X$6752 78 VIA_via2_5
* cell instance $6753 r0 *1 76.285,4.69
X$6753 78 VIA_via2_5
* cell instance $6754 r0 *1 82.175,4.55
X$6754 78 VIA_via2_5
* cell instance $6755 r0 *1 83.125,4.55
X$6755 78 VIA_via2_5
* cell instance $6756 r0 *1 82.935,11.83
X$6756 78 VIA_via2_5
* cell instance $6757 r0 *1 68.495,4.83
X$6757 78 VIA_via2_5
* cell instance $6758 r0 *1 67.735,4.83
X$6758 78 VIA_via2_5
* cell instance $6759 r0 *1 67.355,21.91
X$6759 78 VIA_via2_5
* cell instance $6760 r0 *1 68.305,21.91
X$6760 78 VIA_via2_5
* cell instance $6761 r0 *1 69.825,21.91
X$6761 78 VIA_via2_5
* cell instance $6762 r0 *1 68.115,15.75
X$6762 78 VIA_via2_5
* cell instance $6763 r0 *1 68.495,16.87
X$6763 78 VIA_via2_5
* cell instance $6764 r0 *1 68.115,16.73
X$6764 78 VIA_via2_5
* cell instance $6765 r0 *1 83.125,6.37
X$6765 78 VIA_via1_4
* cell instance $6766 r0 *1 83.125,10.43
X$6766 78 VIA_via1_4
* cell instance $6767 r0 *1 80.845,11.97
X$6767 78 VIA_via1_4
* cell instance $6768 r0 *1 80.845,11.83
X$6768 78 VIA_via2_5
* cell instance $6769 r0 *1 82.175,4.83
X$6769 78 VIA_via1_4
* cell instance $6770 r0 *1 68.495,18.83
X$6770 78 VIA_via1_4
* cell instance $6771 r0 *1 69.825,23.17
X$6771 78 VIA_via1_4
* cell instance $6772 r0 *1 67.355,21.63
X$6772 78 VIA_via1_4
* cell instance $6773 r0 *1 67.165,14.77
X$6773 78 VIA_via1_4
* cell instance $6774 r0 *1 68.115,16.03
X$6774 78 VIA_via1_4
* cell instance $6775 r0 *1 68.495,3.57
X$6775 78 VIA_via1_4
* cell instance $6776 r0 *1 79.895,37.03
X$6776 79 VIA_via1_7
* cell instance $6777 r0 *1 69.635,53.83
X$6777 79 VIA_via1_7
* cell instance $6778 r0 *1 73.245,4.97
X$6778 79 VIA_via1_7
* cell instance $6779 r0 *1 73.245,4.83
X$6779 79 VIA_via2_5
* cell instance $6780 r0 *1 91.485,6.23
X$6780 79 VIA_via1_7
* cell instance $6781 r0 *1 90.155,4.97
X$6781 79 VIA_via1_7
* cell instance $6782 r0 *1 80.845,48.23
X$6782 79 VIA_via1_7
* cell instance $6783 r0 *1 80.845,48.09
X$6783 79 VIA_via2_5
* cell instance $6784 r0 *1 91.485,5.39
X$6784 79 VIA_via2_5
* cell instance $6785 r0 *1 91.295,6.79
X$6785 79 VIA_via2_5
* cell instance $6786 r0 *1 90.155,5.39
X$6786 79 VIA_via2_5
* cell instance $6787 r0 *1 93.575,6.79
X$6787 79 VIA_via2_5
* cell instance $6788 r0 *1 80.465,50.47
X$6788 79 VIA_via2_5
* cell instance $6789 r0 *1 73.245,5.39
X$6789 79 VIA_via2_5
* cell instance $6790 r0 *1 69.635,52.85
X$6790 79 VIA_via2_5
* cell instance $6791 r0 *1 76.855,50.47
X$6791 79 VIA_via2_5
* cell instance $6792 r0 *1 76.855,52.85
X$6792 79 VIA_via2_5
* cell instance $6793 r0 *1 90.345,36.75
X$6793 79 VIA_via2_5
* cell instance $6794 r0 *1 81.225,36.75
X$6794 79 VIA_via2_5
* cell instance $6795 r0 *1 80.085,36.75
X$6795 79 VIA_via2_5
* cell instance $6796 r0 *1 80.465,48.09
X$6796 79 VIA_via2_5
* cell instance $6797 r0 *1 94.145,29.75
X$6797 79 VIA_via2_5
* cell instance $6798 r0 *1 94.335,33.81
X$6798 79 VIA_via2_5
* cell instance $6799 r0 *1 93.955,29.75
X$6799 79 VIA_via2_5
* cell instance $6800 r0 *1 90.345,33.81
X$6800 79 VIA_via2_5
* cell instance $6801 r0 *1 94.715,29.75
X$6801 79 VIA_via2_5
* cell instance $6802 r0 *1 80.845,42.21
X$6802 79 VIA_via2_5
* cell instance $6803 r0 *1 81.225,42.21
X$6803 79 VIA_via2_5
* cell instance $6804 r0 *1 94.715,30.03
X$6804 79 VIA_via1_4
* cell instance $6805 r0 *1 90.345,35.63
X$6805 79 VIA_via1_4
* cell instance $6806 r0 *1 93.575,18.83
X$6806 79 VIA_via1_4
* cell instance $6807 r0 *1 66.975,4.97
X$6807 79 VIA_via1_4
* cell instance $6808 r0 *1 66.975,4.97
X$6808 79 VIA_via2_5
* cell instance $6809 r0 *1 76.855,52.43
X$6809 79 VIA_via1_4
* cell instance $6810 r0 *1 79.705,30.17
X$6810 80 VIA_via1_7
* cell instance $6811 r0 *1 79.705,30.17
X$6811 80 VIA_via2_5
* cell instance $6812 r0 *1 44.745,6.23
X$6812 80 VIA_via1_7
* cell instance $6813 r0 *1 44.745,6.23
X$6813 80 VIA_via2_5
* cell instance $6814 r0 *1 56.525,6.23
X$6814 80 VIA_via1_7
* cell instance $6815 r0 *1 56.525,6.23
X$6815 80 VIA_via2_5
* cell instance $6816 r0 *1 70.015,4.97
X$6816 80 VIA_via1_7
* cell instance $6817 r0 *1 70.015,4.97
X$6817 80 VIA_via2_5
* cell instance $6818 r0 *1 64.695,4.97
X$6818 80 VIA_via1_7
* cell instance $6819 r0 *1 64.695,5.11
X$6819 80 VIA_via2_5
* cell instance $6820 r0 *1 77.425,4.97
X$6820 80 VIA_via1_7
* cell instance $6821 r0 *1 77.425,4.97
X$6821 80 VIA_via2_5
* cell instance $6822 r0 *1 50.445,6.79
X$6822 80 VIA_via2_5
* cell instance $6823 r0 *1 61.085,6.09
X$6823 80 VIA_via2_5
* cell instance $6824 r0 *1 56.525,6.93
X$6824 80 VIA_via2_5
* cell instance $6825 r0 *1 64.695,6.09
X$6825 80 VIA_via2_5
* cell instance $6826 r0 *1 51.015,27.51
X$6826 80 VIA_via2_5
* cell instance $6827 r0 *1 41.705,6.65
X$6827 80 VIA_via2_5
* cell instance $6828 r0 *1 45.315,6.79
X$6828 80 VIA_via2_5
* cell instance $6829 r0 *1 41.705,6.37
X$6829 80 VIA_via2_5
* cell instance $6830 r0 *1 45.315,6.37
X$6830 80 VIA_via2_5
* cell instance $6831 r0 *1 40.755,6.65
X$6831 80 VIA_via2_5
* cell instance $6832 r0 *1 79.705,20.37
X$6832 80 VIA_via1_4
* cell instance $6833 r0 *1 40.755,6.37
X$6833 80 VIA_via1_4
* cell instance $6834 r0 *1 61.085,6.37
X$6834 80 VIA_via1_4
* cell instance $6835 r0 *1 50.445,6.37
X$6835 80 VIA_via1_4
* cell instance $6836 r0 *1 48.545,27.51
X$6836 80 VIA_via1_4
* cell instance $6837 r0 *1 48.545,27.51
X$6837 80 VIA_via2_5
* cell instance $6838 r0 *1 79.895,20.65
X$6838 80 VIA_via3_2
* cell instance $6839 r0 *1 79.895,20.65
X$6839 80 VIA_via2_5
* cell instance $6840 r0 *1 80.175,30.17
X$6840 80 VIA_via3_2
* cell instance $6841 r0 *1 80.175,27.37
X$6841 80 VIA_via3_2
* cell instance $6842 r0 *1 73.815,6.51
X$6842 81 VIA_via2_5
* cell instance $6843 r0 *1 76.285,6.51
X$6843 81 VIA_via1_4
* cell instance $6844 r0 *1 76.285,6.51
X$6844 81 VIA_via2_5
* cell instance $6845 r0 *1 74.005,7.63
X$6845 81 VIA_via1_4
* cell instance $6846 r0 *1 74.005,4.83
X$6846 81 VIA_via1_4
* cell instance $6847 r0 *1 80.275,7.63
X$6847 82 VIA_via1_4
* cell instance $6848 r0 *1 80.085,4.83
X$6848 82 VIA_via1_4
* cell instance $6849 r0 *1 81.225,5.95
X$6849 82 VIA_via1_4
* cell instance $6850 r0 *1 89.965,4.83
X$6850 83 VIA_via2_5
* cell instance $6851 r0 *1 93.005,6.37
X$6851 83 VIA_via2_5
* cell instance $6852 r0 *1 93.195,10.29
X$6852 83 VIA_via2_5
* cell instance $6853 r0 *1 93.005,7.49
X$6853 83 VIA_via2_5
* cell instance $6854 r0 *1 93.005,11.97
X$6854 83 VIA_via1_4
* cell instance $6855 r0 *1 84.265,4.83
X$6855 83 VIA_via1_4
* cell instance $6856 r0 *1 84.265,4.83
X$6856 83 VIA_via2_5
* cell instance $6857 r0 *1 93.005,4.83
X$6857 83 VIA_via1_4
* cell instance $6858 r0 *1 88.445,4.83
X$6858 83 VIA_via1_4
* cell instance $6859 r0 *1 88.445,4.83
X$6859 83 VIA_via2_5
* cell instance $6860 r0 *1 91.105,7.63
X$6860 83 VIA_via1_4
* cell instance $6861 r0 *1 91.105,7.63
X$6861 83 VIA_via2_5
* cell instance $6862 r0 *1 90.155,7.63
X$6862 83 VIA_via1_4
* cell instance $6863 r0 *1 90.155,7.63
X$6863 83 VIA_via2_5
* cell instance $6864 r0 *1 95.095,10.43
X$6864 83 VIA_via1_4
* cell instance $6865 r0 *1 95.095,10.29
X$6865 83 VIA_via2_5
* cell instance $6866 r0 *1 94.335,6.37
X$6866 83 VIA_via1_4
* cell instance $6867 r0 *1 94.335,6.37
X$6867 83 VIA_via2_5
* cell instance $6868 r0 *1 93.195,7.63
X$6868 83 VIA_via1_4
* cell instance $6869 r0 *1 92.245,4.83
X$6869 84 VIA_via1_4
* cell instance $6870 r0 *1 92.245,4.69
X$6870 84 VIA_via2_5
* cell instance $6871 r0 *1 91.295,4.69
X$6871 84 VIA_via1_4
* cell instance $6872 r0 *1 91.295,4.69
X$6872 84 VIA_via2_5
* cell instance $6873 r0 *1 90.915,5.25
X$6873 85 VIA_via2_5
* cell instance $6874 r0 *1 89.395,5.25
X$6874 85 VIA_via2_5
* cell instance $6875 r0 *1 89.395,6.37
X$6875 85 VIA_via1_4
* cell instance $6876 r0 *1 94.525,4.83
X$6876 85 VIA_via1_4
* cell instance $6877 r0 *1 94.525,4.83
X$6877 85 VIA_via2_5
* cell instance $6878 r0 *1 90.915,4.83
X$6878 85 VIA_via1_4
* cell instance $6879 r0 *1 90.915,4.83
X$6879 85 VIA_via2_5
* cell instance $6880 r0 *1 85.405,4.69
X$6880 86 VIA_via2_5
* cell instance $6881 r0 *1 83.695,4.69
X$6881 86 VIA_via2_5
* cell instance $6882 r0 *1 83.505,7.63
X$6882 86 VIA_via1_4
* cell instance $6883 r0 *1 81.605,4.83
X$6883 86 VIA_via1_4
* cell instance $6884 r0 *1 81.605,4.69
X$6884 86 VIA_via2_5
* cell instance $6885 r0 *1 85.405,3.85
X$6885 86 VIA_via1_4
* cell instance $6886 r0 *1 14.725,5.95
X$6886 87 VIA_via2_5
* cell instance $6887 r0 *1 15.675,5.95
X$6887 87 VIA_via1_4
* cell instance $6888 r0 *1 15.675,5.95
X$6888 87 VIA_via2_5
* cell instance $6889 r0 *1 13.395,4.83
X$6889 87 VIA_via1_4
* cell instance $6890 r0 *1 13.395,4.83
X$6890 87 VIA_via2_5
* cell instance $6891 r0 *1 14.725,4.83
X$6891 87 VIA_via1_4
* cell instance $6892 r0 *1 14.725,4.83
X$6892 87 VIA_via2_5
* cell instance $6893 r0 *1 82.365,67.83
X$6893 88 VIA_via1_7
* cell instance $6894 r0 *1 68.305,7.77
X$6894 88 VIA_via1_7
* cell instance $6895 r0 *1 68.305,7.77
X$6895 88 VIA_via2_5
* cell instance $6896 r0 *1 82.555,60.97
X$6896 88 VIA_via1_7
* cell instance $6897 r0 *1 67.545,34.23
X$6897 88 VIA_via1_7
* cell instance $6898 r0 *1 67.545,34.23
X$6898 88 VIA_via2_5
* cell instance $6899 r0 *1 66.975,65.03
X$6899 88 VIA_via1_7
* cell instance $6900 r0 *1 66.975,65.03
X$6900 88 VIA_via2_5
* cell instance $6901 r0 *1 82.365,63.49
X$6901 88 VIA_via2_5
* cell instance $6902 r0 *1 78.565,63.49
X$6902 88 VIA_via2_5
* cell instance $6903 r0 *1 78.565,63.07
X$6903 88 VIA_via2_5
* cell instance $6904 r0 *1 76.285,35.63
X$6904 88 VIA_via2_5
* cell instance $6905 r0 *1 77.045,29.75
X$6905 88 VIA_via2_5
* cell instance $6906 r0 *1 83.315,29.75
X$6906 88 VIA_via2_5
* cell instance $6907 r0 *1 76.095,38.43
X$6907 88 VIA_via1_4
* cell instance $6908 r0 *1 79.895,4.83
X$6908 88 VIA_via1_4
* cell instance $6909 r0 *1 79.895,4.83
X$6909 88 VIA_via3_2
* cell instance $6910 r0 *1 79.895,4.83
X$6910 88 VIA_via2_5
* cell instance $6911 r0 *1 77.045,30.03
X$6911 88 VIA_via1_4
* cell instance $6912 r0 *1 81.415,4.83
X$6912 88 VIA_via1_4
* cell instance $6913 r0 *1 81.415,4.83
X$6913 88 VIA_via2_5
* cell instance $6914 r0 *1 83.505,25.97
X$6914 88 VIA_via1_4
* cell instance $6915 r0 *1 66.595,54.25
X$6915 88 VIA_via1_4
* cell instance $6916 r0 *1 66.595,54.25
X$6916 88 VIA_via2_5
* cell instance $6917 r0 *1 79.895,7.63
X$6917 88 VIA_via4_0
* cell instance $6918 r0 *1 68.695,7.63
X$6918 88 VIA_via4_0
* cell instance $6919 r0 *1 68.695,7.77
X$6919 88 VIA_via3_2
* cell instance $6920 r0 *1 68.415,54.25
X$6920 88 VIA_via3_2
* cell instance $6921 r0 *1 68.415,34.09
X$6921 88 VIA_via3_2
* cell instance $6922 r0 *1 68.415,63.21
X$6922 88 VIA_via3_2
* cell instance $6923 r0 *1 68.415,65.03
X$6923 88 VIA_via3_2
* cell instance $6924 r0 *1 76.535,34.09
X$6924 88 VIA_via3_2
* cell instance $6925 r0 *1 76.535,29.75
X$6925 88 VIA_via3_2
* cell instance $6926 r0 *1 76.535,35.63
X$6926 88 VIA_via3_2
* cell instance $6927 r0 *1 40.375,5.81
X$6927 89 VIA_via1_7
* cell instance $6928 r0 *1 40.375,4.83
X$6928 89 VIA_via2_5
* cell instance $6929 r0 *1 37.525,4.83
X$6929 89 VIA_via1_4
* cell instance $6930 r0 *1 37.525,4.83
X$6930 89 VIA_via2_5
* cell instance $6931 r0 *1 64.885,6.37
X$6931 90 VIA_via2_5
* cell instance $6932 r0 *1 63.555,4.83
X$6932 90 VIA_via1_4
* cell instance $6933 r0 *1 63.555,4.83
X$6933 90 VIA_via2_5
* cell instance $6934 r0 *1 64.885,4.83
X$6934 90 VIA_via1_4
* cell instance $6935 r0 *1 64.885,4.83
X$6935 90 VIA_via2_5
* cell instance $6936 r0 *1 65.645,6.37
X$6936 90 VIA_via1_4
* cell instance $6937 r0 *1 65.645,6.37
X$6937 90 VIA_via2_5
* cell instance $6938 r0 *1 44.555,5.81
X$6938 91 VIA_via1_7
* cell instance $6939 r0 *1 44.555,4.83
X$6939 91 VIA_via2_5
* cell instance $6940 r0 *1 43.035,4.83
X$6940 91 VIA_via1_4
* cell instance $6941 r0 *1 43.035,4.83
X$6941 91 VIA_via2_5
* cell instance $6942 r0 *1 50.255,5.81
X$6942 92 VIA_via1_7
* cell instance $6943 r0 *1 50.255,4.83
X$6943 92 VIA_via2_5
* cell instance $6944 r0 *1 48.735,4.83
X$6944 92 VIA_via1_4
* cell instance $6945 r0 *1 48.735,4.83
X$6945 92 VIA_via2_5
* cell instance $6946 r0 *1 19.855,5.81
X$6946 93 VIA_via1_7
* cell instance $6947 r0 *1 19.285,4.83
X$6947 93 VIA_via1_4
* cell instance $6948 r0 *1 22.515,6.23
X$6948 94 VIA_via1_4
* cell instance $6949 r0 *1 21.945,14.77
X$6949 94 VIA_via1_4
* cell instance $6950 r0 *1 26.885,6.23
X$6950 95 VIA_via1_4
* cell instance $6951 r0 *1 26.505,13.23
X$6951 95 VIA_via1_4
* cell instance $6952 r0 *1 30.305,5.81
X$6952 96 VIA_via1_7
* cell instance $6953 r0 *1 29.735,4.83
X$6953 96 VIA_via1_4
* cell instance $6954 r0 *1 36.575,5.39
X$6954 97 VIA_via1_7
* cell instance $6955 r0 *1 36.765,6.37
X$6955 97 VIA_via1_4
* cell instance $6956 r0 *1 38.475,6.23
X$6956 98 VIA_via2_5
* cell instance $6957 r0 *1 39.425,8.89
X$6957 98 VIA_via2_5
* cell instance $6958 r0 *1 39.425,5.39
X$6958 98 VIA_via2_5
* cell instance $6959 r0 *1 40.185,5.39
X$6959 98 VIA_via2_5
* cell instance $6960 r0 *1 40.565,29.75
X$6960 98 VIA_via2_5
* cell instance $6961 r0 *1 39.235,29.75
X$6961 98 VIA_via2_5
* cell instance $6962 r0 *1 38.855,8.89
X$6962 98 VIA_via2_5
* cell instance $6963 r0 *1 40.375,8.89
X$6963 98 VIA_via2_5
* cell instance $6964 r0 *1 39.425,17.57
X$6964 98 VIA_via1_4
* cell instance $6965 r0 *1 38.855,11.97
X$6965 98 VIA_via1_4
* cell instance $6966 r0 *1 39.425,6.37
X$6966 98 VIA_via1_4
* cell instance $6967 r0 *1 39.425,6.23
X$6967 98 VIA_via2_5
* cell instance $6968 r0 *1 40.375,9.17
X$6968 98 VIA_via1_4
* cell instance $6969 r0 *1 40.185,4.83
X$6969 98 VIA_via1_4
* cell instance $6970 r0 *1 38.475,2.45
X$6970 98 VIA_via1_4
* cell instance $6971 r0 *1 39.235,31.57
X$6971 98 VIA_via1_4
* cell instance $6972 r0 *1 40.565,30.03
X$6972 98 VIA_via1_4
* cell instance $6973 r0 *1 51.015,5.25
X$6973 99 VIA_via1_4
* cell instance $6974 r0 *1 50.635,6.37
X$6974 99 VIA_via1_4
* cell instance $6975 r0 *1 50.635,6.37
X$6975 99 VIA_via2_5
* cell instance $6976 r0 *1 49.875,6.37
X$6976 99 VIA_via1_4
* cell instance $6977 r0 *1 49.875,6.37
X$6977 99 VIA_via2_5
* cell instance $6978 r0 *1 51.585,6.23
X$6978 100 VIA_via1_4
* cell instance $6979 r0 *1 51.585,13.23
X$6979 100 VIA_via1_4
* cell instance $6980 r0 *1 59.185,5.81
X$6980 101 VIA_via1_7
* cell instance $6981 r0 *1 58.805,4.83
X$6981 101 VIA_via1_4
* cell instance $6982 r0 *1 60.705,5.81
X$6982 102 VIA_via1_7
* cell instance $6983 r0 *1 60.325,3.57
X$6983 102 VIA_via1_4
* cell instance $6984 r0 *1 58.805,6.37
X$6984 103 VIA_via1_4
* cell instance $6985 r0 *1 58.805,6.51
X$6985 103 VIA_via2_5
* cell instance $6986 r0 *1 61.275,6.37
X$6986 103 VIA_via1_4
* cell instance $6987 r0 *1 61.275,6.51
X$6987 103 VIA_via2_5
* cell instance $6988 r0 *1 61.085,5.25
X$6988 103 VIA_via1_4
* cell instance $6989 r0 *1 63.935,5.39
X$6989 104 VIA_via1_7
* cell instance $6990 r0 *1 63.365,6.37
X$6990 104 VIA_via1_4
* cell instance $6991 r0 *1 65.835,5.39
X$6991 105 VIA_via1_7
* cell instance $6992 r0 *1 65.645,18.83
X$6992 105 VIA_via1_4
* cell instance $6993 r0 *1 11.685,6.09
X$6993 106 VIA_via2_5
* cell instance $6994 r0 *1 10.735,6.09
X$6994 106 VIA_via1_4
* cell instance $6995 r0 *1 10.735,6.09
X$6995 106 VIA_via2_5
* cell instance $6996 r0 *1 12.065,9.17
X$6996 106 VIA_via1_4
* cell instance $6997 r0 *1 11.685,6.37
X$6997 106 VIA_via1_4
* cell instance $6998 r0 *1 5.415,25.97
X$6998 107 VIA_via2_5
* cell instance $6999 r0 *1 5.415,25.41
X$6999 107 VIA_via2_5
* cell instance $7000 r0 *1 8.455,25.41
X$7000 107 VIA_via2_5
* cell instance $7001 r0 *1 12.825,12.11
X$7001 107 VIA_via2_5
* cell instance $7002 r0 *1 4.465,27.23
X$7002 107 VIA_via2_5
* cell instance $7003 r0 *1 9.595,12.39
X$7003 107 VIA_via2_5
* cell instance $7004 r0 *1 15.675,25.41
X$7004 107 VIA_via2_5
* cell instance $7005 r0 *1 12.825,4.83
X$7005 107 VIA_via1_4
* cell instance $7006 r0 *1 12.825,4.97
X$7006 107 VIA_via2_5
* cell instance $7007 r0 *1 10.925,4.83
X$7007 107 VIA_via1_4
* cell instance $7008 r0 *1 10.925,4.97
X$7008 107 VIA_via2_5
* cell instance $7009 r0 *1 13.965,11.97
X$7009 107 VIA_via1_4
* cell instance $7010 r0 *1 13.965,12.11
X$7010 107 VIA_via2_5
* cell instance $7011 r0 *1 9.595,13.23
X$7011 107 VIA_via1_4
* cell instance $7012 r0 *1 5.415,27.23
X$7012 107 VIA_via1_4
* cell instance $7013 r0 *1 5.415,27.23
X$7013 107 VIA_via2_5
* cell instance $7014 r0 *1 4.085,30.03
X$7014 107 VIA_via1_4
* cell instance $7015 r0 *1 2.185,25.97
X$7015 107 VIA_via1_4
* cell instance $7016 r0 *1 2.185,25.97
X$7016 107 VIA_via2_5
* cell instance $7017 r0 *1 15.865,30.03
X$7017 107 VIA_via1_4
* cell instance $7018 r0 *1 88.445,5.81
X$7018 108 VIA_via1_7
* cell instance $7019 r0 *1 88.445,5.81
X$7019 108 VIA_via2_5
* cell instance $7020 r0 *1 87.685,5.81
X$7020 108 VIA_via2_5
* cell instance $7021 r0 *1 87.685,4.83
X$7021 108 VIA_via1_4
* cell instance $7022 r0 *1 83.505,5.81
X$7022 109 VIA_via1_7
* cell instance $7023 r0 *1 83.505,4.83
X$7023 109 VIA_via1_4
* cell instance $7024 r0 *1 78.565,5.39
X$7024 110 VIA_via1_7
* cell instance $7025 r0 *1 78.565,5.53
X$7025 110 VIA_via2_5
* cell instance $7026 r0 *1 77.805,5.53
X$7026 110 VIA_via2_5
* cell instance $7027 r0 *1 77.805,18.83
X$7027 110 VIA_via1_4
* cell instance $7028 r0 *1 33.725,5.81
X$7028 111 VIA_via1_7
* cell instance $7029 r0 *1 33.725,5.81
X$7029 111 VIA_via2_5
* cell instance $7030 r0 *1 32.965,5.81
X$7030 111 VIA_via2_5
* cell instance $7031 r0 *1 32.965,4.83
X$7031 111 VIA_via1_4
* cell instance $7032 r0 *1 55.195,15.89
X$7032 112 VIA_via2_5
* cell instance $7033 r0 *1 54.435,6.09
X$7033 112 VIA_via2_5
* cell instance $7034 r0 *1 55.765,6.09
X$7034 112 VIA_via2_5
* cell instance $7035 r0 *1 56.715,6.09
X$7035 112 VIA_via2_5
* cell instance $7036 r0 *1 54.625,32.83
X$7036 112 VIA_via2_5
* cell instance $7037 r0 *1 56.905,32.83
X$7037 112 VIA_via1_4
* cell instance $7038 r0 *1 56.905,32.83
X$7038 112 VIA_via2_5
* cell instance $7039 r0 *1 56.905,35.63
X$7039 112 VIA_via1_4
* cell instance $7040 r0 *1 54.435,2.45
X$7040 112 VIA_via1_4
* cell instance $7041 r0 *1 54.435,6.37
X$7041 112 VIA_via1_4
* cell instance $7042 r0 *1 54.625,24.43
X$7042 112 VIA_via1_4
* cell instance $7043 r0 *1 56.145,16.03
X$7043 112 VIA_via1_4
* cell instance $7044 r0 *1 56.145,15.89
X$7044 112 VIA_via2_5
* cell instance $7045 r0 *1 54.815,16.03
X$7045 112 VIA_via1_4
* cell instance $7046 r0 *1 54.815,15.89
X$7046 112 VIA_via2_5
* cell instance $7047 r0 *1 56.715,4.83
X$7047 112 VIA_via1_4
* cell instance $7048 r0 *1 55.385,5.81
X$7048 113 VIA_via1_7
* cell instance $7049 r0 *1 55.385,4.97
X$7049 113 VIA_via2_5
* cell instance $7050 r0 *1 54.055,4.83
X$7050 113 VIA_via1_4
* cell instance $7051 r0 *1 54.055,4.97
X$7051 113 VIA_via2_5
* cell instance $7052 r0 *1 13.775,5.39
X$7052 114 VIA_via1_7
* cell instance $7053 r0 *1 13.395,6.37
X$7053 114 VIA_via1_4
* cell instance $7054 r0 *1 27.455,6.37
X$7054 115 VIA_via2_5
* cell instance $7055 r0 *1 25.365,6.37
X$7055 115 VIA_via2_5
* cell instance $7056 r0 *1 27.455,5.25
X$7056 115 VIA_via1_4
* cell instance $7057 r0 *1 25.175,6.37
X$7057 115 VIA_via1_4
* cell instance $7058 r0 *1 26.505,6.37
X$7058 115 VIA_via1_4
* cell instance $7059 r0 *1 26.505,6.37
X$7059 115 VIA_via2_5
* cell instance $7060 r0 *1 32.015,6.37
X$7060 116 VIA_via2_5
* cell instance $7061 r0 *1 30.875,6.37
X$7061 116 VIA_via1_4
* cell instance $7062 r0 *1 30.875,6.37
X$7062 116 VIA_via2_5
* cell instance $7063 r0 *1 32.015,5.25
X$7063 116 VIA_via1_4
* cell instance $7064 r0 *1 29.925,6.37
X$7064 116 VIA_via1_4
* cell instance $7065 r0 *1 29.925,6.37
X$7065 116 VIA_via2_5
* cell instance $7066 r0 *1 35.245,6.37
X$7066 117 VIA_via2_5
* cell instance $7067 r0 *1 33.345,6.37
X$7067 117 VIA_via1_4
* cell instance $7068 r0 *1 33.345,6.37
X$7068 117 VIA_via2_5
* cell instance $7069 r0 *1 34.105,6.37
X$7069 117 VIA_via1_4
* cell instance $7070 r0 *1 34.105,6.37
X$7070 117 VIA_via2_5
* cell instance $7071 r0 *1 35.245,5.25
X$7071 117 VIA_via1_4
* cell instance $7072 r0 *1 36.195,6.37
X$7072 118 VIA_via2_5
* cell instance $7073 r0 *1 34.675,6.37
X$7073 118 VIA_via1_4
* cell instance $7074 r0 *1 34.675,6.51
X$7074 118 VIA_via2_5
* cell instance $7075 r0 *1 36.195,4.83
X$7075 118 VIA_via1_4
* cell instance $7076 r0 *1 39.045,6.37
X$7076 118 VIA_via1_4
* cell instance $7077 r0 *1 39.045,6.37
X$7077 118 VIA_via2_5
* cell instance $7078 r0 *1 39.995,6.37
X$7078 119 VIA_via1_4
* cell instance $7079 r0 *1 39.995,6.37
X$7079 119 VIA_via2_5
* cell instance $7080 r0 *1 40.945,6.37
X$7080 119 VIA_via1_4
* cell instance $7081 r0 *1 40.945,6.37
X$7081 119 VIA_via2_5
* cell instance $7082 r0 *1 39.805,5.25
X$7082 119 VIA_via1_4
* cell instance $7083 r0 *1 44.935,6.37
X$7083 120 VIA_via1_4
* cell instance $7084 r0 *1 44.175,6.37
X$7084 120 VIA_via1_4
* cell instance $7085 r0 *1 45.315,5.25
X$7085 120 VIA_via1_4
* cell instance $7086 r0 *1 57.475,10.01
X$7086 121 VIA_via2_5
* cell instance $7087 r0 *1 55.575,10.01
X$7087 121 VIA_via2_5
* cell instance $7088 r0 *1 57.095,6.37
X$7088 121 VIA_via2_5
* cell instance $7089 r0 *1 57.095,10.01
X$7089 121 VIA_via2_5
* cell instance $7090 r0 *1 57.665,31.71
X$7090 121 VIA_via2_5
* cell instance $7091 r0 *1 58.615,31.57
X$7091 121 VIA_via1_4
* cell instance $7092 r0 *1 58.615,31.71
X$7092 121 VIA_via2_5
* cell instance $7093 r0 *1 59.375,35.63
X$7093 121 VIA_via1_4
* cell instance $7094 r0 *1 58.235,6.37
X$7094 121 VIA_via1_4
* cell instance $7095 r0 *1 58.235,6.37
X$7095 121 VIA_via2_5
* cell instance $7096 r0 *1 59.755,6.37
X$7096 121 VIA_via1_4
* cell instance $7097 r0 *1 59.755,6.37
X$7097 121 VIA_via2_5
* cell instance $7098 r0 *1 57.095,11.97
X$7098 121 VIA_via1_4
* cell instance $7099 r0 *1 55.575,10.43
X$7099 121 VIA_via1_4
* cell instance $7100 r0 *1 58.995,32.83
X$7100 121 VIA_via1_4
* cell instance $7101 r0 *1 59.945,2.45
X$7101 121 VIA_via1_4
* cell instance $7102 r0 *1 62.605,6.37
X$7102 122 VIA_via2_5
* cell instance $7103 r0 *1 60.325,6.37
X$7103 122 VIA_via1_4
* cell instance $7104 r0 *1 60.325,6.37
X$7104 122 VIA_via2_5
* cell instance $7105 r0 *1 62.605,3.85
X$7105 122 VIA_via1_4
* cell instance $7106 r0 *1 61.845,6.37
X$7106 122 VIA_via1_4
* cell instance $7107 r0 *1 61.845,6.37
X$7107 122 VIA_via2_5
* cell instance $7108 r0 *1 63.175,6.23
X$7108 123 VIA_via2_5
* cell instance $7109 r0 *1 63.175,20.37
X$7109 123 VIA_via1_4
* cell instance $7110 r0 *1 62.225,6.23
X$7110 123 VIA_via1_4
* cell instance $7111 r0 *1 62.225,6.23
X$7111 123 VIA_via2_5
* cell instance $7112 r0 *1 68.495,7.63
X$7112 124 VIA_via1_4
* cell instance $7113 r0 *1 69.065,6.65
X$7113 124 VIA_via1_4
* cell instance $7114 r0 *1 68.305,9.17
X$7114 124 VIA_via1_4
* cell instance $7115 r0 *1 74.385,5.39
X$7115 125 VIA_via1_7
* cell instance $7116 r0 *1 74.005,6.37
X$7116 125 VIA_via1_4
* cell instance $7117 r0 *1 57.285,16.17
X$7117 126 VIA_via1_7
* cell instance $7118 r0 *1 57.285,16.17
X$7118 126 VIA_via2_5
* cell instance $7119 r0 *1 68.305,30.17
X$7119 126 VIA_via1_7
* cell instance $7120 r0 *1 73.245,7.77
X$7120 126 VIA_via1_7
* cell instance $7121 r0 *1 90.725,9.03
X$7121 126 VIA_via1_7
* cell instance $7122 r0 *1 60.325,10.01
X$7122 126 VIA_via2_5
* cell instance $7123 r0 *1 90.725,8.05
X$7123 126 VIA_via2_5
* cell instance $7124 r0 *1 56.905,10.15
X$7124 126 VIA_via2_5
* cell instance $7125 r0 *1 53.105,10.15
X$7125 126 VIA_via2_5
* cell instance $7126 r0 *1 56.715,15.61
X$7126 126 VIA_via2_5
* cell instance $7127 r0 *1 88.445,7.91
X$7127 126 VIA_via2_5
* cell instance $7128 r0 *1 73.245,10.01
X$7128 126 VIA_via2_5
* cell instance $7129 r0 *1 73.245,8.05
X$7129 126 VIA_via2_5
* cell instance $7130 r0 *1 68.305,30.73
X$7130 126 VIA_via2_5
* cell instance $7131 r0 *1 68.305,31.43
X$7131 126 VIA_via2_5
* cell instance $7132 r0 *1 88.635,31.71
X$7132 126 VIA_via2_5
* cell instance $7133 r0 *1 93.575,32.69
X$7133 126 VIA_via2_5
* cell instance $7134 r0 *1 88.635,32.69
X$7134 126 VIA_via2_5
* cell instance $7135 r0 *1 91.675,32.69
X$7135 126 VIA_via2_5
* cell instance $7136 r0 *1 88.635,6.37
X$7136 126 VIA_via1_4
* cell instance $7137 r0 *1 91.675,35.63
X$7137 126 VIA_via1_4
* cell instance $7138 r0 *1 93.575,31.57
X$7138 126 VIA_via1_4
* cell instance $7139 r0 *1 60.325,10.43
X$7139 126 VIA_via1_4
* cell instance $7140 r0 *1 53.105,10.43
X$7140 126 VIA_via1_4
* cell instance $7141 r0 *1 93.575,23.17
X$7141 126 VIA_via1_4
* cell instance $7142 r0 *1 55.005,35.91
X$7142 126 VIA_via1_4
* cell instance $7143 r0 *1 55.005,35.91
X$7143 126 VIA_via2_5
* cell instance $7144 r0 *1 57.495,16.17
X$7144 126 VIA_via3_2
* cell instance $7145 r0 *1 57.495,15.61
X$7145 126 VIA_via3_2
* cell instance $7146 r0 *1 57.495,30.73
X$7146 126 VIA_via3_2
* cell instance $7147 r0 *1 57.495,35.91
X$7147 126 VIA_via3_2
* cell instance $7148 r0 *1 91.485,6.51
X$7148 127 VIA_via2_5
* cell instance $7149 r0 *1 95.855,6.65
X$7149 127 VIA_via1_4
* cell instance $7150 r0 *1 95.855,6.65
X$7150 127 VIA_via2_5
* cell instance $7151 r0 *1 91.485,9.17
X$7151 127 VIA_via1_4
* cell instance $7152 r0 *1 92.245,6.37
X$7152 127 VIA_via1_4
* cell instance $7153 r0 *1 92.245,6.51
X$7153 127 VIA_via2_5
* cell instance $7154 r0 *1 93.575,6.37
X$7154 128 VIA_via1_4
* cell instance $7155 r0 *1 93.575,6.51
X$7155 128 VIA_via2_5
* cell instance $7156 r0 *1 92.625,6.51
X$7156 128 VIA_via1_4
* cell instance $7157 r0 *1 92.625,6.51
X$7157 128 VIA_via2_5
* cell instance $7158 r0 *1 12.065,6.51
X$7158 129 VIA_via1_4
* cell instance $7159 r0 *1 12.065,6.51
X$7159 129 VIA_via2_5
* cell instance $7160 r0 *1 8.455,6.37
X$7160 129 VIA_via1_4
* cell instance $7161 r0 *1 8.455,6.51
X$7161 129 VIA_via2_5
* cell instance $7162 r0 *1 79.895,39.83
X$7162 130 VIA_via1_7
* cell instance $7163 r0 *1 77.425,7.77
X$7163 130 VIA_via1_7
* cell instance $7164 r0 *1 66.215,9.03
X$7164 130 VIA_via1_7
* cell instance $7165 r0 *1 66.215,8.89
X$7165 130 VIA_via2_5
* cell instance $7166 r0 *1 66.215,54.95
X$7166 130 VIA_via2_5
* cell instance $7167 r0 *1 66.595,63.35
X$7167 130 VIA_via2_5
* cell instance $7168 r0 *1 77.425,8.89
X$7168 130 VIA_via2_5
* cell instance $7169 r0 *1 77.425,6.51
X$7169 130 VIA_via2_5
* cell instance $7170 r0 *1 85.025,63.35
X$7170 130 VIA_via2_5
* cell instance $7171 r0 *1 75.145,32.55
X$7171 130 VIA_via2_5
* cell instance $7172 r0 *1 79.895,31.99
X$7172 130 VIA_via2_5
* cell instance $7173 r0 *1 79.895,32.55
X$7173 130 VIA_via2_5
* cell instance $7174 r0 *1 86.355,31.99
X$7174 130 VIA_via2_5
* cell instance $7175 r0 *1 66.595,63.63
X$7175 130 VIA_via1_4
* cell instance $7176 r0 *1 82.365,6.37
X$7176 130 VIA_via1_4
* cell instance $7177 r0 *1 82.365,6.51
X$7177 130 VIA_via2_5
* cell instance $7178 r0 *1 86.735,25.97
X$7178 130 VIA_via1_4
* cell instance $7179 r0 *1 75.145,32.83
X$7179 130 VIA_via1_4
* cell instance $7180 r0 *1 64.695,54.95
X$7180 130 VIA_via1_4
* cell instance $7181 r0 *1 64.695,54.95
X$7181 130 VIA_via2_5
* cell instance $7182 r0 *1 85.595,66.43
X$7182 130 VIA_via1_4
* cell instance $7183 r0 *1 85.405,63.63
X$7183 130 VIA_via1_4
* cell instance $7184 r0 *1 67.545,32.83
X$7184 130 VIA_via1_4
* cell instance $7185 r0 *1 67.575,8.89
X$7185 130 VIA_via3_2
* cell instance $7186 r0 *1 66.735,54.95
X$7186 130 VIA_via3_2
* cell instance $7187 r0 *1 67.575,32.55
X$7187 130 VIA_via3_2
* cell instance $7188 r0 *1 67.545,32.55
X$7188 130 VIA_via2_5
* cell instance $7189 r0 *1 21.565,5.25
X$7189 131 VIA_via1_4
* cell instance $7190 r0 *1 19.475,6.37
X$7190 131 VIA_via1_4
* cell instance $7191 r0 *1 19.475,6.37
X$7191 131 VIA_via2_5
* cell instance $7192 r0 *1 21.565,6.37
X$7192 131 VIA_via1_4
* cell instance $7193 r0 *1 21.565,6.37
X$7193 131 VIA_via2_5
* cell instance $7194 r0 *1 81.035,5.39
X$7194 132 VIA_via1_7
* cell instance $7195 r0 *1 81.035,6.37
X$7195 132 VIA_via2_5
* cell instance $7196 r0 *1 78.945,6.37
X$7196 132 VIA_via1_4
* cell instance $7197 r0 *1 78.945,6.37
X$7197 132 VIA_via2_5
* cell instance $7198 r0 *1 66.405,55.37
X$7198 133 VIA_via1_7
* cell instance $7199 r0 *1 66.405,55.37
X$7199 133 VIA_via2_5
* cell instance $7200 r0 *1 92.055,9.03
X$7200 133 VIA_via1_7
* cell instance $7201 r0 *1 76.665,55.37
X$7201 133 VIA_via1_7
* cell instance $7202 r0 *1 76.665,55.37
X$7202 133 VIA_via2_5
* cell instance $7203 r0 *1 80.655,51.03
X$7203 133 VIA_via1_7
* cell instance $7204 r0 *1 80.655,51.03
X$7204 133 VIA_via2_5
* cell instance $7205 r0 *1 92.055,7.49
X$7205 133 VIA_via2_5
* cell instance $7206 r0 *1 92.055,10.57
X$7206 133 VIA_via2_5
* cell instance $7207 r0 *1 87.305,7.49
X$7207 133 VIA_via2_5
* cell instance $7208 r0 *1 70.585,6.51
X$7208 133 VIA_via2_5
* cell instance $7209 r0 *1 70.585,7.49
X$7209 133 VIA_via2_5
* cell instance $7210 r0 *1 94.905,23.45
X$7210 133 VIA_via2_5
* cell instance $7211 r0 *1 62.225,6.51
X$7211 133 VIA_via2_5
* cell instance $7212 r0 *1 77.615,55.09
X$7212 133 VIA_via2_5
* cell instance $7213 r0 *1 77.615,55.37
X$7213 133 VIA_via2_5
* cell instance $7214 r0 *1 83.505,42.91
X$7214 133 VIA_via2_5
* cell instance $7215 r0 *1 82.365,42.91
X$7215 133 VIA_via2_5
* cell instance $7216 r0 *1 82.175,46.27
X$7216 133 VIA_via2_5
* cell instance $7217 r0 *1 80.655,46.27
X$7217 133 VIA_via2_5
* cell instance $7218 r0 *1 94.525,36.89
X$7218 133 VIA_via2_5
* cell instance $7219 r0 *1 93.195,29.47
X$7219 133 VIA_via2_5
* cell instance $7220 r0 *1 94.905,29.47
X$7220 133 VIA_via2_5
* cell instance $7221 r0 *1 83.125,36.89
X$7221 133 VIA_via2_5
* cell instance $7222 r0 *1 83.125,37.17
X$7222 133 VIA_via1_4
* cell instance $7223 r0 *1 93.195,30.03
X$7223 133 VIA_via1_4
* cell instance $7224 r0 *1 87.305,6.37
X$7224 133 VIA_via1_4
* cell instance $7225 r0 *1 94.335,34.37
X$7225 133 VIA_via1_4
* cell instance $7226 r0 *1 94.905,23.17
X$7226 133 VIA_via1_4
* cell instance $7227 r0 *1 70.205,6.37
X$7227 133 VIA_via1_4
* cell instance $7228 r0 *1 70.205,6.51
X$7228 133 VIA_via2_5
* cell instance $7229 r0 *1 62.225,7.35
X$7229 133 VIA_via1_4
* cell instance $7230 r0 *1 93.615,23.45
X$7230 133 VIA_via3_2
* cell instance $7231 r0 *1 93.615,10.57
X$7231 133 VIA_via3_2
* cell instance $7232 r0 *1 80.455,51.03
X$7232 133 VIA_via3_2
* cell instance $7233 r0 *1 80.455,55.09
X$7233 133 VIA_via3_2
* cell instance $7234 r0 *1 58.805,18.55
X$7234 134 VIA_via2_5
* cell instance $7235 r0 *1 60.895,18.55
X$7235 134 VIA_via2_5
* cell instance $7236 r0 *1 60.895,6.23
X$7236 134 VIA_via2_5
* cell instance $7237 r0 *1 57.665,6.23
X$7237 134 VIA_via1_4
* cell instance $7238 r0 *1 57.665,6.23
X$7238 134 VIA_via2_5
* cell instance $7239 r0 *1 58.805,20.37
X$7239 134 VIA_via1_4
* cell instance $7240 r0 *1 56.335,6.37
X$7240 135 VIA_via2_5
* cell instance $7241 r0 *1 56.715,6.37
X$7241 135 VIA_via1_4
* cell instance $7242 r0 *1 56.715,6.37
X$7242 135 VIA_via2_5
* cell instance $7243 r0 *1 55.005,6.37
X$7243 135 VIA_via1_4
* cell instance $7244 r0 *1 55.005,6.37
X$7244 135 VIA_via2_5
* cell instance $7245 r0 *1 56.335,5.25
X$7245 135 VIA_via1_4
* cell instance $7246 r0 *1 17.575,9.31
X$7246 136 VIA_via2_5
* cell instance $7247 r0 *1 17.575,10.43
X$7247 136 VIA_via1_4
* cell instance $7248 r0 *1 17.955,8.05
X$7248 136 VIA_via1_4
* cell instance $7249 r0 *1 14.915,9.17
X$7249 136 VIA_via1_4
* cell instance $7250 r0 *1 14.915,9.31
X$7250 136 VIA_via2_5
* cell instance $7251 r0 *1 53.295,9.17
X$7251 137 VIA_via2_5
* cell instance $7252 r0 *1 53.295,10.43
X$7252 137 VIA_via1_4
* cell instance $7253 r0 *1 52.915,8.05
X$7253 137 VIA_via1_4
* cell instance $7254 r0 *1 50.255,9.17
X$7254 137 VIA_via1_4
* cell instance $7255 r0 *1 50.255,9.17
X$7255 137 VIA_via2_5
* cell instance $7256 r0 *1 59.375,56.35
X$7256 138 VIA_via1_7
* cell instance $7257 r0 *1 59.375,56.35
X$7257 138 VIA_via2_5
* cell instance $7258 r0 *1 58.045,6.79
X$7258 138 VIA_via2_5
* cell instance $7259 r0 *1 53.295,6.79
X$7259 138 VIA_via2_5
* cell instance $7260 r0 *1 54.245,6.79
X$7260 138 VIA_via2_5
* cell instance $7261 r0 *1 58.045,7.91
X$7261 138 VIA_via2_5
* cell instance $7262 r0 *1 59.375,56.77
X$7262 138 VIA_via2_5
* cell instance $7263 r0 *1 61.275,7.91
X$7263 138 VIA_via2_5
* cell instance $7264 r0 *1 58.045,6.37
X$7264 138 VIA_via1_4
* cell instance $7265 r0 *1 53.295,6.37
X$7265 138 VIA_via1_4
* cell instance $7266 r0 *1 54.245,6.37
X$7266 138 VIA_via1_4
* cell instance $7267 r0 *1 61.275,7.63
X$7267 138 VIA_via1_4
* cell instance $7268 r0 *1 57.095,56.77
X$7268 138 VIA_via1_4
* cell instance $7269 r0 *1 57.095,56.77
X$7269 138 VIA_via2_5
* cell instance $7270 r0 *1 59.735,7.91
X$7270 138 VIA_via4_0
* cell instance $7271 r0 *1 59.735,7.91
X$7271 138 VIA_via5_0
* cell instance $7272 r0 *1 59.735,7.91
X$7272 138 VIA_via3_2
* cell instance $7273 r0 *1 59.735,56.35
X$7273 138 VIA_via3_2
* cell instance $7274 r0 *1 59.735,56.35
X$7274 138 VIA_via4_0
* cell instance $7275 r0 *1 59.735,56.35
X$7275 138 VIA_via5_0
* cell instance $7276 r0 *1 55.765,16.87
X$7276 139 VIA_via2_5
* cell instance $7277 r0 *1 81.035,18.69
X$7277 139 VIA_via2_5
* cell instance $7278 r0 *1 76.475,18.55
X$7278 139 VIA_via2_5
* cell instance $7279 r0 *1 66.405,16.87
X$7279 139 VIA_via2_5
* cell instance $7280 r0 *1 64.505,16.87
X$7280 139 VIA_via2_5
* cell instance $7281 r0 *1 66.405,18.83
X$7281 139 VIA_via2_5
* cell instance $7282 r0 *1 81.035,23.17
X$7282 139 VIA_via1_4
* cell instance $7283 r0 *1 76.095,7.63
X$7283 139 VIA_via1_4
* cell instance $7284 r0 *1 76.095,7.77
X$7284 139 VIA_via2_5
* cell instance $7285 r0 *1 84.645,7.63
X$7285 139 VIA_via1_4
* cell instance $7286 r0 *1 84.645,7.77
X$7286 139 VIA_via2_5
* cell instance $7287 r0 *1 90.725,7.63
X$7287 139 VIA_via1_4
* cell instance $7288 r0 *1 90.725,7.77
X$7288 139 VIA_via2_5
* cell instance $7289 r0 *1 74.575,20.37
X$7289 139 VIA_via1_4
* cell instance $7290 r0 *1 74.765,18.69
X$7290 139 VIA_via1_4
* cell instance $7291 r0 *1 74.765,18.69
X$7291 139 VIA_via2_5
* cell instance $7292 r0 *1 55.955,7.63
X$7292 139 VIA_via1_4
* cell instance $7293 r0 *1 55.955,7.63
X$7293 139 VIA_via2_5
* cell instance $7294 r0 *1 66.405,16.03
X$7294 139 VIA_via1_4
* cell instance $7295 r0 *1 55.765,18.83
X$7295 139 VIA_via1_4
* cell instance $7296 r0 *1 91.865,18.83
X$7296 139 VIA_via1_4
* cell instance $7297 r0 *1 91.865,18.69
X$7297 139 VIA_via2_5
* cell instance $7298 r0 *1 66.595,25.97
X$7298 139 VIA_via1_4
* cell instance $7299 r0 *1 64.125,7.63
X$7299 139 VIA_via1_4
* cell instance $7300 r0 *1 64.125,7.63
X$7300 139 VIA_via2_5
* cell instance $7301 r0 *1 67.925,9.17
X$7301 140 VIA_via2_5
* cell instance $7302 r0 *1 68.875,9.17
X$7302 140 VIA_via1_4
* cell instance $7303 r0 *1 68.875,9.17
X$7303 140 VIA_via2_5
* cell instance $7304 r0 *1 68.115,8.05
X$7304 140 VIA_via1_4
* cell instance $7305 r0 *1 66.405,9.17
X$7305 140 VIA_via1_4
* cell instance $7306 r0 *1 66.405,9.17
X$7306 140 VIA_via2_5
* cell instance $7307 r0 *1 70.965,7.35
X$7307 141 VIA_via2_5
* cell instance $7308 r0 *1 73.435,7.35
X$7308 141 VIA_via2_5
* cell instance $7309 r0 *1 73.055,7.35
X$7309 141 VIA_via1_4
* cell instance $7310 r0 *1 73.055,7.35
X$7310 141 VIA_via2_5
* cell instance $7311 r0 *1 70.965,6.37
X$7311 141 VIA_via1_4
* cell instance $7312 r0 *1 73.435,7.63
X$7312 141 VIA_via1_4
* cell instance $7313 r0 *1 74.385,8.19
X$7313 142 VIA_via1_7
* cell instance $7314 r0 *1 74.005,9.17
X$7314 142 VIA_via1_4
* cell instance $7315 r0 *1 78.565,8.19
X$7315 143 VIA_via1_7
* cell instance $7316 r0 *1 78.375,9.17
X$7316 143 VIA_via1_4
* cell instance $7317 r0 *1 83.315,7.77
X$7317 144 VIA_via1_7
* cell instance $7318 r0 *1 68.115,9.03
X$7318 144 VIA_via1_7
* cell instance $7319 r0 *1 68.115,9.03
X$7319 144 VIA_via2_5
* cell instance $7320 r0 *1 30.875,34.23
X$7320 144 VIA_via1_7
* cell instance $7321 r0 *1 30.875,34.23
X$7321 144 VIA_via2_5
* cell instance $7322 r0 *1 80.085,7.77
X$7322 144 VIA_via1_7
* cell instance $7323 r0 *1 83.315,8.05
X$7323 144 VIA_via2_5
* cell instance $7324 r0 *1 80.275,8.05
X$7324 144 VIA_via2_5
* cell instance $7325 r0 *1 80.275,9.03
X$7325 144 VIA_via2_5
* cell instance $7326 r0 *1 67.925,11.55
X$7326 144 VIA_via2_5
* cell instance $7327 r0 *1 37.715,35.35
X$7327 144 VIA_via2_5
* cell instance $7328 r0 *1 41.325,35.35
X$7328 144 VIA_via2_5
* cell instance $7329 r0 *1 47.215,27.37
X$7329 144 VIA_via2_5
* cell instance $7330 r0 *1 47.215,11.55
X$7330 144 VIA_via2_5
* cell instance $7331 r0 *1 33.915,35.35
X$7331 144 VIA_via2_5
* cell instance $7332 r0 *1 57.285,35.21
X$7332 144 VIA_via2_5
* cell instance $7333 r0 *1 51.395,32.83
X$7333 144 VIA_via2_5
* cell instance $7334 r0 *1 51.395,35.07
X$7334 144 VIA_via2_5
* cell instance $7335 r0 *1 57.285,38.43
X$7335 144 VIA_via2_5
* cell instance $7336 r0 *1 60.515,38.43
X$7336 144 VIA_via1_4
* cell instance $7337 r0 *1 60.515,38.43
X$7337 144 VIA_via2_5
* cell instance $7338 r0 *1 56.715,38.43
X$7338 144 VIA_via1_4
* cell instance $7339 r0 *1 56.715,38.43
X$7339 144 VIA_via2_5
* cell instance $7340 r0 *1 51.395,34.37
X$7340 144 VIA_via1_4
* cell instance $7341 r0 *1 33.915,34.37
X$7341 144 VIA_via1_4
* cell instance $7342 r0 *1 33.915,34.23
X$7342 144 VIA_via2_5
* cell instance $7343 r0 *1 47.025,32.83
X$7343 144 VIA_via1_4
* cell instance $7344 r0 *1 47.025,32.83
X$7344 144 VIA_via2_5
* cell instance $7345 r0 *1 37.715,35.63
X$7345 144 VIA_via1_4
* cell instance $7346 r0 *1 41.705,27.37
X$7346 144 VIA_via1_4
* cell instance $7347 r0 *1 41.705,27.37
X$7347 144 VIA_via2_5
* cell instance $7348 r0 *1 41.325,27.65
X$7348 144 VIA_via1_4
* cell instance $7349 r0 *1 85.785,7.63
X$7349 145 VIA_via2_5
* cell instance $7350 r0 *1 82.555,7.63
X$7350 145 VIA_via2_5
* cell instance $7351 r0 *1 84.075,7.63
X$7351 145 VIA_via1_4
* cell instance $7352 r0 *1 84.075,7.63
X$7352 145 VIA_via2_5
* cell instance $7353 r0 *1 82.555,6.37
X$7353 145 VIA_via1_4
* cell instance $7354 r0 *1 85.785,5.25
X$7354 145 VIA_via1_4
* cell instance $7355 r0 *1 89.775,6.23
X$7355 146 VIA_via1_4
* cell instance $7356 r0 *1 88.635,9.17
X$7356 146 VIA_via1_4
* cell instance $7357 r0 *1 9.595,7.63
X$7357 147 VIA_via1_4
* cell instance $7358 r0 *1 9.595,7.49
X$7358 147 VIA_via2_5
* cell instance $7359 r0 *1 13.205,7.49
X$7359 147 VIA_via1_4
* cell instance $7360 r0 *1 13.205,7.49
X$7360 147 VIA_via2_5
* cell instance $7361 r0 *1 12.825,8.05
X$7361 148 VIA_via2_5
* cell instance $7362 r0 *1 11.875,8.05
X$7362 148 VIA_via1_4
* cell instance $7363 r0 *1 11.875,8.05
X$7363 148 VIA_via2_5
* cell instance $7364 r0 *1 12.825,7.63
X$7364 148 VIA_via1_4
* cell instance $7365 r0 *1 12.635,9.17
X$7365 148 VIA_via1_4
* cell instance $7366 r0 *1 16.055,9.17
X$7366 149 VIA_via2_5
* cell instance $7367 r0 *1 16.055,7.63
X$7367 149 VIA_via2_5
* cell instance $7368 r0 *1 33.535,11.97
X$7368 149 VIA_via2_5
* cell instance $7369 r0 *1 33.535,18.83
X$7369 149 VIA_via2_5
* cell instance $7370 r0 *1 37.335,11.97
X$7370 149 VIA_via2_5
* cell instance $7371 r0 *1 37.335,9.31
X$7371 149 VIA_via2_5
* cell instance $7372 r0 *1 15.105,20.51
X$7372 149 VIA_via2_5
* cell instance $7373 r0 *1 23.465,18.83
X$7373 149 VIA_via2_5
* cell instance $7374 r0 *1 24.415,18.83
X$7374 149 VIA_via2_5
* cell instance $7375 r0 *1 6.555,20.37
X$7375 149 VIA_via1_4
* cell instance $7376 r0 *1 6.555,20.37
X$7376 149 VIA_via2_5
* cell instance $7377 r0 *1 10.355,9.17
X$7377 149 VIA_via1_4
* cell instance $7378 r0 *1 10.355,9.17
X$7378 149 VIA_via2_5
* cell instance $7379 r0 *1 16.055,6.37
X$7379 149 VIA_via1_4
* cell instance $7380 r0 *1 23.275,7.63
X$7380 149 VIA_via1_4
* cell instance $7381 r0 *1 23.275,7.63
X$7381 149 VIA_via2_5
* cell instance $7382 r0 *1 45.695,18.83
X$7382 149 VIA_via1_4
* cell instance $7383 r0 *1 45.695,18.83
X$7383 149 VIA_via2_5
* cell instance $7384 r0 *1 32.205,11.97
X$7384 149 VIA_via1_4
* cell instance $7385 r0 *1 32.205,11.97
X$7385 149 VIA_via2_5
* cell instance $7386 r0 *1 26.505,18.83
X$7386 149 VIA_via1_4
* cell instance $7387 r0 *1 26.505,18.83
X$7387 149 VIA_via2_5
* cell instance $7388 r0 *1 33.345,23.17
X$7388 149 VIA_via1_4
* cell instance $7389 r0 *1 37.335,7.63
X$7389 149 VIA_via1_4
* cell instance $7390 r0 *1 46.455,9.17
X$7390 149 VIA_via1_4
* cell instance $7391 r0 *1 46.455,9.31
X$7391 149 VIA_via2_5
* cell instance $7392 r0 *1 15.105,21.63
X$7392 149 VIA_via1_4
* cell instance $7393 r0 *1 24.415,20.37
X$7393 149 VIA_via1_4
* cell instance $7394 r0 *1 24.415,20.51
X$7394 149 VIA_via2_5
* cell instance $7395 r0 *1 80.655,7.63
X$7395 150 VIA_via2_5
* cell instance $7396 r0 *1 77.615,7.63
X$7396 150 VIA_via1_4
* cell instance $7397 r0 *1 77.615,7.63
X$7397 150 VIA_via2_5
* cell instance $7398 r0 *1 80.655,8.75
X$7398 150 VIA_via1_4
* cell instance $7399 r0 *1 80.845,7.63
X$7399 150 VIA_via1_4
* cell instance $7400 r0 *1 80.845,7.63
X$7400 150 VIA_via2_5
* cell instance $7401 r0 *1 71.345,6.79
X$7401 151 VIA_via1_7
* cell instance $7402 r0 *1 71.345,6.79
X$7402 151 VIA_via2_5
* cell instance $7403 r0 *1 70.775,6.79
X$7403 151 VIA_via2_5
* cell instance $7404 r0 *1 70.775,7.63
X$7404 151 VIA_via1_4
* cell instance $7405 r0 *1 69.445,7.21
X$7405 152 VIA_via1_7
* cell instance $7406 r0 *1 69.445,7.21
X$7406 152 VIA_via2_5
* cell instance $7407 r0 *1 66.785,7.21
X$7407 152 VIA_via2_5
* cell instance $7408 r0 *1 66.785,6.37
X$7408 152 VIA_via1_4
* cell instance $7409 r0 *1 67.165,15.61
X$7409 153 VIA_via1_7
* cell instance $7410 r0 *1 67.165,15.61
X$7410 153 VIA_via2_5
* cell instance $7411 r0 *1 67.545,7.63
X$7411 153 VIA_via2_5
* cell instance $7412 r0 *1 68.305,15.61
X$7412 153 VIA_via2_5
* cell instance $7413 r0 *1 62.795,15.61
X$7413 153 VIA_via2_5
* cell instance $7414 r0 *1 63.745,15.61
X$7414 153 VIA_via2_5
* cell instance $7415 r0 *1 62.795,14.77
X$7415 153 VIA_via1_4
* cell instance $7416 r0 *1 63.745,16.03
X$7416 153 VIA_via1_4
* cell instance $7417 r0 *1 68.115,17.57
X$7417 153 VIA_via1_4
* cell instance $7418 r0 *1 68.305,14.77
X$7418 153 VIA_via1_4
* cell instance $7419 r0 *1 67.735,13.23
X$7419 153 VIA_via1_4
* cell instance $7420 r0 *1 67.355,11.97
X$7420 153 VIA_via1_4
* cell instance $7421 r0 *1 71.535,7.63
X$7421 153 VIA_via1_4
* cell instance $7422 r0 *1 71.535,7.63
X$7422 153 VIA_via2_5
* cell instance $7423 r0 *1 4.275,26.95
X$7423 154 VIA_via2_5
* cell instance $7424 r0 *1 7.505,26.95
X$7424 154 VIA_via2_5
* cell instance $7425 r0 *1 13.585,8.47
X$7425 154 VIA_via2_5
* cell instance $7426 r0 *1 2.755,26.95
X$7426 154 VIA_via2_5
* cell instance $7427 r0 *1 11.115,8.47
X$7427 154 VIA_via2_5
* cell instance $7428 r0 *1 12.255,8.47
X$7428 154 VIA_via2_5
* cell instance $7429 r0 *1 9.025,8.47
X$7429 154 VIA_via2_5
* cell instance $7430 r0 *1 14.155,26.95
X$7430 154 VIA_via2_5
* cell instance $7431 r0 *1 11.115,6.37
X$7431 154 VIA_via1_4
* cell instance $7432 r0 *1 9.025,10.43
X$7432 154 VIA_via1_4
* cell instance $7433 r0 *1 12.255,7.63
X$7433 154 VIA_via1_4
* cell instance $7434 r0 *1 13.585,10.43
X$7434 154 VIA_via1_4
* cell instance $7435 r0 *1 7.505,27.23
X$7435 154 VIA_via1_4
* cell instance $7436 r0 *1 2.755,26.25
X$7436 154 VIA_via1_4
* cell instance $7437 r0 *1 4.275,27.23
X$7437 154 VIA_via1_4
* cell instance $7438 r0 *1 14.155,27.23
X$7438 154 VIA_via1_4
* cell instance $7439 r0 *1 33.725,11.83
X$7439 155 VIA_via1_7
* cell instance $7440 r0 *1 44.365,11.83
X$7440 155 VIA_via1_7
* cell instance $7441 r0 *1 13.775,11.83
X$7441 155 VIA_via1_7
* cell instance $7442 r0 *1 14.155,9.03
X$7442 155 VIA_via1_7
* cell instance $7443 r0 *1 14.155,9.03
X$7443 155 VIA_via2_5
* cell instance $7444 r0 *1 51.205,10.15
X$7444 155 VIA_via2_5
* cell instance $7445 r0 *1 13.775,9.03
X$7445 155 VIA_via2_5
* cell instance $7446 r0 *1 13.775,10.43
X$7446 155 VIA_via2_5
* cell instance $7447 r0 *1 33.725,10.71
X$7447 155 VIA_via2_5
* cell instance $7448 r0 *1 40.185,10.15
X$7448 155 VIA_via2_5
* cell instance $7449 r0 *1 44.365,10.15
X$7449 155 VIA_via2_5
* cell instance $7450 r0 *1 28.215,9.31
X$7450 155 VIA_via2_5
* cell instance $7451 r0 *1 21.375,9.31
X$7451 155 VIA_via2_5
* cell instance $7452 r0 *1 21.375,10.43
X$7452 155 VIA_via1_4
* cell instance $7453 r0 *1 22.705,9.17
X$7453 155 VIA_via1_4
* cell instance $7454 r0 *1 22.705,9.31
X$7454 155 VIA_via2_5
* cell instance $7455 r0 *1 13.395,10.43
X$7455 155 VIA_via1_4
* cell instance $7456 r0 *1 13.395,10.43
X$7456 155 VIA_via2_5
* cell instance $7457 r0 *1 28.215,10.43
X$7457 155 VIA_via1_4
* cell instance $7458 r0 *1 28.215,10.29
X$7458 155 VIA_via2_5
* cell instance $7459 r0 *1 40.185,9.17
X$7459 155 VIA_via1_4
* cell instance $7460 r0 *1 51.205,10.43
X$7460 155 VIA_via1_4
* cell instance $7461 r0 *1 54.815,10.29
X$7461 155 VIA_via1_4
* cell instance $7462 r0 *1 54.815,10.29
X$7462 155 VIA_via2_5
* cell instance $7463 r0 *1 15.295,8.61
X$7463 156 VIA_via1_7
* cell instance $7464 r0 *1 15.675,7.63
X$7464 156 VIA_via1_4
* cell instance $7465 r0 *1 39.995,8.75
X$7465 157 VIA_via1_4
* cell instance $7466 r0 *1 40.945,9.17
X$7466 157 VIA_via1_4
* cell instance $7467 r0 *1 40.755,11.97
X$7467 157 VIA_via1_4
* cell instance $7468 r0 *1 56.525,18.41
X$7468 158 VIA_via1_7
* cell instance $7469 r0 *1 52.155,12.67
X$7469 158 VIA_via2_5
* cell instance $7470 r0 *1 56.525,14.63
X$7470 158 VIA_via2_5
* cell instance $7471 r0 *1 55.385,18.83
X$7471 158 VIA_via2_5
* cell instance $7472 r0 *1 51.965,21.63
X$7472 158 VIA_via2_5
* cell instance $7473 r0 *1 55.385,21.63
X$7473 158 VIA_via2_5
* cell instance $7474 r0 *1 55.575,12.67
X$7474 158 VIA_via2_5
* cell instance $7475 r0 *1 56.525,17.57
X$7475 158 VIA_via2_5
* cell instance $7476 r0 *1 60.705,17.57
X$7476 158 VIA_via1_4
* cell instance $7477 r0 *1 60.705,17.57
X$7477 158 VIA_via2_5
* cell instance $7478 r0 *1 52.345,9.17
X$7478 158 VIA_via1_4
* cell instance $7479 r0 *1 55.005,21.63
X$7479 158 VIA_via1_4
* cell instance $7480 r0 *1 55.005,21.63
X$7480 158 VIA_via2_5
* cell instance $7481 r0 *1 51.775,24.43
X$7481 158 VIA_via1_4
* cell instance $7482 r0 *1 55.385,20.37
X$7482 158 VIA_via1_4
* cell instance $7483 r0 *1 56.715,18.83
X$7483 158 VIA_via1_4
* cell instance $7484 r0 *1 56.715,18.83
X$7484 158 VIA_via2_5
* cell instance $7485 r0 *1 55.575,14.77
X$7485 158 VIA_via1_4
* cell instance $7486 r0 *1 55.575,14.63
X$7486 158 VIA_via2_5
* cell instance $7487 r0 *1 58.995,14.77
X$7487 158 VIA_via1_4
* cell instance $7488 r0 *1 58.995,14.77
X$7488 158 VIA_via2_5
* cell instance $7489 r0 *1 94.715,9.17
X$7489 159 VIA_via2_5
* cell instance $7490 r0 *1 94.715,8.05
X$7490 159 VIA_via1_4
* cell instance $7491 r0 *1 92.815,9.17
X$7491 159 VIA_via1_4
* cell instance $7492 r0 *1 92.815,9.17
X$7492 159 VIA_via2_5
* cell instance $7493 r0 *1 90.915,9.17
X$7493 159 VIA_via1_4
* cell instance $7494 r0 *1 90.915,9.17
X$7494 159 VIA_via2_5
* cell instance $7495 r0 *1 96.045,11.97
X$7495 160 VIA_via1_4
* cell instance $7496 r0 *1 96.045,11.97
X$7496 160 VIA_via2_5
* cell instance $7497 r0 *1 97.255,8.47
X$7497 160 VIA_via4_0
* cell instance $7498 r0 *1 97.255,11.97
X$7498 160 VIA_via3_2
* cell instance $7499 r0 *1 93.195,8.61
X$7499 161 VIA_via1_7
* cell instance $7500 r0 *1 93.195,8.61
X$7500 161 VIA_via2_5
* cell instance $7501 r0 *1 92.435,8.61
X$7501 161 VIA_via2_5
* cell instance $7502 r0 *1 92.435,7.63
X$7502 161 VIA_via1_4
* cell instance $7503 r0 *1 84.455,8.19
X$7503 162 VIA_via1_7
* cell instance $7504 r0 *1 87.685,8.61
X$7504 162 VIA_via2_5
* cell instance $7505 r0 *1 84.455,8.61
X$7505 162 VIA_via2_5
* cell instance $7506 r0 *1 87.685,9.17
X$7506 162 VIA_via1_4
* cell instance $7507 r0 *1 67.355,8.61
X$7507 163 VIA_via1_7
* cell instance $7508 r0 *1 67.355,8.61
X$7508 163 VIA_via2_5
* cell instance $7509 r0 *1 65.835,8.61
X$7509 163 VIA_via2_5
* cell instance $7510 r0 *1 65.835,7.63
X$7510 163 VIA_via1_4
* cell instance $7511 r0 *1 50.635,8.61
X$7511 164 VIA_via1_7
* cell instance $7512 r0 *1 50.635,7.63
X$7512 164 VIA_via1_4
* cell instance $7513 r0 *1 26.505,9.03
X$7513 165 VIA_via2_5
* cell instance $7514 r0 *1 26.505,9.45
X$7514 165 VIA_via2_5
* cell instance $7515 r0 *1 23.465,9.17
X$7515 165 VIA_via1_4
* cell instance $7516 r0 *1 23.465,9.03
X$7516 165 VIA_via2_5
* cell instance $7517 r0 *1 27.075,9.45
X$7517 165 VIA_via1_4
* cell instance $7518 r0 *1 27.075,9.45
X$7518 165 VIA_via2_5
* cell instance $7519 r0 *1 26.505,11.97
X$7519 165 VIA_via1_4
* cell instance $7520 r0 *1 16.625,10.01
X$7520 166 VIA_via1_7
* cell instance $7521 r0 *1 16.245,9.17
X$7521 166 VIA_via1_4
* cell instance $7522 r0 *1 22.705,11.83
X$7522 167 VIA_via2_5
* cell instance $7523 r0 *1 20.995,11.97
X$7523 167 VIA_via1_4
* cell instance $7524 r0 *1 20.995,11.83
X$7524 167 VIA_via2_5
* cell instance $7525 r0 *1 22.515,10.29
X$7525 167 VIA_via1_4
* cell instance $7526 r0 *1 25.555,11.41
X$7526 168 VIA_via1_7
* cell instance $7527 r0 *1 25.175,10.43
X$7527 168 VIA_via1_4
* cell instance $7528 r0 *1 31.635,10.43
X$7528 169 VIA_via2_5
* cell instance $7529 r0 *1 32.015,10.43
X$7529 169 VIA_via2_5
* cell instance $7530 r0 *1 31.635,11.97
X$7530 169 VIA_via1_4
* cell instance $7531 r0 *1 32.015,9.45
X$7531 169 VIA_via1_4
* cell instance $7532 r0 *1 28.975,10.43
X$7532 169 VIA_via1_4
* cell instance $7533 r0 *1 28.975,10.43
X$7533 169 VIA_via2_5
* cell instance $7534 r0 *1 35.245,9.17
X$7534 170 VIA_via2_5
* cell instance $7535 r0 *1 35.245,11.97
X$7535 170 VIA_via1_4
* cell instance $7536 r0 *1 36.195,9.17
X$7536 170 VIA_via1_4
* cell instance $7537 r0 *1 36.195,9.17
X$7537 170 VIA_via2_5
* cell instance $7538 r0 *1 35.245,9.45
X$7538 170 VIA_via1_4
* cell instance $7539 r0 *1 29.545,11.83
X$7539 171 VIA_via1_7
* cell instance $7540 r0 *1 29.545,11.69
X$7540 171 VIA_via2_5
* cell instance $7541 r0 *1 38.665,11.83
X$7541 171 VIA_via1_7
* cell instance $7542 r0 *1 18.525,11.83
X$7542 171 VIA_via1_7
* cell instance $7543 r0 *1 18.525,11.69
X$7543 171 VIA_via2_5
* cell instance $7544 r0 *1 24.415,11.83
X$7544 171 VIA_via1_7
* cell instance $7545 r0 *1 24.415,11.69
X$7545 171 VIA_via2_5
* cell instance $7546 r0 *1 51.585,10.29
X$7546 171 VIA_via2_5
* cell instance $7547 r0 *1 49.495,10.29
X$7547 171 VIA_via2_5
* cell instance $7548 r0 *1 15.485,10.85
X$7548 171 VIA_via2_5
* cell instance $7549 r0 *1 18.525,10.85
X$7549 171 VIA_via2_5
* cell instance $7550 r0 *1 38.665,10.29
X$7550 171 VIA_via2_5
* cell instance $7551 r0 *1 35.625,11.69
X$7551 171 VIA_via2_5
* cell instance $7552 r0 *1 35.625,10.29
X$7552 171 VIA_via2_5
* cell instance $7553 r0 *1 29.545,10.71
X$7553 171 VIA_via2_5
* cell instance $7554 r0 *1 8.835,12.25
X$7554 171 VIA_via2_5
* cell instance $7555 r0 *1 9.405,12.25
X$7555 171 VIA_via2_5
* cell instance $7556 r0 *1 24.415,10.71
X$7556 171 VIA_via2_5
* cell instance $7557 r0 *1 8.835,10.85
X$7557 171 VIA_via2_5
* cell instance $7558 r0 *1 8.835,10.43
X$7558 171 VIA_via1_4
* cell instance $7559 r0 *1 9.405,13.23
X$7559 171 VIA_via1_4
* cell instance $7560 r0 *1 15.485,10.43
X$7560 171 VIA_via1_4
* cell instance $7561 r0 *1 35.435,9.17
X$7561 171 VIA_via1_4
* cell instance $7562 r0 *1 42.655,10.43
X$7562 171 VIA_via1_4
* cell instance $7563 r0 *1 42.655,10.29
X$7563 171 VIA_via2_5
* cell instance $7564 r0 *1 49.495,9.17
X$7564 171 VIA_via1_4
* cell instance $7565 r0 *1 51.585,11.55
X$7565 171 VIA_via1_4
* cell instance $7566 r0 *1 43.415,9.45
X$7566 172 VIA_via2_5
* cell instance $7567 r0 *1 43.225,11.97
X$7567 172 VIA_via1_4
* cell instance $7568 r0 *1 43.415,10.43
X$7568 172 VIA_via1_4
* cell instance $7569 r0 *1 44.745,9.45
X$7569 172 VIA_via1_4
* cell instance $7570 r0 *1 44.745,9.45
X$7570 172 VIA_via2_5
* cell instance $7571 r0 *1 56.145,9.45
X$7571 173 VIA_via2_5
* cell instance $7572 r0 *1 61.085,9.45
X$7572 173 VIA_via2_5
* cell instance $7573 r0 *1 61.085,10.43
X$7573 173 VIA_via1_4
* cell instance $7574 r0 *1 58.805,9.45
X$7574 173 VIA_via1_4
* cell instance $7575 r0 *1 58.805,9.45
X$7575 173 VIA_via2_5
* cell instance $7576 r0 *1 56.145,10.43
X$7576 173 VIA_via1_4
* cell instance $7577 r0 *1 87.685,67.83
X$7577 174 VIA_via1_7
* cell instance $7578 r0 *1 64.695,60.97
X$7578 174 VIA_via1_7
* cell instance $7579 r0 *1 64.775,60.83
X$7579 174 VIA_via3_2
* cell instance $7580 r0 *1 64.695,60.83
X$7580 174 VIA_via2_5
* cell instance $7581 r0 *1 89.015,21.77
X$7581 174 VIA_via1_7
* cell instance $7582 r0 *1 78.375,30.17
X$7582 174 VIA_via1_7
* cell instance $7583 r0 *1 83.885,60.97
X$7583 174 VIA_via1_7
* cell instance $7584 r0 *1 83.885,61.11
X$7584 174 VIA_via2_5
* cell instance $7585 r0 *1 86.355,38.57
X$7585 174 VIA_via1_7
* cell instance $7586 r0 *1 84.645,10.43
X$7586 174 VIA_via2_5
* cell instance $7587 r0 *1 82.175,9.87
X$7587 174 VIA_via2_5
* cell instance $7588 r0 *1 69.255,10.15
X$7588 174 VIA_via2_5
* cell instance $7589 r0 *1 87.495,61.11
X$7589 174 VIA_via2_5
* cell instance $7590 r0 *1 69.255,9.87
X$7590 174 VIA_via2_5
* cell instance $7591 r0 *1 84.645,9.87
X$7591 174 VIA_via2_5
* cell instance $7592 r0 *1 86.165,38.71
X$7592 174 VIA_via2_5
* cell instance $7593 r0 *1 78.375,31.15
X$7593 174 VIA_via2_5
* cell instance $7594 r0 *1 89.015,32.41
X$7594 174 VIA_via2_5
* cell instance $7595 r0 *1 85.595,32.41
X$7595 174 VIA_via2_5
* cell instance $7596 r0 *1 78.375,30.73
X$7596 174 VIA_via2_5
* cell instance $7597 r0 *1 85.595,30.73
X$7597 174 VIA_via2_5
* cell instance $7598 r0 *1 85.595,32.83
X$7598 174 VIA_via1_4
* cell instance $7599 r0 *1 84.265,10.43
X$7599 174 VIA_via1_4
* cell instance $7600 r0 *1 84.265,10.43
X$7600 174 VIA_via2_5
* cell instance $7601 r0 *1 82.365,10.43
X$7601 174 VIA_via1_4
* cell instance $7602 r0 *1 63.935,36.75
X$7602 174 VIA_via1_4
* cell instance $7603 r0 *1 63.935,36.75
X$7603 174 VIA_via2_5
* cell instance $7604 r0 *1 62.985,10.43
X$7604 174 VIA_via1_4
* cell instance $7605 r0 *1 62.985,10.43
X$7605 174 VIA_via2_5
* cell instance $7606 r0 *1 64.775,10.43
X$7606 174 VIA_via3_2
* cell instance $7607 r0 *1 64.775,31.15
X$7607 174 VIA_via3_2
* cell instance $7608 r0 *1 86.335,32.41
X$7608 174 VIA_via3_2
* cell instance $7609 r0 *1 64.775,36.75
X$7609 174 VIA_via3_2
* cell instance $7610 r0 *1 86.335,38.71
X$7610 174 VIA_via3_2
* cell instance $7611 r0 *1 64.775,61.11
X$7611 174 VIA_via3_2
* cell instance $7612 r0 *1 74.195,9.59
X$7612 175 VIA_via1_7
* cell instance $7613 r0 *1 74.195,13.23
X$7613 175 VIA_via1_4
* cell instance $7614 r0 *1 78.565,10.29
X$7614 176 VIA_via1_4
* cell instance $7615 r0 *1 78.565,10.29
X$7615 176 VIA_via2_5
* cell instance $7616 r0 *1 74.955,10.43
X$7616 176 VIA_via1_4
* cell instance $7617 r0 *1 74.955,10.29
X$7617 176 VIA_via2_5
* cell instance $7618 r0 *1 75.145,13.23
X$7618 176 VIA_via1_4
* cell instance $7619 r0 *1 91.865,10.15
X$7619 177 VIA_via2_5
* cell instance $7620 r0 *1 89.015,10.15
X$7620 177 VIA_via2_5
* cell instance $7621 r0 *1 74.385,9.45
X$7621 177 VIA_via2_5
* cell instance $7622 r0 *1 74.005,56.35
X$7622 177 VIA_via2_5
* cell instance $7623 r0 *1 85.595,57.05
X$7623 177 VIA_via2_5
* cell instance $7624 r0 *1 78.565,57.05
X$7624 177 VIA_via2_5
* cell instance $7625 r0 *1 74.765,33.25
X$7625 177 VIA_via2_5
* cell instance $7626 r0 *1 92.815,33.25
X$7626 177 VIA_via2_5
* cell instance $7627 r0 *1 74.385,9.17
X$7627 177 VIA_via1_4
* cell instance $7628 r0 *1 92.625,37.17
X$7628 177 VIA_via1_4
* cell instance $7629 r0 *1 91.865,10.43
X$7629 177 VIA_via1_4
* cell instance $7630 r0 *1 89.015,9.17
X$7630 177 VIA_via1_4
* cell instance $7631 r0 *1 89.015,9.31
X$7631 177 VIA_via2_5
* cell instance $7632 r0 *1 92.815,32.83
X$7632 177 VIA_via1_4
* cell instance $7633 r0 *1 92.815,23.17
X$7633 177 VIA_via1_4
* cell instance $7634 r0 *1 70.585,56.77
X$7634 177 VIA_via1_4
* cell instance $7635 r0 *1 70.585,56.77
X$7635 177 VIA_via2_5
* cell instance $7636 r0 *1 73.245,32.83
X$7636 177 VIA_via1_4
* cell instance $7637 r0 *1 73.245,32.97
X$7637 177 VIA_via2_5
* cell instance $7638 r0 *1 74.765,53.55
X$7638 177 VIA_via1_4
* cell instance $7639 r0 *1 74.385,54.25
X$7639 177 VIA_via1_4
* cell instance $7640 r0 *1 78.565,56.77
X$7640 177 VIA_via1_4
* cell instance $7641 r0 *1 78.565,56.77
X$7641 177 VIA_via2_5
* cell instance $7642 r0 *1 85.595,55.23
X$7642 177 VIA_via1_4
* cell instance $7643 r0 *1 74.855,32.97
X$7643 177 VIA_via3_2
* cell instance $7644 r0 *1 74.765,32.97
X$7644 177 VIA_via2_5
* cell instance $7645 r0 *1 74.855,9.45
X$7645 177 VIA_via3_2
* cell instance $7646 r0 *1 84.265,10.15
X$7646 178 VIA_via2_5
* cell instance $7647 r0 *1 84.265,9.45
X$7647 178 VIA_via1_4
* cell instance $7648 r0 *1 82.555,10.43
X$7648 178 VIA_via1_4
* cell instance $7649 r0 *1 82.555,10.29
X$7649 178 VIA_via2_5
* cell instance $7650 r0 *1 82.745,11.97
X$7650 178 VIA_via1_4
* cell instance $7651 r0 *1 85.405,10.01
X$7651 179 VIA_via1_7
* cell instance $7652 r0 *1 85.215,9.17
X$7652 179 VIA_via1_4
* cell instance $7653 r0 *1 89.585,9.45
X$7653 180 VIA_via2_5
* cell instance $7654 r0 *1 84.455,9.45
X$7654 180 VIA_via2_5
* cell instance $7655 r0 *1 87.495,9.45
X$7655 180 VIA_via1_4
* cell instance $7656 r0 *1 87.495,9.45
X$7656 180 VIA_via2_5
* cell instance $7657 r0 *1 89.585,10.43
X$7657 180 VIA_via1_4
* cell instance $7658 r0 *1 84.455,10.43
X$7658 180 VIA_via1_4
* cell instance $7659 r0 *1 87.875,9.59
X$7659 181 VIA_via1_7
* cell instance $7660 r0 *1 88.065,11.97
X$7660 181 VIA_via1_4
* cell instance $7661 r0 *1 88.825,9.59
X$7661 182 VIA_via1_7
* cell instance $7662 r0 *1 88.825,11.97
X$7662 182 VIA_via1_4
* cell instance $7663 r0 *1 85.975,10.57
X$7663 183 VIA_via2_5
* cell instance $7664 r0 *1 85.975,11.97
X$7664 183 VIA_via1_4
* cell instance $7665 r0 *1 88.635,10.43
X$7665 183 VIA_via1_4
* cell instance $7666 r0 *1 88.635,10.43
X$7666 183 VIA_via2_5
* cell instance $7667 r0 *1 89.015,10.43
X$7667 183 VIA_via1_4
* cell instance $7668 r0 *1 89.015,10.57
X$7668 183 VIA_via2_5
* cell instance $7669 r0 *1 91.865,9.59
X$7669 184 VIA_via1_7
* cell instance $7670 r0 *1 91.485,10.43
X$7670 184 VIA_via1_4
* cell instance $7671 r0 *1 93.955,10.57
X$7671 185 VIA_via2_5
* cell instance $7672 r0 *1 93.955,13.23
X$7672 185 VIA_via1_4
* cell instance $7673 r0 *1 96.615,10.43
X$7673 185 VIA_via1_4
* cell instance $7674 r0 *1 96.615,10.43
X$7674 185 VIA_via2_5
* cell instance $7675 r0 *1 93.005,10.43
X$7675 185 VIA_via1_4
* cell instance $7676 r0 *1 93.005,10.43
X$7676 185 VIA_via2_5
* cell instance $7677 r0 *1 94.335,10.15
X$7677 186 VIA_via2_5
* cell instance $7678 r0 *1 93.385,10.15
X$7678 186 VIA_via1_4
* cell instance $7679 r0 *1 93.385,10.15
X$7679 186 VIA_via2_5
* cell instance $7680 r0 *1 94.335,10.43
X$7680 186 VIA_via1_4
* cell instance $7681 r0 *1 66.975,51.03
X$7681 187 VIA_via1_7
* cell instance $7682 r0 *1 94.905,16.17
X$7682 187 VIA_via1_7
* cell instance $7683 r0 *1 94.335,44.17
X$7683 187 VIA_via1_7
* cell instance $7684 r0 *1 94.335,44.31
X$7684 187 VIA_via2_5
* cell instance $7685 r0 *1 89.205,10.01
X$7685 187 VIA_via2_5
* cell instance $7686 r0 *1 92.245,10.01
X$7686 187 VIA_via2_5
* cell instance $7687 r0 *1 89.205,15.75
X$7687 187 VIA_via2_5
* cell instance $7688 r0 *1 88.445,15.75
X$7688 187 VIA_via2_5
* cell instance $7689 r0 *1 94.525,16.17
X$7689 187 VIA_via2_5
* cell instance $7690 r0 *1 74.195,10.01
X$7690 187 VIA_via2_5
* cell instance $7691 r0 *1 92.815,44.17
X$7691 187 VIA_via2_5
* cell instance $7692 r0 *1 80.085,45.71
X$7692 187 VIA_via2_5
* cell instance $7693 r0 *1 80.085,48.51
X$7693 187 VIA_via2_5
* cell instance $7694 r0 *1 87.495,44.45
X$7694 187 VIA_via2_5
* cell instance $7695 r0 *1 94.525,26.95
X$7695 187 VIA_via2_5
* cell instance $7696 r0 *1 66.975,48.65
X$7696 187 VIA_via2_5
* cell instance $7697 r0 *1 95.475,26.95
X$7697 187 VIA_via2_5
* cell instance $7698 r0 *1 88.445,16.03
X$7698 187 VIA_via1_4
* cell instance $7699 r0 *1 93.195,39.97
X$7699 187 VIA_via1_4
* cell instance $7700 r0 *1 95.475,27.23
X$7700 187 VIA_via1_4
* cell instance $7701 r0 *1 92.245,10.43
X$7701 187 VIA_via1_4
* cell instance $7702 r0 *1 66.785,48.65
X$7702 187 VIA_via1_4
* cell instance $7703 r0 *1 66.785,48.65
X$7703 187 VIA_via2_5
* cell instance $7704 r0 *1 74.195,10.43
X$7704 187 VIA_via1_4
* cell instance $7705 r0 *1 85.405,30.03
X$7705 187 VIA_via1_4
* cell instance $7706 r0 *1 85.405,29.89
X$7706 187 VIA_via2_5
* cell instance $7707 r0 *1 87.495,45.57
X$7707 187 VIA_via1_4
* cell instance $7708 r0 *1 87.495,45.57
X$7708 187 VIA_via2_5
* cell instance $7709 r0 *1 87.735,26.95
X$7709 187 VIA_via3_2
* cell instance $7710 r0 *1 87.735,29.89
X$7710 187 VIA_via3_2
* cell instance $7711 r0 *1 87.735,44.45
X$7711 187 VIA_via3_2
* cell instance $7712 r0 *1 86.925,62.23
X$7712 188 VIA_via1_7
* cell instance $7713 r0 *1 52.915,55.37
X$7713 188 VIA_via1_7
* cell instance $7714 r0 *1 89.585,38.57
X$7714 188 VIA_via1_7
* cell instance $7715 r0 *1 63.365,11.83
X$7715 188 VIA_via1_7
* cell instance $7716 r0 *1 63.365,11.69
X$7716 188 VIA_via2_5
* cell instance $7717 r0 *1 64.125,62.23
X$7717 188 VIA_via1_7
* cell instance $7718 r0 *1 64.125,62.23
X$7718 188 VIA_via2_5
* cell instance $7719 r0 *1 89.395,12.11
X$7719 188 VIA_via2_5
* cell instance $7720 r0 *1 89.395,10.29
X$7720 188 VIA_via2_5
* cell instance $7721 r0 *1 60.515,62.23
X$7721 188 VIA_via2_5
* cell instance $7722 r0 *1 60.515,58.87
X$7722 188 VIA_via2_5
* cell instance $7723 r0 *1 53.295,58.87
X$7723 188 VIA_via2_5
* cell instance $7724 r0 *1 65.075,61.53
X$7724 188 VIA_via2_5
* cell instance $7725 r0 *1 65.075,62.23
X$7725 188 VIA_via2_5
* cell instance $7726 r0 *1 88.065,61.81
X$7726 188 VIA_via2_5
* cell instance $7727 r0 *1 87.305,61.81
X$7727 188 VIA_via2_5
* cell instance $7728 r0 *1 87.685,62.93
X$7728 188 VIA_via2_5
* cell instance $7729 r0 *1 87.305,62.93
X$7729 188 VIA_via2_5
* cell instance $7730 r0 *1 87.685,48.23
X$7730 188 VIA_via2_5
* cell instance $7731 r0 *1 88.065,48.09
X$7731 188 VIA_via2_5
* cell instance $7732 r0 *1 89.585,42.07
X$7732 188 VIA_via2_5
* cell instance $7733 r0 *1 88.065,42.07
X$7733 188 VIA_via2_5
* cell instance $7734 r0 *1 81.985,11.97
X$7734 188 VIA_via1_4
* cell instance $7735 r0 *1 81.985,12.11
X$7735 188 VIA_via2_5
* cell instance $7736 r0 *1 88.825,10.43
X$7736 188 VIA_via1_4
* cell instance $7737 r0 *1 88.825,10.29
X$7737 188 VIA_via2_5
* cell instance $7738 r0 *1 89.775,34.37
X$7738 188 VIA_via1_4
* cell instance $7739 r0 *1 87.495,66.43
X$7739 188 VIA_via1_4
* cell instance $7740 r0 *1 89.205,23.17
X$7740 188 VIA_via1_4
* cell instance $7741 r0 *1 53.295,52.85
X$7741 188 VIA_via1_4
* cell instance $7742 r0 *1 17.005,9.45
X$7742 189 VIA_via2_5
* cell instance $7743 r0 *1 18.525,9.45
X$7743 189 VIA_via1_4
* cell instance $7744 r0 *1 18.525,9.45
X$7744 189 VIA_via2_5
* cell instance $7745 r0 *1 17.005,10.43
X$7745 189 VIA_via1_4
* cell instance $7746 r0 *1 17.005,10.29
X$7746 189 VIA_via2_5
* cell instance $7747 r0 *1 16.245,10.43
X$7747 189 VIA_via1_4
* cell instance $7748 r0 *1 16.245,10.29
X$7748 189 VIA_via2_5
* cell instance $7749 r0 *1 70.965,10.71
X$7749 190 VIA_via2_5
* cell instance $7750 r0 *1 71.345,10.71
X$7750 190 VIA_via2_5
* cell instance $7751 r0 *1 54.055,37.45
X$7751 190 VIA_via2_5
* cell instance $7752 r0 *1 87.685,24.57
X$7752 190 VIA_via2_5
* cell instance $7753 r0 *1 86.545,40.81
X$7753 190 VIA_via2_5
* cell instance $7754 r0 *1 88.065,39.97
X$7754 190 VIA_via2_5
* cell instance $7755 r0 *1 69.635,40.81
X$7755 190 VIA_via2_5
* cell instance $7756 r0 *1 62.985,39.97
X$7756 190 VIA_via2_5
* cell instance $7757 r0 *1 62.985,40.81
X$7757 190 VIA_via2_5
* cell instance $7758 r0 *1 57.855,39.97
X$7758 190 VIA_via1_4
* cell instance $7759 r0 *1 57.855,40.11
X$7759 190 VIA_via2_5
* cell instance $7760 r0 *1 54.055,39.97
X$7760 190 VIA_via1_4
* cell instance $7761 r0 *1 54.055,40.11
X$7761 190 VIA_via2_5
* cell instance $7762 r0 *1 52.535,37.17
X$7762 190 VIA_via1_4
* cell instance $7763 r0 *1 52.535,37.31
X$7763 190 VIA_via2_5
* cell instance $7764 r0 *1 62.605,39.97
X$7764 190 VIA_via1_4
* cell instance $7765 r0 *1 62.605,39.97
X$7765 190 VIA_via2_5
* cell instance $7766 r0 *1 88.065,9.17
X$7766 190 VIA_via1_4
* cell instance $7767 r0 *1 88.065,9.17
X$7767 190 VIA_via2_5
* cell instance $7768 r0 *1 88.015,9.17
X$7768 190 VIA_via3_2
* cell instance $7769 r0 *1 86.545,39.97
X$7769 190 VIA_via1_4
* cell instance $7770 r0 *1 86.545,39.97
X$7770 190 VIA_via2_5
* cell instance $7771 r0 *1 84.075,10.43
X$7771 190 VIA_via1_4
* cell instance $7772 r0 *1 84.075,10.29
X$7772 190 VIA_via2_5
* cell instance $7773 r0 *1 48.355,37.17
X$7773 190 VIA_via1_4
* cell instance $7774 r0 *1 48.355,37.31
X$7774 190 VIA_via2_5
* cell instance $7775 r0 *1 86.925,24.43
X$7775 190 VIA_via1_4
* cell instance $7776 r0 *1 86.925,24.57
X$7776 190 VIA_via2_5
* cell instance $7777 r0 *1 70.965,10.43
X$7777 190 VIA_via1_4
* cell instance $7778 r0 *1 69.825,31.57
X$7778 190 VIA_via1_4
* cell instance $7779 r0 *1 88.015,24.57
X$7779 190 VIA_via3_2
* cell instance $7780 r0 *1 88.015,10.29
X$7780 190 VIA_via3_2
* cell instance $7781 r0 *1 91.865,41.37
X$7781 191 VIA_via1_7
* cell instance $7782 r0 *1 85.975,14.63
X$7782 191 VIA_via1_7
* cell instance $7783 r0 *1 86.165,45.43
X$7783 191 VIA_via1_7
* cell instance $7784 r0 *1 86.165,45.29
X$7784 191 VIA_via2_5
* cell instance $7785 r0 *1 91.865,13.37
X$7785 191 VIA_via1_7
* cell instance $7786 r0 *1 91.865,13.37
X$7786 191 VIA_via2_5
* cell instance $7787 r0 *1 91.865,14.63
X$7787 191 VIA_via1_7
* cell instance $7788 r0 *1 86.165,9.73
X$7788 191 VIA_via2_5
* cell instance $7789 r0 *1 86.165,13.37
X$7789 191 VIA_via2_5
* cell instance $7790 r0 *1 90.725,13.37
X$7790 191 VIA_via2_5
* cell instance $7791 r0 *1 72.865,9.73
X$7791 191 VIA_via2_5
* cell instance $7792 r0 *1 64.885,50.05
X$7792 191 VIA_via2_5
* cell instance $7793 r0 *1 65.265,50.05
X$7793 191 VIA_via2_5
* cell instance $7794 r0 *1 91.865,43.61
X$7794 191 VIA_via2_5
* cell instance $7795 r0 *1 91.675,43.61
X$7795 191 VIA_via2_5
* cell instance $7796 r0 *1 87.685,45.29
X$7796 191 VIA_via2_5
* cell instance $7797 r0 *1 87.685,43.61
X$7797 191 VIA_via2_5
* cell instance $7798 r0 *1 90.915,30.17
X$7798 191 VIA_via2_5
* cell instance $7799 r0 *1 83.885,30.17
X$7799 191 VIA_via2_5
* cell instance $7800 r0 *1 90.915,27.23
X$7800 191 VIA_via2_5
* cell instance $7801 r0 *1 65.265,45.29
X$7801 191 VIA_via2_5
* cell instance $7802 r0 *1 91.295,27.23
X$7802 191 VIA_via1_4
* cell instance $7803 r0 *1 91.295,27.23
X$7803 191 VIA_via2_5
* cell instance $7804 r0 *1 84.075,30.03
X$7804 191 VIA_via1_4
* cell instance $7805 r0 *1 91.865,44.03
X$7805 191 VIA_via1_4
* cell instance $7806 r0 *1 64.885,52.43
X$7806 191 VIA_via1_4
* cell instance $7807 r0 *1 64.315,50.05
X$7807 191 VIA_via1_4
* cell instance $7808 r0 *1 64.315,50.05
X$7808 191 VIA_via2_5
* cell instance $7809 r0 *1 72.865,10.43
X$7809 191 VIA_via1_4
* cell instance $7810 r0 *1 88.015,30.17
X$7810 191 VIA_via3_2
* cell instance $7811 r0 *1 88.015,43.61
X$7811 191 VIA_via3_2
* cell instance $7812 r0 *1 83.505,10.01
X$7812 192 VIA_via1_7
* cell instance $7813 r0 *1 83.505,9.45
X$7813 192 VIA_via2_5
* cell instance $7814 r0 *1 81.985,9.45
X$7814 192 VIA_via2_5
* cell instance $7815 r0 *1 81.985,9.17
X$7815 192 VIA_via1_4
* cell instance $7816 r0 *1 24.795,9.45
X$7816 193 VIA_via2_5
* cell instance $7817 r0 *1 23.845,9.45
X$7817 193 VIA_via1_4
* cell instance $7818 r0 *1 23.845,9.45
X$7818 193 VIA_via2_5
* cell instance $7819 r0 *1 24.795,9.17
X$7819 193 VIA_via1_4
* cell instance $7820 r0 *1 32.965,9.17
X$7820 194 VIA_via1_4
* cell instance $7821 r0 *1 32.965,9.31
X$7821 194 VIA_via2_5
* cell instance $7822 r0 *1 36.575,9.31
X$7822 194 VIA_via1_4
* cell instance $7823 r0 *1 36.575,9.31
X$7823 194 VIA_via2_5
* cell instance $7824 r0 *1 69.255,9.59
X$7824 195 VIA_via1_7
* cell instance $7825 r0 *1 69.255,9.59
X$7825 195 VIA_via2_5
* cell instance $7826 r0 *1 70.585,9.59
X$7826 195 VIA_via2_5
* cell instance $7827 r0 *1 70.585,10.43
X$7827 195 VIA_via1_4
* cell instance $7828 r0 *1 41.325,9.17
X$7828 196 VIA_via1_4
* cell instance $7829 r0 *1 41.325,9.17
X$7829 196 VIA_via2_5
* cell instance $7830 r0 *1 37.715,9.17
X$7830 196 VIA_via1_4
* cell instance $7831 r0 *1 37.715,9.17
X$7831 196 VIA_via2_5
* cell instance $7832 r0 *1 43.795,10.01
X$7832 197 VIA_via1_7
* cell instance $7833 r0 *1 43.795,9.17
X$7833 197 VIA_via2_5
* cell instance $7834 r0 *1 42.465,9.17
X$7834 197 VIA_via1_4
* cell instance $7835 r0 *1 42.465,9.17
X$7835 197 VIA_via2_5
* cell instance $7836 r0 *1 56.525,10.01
X$7836 198 VIA_via1_7
* cell instance $7837 r0 *1 56.525,9.17
X$7837 198 VIA_via1_4
* cell instance $7838 r0 *1 52.345,10.01
X$7838 199 VIA_via1_7
* cell instance $7839 r0 *1 52.345,10.01
X$7839 199 VIA_via2_5
* cell instance $7840 r0 *1 51.585,10.01
X$7840 199 VIA_via2_5
* cell instance $7841 r0 *1 51.585,9.17
X$7841 199 VIA_via1_4
* cell instance $7842 r0 *1 9.975,10.99
X$7842 200 VIA_via1_7
* cell instance $7843 r0 *1 9.025,11.97
X$7843 200 VIA_via1_4
* cell instance $7844 r0 *1 9.595,10.71
X$7844 201 VIA_via2_5
* cell instance $7845 r0 *1 11.305,10.71
X$7845 201 VIA_via2_5
* cell instance $7846 r0 *1 9.595,10.43
X$7846 201 VIA_via1_4
* cell instance $7847 r0 *1 11.305,11.55
X$7847 201 VIA_via1_4
* cell instance $7848 r0 *1 11.685,11.97
X$7848 201 VIA_via1_4
* cell instance $7849 r0 *1 13.205,10.99
X$7849 202 VIA_via2_5
* cell instance $7850 r0 *1 14.155,10.99
X$7850 202 VIA_via2_5
* cell instance $7851 r0 *1 12.255,10.99
X$7851 202 VIA_via2_5
* cell instance $7852 r0 *1 12.255,11.97
X$7852 202 VIA_via1_4
* cell instance $7853 r0 *1 13.205,10.43
X$7853 202 VIA_via1_4
* cell instance $7854 r0 *1 14.155,10.43
X$7854 202 VIA_via1_4
* cell instance $7855 r0 *1 17.955,10.99
X$7855 203 VIA_via1_7
* cell instance $7856 r0 *1 17.955,14.77
X$7856 203 VIA_via1_4
* cell instance $7857 r0 *1 18.335,5.39
X$7857 204 VIA_via1_7
* cell instance $7858 r0 *1 17.955,13.23
X$7858 204 VIA_via1_4
* cell instance $7859 r0 *1 19.665,11.41
X$7859 205 VIA_via1_7
* cell instance $7860 r0 *1 18.905,10.43
X$7860 205 VIA_via1_4
* cell instance $7861 r0 *1 25.365,11.97
X$7861 206 VIA_via2_5
* cell instance $7862 r0 *1 27.455,11.97
X$7862 206 VIA_via2_5
* cell instance $7863 r0 *1 25.175,11.97
X$7863 206 VIA_via1_4
* cell instance $7864 r0 *1 25.935,11.97
X$7864 206 VIA_via1_4
* cell instance $7865 r0 *1 25.935,11.97
X$7865 206 VIA_via2_5
* cell instance $7866 r0 *1 27.455,10.85
X$7866 206 VIA_via1_4
* cell instance $7867 r0 *1 29.735,9.17
X$7867 207 VIA_via1_4
* cell instance $7868 r0 *1 29.355,10.57
X$7868 207 VIA_via1_4
* cell instance $7869 r0 *1 30.685,11.41
X$7869 208 VIA_via1_7
* cell instance $7870 r0 *1 30.305,10.43
X$7870 208 VIA_via1_4
* cell instance $7871 r0 *1 32.395,11.83
X$7871 209 VIA_via2_5
* cell instance $7872 r0 *1 32.585,10.71
X$7872 209 VIA_via1_4
* cell instance $7873 r0 *1 31.065,11.97
X$7873 209 VIA_via1_4
* cell instance $7874 r0 *1 31.065,11.83
X$7874 209 VIA_via2_5
* cell instance $7875 r0 *1 30.305,11.97
X$7875 209 VIA_via1_4
* cell instance $7876 r0 *1 30.305,11.83
X$7876 209 VIA_via2_5
* cell instance $7877 r0 *1 34.865,11.41
X$7877 210 VIA_via1_7
* cell instance $7878 r0 *1 34.675,10.43
X$7878 210 VIA_via1_4
* cell instance $7879 r0 *1 35.055,6.23
X$7879 211 VIA_via1_4
* cell instance $7880 r0 *1 34.865,16.03
X$7880 211 VIA_via1_4
* cell instance $7881 r0 *1 39.995,11.83
X$7881 212 VIA_via1_7
* cell instance $7882 r0 *1 39.995,11.83
X$7882 212 VIA_via2_5
* cell instance $7883 r0 *1 10.545,51.03
X$7883 212 VIA_via1_7
* cell instance $7884 r0 *1 10.545,51.03
X$7884 212 VIA_via2_5
* cell instance $7885 r0 *1 25.745,13.23
X$7885 212 VIA_via2_5
* cell instance $7886 r0 *1 11.495,12.53
X$7886 212 VIA_via2_5
* cell instance $7887 r0 *1 16.815,13.09
X$7887 212 VIA_via2_5
* cell instance $7888 r0 *1 13.965,12.53
X$7888 212 VIA_via2_5
* cell instance $7889 r0 *1 20.805,13.23
X$7889 212 VIA_via1_4
* cell instance $7890 r0 *1 20.805,13.23
X$7890 212 VIA_via2_5
* cell instance $7891 r0 *1 11.495,11.97
X$7891 212 VIA_via1_4
* cell instance $7892 r0 *1 16.815,10.43
X$7892 212 VIA_via1_4
* cell instance $7893 r0 *1 35.055,11.97
X$7893 212 VIA_via1_4
* cell instance $7894 r0 *1 35.055,12.11
X$7894 212 VIA_via2_5
* cell instance $7895 r0 *1 30.875,11.97
X$7895 212 VIA_via1_4
* cell instance $7896 r0 *1 30.875,12.11
X$7896 212 VIA_via2_5
* cell instance $7897 r0 *1 25.745,11.97
X$7897 212 VIA_via1_4
* cell instance $7898 r0 *1 25.745,12.11
X$7898 212 VIA_via2_5
* cell instance $7899 r0 *1 43.035,11.97
X$7899 212 VIA_via1_4
* cell instance $7900 r0 *1 43.035,11.97
X$7900 212 VIA_via2_5
* cell instance $7901 r0 *1 42.845,48.65
X$7901 212 VIA_via1_4
* cell instance $7902 r0 *1 42.845,48.65
X$7902 212 VIA_via2_5
* cell instance $7903 r0 *1 13.965,13.23
X$7903 212 VIA_via1_4
* cell instance $7904 r0 *1 13.965,13.09
X$7904 212 VIA_via2_5
* cell instance $7905 r0 *1 43.215,51.03
X$7905 212 VIA_via4_0
* cell instance $7906 r0 *1 43.215,48.65
X$7906 212 VIA_via3_2
* cell instance $7907 r0 *1 12.415,51.03
X$7907 212 VIA_via3_2
* cell instance $7908 r0 *1 12.415,51.03
X$7908 212 VIA_via4_0
* cell instance $7909 r0 *1 43.215,11.97
X$7909 212 VIA_via3_2
* cell instance $7910 r0 *1 39.805,11.41
X$7910 213 VIA_via1_7
* cell instance $7911 r0 *1 39.425,10.43
X$7911 213 VIA_via1_4
* cell instance $7912 r0 *1 41.705,11.97
X$7912 214 VIA_via2_5
* cell instance $7913 r0 *1 40.185,11.97
X$7913 214 VIA_via1_4
* cell instance $7914 r0 *1 40.185,11.97
X$7914 214 VIA_via2_5
* cell instance $7915 r0 *1 39.425,11.97
X$7915 214 VIA_via1_4
* cell instance $7916 r0 *1 39.425,11.97
X$7916 214 VIA_via2_5
* cell instance $7917 r0 *1 41.705,10.85
X$7917 214 VIA_via1_4
* cell instance $7918 r0 *1 45.505,11.41
X$7918 215 VIA_via1_7
* cell instance $7919 r0 *1 44.745,10.43
X$7919 215 VIA_via1_4
* cell instance $7920 r0 *1 47.025,11.97
X$7920 216 VIA_via2_5
* cell instance $7921 r0 *1 43.795,11.97
X$7921 216 VIA_via1_4
* cell instance $7922 r0 *1 43.795,11.97
X$7922 216 VIA_via2_5
* cell instance $7923 r0 *1 47.025,10.85
X$7923 216 VIA_via1_4
* cell instance $7924 r0 *1 45.125,11.97
X$7924 216 VIA_via1_4
* cell instance $7925 r0 *1 45.125,11.97
X$7925 216 VIA_via2_5
* cell instance $7926 r0 *1 58.045,11.41
X$7926 217 VIA_via1_7
* cell instance $7927 r0 *1 57.855,10.43
X$7927 217 VIA_via1_4
* cell instance $7928 r0 *1 60.135,11.97
X$7928 218 VIA_via2_5
* cell instance $7929 r0 *1 60.135,10.43
X$7929 218 VIA_via1_4
* cell instance $7930 r0 *1 60.515,10.43
X$7930 218 VIA_via1_4
* cell instance $7931 r0 *1 57.665,11.97
X$7931 218 VIA_via1_4
* cell instance $7932 r0 *1 57.665,11.97
X$7932 218 VIA_via2_5
* cell instance $7933 r0 *1 61.275,11.97
X$7933 219 VIA_via1_4
* cell instance $7934 r0 *1 61.275,11.97
X$7934 219 VIA_via2_5
* cell instance $7935 r0 *1 62.225,11.97
X$7935 219 VIA_via1_4
* cell instance $7936 r0 *1 62.225,11.97
X$7936 219 VIA_via2_5
* cell instance $7937 r0 *1 63.555,11.97
X$7937 219 VIA_via1_4
* cell instance $7938 r0 *1 63.555,11.97
X$7938 219 VIA_via2_5
* cell instance $7939 r0 *1 63.555,10.71
X$7939 220 VIA_via2_5
* cell instance $7940 r0 *1 63.175,10.71
X$7940 220 VIA_via2_5
* cell instance $7941 r0 *1 63.555,9.45
X$7941 220 VIA_via1_4
* cell instance $7942 r0 *1 63.175,10.43
X$7942 220 VIA_via1_4
* cell instance $7943 r0 *1 64.125,11.97
X$7943 220 VIA_via1_4
* cell instance $7944 r0 *1 75.525,12.81
X$7944 221 VIA_via1_7
* cell instance $7945 r0 *1 75.335,11.97
X$7945 221 VIA_via1_4
* cell instance $7946 r0 *1 75.905,13.23
X$7946 222 VIA_via2_5
* cell instance $7947 r0 *1 75.715,11.55
X$7947 222 VIA_via1_4
* cell instance $7948 r0 *1 74.005,13.23
X$7948 222 VIA_via1_4
* cell instance $7949 r0 *1 74.005,13.23
X$7949 222 VIA_via2_5
* cell instance $7950 r0 *1 84.835,59.43
X$7950 223 VIA_via1_7
* cell instance $7951 r0 *1 84.835,59.43
X$7951 223 VIA_via2_5
* cell instance $7952 r0 *1 84.935,59.43
X$7952 223 VIA_via3_2
* cell instance $7953 r0 *1 87.685,38.57
X$7953 223 VIA_via1_7
* cell instance $7954 r0 *1 87.685,38.57
X$7954 223 VIA_via2_5
* cell instance $7955 r0 *1 80.085,11.83
X$7955 223 VIA_via1_7
* cell instance $7956 r0 *1 80.085,11.83
X$7956 223 VIA_via2_5
* cell instance $7957 r0 *1 61.975,40.95
X$7957 223 VIA_via5_0
* cell instance $7958 r0 *1 85.785,11.69
X$7958 223 VIA_via2_5
* cell instance $7959 r0 *1 85.785,23.45
X$7959 223 VIA_via2_5
* cell instance $7960 r0 *1 86.545,23.45
X$7960 223 VIA_via2_5
* cell instance $7961 r0 *1 84.835,23.45
X$7961 223 VIA_via2_5
* cell instance $7962 r0 *1 86.355,67.83
X$7962 223 VIA_via2_5
* cell instance $7963 r0 *1 86.335,67.83
X$7963 223 VIA_via3_2
* cell instance $7964 r0 *1 86.355,67.83
X$7964 223 VIA_via1_7
* cell instance $7965 r0 *1 62.035,12.25
X$7965 223 VIA_via2_5
* cell instance $7966 r0 *1 76.285,29.05
X$7966 223 VIA_via2_5
* cell instance $7967 r0 *1 84.645,29.05
X$7967 223 VIA_via2_5
* cell instance $7968 r0 *1 85.215,38.57
X$7968 223 VIA_via2_5
* cell instance $7969 r0 *1 85.215,34.37
X$7969 223 VIA_via1_4
* cell instance $7970 r0 *1 85.785,11.97
X$7970 223 VIA_via1_4
* cell instance $7971 r0 *1 76.285,28.77
X$7971 223 VIA_via1_4
* cell instance $7972 r0 *1 86.545,23.17
X$7972 223 VIA_via1_4
* cell instance $7973 r0 *1 62.035,11.97
X$7973 223 VIA_via1_4
* cell instance $7974 r0 *1 61.975,63.63
X$7974 223 VIA_via4_0
* cell instance $7975 r0 *1 61.975,63.63
X$7975 223 VIA_via3_2
* cell instance $7976 r0 *1 61.975,63.63
X$7976 223 VIA_via5_0
* cell instance $7977 r0 *1 62.035,63.63
X$7977 223 VIA_via2_5
* cell instance $7978 r0 *1 62.035,63.63
X$7978 223 VIA_via1_4
* cell instance $7979 r0 *1 84.935,40.95
X$7979 223 VIA_via4_0
* cell instance $7980 r0 *1 84.935,38.57
X$7980 223 VIA_via3_2
* cell instance $7981 r0 *1 86.335,59.43
X$7981 223 VIA_via3_2
* cell instance $7982 r0 *1 62.255,12.25
X$7982 223 VIA_via3_2
* cell instance $7983 r0 *1 62.255,40.95
X$7983 223 VIA_via3_2
* cell instance $7984 r0 *1 62.225,40.95
X$7984 223 VIA_via2_5
* cell instance $7985 r0 *1 62.255,40.95
X$7985 223 VIA_via4_0
* cell instance $7986 r0 *1 62.225,40.95
X$7986 223 VIA_via1_4
* cell instance $7987 r0 *1 86.925,11.41
X$7987 224 VIA_via1_7
* cell instance $7988 r0 *1 86.355,10.43
X$7988 224 VIA_via1_4
* cell instance $7989 r0 *1 73.815,13.51
X$7989 225 VIA_via2_5
* cell instance $7990 r0 *1 55.575,65.45
X$7990 225 VIA_via2_5
* cell instance $7991 r0 *1 90.915,12.67
X$7991 225 VIA_via2_5
* cell instance $7992 r0 *1 88.255,13.51
X$7992 225 VIA_via2_5
* cell instance $7993 r0 *1 88.255,12.67
X$7993 225 VIA_via2_5
* cell instance $7994 r0 *1 90.915,14.07
X$7994 225 VIA_via2_5
* cell instance $7995 r0 *1 67.165,60.41
X$7995 225 VIA_via2_5
* cell instance $7996 r0 *1 67.165,59.85
X$7996 225 VIA_via2_5
* cell instance $7997 r0 *1 61.465,50.33
X$7997 225 VIA_via2_5
* cell instance $7998 r0 *1 92.245,14.07
X$7998 225 VIA_via2_5
* cell instance $7999 r0 *1 89.205,60.55
X$7999 225 VIA_via2_5
* cell instance $8000 r0 *1 88.635,59.85
X$8000 225 VIA_via2_5
* cell instance $8001 r0 *1 88.635,60.55
X$8001 225 VIA_via2_5
* cell instance $8002 r0 *1 89.015,49.63
X$8002 225 VIA_via2_5
* cell instance $8003 r0 *1 88.635,49.63
X$8003 225 VIA_via2_5
* cell instance $8004 r0 *1 89.015,42.21
X$8004 225 VIA_via2_5
* cell instance $8005 r0 *1 91.865,24.99
X$8005 225 VIA_via2_5
* cell instance $8006 r0 *1 91.865,28.07
X$8006 225 VIA_via2_5
* cell instance $8007 r0 *1 91.295,28.07
X$8007 225 VIA_via2_5
* cell instance $8008 r0 *1 91.295,31.57
X$8008 225 VIA_via1_4
* cell instance $8009 r0 *1 91.295,31.57
X$8009 225 VIA_via2_5
* cell instance $8010 r0 *1 88.445,11.97
X$8010 225 VIA_via1_4
* cell instance $8011 r0 *1 61.275,47.25
X$8011 225 VIA_via1_4
* cell instance $8012 r0 *1 90.915,11.97
X$8012 225 VIA_via1_4
* cell instance $8013 r0 *1 91.675,38.43
X$8013 225 VIA_via1_4
* cell instance $8014 r0 *1 91.675,38.57
X$8014 225 VIA_via2_5
* cell instance $8015 r0 *1 91.655,38.57
X$8015 225 VIA_via3_2
* cell instance $8016 r0 *1 73.815,13.23
X$8016 225 VIA_via1_4
* cell instance $8017 r0 *1 89.585,62.37
X$8017 225 VIA_via1_4
* cell instance $8018 r0 *1 55.575,65.17
X$8018 225 VIA_via1_4
* cell instance $8019 r0 *1 67.165,60.83
X$8019 225 VIA_via1_4
* cell instance $8020 r0 *1 92.055,24.43
X$8020 225 VIA_via1_4
* cell instance $8021 r0 *1 92.055,24.43
X$8021 225 VIA_via2_5
* cell instance $8022 r0 *1 89.205,60.83
X$8022 225 VIA_via1_4
* cell instance $8023 r0 *1 62.535,60.55
X$8023 225 VIA_via3_2
* cell instance $8024 r0 *1 62.535,50.33
X$8024 225 VIA_via3_2
* cell instance $8025 r0 *1 91.095,38.57
X$8025 225 VIA_via3_2
* cell instance $8026 r0 *1 91.095,42.21
X$8026 225 VIA_via3_2
* cell instance $8027 r0 *1 91.655,31.57
X$8027 225 VIA_via3_2
* cell instance $8028 r0 *1 62.815,65.45
X$8028 225 VIA_via3_2
* cell instance $8029 r0 *1 89.965,10.99
X$8029 226 VIA_via1_7
* cell instance $8030 r0 *1 89.585,11.97
X$8030 226 VIA_via1_4
* cell instance $8031 r0 *1 66.405,60.27
X$8031 227 VIA_via2_5
* cell instance $8032 r0 *1 68.305,60.27
X$8032 227 VIA_via2_5
* cell instance $8033 r0 *1 88.445,60.41
X$8033 227 VIA_via2_5
* cell instance $8034 r0 *1 71.915,33.81
X$8034 227 VIA_via2_5
* cell instance $8035 r0 *1 90.535,31.85
X$8035 227 VIA_via2_5
* cell instance $8036 r0 *1 79.135,35.21
X$8036 227 VIA_via2_5
* cell instance $8037 r0 *1 79.135,35.63
X$8037 227 VIA_via1_4
* cell instance $8038 r0 *1 79.135,35.49
X$8038 227 VIA_via2_5
* cell instance $8039 r0 *1 87.685,11.97
X$8039 227 VIA_via1_4
* cell instance $8040 r0 *1 87.685,11.97
X$8040 227 VIA_via2_5
* cell instance $8041 r0 *1 90.155,11.97
X$8041 227 VIA_via1_4
* cell instance $8042 r0 *1 90.155,11.97
X$8042 227 VIA_via2_5
* cell instance $8043 r0 *1 90.535,31.57
X$8043 227 VIA_via1_4
* cell instance $8044 r0 *1 90.915,38.43
X$8044 227 VIA_via1_4
* cell instance $8045 r0 *1 90.915,38.29
X$8045 227 VIA_via2_5
* cell instance $8046 r0 *1 73.055,13.23
X$8046 227 VIA_via1_4
* cell instance $8047 r0 *1 88.825,62.37
X$8047 227 VIA_via1_4
* cell instance $8048 r0 *1 69.065,49.35
X$8048 227 VIA_via1_4
* cell instance $8049 r0 *1 69.065,49.35
X$8049 227 VIA_via2_5
* cell instance $8050 r0 *1 68.685,50.05
X$8050 227 VIA_via1_4
* cell instance $8051 r0 *1 91.295,24.43
X$8051 227 VIA_via1_4
* cell instance $8052 r0 *1 91.295,24.29
X$8052 227 VIA_via2_5
* cell instance $8053 r0 *1 66.405,60.83
X$8053 227 VIA_via1_4
* cell instance $8054 r0 *1 88.445,60.83
X$8054 227 VIA_via1_4
* cell instance $8055 r0 *1 72.335,49.35
X$8055 227 VIA_via3_2
* cell instance $8056 r0 *1 91.095,31.85
X$8056 227 VIA_via3_2
* cell instance $8057 r0 *1 91.095,35.49
X$8057 227 VIA_via3_2
* cell instance $8058 r0 *1 72.335,35.21
X$8058 227 VIA_via3_2
* cell instance $8059 r0 *1 72.335,33.81
X$8059 227 VIA_via3_2
* cell instance $8060 r0 *1 91.095,24.29
X$8060 227 VIA_via3_2
* cell instance $8061 r0 *1 91.095,38.29
X$8061 227 VIA_via3_2
* cell instance $8062 r0 *1 91.095,11.97
X$8062 227 VIA_via3_2
* cell instance $8063 r0 *1 90.345,11.97
X$8063 228 VIA_via1_4
* cell instance $8064 r0 *1 89.965,11.55
X$8064 228 VIA_via1_4
* cell instance $8065 r0 *1 91.295,11.97
X$8065 229 VIA_via1_4
* cell instance $8066 r0 *1 91.675,10.71
X$8066 229 VIA_via1_4
* cell instance $8067 r0 *1 10.925,10.43
X$8067 230 VIA_via1_4
* cell instance $8068 r0 *1 10.925,10.57
X$8068 230 VIA_via2_5
* cell instance $8069 r0 *1 14.535,10.57
X$8069 230 VIA_via1_4
* cell instance $8070 r0 *1 14.535,10.57
X$8070 230 VIA_via2_5
* cell instance $8071 r0 *1 84.075,10.99
X$8071 231 VIA_via1_7
* cell instance $8072 r0 *1 84.075,10.99
X$8072 231 VIA_via2_5
* cell instance $8073 r0 *1 90.535,10.99
X$8073 231 VIA_via2_5
* cell instance $8074 r0 *1 90.535,11.97
X$8074 231 VIA_via1_4
* cell instance $8075 r0 *1 85.025,11.83
X$8075 232 VIA_via1_4
* cell instance $8076 r0 *1 85.025,11.83
X$8076 232 VIA_via2_5
* cell instance $8077 r0 *1 87.875,11.97
X$8077 232 VIA_via1_4
* cell instance $8078 r0 *1 87.875,11.83
X$8078 232 VIA_via2_5
* cell instance $8079 r0 *1 81.225,8.19
X$8079 233 VIA_via1_7
* cell instance $8080 r0 *1 81.225,10.43
X$8080 233 VIA_via2_5
* cell instance $8081 r0 *1 83.695,10.43
X$8081 233 VIA_via1_4
* cell instance $8082 r0 *1 83.695,10.43
X$8082 233 VIA_via2_5
* cell instance $8083 r0 *1 81.225,11.41
X$8083 234 VIA_via1_7
* cell instance $8084 r0 *1 79.895,10.71
X$8084 234 VIA_via2_5
* cell instance $8085 r0 *1 81.225,10.71
X$8085 234 VIA_via2_5
* cell instance $8086 r0 *1 79.895,10.43
X$8086 234 VIA_via1_4
* cell instance $8087 r0 *1 35.815,10.85
X$8087 235 VIA_via2_5
* cell instance $8088 r0 *1 35.815,11.97
X$8088 235 VIA_via1_4
* cell instance $8089 r0 *1 35.815,11.83
X$8089 235 VIA_via2_5
* cell instance $8090 r0 *1 34.485,11.97
X$8090 235 VIA_via1_4
* cell instance $8091 r0 *1 34.485,11.83
X$8091 235 VIA_via2_5
* cell instance $8092 r0 *1 36.955,10.85
X$8092 235 VIA_via1_4
* cell instance $8093 r0 *1 36.955,10.85
X$8093 235 VIA_via2_5
* cell instance $8094 r0 *1 75.335,10.57
X$8094 236 VIA_via1_4
* cell instance $8095 r0 *1 75.335,10.57
X$8095 236 VIA_via2_5
* cell instance $8096 r0 *1 76.285,10.43
X$8096 236 VIA_via1_4
* cell instance $8097 r0 *1 76.285,10.57
X$8097 236 VIA_via2_5
* cell instance $8098 r0 *1 74.575,11.55
X$8098 237 VIA_via2_5
* cell instance $8099 r0 *1 73.625,11.55
X$8099 237 VIA_via2_5
* cell instance $8100 r0 *1 75.145,11.55
X$8100 237 VIA_via1_4
* cell instance $8101 r0 *1 75.145,11.55
X$8101 237 VIA_via2_5
* cell instance $8102 r0 *1 73.625,10.43
X$8102 237 VIA_via1_4
* cell instance $8103 r0 *1 74.575,13.23
X$8103 237 VIA_via1_4
* cell instance $8104 r0 *1 74.005,10.99
X$8104 238 VIA_via1_7
* cell instance $8105 r0 *1 74.005,10.99
X$8105 238 VIA_via2_5
* cell instance $8106 r0 *1 72.865,10.99
X$8106 238 VIA_via2_5
* cell instance $8107 r0 *1 72.865,11.97
X$8107 238 VIA_via1_4
* cell instance $8108 r0 *1 73.245,11.55
X$8108 239 VIA_via2_5
* cell instance $8109 r0 *1 73.245,13.23
X$8109 239 VIA_via1_4
* cell instance $8110 r0 *1 70.205,11.55
X$8110 239 VIA_via1_4
* cell instance $8111 r0 *1 70.205,11.55
X$8111 239 VIA_via2_5
* cell instance $8112 r0 *1 84.645,70.63
X$8112 240 VIA_via1_7
* cell instance $8113 r0 *1 69.825,13.37
X$8113 240 VIA_via1_7
* cell instance $8114 r0 *1 69.825,13.37
X$8114 240 VIA_via2_5
* cell instance $8115 r0 *1 79.895,13.37
X$8115 240 VIA_via1_7
* cell instance $8116 r0 *1 79.895,13.37
X$8116 240 VIA_via2_5
* cell instance $8117 r0 *1 82.175,20.23
X$8117 240 VIA_via1_7
* cell instance $8118 r0 *1 82.175,13.37
X$8118 240 VIA_via2_5
* cell instance $8119 r0 *1 70.395,69.79
X$8119 240 VIA_via2_5
* cell instance $8120 r0 *1 79.325,60.27
X$8120 240 VIA_via2_5
* cell instance $8121 r0 *1 84.265,60.27
X$8121 240 VIA_via2_5
* cell instance $8122 r0 *1 82.745,43.89
X$8122 240 VIA_via2_5
* cell instance $8123 r0 *1 83.505,29.61
X$8123 240 VIA_via2_5
* cell instance $8124 r0 *1 82.555,29.61
X$8124 240 VIA_via2_5
* cell instance $8125 r0 *1 82.745,32.97
X$8125 240 VIA_via2_5
* cell instance $8126 r0 *1 82.555,33.81
X$8126 240 VIA_via2_5
* cell instance $8127 r0 *1 70.395,70.7
X$8127 240 VIA_via1_4
* cell instance $8128 r0 *1 83.505,32.83
X$8128 240 VIA_via1_4
* cell instance $8129 r0 *1 83.505,32.97
X$8129 240 VIA_via2_5
* cell instance $8130 r0 *1 83.505,44.03
X$8130 240 VIA_via1_4
* cell instance $8131 r0 *1 83.535,43.89
X$8131 240 VIA_via3_2
* cell instance $8132 r0 *1 83.505,43.89
X$8132 240 VIA_via2_5
* cell instance $8133 r0 *1 70.775,39.97
X$8133 240 VIA_via1_4
* cell instance $8134 r0 *1 70.775,39.97
X$8134 240 VIA_via2_5
* cell instance $8135 r0 *1 70.655,39.97
X$8135 240 VIA_via3_2
* cell instance $8136 r0 *1 68.115,10.43
X$8136 240 VIA_via1_4
* cell instance $8137 r0 *1 68.115,10.43
X$8137 240 VIA_via2_5
* cell instance $8138 r0 *1 79.325,59.57
X$8138 240 VIA_via1_4
* cell instance $8139 r0 *1 69.825,33.95
X$8139 240 VIA_via1_4
* cell instance $8140 r0 *1 69.825,33.95
X$8140 240 VIA_via2_5
* cell instance $8141 r0 *1 70.655,10.43
X$8141 240 VIA_via3_2
* cell instance $8142 r0 *1 70.655,69.79
X$8142 240 VIA_via3_2
* cell instance $8143 r0 *1 83.535,60.27
X$8143 240 VIA_via3_2
* cell instance $8144 r0 *1 70.655,33.95
X$8144 240 VIA_via3_2
* cell instance $8145 r0 *1 70.655,13.37
X$8145 240 VIA_via3_2
* cell instance $8146 r0 *1 69.255,10.99
X$8146 241 VIA_via1_7
* cell instance $8147 r0 *1 69.255,10.99
X$8147 241 VIA_via2_5
* cell instance $8148 r0 *1 66.595,10.99
X$8148 241 VIA_via2_5
* cell instance $8149 r0 *1 66.595,11.97
X$8149 241 VIA_via1_4
* cell instance $8150 r0 *1 53.865,10.43
X$8150 242 VIA_via1_4
* cell instance $8151 r0 *1 53.865,10.43
X$8151 242 VIA_via2_5
* cell instance $8152 r0 *1 53.865,9.45
X$8152 242 VIA_via1_4
* cell instance $8153 r0 *1 51.965,10.43
X$8153 242 VIA_via1_4
* cell instance $8154 r0 *1 51.965,10.43
X$8154 242 VIA_via2_5
* cell instance $8155 r0 *1 55.955,16.17
X$8155 243 VIA_via1_7
* cell instance $8156 r0 *1 55.955,16.17
X$8156 243 VIA_via2_5
* cell instance $8157 r0 *1 56.095,16.17
X$8157 243 VIA_via3_2
* cell instance $8158 r0 *1 55.385,15.33
X$8158 243 VIA_via2_5
* cell instance $8159 r0 *1 55.955,15.33
X$8159 243 VIA_via2_5
* cell instance $8160 r0 *1 65.835,48.37
X$8160 243 VIA_via1_4
* cell instance $8161 r0 *1 65.835,48.37
X$8161 243 VIA_via2_5
* cell instance $8162 r0 *1 55.385,10.43
X$8162 243 VIA_via1_4
* cell instance $8163 r0 *1 55.385,10.43
X$8163 243 VIA_via2_5
* cell instance $8164 r0 *1 54.435,10.43
X$8164 243 VIA_via1_4
* cell instance $8165 r0 *1 54.435,10.43
X$8165 243 VIA_via2_5
* cell instance $8166 r0 *1 56.905,58.03
X$8166 243 VIA_via1_4
* cell instance $8167 r0 *1 56.905,58.03
X$8167 243 VIA_via2_5
* cell instance $8168 r0 *1 63.555,56.49
X$8168 243 VIA_via1_4
* cell instance $8169 r0 *1 63.555,56.49
X$8169 243 VIA_via2_5
* cell instance $8170 r0 *1 58.615,58.03
X$8170 243 VIA_via4_0
* cell instance $8171 r0 *1 58.615,58.03
X$8171 243 VIA_via3_2
* cell instance $8172 r0 *1 63.375,58.03
X$8172 243 VIA_via4_0
* cell instance $8173 r0 *1 65.055,56.49
X$8173 243 VIA_via3_2
* cell instance $8174 r0 *1 63.375,56.49
X$8174 243 VIA_via3_2
* cell instance $8175 r0 *1 65.055,48.37
X$8175 243 VIA_via3_2
* cell instance $8176 r0 *1 56.095,45.99
X$8176 243 VIA_via3_2
* cell instance $8177 r0 *1 65.055,45.99
X$8177 243 VIA_via3_2
* cell instance $8178 r0 *1 61.275,10.57
X$8178 244 VIA_via2_5
* cell instance $8179 r0 *1 61.275,9.17
X$8179 244 VIA_via1_4
* cell instance $8180 r0 *1 64.125,10.57
X$8180 244 VIA_via1_4
* cell instance $8181 r0 *1 64.125,10.57
X$8181 244 VIA_via2_5
* cell instance $8182 r0 *1 12.635,12.39
X$8182 245 VIA_via1_7
* cell instance $8183 r0 *1 12.825,16.03
X$8183 245 VIA_via1_4
* cell instance $8184 r0 *1 10.165,13.23
X$8184 246 VIA_via1_4
* cell instance $8185 r0 *1 10.165,13.23
X$8185 246 VIA_via2_5
* cell instance $8186 r0 *1 13.775,13.23
X$8186 246 VIA_via1_4
* cell instance $8187 r0 *1 13.775,13.23
X$8187 246 VIA_via2_5
* cell instance $8188 r0 *1 14.155,13.23
X$8188 246 VIA_via1_4
* cell instance $8189 r0 *1 14.155,13.23
X$8189 246 VIA_via2_5
* cell instance $8190 r0 *1 15.105,5.39
X$8190 247 VIA_via1_7
* cell instance $8191 r0 *1 15.485,14.77
X$8191 247 VIA_via1_4
* cell instance $8192 r0 *1 51.585,15.89
X$8192 248 VIA_via2_5
* cell instance $8193 r0 *1 35.245,13.79
X$8193 248 VIA_via2_5
* cell instance $8194 r0 *1 35.245,15.75
X$8194 248 VIA_via2_5
* cell instance $8195 r0 *1 32.395,13.79
X$8195 248 VIA_via2_5
* cell instance $8196 r0 *1 41.515,15.89
X$8196 248 VIA_via2_5
* cell instance $8197 r0 *1 22.325,13.37
X$8197 248 VIA_via2_5
* cell instance $8198 r0 *1 16.815,14.91
X$8198 248 VIA_via2_5
* cell instance $8199 r0 *1 16.815,13.37
X$8199 248 VIA_via2_5
* cell instance $8200 r0 *1 41.515,14.77
X$8200 248 VIA_via1_4
* cell instance $8201 r0 *1 22.325,14.77
X$8201 248 VIA_via1_4
* cell instance $8202 r0 *1 46.265,16.03
X$8202 248 VIA_via1_4
* cell instance $8203 r0 *1 46.265,15.89
X$8203 248 VIA_via2_5
* cell instance $8204 r0 *1 35.245,16.03
X$8204 248 VIA_via1_4
* cell instance $8205 r0 *1 32.205,13.23
X$8205 248 VIA_via1_4
* cell instance $8206 r0 *1 32.205,13.23
X$8206 248 VIA_via2_5
* cell instance $8207 r0 *1 26.885,13.23
X$8207 248 VIA_via1_4
* cell instance $8208 r0 *1 26.885,13.23
X$8208 248 VIA_via2_5
* cell instance $8209 r0 *1 51.585,17.15
X$8209 248 VIA_via1_4
* cell instance $8210 r0 *1 51.965,13.23
X$8210 248 VIA_via1_4
* cell instance $8211 r0 *1 18.335,13.23
X$8211 248 VIA_via1_4
* cell instance $8212 r0 *1 18.335,13.37
X$8212 248 VIA_via2_5
* cell instance $8213 r0 *1 15.865,14.77
X$8213 248 VIA_via1_4
* cell instance $8214 r0 *1 15.865,14.91
X$8214 248 VIA_via2_5
* cell instance $8215 r0 *1 13.775,14.77
X$8215 248 VIA_via1_4
* cell instance $8216 r0 *1 13.775,14.77
X$8216 248 VIA_via2_5
* cell instance $8217 r0 *1 18.335,14.35
X$8217 249 VIA_via1_4
* cell instance $8218 r0 *1 17.765,16.03
X$8218 249 VIA_via1_4
* cell instance $8219 r0 *1 21.185,11.97
X$8219 250 VIA_via2_5
* cell instance $8220 r0 *1 20.995,13.23
X$8220 250 VIA_via1_4
* cell instance $8221 r0 *1 19.285,11.97
X$8221 250 VIA_via1_4
* cell instance $8222 r0 *1 19.285,11.97
X$8222 250 VIA_via2_5
* cell instance $8223 r0 *1 21.185,10.85
X$8223 250 VIA_via1_4
* cell instance $8224 r0 *1 21.945,13.79
X$8224 251 VIA_via1_7
* cell instance $8225 r0 *1 21.375,14.77
X$8225 251 VIA_via1_4
* cell instance $8226 r0 *1 32.015,12.39
X$8226 252 VIA_via1_7
* cell instance $8227 r0 *1 32.395,13.23
X$8227 252 VIA_via1_4
* cell instance $8228 r0 *1 35.055,18.83
X$8228 253 VIA_via1_4
* cell instance $8229 r0 *1 35.245,13.51
X$8229 253 VIA_via1_4
* cell instance $8230 r0 *1 39.805,49.35
X$8230 254 VIA_via2_5
* cell instance $8231 r0 *1 43.795,49.35
X$8231 254 VIA_via2_5
* cell instance $8232 r0 *1 39.805,50.89
X$8232 254 VIA_via2_5
* cell instance $8233 r0 *1 32.775,14.91
X$8233 254 VIA_via2_5
* cell instance $8234 r0 *1 25.175,14.91
X$8234 254 VIA_via2_5
* cell instance $8235 r0 *1 25.935,14.91
X$8235 254 VIA_via2_5
* cell instance $8236 r0 *1 25.935,15.75
X$8236 254 VIA_via2_5
* cell instance $8237 r0 *1 25.175,15.75
X$8237 254 VIA_via2_5
* cell instance $8238 r0 *1 18.335,16.03
X$8238 254 VIA_via2_5
* cell instance $8239 r0 *1 12.255,50.89
X$8239 254 VIA_via2_5
* cell instance $8240 r0 *1 21.755,14.77
X$8240 254 VIA_via1_4
* cell instance $8241 r0 *1 21.755,14.91
X$8241 254 VIA_via2_5
* cell instance $8242 r0 *1 44.555,13.23
X$8242 254 VIA_via1_4
* cell instance $8243 r0 *1 44.555,13.23
X$8243 254 VIA_via2_5
* cell instance $8244 r0 *1 41.135,13.23
X$8244 254 VIA_via1_4
* cell instance $8245 r0 *1 41.135,13.23
X$8245 254 VIA_via2_5
* cell instance $8246 r0 *1 35.435,13.23
X$8246 254 VIA_via1_4
* cell instance $8247 r0 *1 35.435,13.23
X$8247 254 VIA_via2_5
* cell instance $8248 r0 *1 32.775,13.23
X$8248 254 VIA_via1_4
* cell instance $8249 r0 *1 32.775,13.23
X$8249 254 VIA_via2_5
* cell instance $8250 r0 *1 26.505,14.77
X$8250 254 VIA_via1_4
* cell instance $8251 r0 *1 26.505,14.91
X$8251 254 VIA_via2_5
* cell instance $8252 r0 *1 43.795,48.65
X$8252 254 VIA_via1_4
* cell instance $8253 r0 *1 43.795,48.51
X$8253 254 VIA_via2_5
* cell instance $8254 r0 *1 12.255,51.17
X$8254 254 VIA_via1_4
* cell instance $8255 r0 *1 18.335,14.77
X$8255 254 VIA_via1_4
* cell instance $8256 r0 *1 18.335,14.91
X$8256 254 VIA_via2_5
* cell instance $8257 r0 *1 13.205,16.03
X$8257 254 VIA_via1_4
* cell instance $8258 r0 *1 13.205,16.03
X$8258 254 VIA_via2_5
* cell instance $8259 r0 *1 16.055,16.03
X$8259 254 VIA_via1_4
* cell instance $8260 r0 *1 16.055,16.03
X$8260 254 VIA_via2_5
* cell instance $8261 r0 *1 44.055,48.51
X$8261 254 VIA_via3_2
* cell instance $8262 r0 *1 44.055,13.23
X$8262 254 VIA_via3_2
* cell instance $8263 r0 *1 41.135,12.39
X$8263 255 VIA_via1_7
* cell instance $8264 r0 *1 40.755,13.23
X$8264 255 VIA_via1_4
* cell instance $8265 r0 *1 41.135,14.77
X$8265 256 VIA_via1_4
* cell instance $8266 r0 *1 41.895,6.23
X$8266 256 VIA_via1_4
* cell instance $8267 r0 *1 30.115,17.43
X$8267 257 VIA_via1_7
* cell instance $8268 r0 *1 46.645,23.59
X$8268 257 VIA_via2_5
* cell instance $8269 r0 *1 46.645,23.17
X$8269 257 VIA_via2_5
* cell instance $8270 r0 *1 46.835,15.05
X$8270 257 VIA_via2_5
* cell instance $8271 r0 *1 45.315,15.05
X$8271 257 VIA_via2_5
* cell instance $8272 r0 *1 30.115,15.19
X$8272 257 VIA_via2_5
* cell instance $8273 r0 *1 31.825,23.45
X$8273 257 VIA_via2_5
* cell instance $8274 r0 *1 38.665,15.33
X$8274 257 VIA_via2_5
* cell instance $8275 r0 *1 6.745,18.69
X$8275 257 VIA_via2_5
* cell instance $8276 r0 *1 6.745,21.63
X$8276 257 VIA_via2_5
* cell instance $8277 r0 *1 8.645,15.05
X$8277 257 VIA_via2_5
* cell instance $8278 r0 *1 5.985,23.45
X$8278 257 VIA_via2_5
* cell instance $8279 r0 *1 6.175,15.05
X$8279 257 VIA_via2_5
* cell instance $8280 r0 *1 6.365,21.63
X$8280 257 VIA_via2_5
* cell instance $8281 r0 *1 6.365,23.45
X$8281 257 VIA_via2_5
* cell instance $8282 r0 *1 19.855,15.05
X$8282 257 VIA_via2_5
* cell instance $8283 r0 *1 8.645,18.83
X$8283 257 VIA_via1_4
* cell instance $8284 r0 *1 8.645,18.69
X$8284 257 VIA_via2_5
* cell instance $8285 r0 *1 31.825,23.17
X$8285 257 VIA_via1_4
* cell instance $8286 r0 *1 44.935,14.77
X$8286 257 VIA_via1_4
* cell instance $8287 r0 *1 46.835,14.77
X$8287 257 VIA_via1_4
* cell instance $8288 r0 *1 5.985,24.43
X$8288 257 VIA_via1_4
* cell instance $8289 r0 *1 5.035,21.63
X$8289 257 VIA_via1_4
* cell instance $8290 r0 *1 5.035,21.63
X$8290 257 VIA_via2_5
* cell instance $8291 r0 *1 38.665,14.77
X$8291 257 VIA_via1_4
* cell instance $8292 r0 *1 6.175,14.77
X$8292 257 VIA_via1_4
* cell instance $8293 r0 *1 49.495,23.17
X$8293 257 VIA_via1_4
* cell instance $8294 r0 *1 49.495,23.17
X$8294 257 VIA_via2_5
* cell instance $8295 r0 *1 19.855,16.03
X$8295 257 VIA_via1_4
* cell instance $8296 r0 *1 49.305,14.21
X$8296 258 VIA_via1_7
* cell instance $8297 r0 *1 48.355,11.97
X$8297 258 VIA_via1_4
* cell instance $8298 r0 *1 48.355,14.77
X$8298 259 VIA_via1_4
* cell instance $8299 r0 *1 48.355,14.77
X$8299 259 VIA_via2_5
* cell instance $8300 r0 *1 50.635,12.25
X$8300 259 VIA_via1_4
* cell instance $8301 r0 *1 50.825,14.77
X$8301 259 VIA_via1_4
* cell instance $8302 r0 *1 50.825,14.77
X$8302 259 VIA_via2_5
* cell instance $8303 r0 *1 81.035,42.63
X$8303 260 VIA_via1_7
* cell instance $8304 r0 *1 79.705,70.63
X$8304 260 VIA_via1_7
* cell instance $8305 r0 *1 79.705,70.63
X$8305 260 VIA_via2_5
* cell instance $8306 r0 *1 78.755,63.77
X$8306 260 VIA_via1_7
* cell instance $8307 r0 *1 78.755,63.77
X$8307 260 VIA_via2_5
* cell instance $8308 r0 *1 77.425,17.43
X$8308 260 VIA_via1_7
* cell instance $8309 r0 *1 68.115,70.63
X$8309 260 VIA_via1_7
* cell instance $8310 r0 *1 68.115,70.49
X$8310 260 VIA_via2_5
* cell instance $8311 r0 *1 63.935,13.37
X$8311 260 VIA_via1_7
* cell instance $8312 r0 *1 66.975,14.63
X$8312 260 VIA_via1_7
* cell instance $8313 r0 *1 66.975,14.49
X$8313 260 VIA_via2_5
* cell instance $8314 r0 *1 81.985,23.24
X$8314 260 VIA_via1_7
* cell instance $8315 r0 *1 81.985,23.17
X$8315 260 VIA_via2_5
* cell instance $8316 r0 *1 77.425,13.65
X$8316 260 VIA_via2_5
* cell instance $8317 r0 *1 80.845,23.17
X$8317 260 VIA_via2_5
* cell instance $8318 r0 *1 77.425,18.41
X$8318 260 VIA_via2_5
* cell instance $8319 r0 *1 67.355,14.49
X$8319 260 VIA_via2_5
* cell instance $8320 r0 *1 67.355,13.37
X$8320 260 VIA_via2_5
* cell instance $8321 r0 *1 68.685,40.25
X$8321 260 VIA_via2_5
* cell instance $8322 r0 *1 63.935,14.35
X$8322 260 VIA_via2_5
* cell instance $8323 r0 *1 80.465,41.65
X$8323 260 VIA_via2_5
* cell instance $8324 r0 *1 80.465,40.39
X$8324 260 VIA_via2_5
* cell instance $8325 r0 *1 81.035,41.65
X$8325 260 VIA_via2_5
* cell instance $8326 r0 *1 80.465,31.57
X$8326 260 VIA_via1_4
* cell instance $8327 r0 *1 63.745,48.51
X$8327 260 VIA_via1_4
* cell instance $8328 r0 *1 63.745,48.51
X$8328 260 VIA_via2_5
* cell instance $8329 r0 *1 68.685,39.97
X$8329 260 VIA_via1_4
* cell instance $8330 r0 *1 68.695,39.97
X$8330 260 VIA_via3_2
* cell instance $8331 r0 *1 68.685,39.97
X$8331 260 VIA_via2_5
* cell instance $8332 r0 *1 80.175,18.41
X$8332 260 VIA_via3_2
* cell instance $8333 r0 *1 68.695,70.49
X$8333 260 VIA_via3_2
* cell instance $8334 r0 *1 80.175,23.17
X$8334 260 VIA_via3_2
* cell instance $8335 r0 *1 79.335,70.63
X$8335 260 VIA_via3_2
* cell instance $8336 r0 *1 68.695,48.51
X$8336 260 VIA_via3_2
* cell instance $8337 r0 *1 79.335,63.77
X$8337 260 VIA_via3_2
* cell instance $8338 r0 *1 53.485,13.79
X$8338 261 VIA_via2_5
* cell instance $8339 r0 *1 85.215,12.39
X$8339 261 VIA_via2_5
* cell instance $8340 r0 *1 89.965,12.39
X$8340 261 VIA_via2_5
* cell instance $8341 r0 *1 53.485,29.89
X$8341 261 VIA_via2_5
* cell instance $8342 r0 *1 62.795,34.51
X$8342 261 VIA_via2_5
* cell instance $8343 r0 *1 70.205,12.39
X$8343 261 VIA_via2_5
* cell instance $8344 r0 *1 70.205,13.65
X$8344 261 VIA_via2_5
* cell instance $8345 r0 *1 53.485,34.51
X$8345 261 VIA_via2_5
* cell instance $8346 r0 *1 52.915,34.51
X$8346 261 VIA_via2_5
* cell instance $8347 r0 *1 89.965,11.97
X$8347 261 VIA_via1_4
* cell instance $8348 r0 *1 91.105,32.83
X$8348 261 VIA_via1_4
* cell instance $8349 r0 *1 91.105,32.83
X$8349 261 VIA_via2_5
* cell instance $8350 r0 *1 85.215,11.97
X$8350 261 VIA_via1_4
* cell instance $8351 r0 *1 90.915,37.17
X$8351 261 VIA_via1_4
* cell instance $8352 r0 *1 90.915,37.17
X$8352 261 VIA_via2_5
* cell instance $8353 r0 *1 90.815,37.17
X$8353 261 VIA_via3_2
* cell instance $8354 r0 *1 53.485,20.65
X$8354 261 VIA_via1_4
* cell instance $8355 r0 *1 90.915,23.1
X$8355 261 VIA_via1_4
* cell instance $8356 r0 *1 90.915,23.03
X$8356 261 VIA_via2_5
* cell instance $8357 r0 *1 52.915,35.63
X$8357 261 VIA_via1_4
* cell instance $8358 r0 *1 57.095,34.37
X$8358 261 VIA_via1_4
* cell instance $8359 r0 *1 57.095,34.51
X$8359 261 VIA_via2_5
* cell instance $8360 r0 *1 62.795,35.63
X$8360 261 VIA_via1_4
* cell instance $8361 r0 *1 70.205,11.97
X$8361 261 VIA_via1_4
* cell instance $8362 r0 *1 46.645,30.03
X$8362 261 VIA_via1_4
* cell instance $8363 r0 *1 46.645,29.89
X$8363 261 VIA_via2_5
* cell instance $8364 r0 *1 90.815,32.83
X$8364 261 VIA_via3_2
* cell instance $8365 r0 *1 90.815,23.17
X$8365 261 VIA_via3_2
* cell instance $8366 r0 *1 90.815,12.39
X$8366 261 VIA_via3_2
* cell instance $8367 r0 *1 71.155,5.39
X$8367 262 VIA_via1_7
* cell instance $8368 r0 *1 70.585,17.57
X$8368 262 VIA_via1_4
* cell instance $8369 r0 *1 93.195,13.37
X$8369 263 VIA_via1_7
* cell instance $8370 r0 *1 74.195,14.91
X$8370 263 VIA_via2_5
* cell instance $8371 r0 *1 93.195,15.05
X$8371 263 VIA_via2_5
* cell instance $8372 r0 *1 73.435,38.01
X$8372 263 VIA_via2_5
* cell instance $8373 r0 *1 90.155,39.83
X$8373 263 VIA_via2_5
* cell instance $8374 r0 *1 90.535,39.97
X$8374 263 VIA_via2_5
* cell instance $8375 r0 *1 90.155,38.01
X$8375 263 VIA_via2_5
* cell instance $8376 r0 *1 73.055,31.99
X$8376 263 VIA_via2_5
* cell instance $8377 r0 *1 72.295,31.99
X$8377 263 VIA_via2_5
* cell instance $8378 r0 *1 77.045,31.99
X$8378 263 VIA_via2_5
* cell instance $8379 r0 *1 73.815,31.99
X$8379 263 VIA_via2_5
* cell instance $8380 r0 *1 93.005,17.57
X$8380 263 VIA_via1_4
* cell instance $8381 r0 *1 87.685,14.77
X$8381 263 VIA_via1_4
* cell instance $8382 r0 *1 87.685,14.91
X$8382 263 VIA_via2_5
* cell instance $8383 r0 *1 73.245,38.15
X$8383 263 VIA_via1_4
* cell instance $8384 r0 *1 73.245,38.01
X$8384 263 VIA_via2_5
* cell instance $8385 r0 *1 93.385,27.23
X$8385 263 VIA_via1_4
* cell instance $8386 r0 *1 77.045,32.83
X$8386 263 VIA_via1_4
* cell instance $8387 r0 *1 90.535,44.03
X$8387 263 VIA_via1_4
* cell instance $8388 r0 *1 90.535,43.89
X$8388 263 VIA_via2_5
* cell instance $8389 r0 *1 88.635,44.03
X$8389 263 VIA_via1_4
* cell instance $8390 r0 *1 88.635,43.89
X$8390 263 VIA_via2_5
* cell instance $8391 r0 *1 91.295,39.97
X$8391 263 VIA_via1_4
* cell instance $8392 r0 *1 91.295,39.97
X$8392 263 VIA_via2_5
* cell instance $8393 r0 *1 74.385,13.23
X$8393 263 VIA_via1_4
* cell instance $8394 r0 *1 72.295,31.57
X$8394 263 VIA_via1_4
* cell instance $8395 r0 *1 88.825,14.21
X$8395 264 VIA_via1_7
* cell instance $8396 r0 *1 88.445,13.23
X$8396 264 VIA_via1_4
* cell instance $8397 r0 *1 89.585,44.31
X$8397 265 VIA_via2_5
* cell instance $8398 r0 *1 88.255,44.31
X$8398 265 VIA_via2_5
* cell instance $8399 r0 *1 88.825,12.25
X$8399 265 VIA_via1_4
* cell instance $8400 r0 *1 89.965,51.17
X$8400 265 VIA_via1_4
* cell instance $8401 r0 *1 89.965,49.63
X$8401 265 VIA_via1_4
* cell instance $8402 r0 *1 91.485,12.81
X$8402 266 VIA_via1_7
* cell instance $8403 r0 *1 91.105,11.97
X$8403 266 VIA_via1_4
* cell instance $8404 r0 *1 94.525,13.23
X$8404 267 VIA_via2_5
* cell instance $8405 r0 *1 92.625,13.23
X$8405 267 VIA_via1_4
* cell instance $8406 r0 *1 92.625,13.23
X$8406 267 VIA_via2_5
* cell instance $8407 r0 *1 93.385,13.23
X$8407 267 VIA_via1_4
* cell instance $8408 r0 *1 93.385,13.23
X$8408 267 VIA_via2_5
* cell instance $8409 r0 *1 94.525,12.25
X$8409 267 VIA_via1_4
* cell instance $8410 r0 *1 7.315,14.21
X$8410 268 VIA_via1_7
* cell instance $8411 r0 *1 7.315,13.23
X$8411 268 VIA_via2_5
* cell instance $8412 r0 *1 4.275,13.23
X$8412 268 VIA_via1_4
* cell instance $8413 r0 *1 4.275,13.23
X$8413 268 VIA_via2_5
* cell instance $8414 r0 *1 11.495,13.23
X$8414 269 VIA_via1_4
* cell instance $8415 r0 *1 10.545,13.23
X$8415 269 VIA_via1_4
* cell instance $8416 r0 *1 14.725,12.11
X$8416 270 VIA_via2_5
* cell instance $8417 r0 *1 14.535,11.97
X$8417 270 VIA_via1_4
* cell instance $8418 r0 *1 14.535,12.11
X$8418 270 VIA_via2_5
* cell instance $8419 r0 *1 18.145,12.11
X$8419 270 VIA_via1_4
* cell instance $8420 r0 *1 18.145,12.11
X$8420 270 VIA_via2_5
* cell instance $8421 r0 *1 14.725,13.23
X$8421 270 VIA_via1_4
* cell instance $8422 r0 *1 14.915,11.97
X$8422 271 VIA_via1_4
* cell instance $8423 r0 *1 14.915,11.97
X$8423 271 VIA_via2_5
* cell instance $8424 r0 *1 15.865,11.97
X$8424 271 VIA_via1_4
* cell instance $8425 r0 *1 15.865,11.97
X$8425 271 VIA_via2_5
* cell instance $8426 r0 *1 94.335,13.09
X$8426 272 VIA_via1_4
* cell instance $8427 r0 *1 94.335,13.09
X$8427 272 VIA_via2_5
* cell instance $8428 r0 *1 91.295,13.23
X$8428 272 VIA_via1_4
* cell instance $8429 r0 *1 91.295,13.09
X$8429 272 VIA_via2_5
* cell instance $8430 r0 *1 22.135,12.25
X$8430 273 VIA_via2_5
* cell instance $8431 r0 *1 21.565,12.25
X$8431 273 VIA_via2_5
* cell instance $8432 r0 *1 21.565,13.23
X$8432 273 VIA_via1_4
* cell instance $8433 r0 *1 22.135,10.43
X$8433 273 VIA_via1_4
* cell instance $8434 r0 *1 23.275,12.25
X$8434 273 VIA_via1_4
* cell instance $8435 r0 *1 23.275,12.25
X$8435 273 VIA_via2_5
* cell instance $8436 r0 *1 76.475,35.49
X$8436 274 VIA_via1_7
* cell instance $8437 r0 *1 91.675,21.77
X$8437 274 VIA_via2_5
* cell instance $8438 r0 *1 91.105,21.77
X$8438 274 VIA_via2_5
* cell instance $8439 r0 *1 93.005,37.87
X$8439 274 VIA_via2_5
* cell instance $8440 r0 *1 90.535,38.29
X$8440 274 VIA_via2_5
* cell instance $8441 r0 *1 91.295,37.87
X$8441 274 VIA_via2_5
* cell instance $8442 r0 *1 91.105,28.77
X$8442 274 VIA_via2_5
* cell instance $8443 r0 *1 75.715,32.69
X$8443 274 VIA_via2_5
* cell instance $8444 r0 *1 76.475,34.79
X$8444 274 VIA_via2_5
* cell instance $8445 r0 *1 91.295,34.23
X$8445 274 VIA_via2_5
* cell instance $8446 r0 *1 75.715,34.79
X$8446 274 VIA_via2_5
* cell instance $8447 r0 *1 79.135,34.79
X$8447 274 VIA_via2_5
* cell instance $8448 r0 *1 91.865,34.09
X$8448 274 VIA_via2_5
* cell instance $8449 r0 *1 91.675,13.23
X$8449 274 VIA_via1_4
* cell instance $8450 r0 *1 91.675,13.23
X$8450 274 VIA_via2_5
* cell instance $8451 r0 *1 88.825,13.23
X$8451 274 VIA_via1_4
* cell instance $8452 r0 *1 88.825,13.23
X$8452 274 VIA_via2_5
* cell instance $8453 r0 *1 73.815,32.83
X$8453 274 VIA_via1_4
* cell instance $8454 r0 *1 73.815,32.69
X$8454 274 VIA_via2_5
* cell instance $8455 r0 *1 75.715,11.97
X$8455 274 VIA_via1_4
* cell instance $8456 r0 *1 79.135,34.37
X$8456 274 VIA_via1_4
* cell instance $8457 r0 *1 79.135,34.23
X$8457 274 VIA_via2_5
* cell instance $8458 r0 *1 93.005,38.43
X$8458 274 VIA_via1_4
* cell instance $8459 r0 *1 91.865,28.77
X$8459 274 VIA_via1_4
* cell instance $8460 r0 *1 91.865,28.77
X$8460 274 VIA_via2_5
* cell instance $8461 r0 *1 91.865,45.57
X$8461 274 VIA_via1_4
* cell instance $8462 r0 *1 91.865,45.57
X$8462 274 VIA_via2_5
* cell instance $8463 r0 *1 90.535,45.57
X$8463 274 VIA_via1_4
* cell instance $8464 r0 *1 90.535,45.57
X$8464 274 VIA_via2_5
* cell instance $8465 r0 *1 92.625,21.63
X$8465 274 VIA_via1_4
* cell instance $8466 r0 *1 92.625,21.77
X$8466 274 VIA_via2_5
* cell instance $8467 r0 *1 93.005,12.81
X$8467 275 VIA_via1_7
* cell instance $8468 r0 *1 93.005,12.81
X$8468 275 VIA_via2_5
* cell instance $8469 r0 *1 92.245,12.81
X$8469 275 VIA_via2_5
* cell instance $8470 r0 *1 92.245,11.97
X$8470 275 VIA_via1_4
* cell instance $8471 r0 *1 26.885,12.39
X$8471 276 VIA_via1_7
* cell instance $8472 r0 *1 26.885,12.39
X$8472 276 VIA_via2_5
* cell instance $8473 r0 *1 26.125,12.39
X$8473 276 VIA_via2_5
* cell instance $8474 r0 *1 26.125,14.77
X$8474 276 VIA_via1_4
* cell instance $8475 r0 *1 89.965,52.15
X$8475 277 VIA_via2_5
* cell instance $8476 r0 *1 90.725,12.11
X$8476 277 VIA_via1_4
* cell instance $8477 r0 *1 90.725,12.11
X$8477 277 VIA_via2_5
* cell instance $8478 r0 *1 90.815,12.11
X$8478 277 VIA_via3_2
* cell instance $8479 r0 *1 90.815,12.11
X$8479 277 VIA_via4_0
* cell instance $8480 r0 *1 90.815,12.11
X$8480 277 VIA_via5_0
* cell instance $8481 r0 *1 90.915,52.43
X$8481 277 VIA_via1_4
* cell instance $8482 r0 *1 89.965,52.43
X$8482 277 VIA_via1_4
* cell instance $8483 r0 *1 90.815,52.15
X$8483 277 VIA_via4_0
* cell instance $8484 r0 *1 90.815,52.15
X$8484 277 VIA_via5_0
* cell instance $8485 r0 *1 90.815,52.15
X$8485 277 VIA_via3_2
* cell instance $8486 r0 *1 90.915,52.15
X$8486 277 VIA_via2_5
* cell instance $8487 r0 *1 31.825,6.23
X$8487 278 VIA_via1_4
* cell instance $8488 r0 *1 31.825,13.23
X$8488 278 VIA_via1_4
* cell instance $8489 r0 *1 36.195,12.39
X$8489 279 VIA_via1_7
* cell instance $8490 r0 *1 36.195,12.39
X$8490 279 VIA_via2_5
* cell instance $8491 r0 *1 35.055,12.39
X$8491 279 VIA_via2_5
* cell instance $8492 r0 *1 35.055,13.23
X$8492 279 VIA_via1_4
* cell instance $8493 r0 *1 44.175,12.39
X$8493 280 VIA_via1_7
* cell instance $8494 r0 *1 44.175,13.23
X$8494 280 VIA_via1_4
* cell instance $8495 r0 *1 88.635,12.81
X$8495 281 VIA_via1_7
* cell instance $8496 r0 *1 88.635,11.97
X$8496 281 VIA_via1_4
* cell instance $8497 r0 *1 47.975,14.21
X$8497 282 VIA_via1_7
* cell instance $8498 r0 *1 47.975,13.23
X$8498 282 VIA_via1_4
* cell instance $8499 r0 *1 84.835,11.97
X$8499 283 VIA_via1_4
* cell instance $8500 r0 *1 84.835,11.97
X$8500 283 VIA_via2_5
* cell instance $8501 r0 *1 83.125,11.97
X$8501 283 VIA_via1_4
* cell instance $8502 r0 *1 83.125,11.97
X$8502 283 VIA_via2_5
* cell instance $8503 r0 *1 80.275,11.97
X$8503 284 VIA_via1_4
* cell instance $8504 r0 *1 80.275,11.97
X$8504 284 VIA_via2_5
* cell instance $8505 r0 *1 82.175,10.85
X$8505 284 VIA_via1_4
* cell instance $8506 r0 *1 82.175,11.97
X$8506 284 VIA_via1_4
* cell instance $8507 r0 *1 82.175,11.97
X$8507 284 VIA_via2_5
* cell instance $8508 r0 *1 73.625,13.79
X$8508 285 VIA_via2_5
* cell instance $8509 r0 *1 84.455,13.79
X$8509 285 VIA_via2_5
* cell instance $8510 r0 *1 85.405,48.37
X$8510 285 VIA_via1_4
* cell instance $8511 r0 *1 73.625,13.51
X$8511 285 VIA_via1_4
* cell instance $8512 r0 *1 85.215,51.17
X$8512 285 VIA_via1_4
* cell instance $8513 r0 *1 62.605,54.95
X$8513 286 VIA_via1_7
* cell instance $8514 r0 *1 62.605,54.95
X$8514 286 VIA_via2_5
* cell instance $8515 r0 *1 61.465,55.51
X$8515 286 VIA_via1_4
* cell instance $8516 r0 *1 54.625,16.17
X$8516 286 VIA_via1_7
* cell instance $8517 r0 *1 54.625,16.45
X$8517 286 VIA_via2_5
* cell instance $8518 r0 *1 57.095,16.45
X$8518 286 VIA_via2_5
* cell instance $8519 r0 *1 61.465,55.09
X$8519 286 VIA_via2_5
* cell instance $8520 r0 *1 62.985,49.63
X$8520 286 VIA_via2_5
* cell instance $8521 r0 *1 62.985,54.95
X$8521 286 VIA_via2_5
* cell instance $8522 r0 *1 56.905,11.97
X$8522 286 VIA_via1_4
* cell instance $8523 r0 *1 56.905,11.97
X$8523 286 VIA_via2_5
* cell instance $8524 r0 *1 51.205,11.97
X$8524 286 VIA_via1_4
* cell instance $8525 r0 *1 51.205,11.97
X$8525 286 VIA_via2_5
* cell instance $8526 r0 *1 63.365,49.63
X$8526 286 VIA_via1_4
* cell instance $8527 r0 *1 63.365,49.63
X$8527 286 VIA_via2_5
* cell instance $8528 r0 *1 54.245,55.23
X$8528 286 VIA_via1_4
* cell instance $8529 r0 *1 54.245,55.09
X$8529 286 VIA_via2_5
* cell instance $8530 r0 *1 58.335,16.45
X$8530 286 VIA_via3_2
* cell instance $8531 r0 *1 62.255,49.63
X$8531 286 VIA_via3_2
* cell instance $8532 r0 *1 62.255,42.07
X$8532 286 VIA_via3_2
* cell instance $8533 r0 *1 58.335,42.07
X$8533 286 VIA_via3_2
* cell instance $8534 r0 *1 58.995,11.97
X$8534 287 VIA_via1_4
* cell instance $8535 r0 *1 58.995,12.11
X$8535 287 VIA_via2_5
* cell instance $8536 r0 *1 63.175,12.11
X$8536 287 VIA_via1_4
* cell instance $8537 r0 *1 63.175,12.11
X$8537 287 VIA_via2_5
* cell instance $8538 r0 *1 68.115,14.21
X$8538 288 VIA_via1_7
* cell instance $8539 r0 *1 68.115,14.21
X$8539 288 VIA_via2_5
* cell instance $8540 r0 *1 66.975,14.21
X$8540 288 VIA_via2_5
* cell instance $8541 r0 *1 66.975,13.23
X$8541 288 VIA_via1_4
* cell instance $8542 r0 *1 70.965,10.99
X$8542 289 VIA_via1_7
* cell instance $8543 r0 *1 70.965,13.23
X$8543 289 VIA_via2_5
* cell instance $8544 r0 *1 73.435,13.23
X$8544 289 VIA_via1_4
* cell instance $8545 r0 *1 73.435,13.23
X$8545 289 VIA_via2_5
* cell instance $8546 r0 *1 65.645,12.25
X$8546 290 VIA_via2_5
* cell instance $8547 r0 *1 68.875,12.25
X$8547 290 VIA_via1_4
* cell instance $8548 r0 *1 68.875,12.25
X$8548 290 VIA_via2_5
* cell instance $8549 r0 *1 65.645,14.77
X$8549 290 VIA_via1_4
* cell instance $8550 r0 *1 68.875,10.43
X$8550 290 VIA_via1_4
* cell instance $8551 r0 *1 69.825,11.97
X$8551 291 VIA_via1_4
* cell instance $8552 r0 *1 69.825,11.97
X$8552 291 VIA_via2_5
* cell instance $8553 r0 *1 64.505,11.97
X$8553 291 VIA_via1_4
* cell instance $8554 r0 *1 64.505,11.97
X$8554 291 VIA_via2_5
* cell instance $8555 r0 *1 70.965,13.79
X$8555 292 VIA_via1_7
* cell instance $8556 r0 *1 70.965,13.79
X$8556 292 VIA_via2_5
* cell instance $8557 r0 *1 69.635,13.79
X$8557 292 VIA_via2_5
* cell instance $8558 r0 *1 69.635,14.77
X$8558 292 VIA_via1_4
* cell instance $8559 r0 *1 5.605,16.03
X$8559 293 VIA_via1_4
* cell instance $8560 r0 *1 5.605,16.03
X$8560 293 VIA_via2_5
* cell instance $8561 r0 *1 5.985,15.05
X$8561 293 VIA_via1_4
* cell instance $8562 r0 *1 4.275,16.03
X$8562 293 VIA_via1_4
* cell instance $8563 r0 *1 4.275,16.03
X$8563 293 VIA_via2_5
* cell instance $8564 r0 *1 6.555,13.65
X$8564 294 VIA_via1_4
* cell instance $8565 r0 *1 6.365,14.77
X$8565 294 VIA_via1_4
* cell instance $8566 r0 *1 6.175,16.03
X$8566 294 VIA_via1_4
* cell instance $8567 r0 *1 12.445,15.61
X$8567 295 VIA_via1_7
* cell instance $8568 r0 *1 12.445,16.59
X$8568 295 VIA_via1_7
* cell instance $8569 r0 *1 5.985,37.87
X$8569 295 VIA_via2_5
* cell instance $8570 r0 *1 13.015,37.87
X$8570 295 VIA_via2_5
* cell instance $8571 r0 *1 13.205,38.43
X$8571 295 VIA_via2_5
* cell instance $8572 r0 *1 12.445,14.91
X$8572 295 VIA_via2_5
* cell instance $8573 r0 *1 4.845,14.91
X$8573 295 VIA_via2_5
* cell instance $8574 r0 *1 14.915,18.55
X$8574 295 VIA_via2_5
* cell instance $8575 r0 *1 12.635,18.69
X$8575 295 VIA_via2_5
* cell instance $8576 r0 *1 14.155,18.69
X$8576 295 VIA_via2_5
* cell instance $8577 r0 *1 13.015,35.91
X$8577 295 VIA_via2_5
* cell instance $8578 r0 *1 13.775,35.91
X$8578 295 VIA_via2_5
* cell instance $8579 r0 *1 6.935,14.77
X$8579 295 VIA_via1_4
* cell instance $8580 r0 *1 6.935,14.91
X$8580 295 VIA_via2_5
* cell instance $8581 r0 *1 4.845,16.03
X$8581 295 VIA_via1_4
* cell instance $8582 r0 *1 6.175,32.83
X$8582 295 VIA_via1_4
* cell instance $8583 r0 *1 5.985,41.23
X$8583 295 VIA_via1_4
* cell instance $8584 r0 *1 5.795,38.43
X$8584 295 VIA_via1_4
* cell instance $8585 r0 *1 13.585,18.83
X$8585 295 VIA_via1_4
* cell instance $8586 r0 *1 13.585,18.69
X$8586 295 VIA_via2_5
* cell instance $8587 r0 *1 14.915,17.57
X$8587 295 VIA_via1_4
* cell instance $8588 r0 *1 13.015,35.63
X$8588 295 VIA_via1_4
* cell instance $8589 r0 *1 15.105,38.43
X$8589 295 VIA_via1_4
* cell instance $8590 r0 *1 15.105,38.43
X$8590 295 VIA_via2_5
* cell instance $8591 r0 *1 13.205,39.97
X$8591 295 VIA_via1_4
* cell instance $8592 r0 *1 13.015,9.59
X$8592 296 VIA_via1_7
* cell instance $8593 r0 *1 13.395,14.77
X$8593 296 VIA_via1_4
* cell instance $8594 r0 *1 13.775,23.17
X$8594 297 VIA_via1_4
* cell instance $8595 r0 *1 13.585,14.63
X$8595 297 VIA_via1_4
* cell instance $8596 r0 *1 25.745,16.03
X$8596 298 VIA_via2_5
* cell instance $8597 r0 *1 26.125,16.03
X$8597 298 VIA_via1_4
* cell instance $8598 r0 *1 26.125,16.03
X$8598 298 VIA_via2_5
* cell instance $8599 r0 *1 25.555,15.05
X$8599 298 VIA_via1_4
* cell instance $8600 r0 *1 24.605,16.03
X$8600 298 VIA_via1_4
* cell instance $8601 r0 *1 24.605,16.03
X$8601 298 VIA_via2_5
* cell instance $8602 r0 *1 46.455,18.41
X$8602 299 VIA_via1_7
* cell instance $8603 r0 *1 46.455,18.41
X$8603 299 VIA_via2_5
* cell instance $8604 r0 *1 46.075,19.25
X$8604 299 VIA_via1_4
* cell instance $8605 r0 *1 49.115,18.41
X$8605 299 VIA_via2_5
* cell instance $8606 r0 *1 44.365,21.63
X$8606 299 VIA_via2_5
* cell instance $8607 r0 *1 48.355,18.41
X$8607 299 VIA_via2_5
* cell instance $8608 r0 *1 43.035,18.41
X$8608 299 VIA_via2_5
* cell instance $8609 r0 *1 42.655,18.41
X$8609 299 VIA_via2_5
* cell instance $8610 r0 *1 43.035,21.63
X$8610 299 VIA_via2_5
* cell instance $8611 r0 *1 48.735,16.03
X$8611 299 VIA_via1_4
* cell instance $8612 r0 *1 43.225,14.77
X$8612 299 VIA_via1_4
* cell instance $8613 r0 *1 48.355,17.57
X$8613 299 VIA_via1_4
* cell instance $8614 r0 *1 42.845,21.63
X$8614 299 VIA_via1_4
* cell instance $8615 r0 *1 42.465,16.03
X$8615 299 VIA_via1_4
* cell instance $8616 r0 *1 44.365,23.17
X$8616 299 VIA_via1_4
* cell instance $8617 r0 *1 45.885,20.37
X$8617 299 VIA_via1_4
* cell instance $8618 r0 *1 49.305,21.63
X$8618 299 VIA_via1_4
* cell instance $8619 r0 *1 45.125,14.77
X$8619 300 VIA_via1_4
* cell instance $8620 r0 *1 44.745,15.05
X$8620 300 VIA_via1_4
* cell instance $8621 r0 *1 44.935,16.03
X$8621 300 VIA_via1_4
* cell instance $8622 r0 *1 49.875,15.19
X$8622 301 VIA_via1_7
* cell instance $8623 r0 *1 49.115,38.15
X$8623 301 VIA_via2_5
* cell instance $8624 r0 *1 49.115,28.77
X$8624 301 VIA_via2_5
* cell instance $8625 r0 *1 47.785,42.91
X$8625 301 VIA_via2_5
* cell instance $8626 r0 *1 47.405,18.55
X$8626 301 VIA_via2_5
* cell instance $8627 r0 *1 48.925,18.55
X$8627 301 VIA_via2_5
* cell instance $8628 r0 *1 48.735,38.15
X$8628 301 VIA_via2_5
* cell instance $8629 r0 *1 48.735,34.23
X$8629 301 VIA_via2_5
* cell instance $8630 r0 *1 48.355,28.77
X$8630 301 VIA_via2_5
* cell instance $8631 r0 *1 47.595,14.77
X$8631 301 VIA_via1_4
* cell instance $8632 r0 *1 48.925,14.77
X$8632 301 VIA_via1_4
* cell instance $8633 r0 *1 47.595,18.83
X$8633 301 VIA_via1_4
* cell instance $8634 r0 *1 48.925,18.83
X$8634 301 VIA_via1_4
* cell instance $8635 r0 *1 49.115,42.77
X$8635 301 VIA_via1_4
* cell instance $8636 r0 *1 49.115,42.91
X$8636 301 VIA_via2_5
* cell instance $8637 r0 *1 49.115,41.23
X$8637 301 VIA_via1_4
* cell instance $8638 r0 *1 47.405,38.43
X$8638 301 VIA_via1_4
* cell instance $8639 r0 *1 47.405,38.29
X$8639 301 VIA_via2_5
* cell instance $8640 r0 *1 47.785,44.03
X$8640 301 VIA_via1_4
* cell instance $8641 r0 *1 50.065,28.77
X$8641 301 VIA_via1_4
* cell instance $8642 r0 *1 50.065,28.77
X$8642 301 VIA_via2_5
* cell instance $8643 r0 *1 48.355,34.37
X$8643 301 VIA_via1_4
* cell instance $8644 r0 *1 48.355,34.23
X$8644 301 VIA_via2_5
* cell instance $8645 r0 *1 50.255,14.91
X$8645 302 VIA_via2_5
* cell instance $8646 r0 *1 47.025,14.77
X$8646 302 VIA_via1_4
* cell instance $8647 r0 *1 47.025,14.91
X$8647 302 VIA_via2_5
* cell instance $8648 r0 *1 50.255,13.65
X$8648 302 VIA_via1_4
* cell instance $8649 r0 *1 51.395,14.77
X$8649 302 VIA_via1_4
* cell instance $8650 r0 *1 51.395,14.91
X$8650 302 VIA_via2_5
* cell instance $8651 r0 *1 56.905,16.03
X$8651 303 VIA_via2_5
* cell instance $8652 r0 *1 57.475,16.03
X$8652 303 VIA_via1_4
* cell instance $8653 r0 *1 57.475,16.03
X$8653 303 VIA_via2_5
* cell instance $8654 r0 *1 55.385,16.03
X$8654 303 VIA_via1_4
* cell instance $8655 r0 *1 55.385,16.03
X$8655 303 VIA_via2_5
* cell instance $8656 r0 *1 57.095,15.05
X$8656 303 VIA_via1_4
* cell instance $8657 r0 *1 65.075,13.79
X$8657 304 VIA_via1_7
* cell instance $8658 r0 *1 65.075,14.49
X$8658 304 VIA_via2_5
* cell instance $8659 r0 *1 62.035,14.77
X$8659 304 VIA_via1_4
* cell instance $8660 r0 *1 62.035,14.77
X$8660 304 VIA_via2_5
* cell instance $8661 r0 *1 44.175,16.17
X$8661 305 VIA_via1_7
* cell instance $8662 r0 *1 44.175,16.17
X$8662 305 VIA_via2_5
* cell instance $8663 r0 *1 29.545,16.17
X$8663 305 VIA_via1_7
* cell instance $8664 r0 *1 29.545,16.17
X$8664 305 VIA_via2_5
* cell instance $8665 r0 *1 39.045,16.17
X$8665 305 VIA_via1_7
* cell instance $8666 r0 *1 39.045,16.17
X$8666 305 VIA_via2_5
* cell instance $8667 r0 *1 50.635,16.17
X$8667 305 VIA_via2_5
* cell instance $8668 r0 *1 56.145,16.31
X$8668 305 VIA_via2_5
* cell instance $8669 r0 *1 56.335,14.91
X$8669 305 VIA_via2_5
* cell instance $8670 r0 *1 56.335,16.31
X$8670 305 VIA_via2_5
* cell instance $8671 r0 *1 56.145,25.27
X$8671 305 VIA_via2_5
* cell instance $8672 r0 *1 57.855,25.27
X$8672 305 VIA_via2_5
* cell instance $8673 r0 *1 31.635,25.55
X$8673 305 VIA_via2_5
* cell instance $8674 r0 *1 29.545,16.45
X$8674 305 VIA_via2_5
* cell instance $8675 r0 *1 30.495,16.17
X$8675 305 VIA_via2_5
* cell instance $8676 r0 *1 25.745,16.45
X$8676 305 VIA_via2_5
* cell instance $8677 r0 *1 68.685,14.91
X$8677 305 VIA_via2_5
* cell instance $8678 r0 *1 25.935,16.03
X$8678 305 VIA_via1_4
* cell instance $8679 r0 *1 31.065,21.63
X$8679 305 VIA_via1_4
* cell instance $8680 r0 *1 55.955,23.17
X$8680 305 VIA_via1_4
* cell instance $8681 r0 *1 64.885,14.77
X$8681 305 VIA_via1_4
* cell instance $8682 r0 *1 64.885,14.91
X$8682 305 VIA_via2_5
* cell instance $8683 r0 *1 68.685,16.03
X$8683 305 VIA_via1_4
* cell instance $8684 r0 *1 50.635,14.77
X$8684 305 VIA_via1_4
* cell instance $8685 r0 *1 57.855,27.23
X$8685 305 VIA_via1_4
* cell instance $8686 r0 *1 33.345,25.55
X$8686 305 VIA_via1_4
* cell instance $8687 r0 *1 33.345,25.55
X$8687 305 VIA_via2_5
* cell instance $8688 r0 *1 66.025,14.63
X$8688 306 VIA_via1_4
* cell instance $8689 r0 *1 65.835,17.57
X$8689 306 VIA_via1_4
* cell instance $8690 r0 *1 80.845,15.05
X$8690 307 VIA_via2_5
* cell instance $8691 r0 *1 81.985,15.05
X$8691 307 VIA_via1_4
* cell instance $8692 r0 *1 81.985,15.05
X$8692 307 VIA_via2_5
* cell instance $8693 r0 *1 80.655,13.23
X$8693 307 VIA_via1_4
* cell instance $8694 r0 *1 80.845,17.57
X$8694 307 VIA_via1_4
* cell instance $8695 r0 *1 86.735,14.77
X$8695 308 VIA_via1_4
* cell instance $8696 r0 *1 86.735,14.77
X$8696 308 VIA_via2_5
* cell instance $8697 r0 *1 88.255,15.75
X$8697 308 VIA_via1_4
* cell instance $8698 r0 *1 87.875,14.77
X$8698 308 VIA_via1_4
* cell instance $8699 r0 *1 87.875,14.77
X$8699 308 VIA_via2_5
* cell instance $8700 r0 *1 90.155,16.03
X$8700 309 VIA_via2_5
* cell instance $8701 r0 *1 88.825,16.03
X$8701 309 VIA_via2_5
* cell instance $8702 r0 *1 88.445,14.77
X$8702 309 VIA_via1_4
* cell instance $8703 r0 *1 90.155,17.15
X$8703 309 VIA_via1_4
* cell instance $8704 r0 *1 89.205,16.03
X$8704 309 VIA_via1_4
* cell instance $8705 r0 *1 89.205,16.03
X$8705 309 VIA_via2_5
* cell instance $8706 r0 *1 92.435,18.69
X$8706 310 VIA_via1_7
* cell instance $8707 r0 *1 92.435,18.83
X$8707 310 VIA_via2_5
* cell instance $8708 r0 *1 86.735,17.57
X$8708 310 VIA_via2_5
* cell instance $8709 r0 *1 89.775,18.83
X$8709 310 VIA_via2_5
* cell instance $8710 r0 *1 89.775,17.57
X$8710 310 VIA_via2_5
* cell instance $8711 r0 *1 95.285,17.01
X$8711 310 VIA_via2_5
* cell instance $8712 r0 *1 93.195,17.01
X$8712 310 VIA_via2_5
* cell instance $8713 r0 *1 92.815,17.01
X$8713 310 VIA_via2_5
* cell instance $8714 r0 *1 94.905,18.83
X$8714 310 VIA_via2_5
* cell instance $8715 r0 *1 88.635,17.57
X$8715 310 VIA_via1_4
* cell instance $8716 r0 *1 88.635,17.57
X$8716 310 VIA_via2_5
* cell instance $8717 r0 *1 95.095,14.77
X$8717 310 VIA_via1_4
* cell instance $8718 r0 *1 93.195,16.03
X$8718 310 VIA_via1_4
* cell instance $8719 r0 *1 94.905,20.37
X$8719 310 VIA_via1_4
* cell instance $8720 r0 *1 94.715,21.63
X$8720 310 VIA_via1_4
* cell instance $8721 r0 *1 92.815,18.83
X$8721 310 VIA_via1_4
* cell instance $8722 r0 *1 92.815,18.83
X$8722 310 VIA_via2_5
* cell instance $8723 r0 *1 89.775,20.37
X$8723 310 VIA_via1_4
* cell instance $8724 r0 *1 86.735,16.03
X$8724 310 VIA_via1_4
* cell instance $8725 r0 *1 96.045,15.61
X$8725 311 VIA_via1_7
* cell instance $8726 r0 *1 96.045,14.77
X$8726 311 VIA_via2_5
* cell instance $8727 r0 *1 94.335,14.77
X$8727 311 VIA_via1_4
* cell instance $8728 r0 *1 94.335,14.77
X$8728 311 VIA_via2_5
* cell instance $8729 r0 *1 5.225,15.61
X$8729 312 VIA_via1_7
* cell instance $8730 r0 *1 5.225,14.77
X$8730 312 VIA_via2_5
* cell instance $8731 r0 *1 3.705,14.77
X$8731 312 VIA_via1_4
* cell instance $8732 r0 *1 3.705,14.77
X$8732 312 VIA_via2_5
* cell instance $8733 r0 *1 93.385,14.91
X$8733 313 VIA_via2_5
* cell instance $8734 r0 *1 94.715,14.91
X$8734 313 VIA_via2_5
* cell instance $8735 r0 *1 93.195,17.57
X$8735 313 VIA_via1_4
* cell instance $8736 r0 *1 92.625,14.77
X$8736 313 VIA_via1_4
* cell instance $8737 r0 *1 92.625,14.91
X$8737 313 VIA_via2_5
* cell instance $8738 r0 *1 94.715,15.75
X$8738 313 VIA_via1_4
* cell instance $8739 r0 *1 81.035,13.79
X$8739 314 VIA_via1_7
* cell instance $8740 r0 *1 81.035,14.77
X$8740 314 VIA_via2_5
* cell instance $8741 r0 *1 79.705,14.77
X$8741 314 VIA_via1_4
* cell instance $8742 r0 *1 79.705,14.77
X$8742 314 VIA_via2_5
* cell instance $8743 r0 *1 69.255,14.77
X$8743 315 VIA_via2_5
* cell instance $8744 r0 *1 67.735,14.77
X$8744 315 VIA_via1_4
* cell instance $8745 r0 *1 67.735,14.77
X$8745 315 VIA_via2_5
* cell instance $8746 r0 *1 69.255,13.65
X$8746 315 VIA_via1_4
* cell instance $8747 r0 *1 68.875,16.03
X$8747 315 VIA_via1_4
* cell instance $8748 r0 *1 64.695,14.77
X$8748 316 VIA_via2_5
* cell instance $8749 r0 *1 64.315,14.77
X$8749 316 VIA_via1_4
* cell instance $8750 r0 *1 64.315,14.77
X$8750 316 VIA_via2_5
* cell instance $8751 r0 *1 65.075,14.77
X$8751 316 VIA_via1_4
* cell instance $8752 r0 *1 65.075,14.77
X$8752 316 VIA_via2_5
* cell instance $8753 r0 *1 64.695,13.23
X$8753 316 VIA_via1_4
* cell instance $8754 r0 *1 39.805,14.91
X$8754 317 VIA_via1_4
* cell instance $8755 r0 *1 39.805,14.91
X$8755 317 VIA_via2_5
* cell instance $8756 r0 *1 35.815,14.77
X$8756 317 VIA_via1_4
* cell instance $8757 r0 *1 35.815,14.91
X$8757 317 VIA_via2_5
* cell instance $8758 r0 *1 24.415,16.17
X$8758 318 VIA_via1_7
* cell instance $8759 r0 *1 24.415,16.17
X$8759 318 VIA_via2_5
* cell instance $8760 r0 *1 4.085,16.17
X$8760 318 VIA_via1_7
* cell instance $8761 r0 *1 8.645,20.23
X$8761 318 VIA_via1_7
* cell instance $8762 r0 *1 8.645,20.09
X$8762 318 VIA_via2_5
* cell instance $8763 r0 *1 48.165,14.63
X$8763 318 VIA_via1_7
* cell instance $8764 r0 *1 48.165,14.63
X$8764 318 VIA_via2_5
* cell instance $8765 r0 *1 28.215,16.17
X$8765 318 VIA_via1_7
* cell instance $8766 r0 *1 28.215,16.17
X$8766 318 VIA_via2_5
* cell instance $8767 r0 *1 29.735,16.31
X$8767 318 VIA_via2_5
* cell instance $8768 r0 *1 29.735,17.85
X$8768 318 VIA_via2_5
* cell instance $8769 r0 *1 37.525,17.85
X$8769 318 VIA_via2_5
* cell instance $8770 r0 *1 4.275,21.63
X$8770 318 VIA_via2_5
* cell instance $8771 r0 *1 4.275,20.09
X$8771 318 VIA_via2_5
* cell instance $8772 r0 *1 23.275,19.25
X$8772 318 VIA_via2_5
* cell instance $8773 r0 *1 23.275,16.17
X$8773 318 VIA_via2_5
* cell instance $8774 r0 *1 8.645,19.39
X$8774 318 VIA_via2_5
* cell instance $8775 r0 *1 43.605,17.57
X$8775 318 VIA_via1_4
* cell instance $8776 r0 *1 43.605,17.71
X$8776 318 VIA_via2_5
* cell instance $8777 r0 *1 4.085,24.43
X$8777 318 VIA_via1_4
* cell instance $8778 r0 *1 37.525,17.57
X$8778 318 VIA_via1_4
* cell instance $8779 r0 *1 3.705,21.63
X$8779 318 VIA_via1_4
* cell instance $8780 r0 *1 3.705,21.63
X$8780 318 VIA_via2_5
* cell instance $8781 r0 *1 48.925,24.15
X$8781 318 VIA_via1_4
* cell instance $8782 r0 *1 48.925,24.15
X$8782 318 VIA_via2_5
* cell instance $8783 r0 *1 29.735,21.63
X$8783 318 VIA_via1_4
* cell instance $8784 r0 *1 48.535,14.63
X$8784 318 VIA_via3_2
* cell instance $8785 r0 *1 48.535,24.15
X$8785 318 VIA_via3_2
* cell instance $8786 r0 *1 48.535,17.71
X$8786 318 VIA_via3_2
* cell instance $8787 r0 *1 39.805,17.99
X$8787 319 VIA_via1_7
* cell instance $8788 r0 *1 37.525,45.57
X$8788 319 VIA_via2_5
* cell instance $8789 r0 *1 36.765,23.17
X$8789 319 VIA_via2_5
* cell instance $8790 r0 *1 38.285,23.45
X$8790 319 VIA_via2_5
* cell instance $8791 r0 *1 36.575,45.43
X$8791 319 VIA_via2_5
* cell instance $8792 r0 *1 38.285,17.99
X$8792 319 VIA_via2_5
* cell instance $8793 r0 *1 39.615,17.99
X$8793 319 VIA_via2_5
* cell instance $8794 r0 *1 38.285,14.77
X$8794 319 VIA_via2_5
* cell instance $8795 r0 *1 39.615,23.45
X$8795 319 VIA_via2_5
* cell instance $8796 r0 *1 39.615,23.17
X$8796 319 VIA_via1_4
* cell instance $8797 r0 *1 39.425,14.77
X$8797 319 VIA_via1_4
* cell instance $8798 r0 *1 39.425,14.77
X$8798 319 VIA_via2_5
* cell instance $8799 r0 *1 38.285,23.17
X$8799 319 VIA_via1_4
* cell instance $8800 r0 *1 38.285,23.17
X$8800 319 VIA_via2_5
* cell instance $8801 r0 *1 38.285,17.57
X$8801 319 VIA_via1_4
* cell instance $8802 r0 *1 38.475,45.57
X$8802 319 VIA_via1_4
* cell instance $8803 r0 *1 38.475,45.57
X$8803 319 VIA_via2_5
* cell instance $8804 r0 *1 36.575,46.83
X$8804 319 VIA_via1_4
* cell instance $8805 r0 *1 41.705,45.57
X$8805 319 VIA_via1_4
* cell instance $8806 r0 *1 41.705,45.57
X$8806 319 VIA_via2_5
* cell instance $8807 r0 *1 40.185,45.57
X$8807 319 VIA_via1_4
* cell instance $8808 r0 *1 40.185,45.57
X$8808 319 VIA_via2_5
* cell instance $8809 r0 *1 36.575,35.63
X$8809 319 VIA_via1_4
* cell instance $8810 r0 *1 36.765,28.77
X$8810 319 VIA_via1_4
* cell instance $8811 r0 *1 42.465,14.77
X$8811 320 VIA_via1_4
* cell instance $8812 r0 *1 42.465,14.77
X$8812 320 VIA_via2_5
* cell instance $8813 r0 *1 46.075,14.77
X$8813 320 VIA_via1_4
* cell instance $8814 r0 *1 46.075,14.77
X$8814 320 VIA_via2_5
* cell instance $8815 r0 *1 15.105,13.79
X$8815 321 VIA_via1_7
* cell instance $8816 r0 *1 15.675,16.03
X$8816 321 VIA_via1_4
* cell instance $8817 r0 *1 16.815,20.37
X$8817 322 VIA_via1_4
* cell instance $8818 r0 *1 15.865,15.75
X$8818 322 VIA_via1_4
* cell instance $8819 r0 *1 18.145,13.51
X$8819 323 VIA_via1_4
* cell instance $8820 r0 *1 17.955,16.03
X$8820 323 VIA_via1_4
* cell instance $8821 r0 *1 27.265,20.37
X$8821 324 VIA_via2_5
* cell instance $8822 r0 *1 22.515,20.37
X$8822 324 VIA_via2_5
* cell instance $8823 r0 *1 24.035,20.37
X$8823 324 VIA_via2_5
* cell instance $8824 r0 *1 24.035,16.03
X$8824 324 VIA_via2_5
* cell instance $8825 r0 *1 27.265,21.63
X$8825 324 VIA_via1_4
* cell instance $8826 r0 *1 25.175,20.37
X$8826 324 VIA_via1_4
* cell instance $8827 r0 *1 25.365,20.37
X$8827 324 VIA_via1_4
* cell instance $8828 r0 *1 25.365,20.37
X$8828 324 VIA_via2_5
* cell instance $8829 r0 *1 27.645,20.37
X$8829 324 VIA_via1_4
* cell instance $8830 r0 *1 22.515,21.63
X$8830 324 VIA_via1_4
* cell instance $8831 r0 *1 21.945,20.37
X$8831 324 VIA_via1_4
* cell instance $8832 r0 *1 21.945,20.37
X$8832 324 VIA_via2_5
* cell instance $8833 r0 *1 22.705,16.03
X$8833 324 VIA_via1_4
* cell instance $8834 r0 *1 22.705,16.03
X$8834 324 VIA_via2_5
* cell instance $8835 r0 *1 24.035,14.77
X$8835 324 VIA_via1_4
* cell instance $8836 r0 *1 20.045,16.03
X$8836 325 VIA_via1_4
* cell instance $8837 r0 *1 20.045,15.89
X$8837 325 VIA_via2_5
* cell instance $8838 r0 *1 24.225,15.89
X$8838 325 VIA_via1_4
* cell instance $8839 r0 *1 24.225,15.89
X$8839 325 VIA_via2_5
* cell instance $8840 r0 *1 26.695,16.03
X$8840 325 VIA_via1_4
* cell instance $8841 r0 *1 26.695,15.89
X$8841 325 VIA_via2_5
* cell instance $8842 r0 *1 25.555,15.61
X$8842 326 VIA_via1_7
* cell instance $8843 r0 *1 25.555,15.61
X$8843 326 VIA_via2_5
* cell instance $8844 r0 *1 23.275,15.33
X$8844 326 VIA_via2_5
* cell instance $8845 r0 *1 23.275,14.77
X$8845 326 VIA_via1_4
* cell instance $8846 r0 *1 26.125,17.57
X$8846 327 VIA_via1_4
* cell instance $8847 r0 *1 26.695,13.51
X$8847 327 VIA_via1_4
* cell instance $8848 r0 *1 30.305,15.75
X$8848 328 VIA_via2_5
* cell instance $8849 r0 *1 34.675,15.75
X$8849 328 VIA_via1_4
* cell instance $8850 r0 *1 34.675,15.75
X$8850 328 VIA_via2_5
* cell instance $8851 r0 *1 30.305,17.57
X$8851 328 VIA_via1_4
* cell instance $8852 r0 *1 30.305,16.03
X$8852 328 VIA_via1_4
* cell instance $8853 r0 *1 35.815,20.37
X$8853 329 VIA_via2_5
* cell instance $8854 r0 *1 33.725,24.43
X$8854 329 VIA_via2_5
* cell instance $8855 r0 *1 33.725,23.17
X$8855 329 VIA_via2_5
* cell instance $8856 r0 *1 29.545,24.43
X$8856 329 VIA_via2_5
* cell instance $8857 r0 *1 37.335,20.37
X$8857 329 VIA_via2_5
* cell instance $8858 r0 *1 39.425,20.37
X$8858 329 VIA_via2_5
* cell instance $8859 r0 *1 37.145,16.03
X$8859 329 VIA_via1_4
* cell instance $8860 r0 *1 33.725,23.45
X$8860 329 VIA_via1_4
* cell instance $8861 r0 *1 33.345,24.43
X$8861 329 VIA_via1_4
* cell instance $8862 r0 *1 33.345,24.43
X$8862 329 VIA_via2_5
* cell instance $8863 r0 *1 35.815,23.17
X$8863 329 VIA_via1_4
* cell instance $8864 r0 *1 35.815,23.17
X$8864 329 VIA_via2_5
* cell instance $8865 r0 *1 39.425,21.63
X$8865 329 VIA_via1_4
* cell instance $8866 r0 *1 39.045,20.37
X$8866 329 VIA_via1_4
* cell instance $8867 r0 *1 39.045,20.37
X$8867 329 VIA_via2_5
* cell instance $8868 r0 *1 29.545,23.17
X$8868 329 VIA_via1_4
* cell instance $8869 r0 *1 34.295,20.37
X$8869 329 VIA_via1_4
* cell instance $8870 r0 *1 34.295,20.37
X$8870 329 VIA_via2_5
* cell instance $8871 r0 *1 29.355,27.23
X$8871 329 VIA_via1_4
* cell instance $8872 r0 *1 38.095,16.03
X$8872 330 VIA_via2_5
* cell instance $8873 r0 *1 38.855,16.03
X$8873 330 VIA_via2_5
* cell instance $8874 r0 *1 38.095,15.05
X$8874 330 VIA_via1_4
* cell instance $8875 r0 *1 39.805,16.03
X$8875 330 VIA_via1_4
* cell instance $8876 r0 *1 39.805,16.03
X$8876 330 VIA_via2_5
* cell instance $8877 r0 *1 38.855,14.77
X$8877 330 VIA_via1_4
* cell instance $8878 r0 *1 40.945,13.51
X$8878 331 VIA_via1_4
* cell instance $8879 r0 *1 41.135,17.57
X$8879 331 VIA_via1_4
* cell instance $8880 r0 *1 55.765,15.61
X$8880 332 VIA_via1_7
* cell instance $8881 r0 *1 54.815,14.77
X$8881 332 VIA_via1_4
* cell instance $8882 r0 *1 60.515,16.03
X$8882 333 VIA_via2_5
* cell instance $8883 r0 *1 60.515,15.05
X$8883 333 VIA_via1_4
* cell instance $8884 r0 *1 58.045,16.03
X$8884 333 VIA_via1_4
* cell instance $8885 r0 *1 58.045,16.03
X$8885 333 VIA_via2_5
* cell instance $8886 r0 *1 56.715,16.03
X$8886 333 VIA_via1_4
* cell instance $8887 r0 *1 56.715,15.89
X$8887 333 VIA_via2_5
* cell instance $8888 r0 *1 73.625,16.03
X$8888 334 VIA_via2_5
* cell instance $8889 r0 *1 74.955,16.03
X$8889 334 VIA_via2_5
* cell instance $8890 r0 *1 80.465,16.03
X$8890 334 VIA_via2_5
* cell instance $8891 r0 *1 72.295,20.37
X$8891 334 VIA_via2_5
* cell instance $8892 r0 *1 70.395,16.03
X$8892 334 VIA_via2_5
* cell instance $8893 r0 *1 74.955,20.37
X$8893 334 VIA_via1_4
* cell instance $8894 r0 *1 74.955,20.37
X$8894 334 VIA_via2_5
* cell instance $8895 r0 *1 80.465,14.77
X$8895 334 VIA_via1_4
* cell instance $8896 r0 *1 74.765,16.03
X$8896 334 VIA_via1_4
* cell instance $8897 r0 *1 74.765,16.03
X$8897 334 VIA_via2_5
* cell instance $8898 r0 *1 77.995,16.03
X$8898 334 VIA_via1_4
* cell instance $8899 r0 *1 77.995,16.03
X$8899 334 VIA_via2_5
* cell instance $8900 r0 *1 73.625,17.57
X$8900 334 VIA_via1_4
* cell instance $8901 r0 *1 67.735,20.37
X$8901 334 VIA_via1_4
* cell instance $8902 r0 *1 67.735,20.37
X$8902 334 VIA_via2_5
* cell instance $8903 r0 *1 72.865,20.37
X$8903 334 VIA_via1_4
* cell instance $8904 r0 *1 72.865,20.37
X$8904 334 VIA_via2_5
* cell instance $8905 r0 *1 72.295,21.63
X$8905 334 VIA_via1_4
* cell instance $8906 r0 *1 70.395,14.77
X$8906 334 VIA_via1_4
* cell instance $8907 r0 *1 93.005,15.19
X$8907 335 VIA_via1_7
* cell instance $8908 r0 *1 92.435,16.03
X$8908 335 VIA_via1_4
* cell instance $8909 r0 *1 96.615,16.03
X$8909 336 VIA_via2_5
* cell instance $8910 r0 *1 93.765,16.03
X$8910 336 VIA_via2_5
* cell instance $8911 r0 *1 95.665,16.03
X$8911 336 VIA_via1_4
* cell instance $8912 r0 *1 95.665,16.03
X$8912 336 VIA_via2_5
* cell instance $8913 r0 *1 93.765,17.57
X$8913 336 VIA_via1_4
* cell instance $8914 r0 *1 96.615,15.05
X$8914 336 VIA_via1_4
* cell instance $8915 r0 *1 6.555,16.03
X$8915 337 VIA_via1_4
* cell instance $8916 r0 *1 6.555,16.03
X$8916 337 VIA_via2_5
* cell instance $8917 r0 *1 10.545,16.03
X$8917 337 VIA_via1_4
* cell instance $8918 r0 *1 10.545,16.03
X$8918 337 VIA_via2_5
* cell instance $8919 r0 *1 16.815,16.87
X$8919 338 VIA_via2_5
* cell instance $8920 r0 *1 17.385,16.73
X$8920 338 VIA_via2_5
* cell instance $8921 r0 *1 15.675,15.19
X$8921 338 VIA_via2_5
* cell instance $8922 r0 *1 17.385,15.19
X$8922 338 VIA_via2_5
* cell instance $8923 r0 *1 15.675,14.63
X$8923 338 VIA_via1_4
* cell instance $8924 r0 *1 17.005,20.37
X$8924 338 VIA_via1_4
* cell instance $8925 r0 *1 10.735,15.89
X$8925 339 VIA_via1_4
* cell instance $8926 r0 *1 10.735,15.89
X$8926 339 VIA_via2_5
* cell instance $8927 r0 *1 17.195,16.03
X$8927 339 VIA_via1_4
* cell instance $8928 r0 *1 17.195,15.89
X$8928 339 VIA_via2_5
* cell instance $8929 r0 *1 20.235,51.59
X$8929 340 VIA_via2_5
* cell instance $8930 r0 *1 20.045,53.97
X$8930 340 VIA_via1_4
* cell instance $8931 r0 *1 15.865,51.17
X$8931 340 VIA_via1_4
* cell instance $8932 r0 *1 15.865,51.03
X$8932 340 VIA_via2_5
* cell instance $8933 r0 *1 17.955,15.75
X$8933 340 VIA_via1_4
* cell instance $8934 r0 *1 17.955,15.75
X$8934 340 VIA_via2_5
* cell instance $8935 r0 *1 18.015,15.75
X$8935 340 VIA_via3_2
* cell instance $8936 r0 *1 18.015,51.03
X$8936 340 VIA_via3_2
* cell instance $8937 r0 *1 21.945,16.03
X$8937 341 VIA_via1_4
* cell instance $8938 r0 *1 21.945,16.03
X$8938 341 VIA_via2_5
* cell instance $8939 r0 *1 20.995,16.03
X$8939 341 VIA_via1_4
* cell instance $8940 r0 *1 20.995,16.03
X$8940 341 VIA_via2_5
* cell instance $8941 r0 *1 87.115,16.03
X$8941 342 VIA_via2_5
* cell instance $8942 r0 *1 85.975,16.03
X$8942 342 VIA_via1_4
* cell instance $8943 r0 *1 85.975,16.03
X$8943 342 VIA_via2_5
* cell instance $8944 r0 *1 87.115,14.63
X$8944 342 VIA_via1_4
* cell instance $8945 r0 *1 29.355,15.61
X$8945 343 VIA_via1_7
* cell instance $8946 r0 *1 29.355,15.61
X$8946 343 VIA_via2_5
* cell instance $8947 r0 *1 27.455,15.61
X$8947 343 VIA_via2_5
* cell instance $8948 r0 *1 27.455,14.77
X$8948 343 VIA_via1_4
* cell instance $8949 r0 *1 28.405,16.03
X$8949 344 VIA_via1_4
* cell instance $8950 r0 *1 28.405,16.03
X$8950 344 VIA_via2_5
* cell instance $8951 r0 *1 29.735,16.03
X$8951 344 VIA_via1_4
* cell instance $8952 r0 *1 29.735,16.03
X$8952 344 VIA_via2_5
* cell instance $8953 r0 *1 29.735,15.05
X$8953 344 VIA_via1_4
* cell instance $8954 r0 *1 69.445,15.05
X$8954 345 VIA_via2_5
* cell instance $8955 r0 *1 70.585,15.05
X$8955 345 VIA_via2_5
* cell instance $8956 r0 *1 70.585,13.23
X$8956 345 VIA_via1_4
* cell instance $8957 r0 *1 71.915,15.05
X$8957 345 VIA_via1_4
* cell instance $8958 r0 *1 71.915,15.05
X$8958 345 VIA_via2_5
* cell instance $8959 r0 *1 69.445,16.03
X$8959 345 VIA_via1_4
* cell instance $8960 r0 *1 31.065,16.03
X$8960 346 VIA_via1_4
* cell instance $8961 r0 *1 30.685,16.03
X$8961 346 VIA_via1_4
* cell instance $8962 r0 *1 63.555,17.01
X$8962 347 VIA_via1_7
* cell instance $8963 r0 *1 63.175,16.03
X$8963 347 VIA_via2_5
* cell instance $8964 r0 *1 63.555,16.03
X$8964 347 VIA_via2_5
* cell instance $8965 r0 *1 62.985,16.03
X$8965 347 VIA_via1_4
* cell instance $8966 r0 *1 40.185,16.03
X$8966 348 VIA_via1_4
* cell instance $8967 r0 *1 40.375,16.03
X$8967 348 VIA_via1_4
* cell instance $8968 r0 *1 57.095,15.61
X$8968 349 VIA_via1_7
* cell instance $8969 r0 *1 58.235,15.33
X$8969 349 VIA_via2_5
* cell instance $8970 r0 *1 57.095,15.33
X$8970 349 VIA_via2_5
* cell instance $8971 r0 *1 58.235,14.77
X$8971 349 VIA_via1_4
* cell instance $8972 r0 *1 44.745,17.01
X$8972 350 VIA_via1_7
* cell instance $8973 r0 *1 44.745,16.03
X$8973 350 VIA_via2_5
* cell instance $8974 r0 *1 41.705,16.03
X$8974 350 VIA_via1_4
* cell instance $8975 r0 *1 41.705,16.03
X$8975 350 VIA_via2_5
* cell instance $8976 r0 *1 45.885,16.03
X$8976 351 VIA_via1_4
* cell instance $8977 r0 *1 45.885,6.23
X$8977 351 VIA_via1_4
* cell instance $8978 r0 *1 49.305,18.41
X$8978 352 VIA_via1_7
* cell instance $8979 r0 *1 49.305,16.03
X$8979 352 VIA_via2_5
* cell instance $8980 r0 *1 47.975,16.03
X$8980 352 VIA_via1_4
* cell instance $8981 r0 *1 47.975,16.03
X$8981 352 VIA_via2_5
* cell instance $8982 r0 *1 51.775,15.19
X$8982 353 VIA_via1_7
* cell instance $8983 r0 *1 51.775,16.03
X$8983 353 VIA_via1_4
* cell instance $8984 r0 *1 11.305,61.95
X$8984 354 VIA_via2_5
* cell instance $8985 r0 *1 11.115,69.51
X$8985 354 VIA_via2_5
* cell instance $8986 r0 *1 11.875,69.51
X$8986 354 VIA_via2_5
* cell instance $8987 r0 *1 10.545,69.51
X$8987 354 VIA_via2_5
* cell instance $8988 r0 *1 32.775,16.87
X$8988 354 VIA_via2_5
* cell instance $8989 r0 *1 31.445,16.31
X$8989 354 VIA_via2_5
* cell instance $8990 r0 *1 27.075,16.87
X$8990 354 VIA_via2_5
* cell instance $8991 r0 *1 11.305,20.23
X$8991 354 VIA_via2_5
* cell instance $8992 r0 *1 15.675,16.87
X$8992 354 VIA_via2_5
* cell instance $8993 r0 *1 10.925,16.73
X$8993 354 VIA_via2_5
* cell instance $8994 r0 *1 15.675,17.71
X$8994 354 VIA_via2_5
* cell instance $8995 r0 *1 10.355,20.37
X$8995 354 VIA_via1_4
* cell instance $8996 r0 *1 10.355,20.23
X$8996 354 VIA_via2_5
* cell instance $8997 r0 *1 11.305,21.63
X$8997 354 VIA_via1_4
* cell instance $8998 r0 *1 10.925,16.03
X$8998 354 VIA_via1_4
* cell instance $8999 r0 *1 31.445,16.03
X$8999 354 VIA_via1_4
* cell instance $9000 r0 *1 32.585,20.37
X$9000 354 VIA_via1_4
* cell instance $9001 r0 *1 32.585,20.37
X$9001 354 VIA_via2_5
* cell instance $9002 r0 *1 27.075,17.57
X$9002 354 VIA_via1_4
* cell instance $9003 r0 *1 27.075,17.71
X$9003 354 VIA_via2_5
* cell instance $9004 r0 *1 11.305,53.97
X$9004 354 VIA_via1_4
* cell instance $9005 r0 *1 11.875,70.77
X$9005 354 VIA_via1_4
* cell instance $9006 r0 *1 11.115,69.23
X$9006 354 VIA_via1_4
* cell instance $9007 r0 *1 32.015,61.95
X$9007 354 VIA_via1_4
* cell instance $9008 r0 *1 32.015,61.95
X$9008 354 VIA_via2_5
* cell instance $9009 r0 *1 16.245,17.57
X$9009 354 VIA_via1_4
* cell instance $9010 r0 *1 16.245,17.71
X$9010 354 VIA_via2_5
* cell instance $9011 r0 *1 32.855,61.95
X$9011 354 VIA_via3_2
* cell instance $9012 r0 *1 10.735,20.23
X$9012 354 VIA_via3_2
* cell instance $9013 r0 *1 10.735,16.73
X$9013 354 VIA_via3_2
* cell instance $9014 r0 *1 32.855,20.37
X$9014 354 VIA_via3_2
* cell instance $9015 r0 *1 32.775,20.37
X$9015 354 VIA_via2_5
* cell instance $9016 r0 *1 16.055,18.41
X$9016 355 VIA_via1_7
* cell instance $9017 r0 *1 16.245,16.03
X$9017 355 VIA_via1_4
* cell instance $9018 r0 *1 53.295,21.21
X$9018 356 VIA_via1_7
* cell instance $9019 r0 *1 52.155,18.13
X$9019 356 VIA_via2_5
* cell instance $9020 r0 *1 53.295,18.13
X$9020 356 VIA_via2_5
* cell instance $9021 r0 *1 34.105,17.99
X$9021 356 VIA_via2_5
* cell instance $9022 r0 *1 40.185,18.13
X$9022 356 VIA_via2_5
* cell instance $9023 r0 *1 31.445,17.99
X$9023 356 VIA_via2_5
* cell instance $9024 r0 *1 24.985,17.99
X$9024 356 VIA_via2_5
* cell instance $9025 r0 *1 44.365,18.13
X$9025 356 VIA_via2_5
* cell instance $9026 r0 *1 24.985,17.29
X$9026 356 VIA_via2_5
* cell instance $9027 r0 *1 15.865,20.65
X$9027 356 VIA_via2_5
* cell instance $9028 r0 *1 17.005,17.43
X$9028 356 VIA_via2_5
* cell instance $9029 r0 *1 17.005,18.41
X$9029 356 VIA_via2_5
* cell instance $9030 r0 *1 15.865,18.41
X$9030 356 VIA_via2_5
* cell instance $9031 r0 *1 12.635,20.65
X$9031 356 VIA_via2_5
* cell instance $9032 r0 *1 40.185,17.57
X$9032 356 VIA_via1_4
* cell instance $9033 r0 *1 44.365,18.83
X$9033 356 VIA_via1_4
* cell instance $9034 r0 *1 34.105,18.83
X$9034 356 VIA_via1_4
* cell instance $9035 r0 *1 31.445,17.57
X$9035 356 VIA_via1_4
* cell instance $9036 r0 *1 24.985,17.57
X$9036 356 VIA_via1_4
* cell instance $9037 r0 *1 52.155,17.57
X$9037 356 VIA_via1_4
* cell instance $9038 r0 *1 12.635,23.17
X$9038 356 VIA_via1_4
* cell instance $9039 r0 *1 20.615,17.57
X$9039 356 VIA_via1_4
* cell instance $9040 r0 *1 20.615,17.43
X$9040 356 VIA_via2_5
* cell instance $9041 r0 *1 15.865,20.37
X$9041 356 VIA_via1_4
* cell instance $9042 r0 *1 16.815,16.03
X$9042 356 VIA_via1_4
* cell instance $9043 r0 *1 17.005,16.31
X$9043 357 VIA_via2_5
* cell instance $9044 r0 *1 17.005,16.03
X$9044 357 VIA_via1_4
* cell instance $9045 r0 *1 16.625,16.45
X$9045 357 VIA_via1_4
* cell instance $9046 r0 *1 16.625,16.45
X$9046 357 VIA_via2_5
* cell instance $9047 r0 *1 25.175,16.45
X$9047 358 VIA_via2_5
* cell instance $9048 r0 *1 23.275,42.49
X$9048 358 VIA_via2_5
* cell instance $9049 r0 *1 22.135,42.49
X$9049 358 VIA_via2_5
* cell instance $9050 r0 *1 23.655,26.11
X$9050 358 VIA_via2_5
* cell instance $9051 r0 *1 24.415,26.11
X$9051 358 VIA_via2_5
* cell instance $9052 r0 *1 20.425,26.11
X$9052 358 VIA_via2_5
* cell instance $9053 r0 *1 20.615,16.45
X$9053 358 VIA_via2_5
* cell instance $9054 r0 *1 20.425,34.37
X$9054 358 VIA_via2_5
* cell instance $9055 r0 *1 22.325,34.37
X$9055 358 VIA_via2_5
* cell instance $9056 r0 *1 20.235,16.45
X$9056 358 VIA_via2_5
* cell instance $9057 r0 *1 20.615,16.03
X$9057 358 VIA_via1_4
* cell instance $9058 r0 *1 25.175,16.03
X$9058 358 VIA_via1_4
* cell instance $9059 r0 *1 20.425,35.63
X$9059 358 VIA_via1_4
* cell instance $9060 r0 *1 22.515,38.43
X$9060 358 VIA_via1_4
* cell instance $9061 r0 *1 21.945,42.77
X$9061 358 VIA_via1_4
* cell instance $9062 r0 *1 23.275,42.77
X$9062 358 VIA_via1_4
* cell instance $9063 r0 *1 24.415,23.17
X$9063 358 VIA_via1_4
* cell instance $9064 r0 *1 20.425,21.63
X$9064 358 VIA_via1_4
* cell instance $9065 r0 *1 23.655,34.37
X$9065 358 VIA_via1_4
* cell instance $9066 r0 *1 23.655,34.37
X$9066 358 VIA_via2_5
* cell instance $9067 r0 *1 22.135,25.97
X$9067 358 VIA_via1_4
* cell instance $9068 r0 *1 22.135,26.11
X$9068 358 VIA_via2_5
* cell instance $9069 r0 *1 23.655,28.77
X$9069 358 VIA_via1_4
* cell instance $9070 r0 *1 20.805,17.57
X$9070 359 VIA_via1_4
* cell instance $9071 r0 *1 20.425,17.15
X$9071 359 VIA_via1_4
* cell instance $9072 r0 *1 58.615,21.49
X$9072 360 VIA_via2_5
* cell instance $9073 r0 *1 57.665,21.49
X$9073 360 VIA_via2_5
* cell instance $9074 r0 *1 52.915,18.27
X$9074 360 VIA_via2_5
* cell instance $9075 r0 *1 57.665,17.71
X$9075 360 VIA_via2_5
* cell instance $9076 r0 *1 45.125,18.27
X$9076 360 VIA_via2_5
* cell instance $9077 r0 *1 32.205,18.55
X$9077 360 VIA_via2_5
* cell instance $9078 r0 *1 40.945,18.69
X$9078 360 VIA_via2_5
* cell instance $9079 r0 *1 40.945,18.27
X$9079 360 VIA_via2_5
* cell instance $9080 r0 *1 17.575,17.57
X$9080 360 VIA_via2_5
* cell instance $9081 r0 *1 16.435,19.11
X$9081 360 VIA_via2_5
* cell instance $9082 r0 *1 17.575,19.11
X$9082 360 VIA_via2_5
* cell instance $9083 r0 *1 40.945,17.57
X$9083 360 VIA_via1_4
* cell instance $9084 r0 *1 21.375,17.57
X$9084 360 VIA_via1_4
* cell instance $9085 r0 *1 21.375,17.57
X$9085 360 VIA_via2_5
* cell instance $9086 r0 *1 45.125,18.83
X$9086 360 VIA_via1_4
* cell instance $9087 r0 *1 34.865,18.83
X$9087 360 VIA_via1_4
* cell instance $9088 r0 *1 34.865,18.69
X$9088 360 VIA_via2_5
* cell instance $9089 r0 *1 32.205,17.57
X$9089 360 VIA_via1_4
* cell instance $9090 r0 *1 32.205,17.57
X$9090 360 VIA_via2_5
* cell instance $9091 r0 *1 25.745,17.57
X$9091 360 VIA_via1_4
* cell instance $9092 r0 *1 25.745,17.43
X$9092 360 VIA_via2_5
* cell instance $9093 r0 *1 58.805,21.63
X$9093 360 VIA_via1_4
* cell instance $9094 r0 *1 58.425,22.75
X$9094 360 VIA_via1_4
* cell instance $9095 r0 *1 52.915,17.57
X$9095 360 VIA_via1_4
* cell instance $9096 r0 *1 52.915,17.71
X$9096 360 VIA_via2_5
* cell instance $9097 r0 *1 16.625,20.37
X$9097 360 VIA_via1_4
* cell instance $9098 r0 *1 17.575,16.03
X$9098 360 VIA_via1_4
* cell instance $9099 r0 *1 25.935,17.57
X$9099 361 VIA_via1_4
* cell instance $9100 r0 *1 26.315,14.63
X$9100 361 VIA_via1_4
* cell instance $9101 r0 *1 27.075,16.59
X$9101 362 VIA_via1_7
* cell instance $9102 r0 *1 26.695,17.57
X$9102 362 VIA_via1_4
* cell instance $9103 r0 *1 31.445,16.59
X$9103 363 VIA_via1_7
* cell instance $9104 r0 *1 31.825,17.57
X$9104 363 VIA_via1_4
* cell instance $9105 r0 *1 32.395,17.57
X$9105 364 VIA_via1_4
* cell instance $9106 r0 *1 32.585,13.51
X$9106 364 VIA_via1_4
* cell instance $9107 r0 *1 32.205,13.79
X$9107 365 VIA_via1_7
* cell instance $9108 r0 *1 32.205,17.29
X$9108 365 VIA_via2_5
* cell instance $9109 r0 *1 32.585,17.57
X$9109 365 VIA_via1_4
* cell instance $9110 r0 *1 32.585,17.57
X$9110 365 VIA_via2_5
* cell instance $9111 r0 *1 38.475,17.57
X$9111 366 VIA_via2_5
* cell instance $9112 r0 *1 38.665,16.45
X$9112 366 VIA_via1_4
* cell instance $9113 r0 *1 39.235,16.03
X$9113 366 VIA_via1_4
* cell instance $9114 r0 *1 37.715,17.57
X$9114 366 VIA_via1_4
* cell instance $9115 r0 *1 37.715,17.57
X$9115 366 VIA_via2_5
* cell instance $9116 r0 *1 55.765,40.39
X$9116 367 VIA_via1_7
* cell instance $9117 r0 *1 55.765,40.39
X$9117 367 VIA_via2_5
* cell instance $9118 r0 *1 58.235,18.41
X$9118 367 VIA_via2_5
* cell instance $9119 r0 *1 60.135,20.37
X$9119 367 VIA_via2_5
* cell instance $9120 r0 *1 60.135,24.01
X$9120 367 VIA_via2_5
* cell instance $9121 r0 *1 76.095,22.89
X$9121 367 VIA_via2_5
* cell instance $9122 r0 *1 68.495,40.39
X$9122 367 VIA_via2_5
* cell instance $9123 r0 *1 70.205,23.03
X$9123 367 VIA_via2_5
* cell instance $9124 r0 *1 70.205,23.31
X$9124 367 VIA_via2_5
* cell instance $9125 r0 *1 45.315,16.87
X$9125 367 VIA_via2_5
* cell instance $9126 r0 *1 40.755,16.73
X$9126 367 VIA_via2_5
* cell instance $9127 r0 *1 59.375,40.39
X$9127 367 VIA_via2_5
* cell instance $9128 r0 *1 65.075,24.01
X$9128 367 VIA_via2_5
* cell instance $9129 r0 *1 45.315,17.57
X$9129 367 VIA_via1_4
* cell instance $9130 r0 *1 40.755,16.03
X$9130 367 VIA_via1_4
* cell instance $9131 r0 *1 75.525,23.17
X$9131 367 VIA_via1_4
* cell instance $9132 r0 *1 75.525,23.03
X$9132 367 VIA_via2_5
* cell instance $9133 r0 *1 75.905,20.37
X$9133 367 VIA_via1_4
* cell instance $9134 r0 *1 68.495,39.97
X$9134 367 VIA_via1_4
* cell instance $9135 r0 *1 70.205,21.63
X$9135 367 VIA_via1_4
* cell instance $9136 r0 *1 65.075,23.17
X$9136 367 VIA_via1_4
* cell instance $9137 r0 *1 65.075,23.31
X$9137 367 VIA_via2_5
* cell instance $9138 r0 *1 59.945,24.43
X$9138 367 VIA_via1_4
* cell instance $9139 r0 *1 58.235,20.37
X$9139 367 VIA_via1_4
* cell instance $9140 r0 *1 58.235,20.37
X$9140 367 VIA_via2_5
* cell instance $9141 r0 *1 52.155,16.03
X$9141 367 VIA_via1_4
* cell instance $9142 r0 *1 52.175,16.87
X$9142 367 VIA_via4_0
* cell instance $9143 r0 *1 46.015,16.87
X$9143 367 VIA_via3_2
* cell instance $9144 r0 *1 46.015,16.87
X$9144 367 VIA_via4_0
* cell instance $9145 r0 *1 52.175,18.41
X$9145 367 VIA_via3_2
* cell instance $9146 r0 *1 52.175,16.31
X$9146 367 VIA_via3_2
* cell instance $9147 r0 *1 52.155,16.31
X$9147 367 VIA_via2_5
* cell instance $9148 r0 *1 43.985,16.45
X$9148 368 VIA_via1_4
* cell instance $9149 r0 *1 43.795,17.57
X$9149 368 VIA_via1_4
* cell instance $9150 r0 *1 44.365,16.03
X$9150 368 VIA_via1_4
* cell instance $9151 r0 *1 45.315,16.59
X$9151 369 VIA_via1_7
* cell instance $9152 r0 *1 44.935,17.57
X$9152 369 VIA_via1_4
* cell instance $9153 r0 *1 77.045,18.27
X$9153 370 VIA_via2_5
* cell instance $9154 r0 *1 51.965,17.15
X$9154 370 VIA_via2_5
* cell instance $9155 r0 *1 57.095,17.01
X$9155 370 VIA_via2_5
* cell instance $9156 r0 *1 51.965,18.55
X$9156 370 VIA_via2_5
* cell instance $9157 r0 *1 57.095,17.99
X$9157 370 VIA_via2_5
* cell instance $9158 r0 *1 70.775,18.41
X$9158 370 VIA_via2_5
* cell instance $9159 r0 *1 64.885,18.41
X$9159 370 VIA_via2_5
* cell instance $9160 r0 *1 46.265,20.51
X$9160 370 VIA_via2_5
* cell instance $9161 r0 *1 75.525,25.27
X$9161 370 VIA_via2_5
* cell instance $9162 r0 *1 77.425,25.27
X$9162 370 VIA_via2_5
* cell instance $9163 r0 *1 64.885,17.99
X$9163 370 VIA_via2_5
* cell instance $9164 r0 *1 80.085,25.27
X$9164 370 VIA_via2_5
* cell instance $9165 r0 *1 62.035,21.77
X$9165 370 VIA_via2_5
* cell instance $9166 r0 *1 46.645,17.15
X$9166 370 VIA_via1_4
* cell instance $9167 r0 *1 46.645,17.15
X$9167 370 VIA_via2_5
* cell instance $9168 r0 *1 46.265,17.85
X$9168 370 VIA_via1_4
* cell instance $9169 r0 *1 41.705,20.37
X$9169 370 VIA_via1_4
* cell instance $9170 r0 *1 41.705,20.51
X$9170 370 VIA_via2_5
* cell instance $9171 r0 *1 80.085,24.43
X$9171 370 VIA_via1_4
* cell instance $9172 r0 *1 45.695,20.37
X$9172 370 VIA_via1_4
* cell instance $9173 r0 *1 45.695,20.51
X$9173 370 VIA_via2_5
* cell instance $9174 r0 *1 75.335,30.03
X$9174 370 VIA_via1_4
* cell instance $9175 r0 *1 77.045,18.83
X$9175 370 VIA_via1_4
* cell instance $9176 r0 *1 70.775,18.83
X$9176 370 VIA_via1_4
* cell instance $9177 r0 *1 57.095,21.63
X$9177 370 VIA_via1_4
* cell instance $9178 r0 *1 57.095,21.77
X$9178 370 VIA_via2_5
* cell instance $9179 r0 *1 62.035,24.43
X$9179 370 VIA_via1_4
* cell instance $9180 r0 *1 64.885,18.83
X$9180 370 VIA_via1_4
* cell instance $9181 r0 *1 52.345,18.83
X$9181 370 VIA_via1_4
* cell instance $9182 r0 *1 52.345,18.69
X$9182 370 VIA_via2_5
* cell instance $9183 r0 *1 52.155,16.59
X$9183 371 VIA_via1_7
* cell instance $9184 r0 *1 52.535,17.57
X$9184 371 VIA_via1_4
* cell instance $9185 r0 *1 56.715,41.23
X$9185 372 VIA_via1_7
* cell instance $9186 r0 *1 60.325,18.27
X$9186 372 VIA_via2_5
* cell instance $9187 r0 *1 60.895,23.45
X$9187 372 VIA_via2_5
* cell instance $9188 r0 *1 60.855,23.45
X$9188 372 VIA_via3_2
* cell instance $9189 r0 *1 60.325,17.43
X$9189 372 VIA_via2_5
* cell instance $9190 r0 *1 78.185,17.99
X$9190 372 VIA_via2_5
* cell instance $9191 r0 *1 80.085,18.97
X$9191 372 VIA_via2_5
* cell instance $9192 r0 *1 71.155,41.51
X$9192 372 VIA_via2_5
* cell instance $9193 r0 *1 66.025,18.27
X$9193 372 VIA_via2_5
* cell instance $9194 r0 *1 56.715,41.51
X$9194 372 VIA_via2_5
* cell instance $9195 r0 *1 78.185,45.15
X$9195 372 VIA_via2_5
* cell instance $9196 r0 *1 79.515,45.15
X$9196 372 VIA_via2_5
* cell instance $9197 r0 *1 71.155,45.15
X$9197 372 VIA_via2_5
* cell instance $9198 r0 *1 80.085,21.63
X$9198 372 VIA_via1_4
* cell instance $9199 r0 *1 79.515,45.57
X$9199 372 VIA_via1_4
* cell instance $9200 r0 *1 71.155,45.57
X$9200 372 VIA_via1_4
* cell instance $9201 r0 *1 78.185,18.83
X$9201 372 VIA_via1_4
* cell instance $9202 r0 *1 78.185,18.83
X$9202 372 VIA_via2_5
* cell instance $9203 r0 *1 58.805,17.57
X$9203 372 VIA_via1_4
* cell instance $9204 r0 *1 58.805,17.43
X$9204 372 VIA_via2_5
* cell instance $9205 r0 *1 70.965,17.57
X$9205 372 VIA_via1_4
* cell instance $9206 r0 *1 70.965,17.71
X$9206 372 VIA_via2_5
* cell instance $9207 r0 *1 60.895,23.17
X$9207 372 VIA_via1_4
* cell instance $9208 r0 *1 55.005,17.57
X$9208 372 VIA_via1_4
* cell instance $9209 r0 *1 55.005,17.43
X$9209 372 VIA_via2_5
* cell instance $9210 r0 *1 66.025,18.83
X$9210 372 VIA_via1_4
* cell instance $9211 r0 *1 78.375,58.03
X$9211 372 VIA_via1_4
* cell instance $9212 r0 *1 60.855,41.51
X$9212 372 VIA_via3_2
* cell instance $9213 r0 *1 67.355,16.17
X$9213 373 VIA_via1_7
* cell instance $9214 r0 *1 66.975,30.17
X$9214 373 VIA_via1_7
* cell instance $9215 r0 *1 66.975,30.17
X$9215 373 VIA_via2_5
* cell instance $9216 r0 *1 75.525,63.77
X$9216 373 VIA_via1_7
* cell instance $9217 r0 *1 75.525,63.77
X$9217 373 VIA_via2_5
* cell instance $9218 r0 *1 62.415,17.43
X$9218 373 VIA_via1_7
* cell instance $9219 r0 *1 61.275,73.43
X$9219 373 VIA_via1_7
* cell instance $9220 r0 *1 61.275,73.43
X$9220 373 VIA_via2_5
* cell instance $9221 r0 *1 75.905,23.73
X$9221 373 VIA_via2_5
* cell instance $9222 r0 *1 75.715,72.17
X$9222 373 VIA_via2_5
* cell instance $9223 r0 *1 75.695,72.17
X$9223 373 VIA_via3_2
* cell instance $9224 r0 *1 75.715,72.17
X$9224 373 VIA_via1_7
* cell instance $9225 r0 *1 69.065,30.45
X$9225 373 VIA_via2_5
* cell instance $9226 r0 *1 68.685,40.95
X$9226 373 VIA_via2_5
* cell instance $9227 r0 *1 62.035,48.79
X$9227 373 VIA_via2_5
* cell instance $9228 r0 *1 62.415,17.01
X$9228 373 VIA_via2_5
* cell instance $9229 r0 *1 69.065,40.95
X$9229 373 VIA_via2_5
* cell instance $9230 r0 *1 64.885,48.79
X$9230 373 VIA_via2_5
* cell instance $9231 r0 *1 68.685,42.91
X$9231 373 VIA_via2_5
* cell instance $9232 r0 *1 67.545,42.91
X$9232 373 VIA_via2_5
* cell instance $9233 r0 *1 64.885,43.47
X$9233 373 VIA_via2_5
* cell instance $9234 r0 *1 67.545,43.47
X$9234 373 VIA_via2_5
* cell instance $9235 r0 *1 76.285,42.77
X$9235 373 VIA_via1_4
* cell instance $9236 r0 *1 76.285,42.91
X$9236 373 VIA_via2_5
* cell instance $9237 r0 *1 67.545,44.03
X$9237 373 VIA_via1_4
* cell instance $9238 r0 *1 75.905,23.17
X$9238 373 VIA_via1_4
* cell instance $9239 r0 *1 75.905,23.31
X$9239 373 VIA_via2_5
* cell instance $9240 r0 *1 75.905,17.57
X$9240 373 VIA_via1_4
* cell instance $9241 r0 *1 75.905,17.57
X$9241 373 VIA_via2_5
* cell instance $9242 r0 *1 62.035,50.75
X$9242 373 VIA_via1_4
* cell instance $9243 r0 *1 61.655,51.45
X$9243 373 VIA_via1_4
* cell instance $9244 r0 *1 61.975,71.47
X$9244 373 VIA_via3_2
* cell instance $9245 r0 *1 61.975,73.43
X$9245 373 VIA_via3_2
* cell instance $9246 r0 *1 61.695,51.73
X$9246 373 VIA_via3_2
* cell instance $9247 r0 *1 61.655,51.73
X$9247 373 VIA_via2_5
* cell instance $9248 r0 *1 67.295,17.01
X$9248 373 VIA_via3_2
* cell instance $9249 r0 *1 67.165,17.01
X$9249 373 VIA_via2_5
* cell instance $9250 r0 *1 75.695,71.61
X$9250 373 VIA_via3_2
* cell instance $9251 r0 *1 67.295,23.73
X$9251 373 VIA_via3_2
* cell instance $9252 r0 *1 75.695,17.57
X$9252 373 VIA_via3_2
* cell instance $9253 r0 *1 67.295,30.45
X$9253 373 VIA_via3_2
* cell instance $9254 r0 *1 75.695,23.31
X$9254 373 VIA_via3_2
* cell instance $9255 r0 *1 67.295,30.17
X$9255 373 VIA_via3_2
* cell instance $9256 r0 *1 75.695,63.77
X$9256 373 VIA_via3_2
* cell instance $9257 r0 *1 80.655,17.43
X$9257 374 VIA_via2_5
* cell instance $9258 r0 *1 79.135,59.15
X$9258 374 VIA_via2_5
* cell instance $9259 r0 *1 63.555,20.09
X$9259 374 VIA_via2_5
* cell instance $9260 r0 *1 65.265,20.09
X$9260 374 VIA_via2_5
* cell instance $9261 r0 *1 65.265,17.57
X$9261 374 VIA_via2_5
* cell instance $9262 r0 *1 78.755,42.63
X$9262 374 VIA_via2_5
* cell instance $9263 r0 *1 79.895,42.63
X$9263 374 VIA_via2_5
* cell instance $9264 r0 *1 80.465,23.17
X$9264 374 VIA_via1_4
* cell instance $9265 r0 *1 80.085,32.83
X$9265 374 VIA_via1_4
* cell instance $9266 r0 *1 79.895,44.03
X$9266 374 VIA_via1_4
* cell instance $9267 r0 *1 71.915,42.77
X$9267 374 VIA_via1_4
* cell instance $9268 r0 *1 71.915,42.63
X$9268 374 VIA_via2_5
* cell instance $9269 r0 *1 79.895,17.57
X$9269 374 VIA_via1_4
* cell instance $9270 r0 *1 79.895,17.43
X$9270 374 VIA_via2_5
* cell instance $9271 r0 *1 66.215,17.57
X$9271 374 VIA_via1_4
* cell instance $9272 r0 *1 66.215,17.57
X$9272 374 VIA_via2_5
* cell instance $9273 r0 *1 59.185,20.37
X$9273 374 VIA_via1_4
* cell instance $9274 r0 *1 59.185,20.51
X$9274 374 VIA_via2_5
* cell instance $9275 r0 *1 70.205,17.57
X$9275 374 VIA_via1_4
* cell instance $9276 r0 *1 70.205,17.57
X$9276 374 VIA_via2_5
* cell instance $9277 r0 *1 63.555,20.37
X$9277 374 VIA_via1_4
* cell instance $9278 r0 *1 63.555,20.51
X$9278 374 VIA_via2_5
* cell instance $9279 r0 *1 59.375,59.15
X$9279 374 VIA_via1_4
* cell instance $9280 r0 *1 59.375,59.15
X$9280 374 VIA_via2_5
* cell instance $9281 r0 *1 79.135,60.83
X$9281 374 VIA_via1_4
* cell instance $9282 r0 *1 76.095,18.83
X$9282 375 VIA_via1_4
* cell instance $9283 r0 *1 76.095,17.57
X$9283 375 VIA_via1_4
* cell instance $9284 r0 *1 76.285,16.45
X$9284 375 VIA_via1_4
* cell instance $9285 r0 *1 79.325,17.71
X$9285 376 VIA_via2_5
* cell instance $9286 r0 *1 80.275,17.57
X$9286 376 VIA_via1_4
* cell instance $9287 r0 *1 80.275,17.71
X$9287 376 VIA_via2_5
* cell instance $9288 r0 *1 79.515,16.45
X$9288 376 VIA_via1_4
* cell instance $9289 r0 *1 78.185,17.57
X$9289 376 VIA_via1_4
* cell instance $9290 r0 *1 78.185,17.71
X$9290 376 VIA_via2_5
* cell instance $9291 r0 *1 96.425,12.39
X$9291 377 VIA_via1_7
* cell instance $9292 r0 *1 85.215,17.43
X$9292 377 VIA_via2_5
* cell instance $9293 r0 *1 82.555,17.43
X$9293 377 VIA_via2_5
* cell instance $9294 r0 *1 92.055,16.87
X$9294 377 VIA_via2_5
* cell instance $9295 r0 *1 93.955,16.87
X$9295 377 VIA_via2_5
* cell instance $9296 r0 *1 95.095,16.87
X$9296 377 VIA_via2_5
* cell instance $9297 r0 *1 92.055,17.43
X$9297 377 VIA_via2_5
* cell instance $9298 r0 *1 96.425,16.87
X$9298 377 VIA_via2_5
* cell instance $9299 r0 *1 85.025,21.63
X$9299 377 VIA_via1_4
* cell instance $9300 r0 *1 92.055,14.77
X$9300 377 VIA_via1_4
* cell instance $9301 r0 *1 95.095,16.03
X$9301 377 VIA_via1_4
* cell instance $9302 r0 *1 82.365,20.37
X$9302 377 VIA_via1_4
* cell instance $9303 r0 *1 82.555,16.03
X$9303 377 VIA_via1_4
* cell instance $9304 r0 *1 95.095,23.17
X$9304 377 VIA_via1_4
* cell instance $9305 r0 *1 93.765,18.83
X$9305 377 VIA_via1_4
* cell instance $9306 r0 *1 80.465,17.01
X$9306 378 VIA_via2_5
* cell instance $9307 r0 *1 83.125,17.01
X$9307 378 VIA_via2_5
* cell instance $9308 r0 *1 80.465,20.37
X$9308 378 VIA_via1_4
* cell instance $9309 r0 *1 83.125,16.03
X$9309 378 VIA_via1_4
* cell instance $9310 r0 *1 85.215,17.15
X$9310 378 VIA_via1_4
* cell instance $9311 r0 *1 85.215,17.01
X$9311 378 VIA_via2_5
* cell instance $9312 r0 *1 89.585,16.59
X$9312 379 VIA_via1_7
* cell instance $9313 r0 *1 89.585,16.87
X$9313 379 VIA_via2_5
* cell instance $9314 r0 *1 87.875,16.87
X$9314 379 VIA_via2_5
* cell instance $9315 r0 *1 87.875,17.57
X$9315 379 VIA_via1_4
* cell instance $9316 r0 *1 20.995,17.29
X$9316 380 VIA_via2_5
* cell instance $9317 r0 *1 20.995,17.57
X$9317 380 VIA_via1_4
* cell instance $9318 r0 *1 16.245,17.15
X$9318 380 VIA_via1_4
* cell instance $9319 r0 *1 16.245,17.29
X$9319 380 VIA_via2_5
* cell instance $9320 r0 *1 13.395,66.29
X$9320 381 VIA_via2_5
* cell instance $9321 r0 *1 12.825,63.35
X$9321 381 VIA_via2_5
* cell instance $9322 r0 *1 13.395,63.35
X$9322 381 VIA_via2_5
* cell instance $9323 r0 *1 30.685,18.41
X$9323 381 VIA_via2_5
* cell instance $9324 r0 *1 25.365,18.41
X$9324 381 VIA_via2_5
* cell instance $9325 r0 *1 35.815,18.41
X$9325 381 VIA_via2_5
* cell instance $9326 r0 *1 17.575,20.65
X$9326 381 VIA_via2_5
* cell instance $9327 r0 *1 17.455,20.65
X$9327 381 VIA_via3_2
* cell instance $9328 r0 *1 20.425,18.69
X$9328 381 VIA_via2_5
* cell instance $9329 r0 *1 20.425,17.85
X$9329 381 VIA_via2_5
* cell instance $9330 r0 *1 13.015,54.11
X$9330 381 VIA_via2_5
* cell instance $9331 r0 *1 14.155,24.71
X$9331 381 VIA_via2_5
* cell instance $9332 r0 *1 12.825,24.71
X$9332 381 VIA_via2_5
* cell instance $9333 r0 *1 25.365,18.83
X$9333 381 VIA_via1_4
* cell instance $9334 r0 *1 25.365,18.69
X$9334 381 VIA_via2_5
* cell instance $9335 r0 *1 31.255,20.37
X$9335 381 VIA_via1_4
* cell instance $9336 r0 *1 35.815,18.83
X$9336 381 VIA_via1_4
* cell instance $9337 r0 *1 35.245,54.11
X$9337 381 VIA_via1_4
* cell instance $9338 r0 *1 35.245,54.11
X$9338 381 VIA_via2_5
* cell instance $9339 r0 *1 14.155,24.5
X$9339 381 VIA_via1_4
* cell instance $9340 r0 *1 13.965,66.43
X$9340 381 VIA_via1_4
* cell instance $9341 r0 *1 13.965,66.29
X$9341 381 VIA_via2_5
* cell instance $9342 r0 *1 14.155,53.97
X$9342 381 VIA_via1_4
* cell instance $9343 r0 *1 14.155,54.11
X$9343 381 VIA_via2_5
* cell instance $9344 r0 *1 20.425,17.57
X$9344 381 VIA_via1_4
* cell instance $9345 r0 *1 17.575,20.37
X$9345 381 VIA_via1_4
* cell instance $9346 r0 *1 16.625,16.03
X$9346 381 VIA_via1_4
* cell instance $9347 r0 *1 16.625,16.17
X$9347 381 VIA_via2_5
* cell instance $9348 r0 *1 13.395,73.57
X$9348 381 VIA_via1_4
* cell instance $9349 r0 *1 14.375,54.11
X$9349 381 VIA_via4_0
* cell instance $9350 r0 *1 14.375,54.11
X$9350 381 VIA_via3_2
* cell instance $9351 r0 *1 34.535,54.11
X$9351 381 VIA_via3_2
* cell instance $9352 r0 *1 34.535,54.11
X$9352 381 VIA_via4_0
* cell instance $9353 r0 *1 17.455,16.17
X$9353 381 VIA_via3_2
* cell instance $9354 r0 *1 17.455,17.85
X$9354 381 VIA_via3_2
* cell instance $9355 r0 *1 17.455,24.71
X$9355 381 VIA_via3_2
* cell instance $9356 r0 *1 78.565,17.01
X$9356 382 VIA_via1_7
* cell instance $9357 r0 *1 78.565,17.01
X$9357 382 VIA_via2_5
* cell instance $9358 r0 *1 77.235,17.01
X$9358 382 VIA_via2_5
* cell instance $9359 r0 *1 77.235,16.03
X$9359 382 VIA_via1_4
* cell instance $9360 r0 *1 77.045,17.01
X$9360 383 VIA_via1_7
* cell instance $9361 r0 *1 77.045,16.87
X$9361 383 VIA_via2_5
* cell instance $9362 r0 *1 74.005,16.87
X$9362 383 VIA_via2_5
* cell instance $9363 r0 *1 74.005,16.03
X$9363 383 VIA_via1_4
* cell instance $9364 r0 *1 69.635,17.15
X$9364 384 VIA_via2_5
* cell instance $9365 r0 *1 67.545,17.15
X$9365 384 VIA_via2_5
* cell instance $9366 r0 *1 69.825,18.83
X$9366 384 VIA_via1_4
* cell instance $9367 r0 *1 69.635,17.85
X$9367 384 VIA_via1_4
* cell instance $9368 r0 *1 67.545,16.03
X$9368 384 VIA_via1_4
* cell instance $9369 r0 *1 68.495,16.59
X$9369 385 VIA_via1_7
* cell instance $9370 r0 *1 68.495,16.59
X$9370 385 VIA_via2_5
* cell instance $9371 r0 *1 67.355,16.59
X$9371 385 VIA_via2_5
* cell instance $9372 r0 *1 67.355,17.57
X$9372 385 VIA_via1_4
* cell instance $9373 r0 *1 62.605,16.45
X$9373 386 VIA_via2_5
* cell instance $9374 r0 *1 65.265,16.45
X$9374 386 VIA_via1_4
* cell instance $9375 r0 *1 65.265,16.45
X$9375 386 VIA_via2_5
* cell instance $9376 r0 *1 62.605,17.57
X$9376 386 VIA_via1_4
* cell instance $9377 r0 *1 62.605,18.83
X$9377 386 VIA_via1_4
* cell instance $9378 r0 *1 31.255,17.01
X$9378 387 VIA_via1_7
* cell instance $9379 r0 *1 31.255,17.01
X$9379 387 VIA_via2_5
* cell instance $9380 r0 *1 32.395,17.01
X$9380 387 VIA_via2_5
* cell instance $9381 r0 *1 32.395,16.03
X$9381 387 VIA_via1_4
* cell instance $9382 r0 *1 35.245,16.59
X$9382 388 VIA_via1_7
* cell instance $9383 r0 *1 35.245,16.59
X$9383 388 VIA_via2_5
* cell instance $9384 r0 *1 35.245,19.11
X$9384 388 VIA_via2_5
* cell instance $9385 r0 *1 35.245,18.83
X$9385 388 VIA_via1_4
* cell instance $9386 r0 *1 35.095,16.59
X$9386 388 VIA_via3_2
* cell instance $9387 r0 *1 35.095,19.11
X$9387 388 VIA_via3_2
* cell instance $9388 r0 *1 38.665,17.01
X$9388 389 VIA_via1_7
* cell instance $9389 r0 *1 38.665,17.01
X$9389 389 VIA_via2_5
* cell instance $9390 r0 *1 36.385,17.01
X$9390 389 VIA_via2_5
* cell instance $9391 r0 *1 36.385,16.03
X$9391 389 VIA_via1_4
* cell instance $9392 r0 *1 51.965,13.79
X$9392 390 VIA_via1_7
* cell instance $9393 r0 *1 51.965,16.87
X$9393 390 VIA_via2_5
* cell instance $9394 r0 *1 53.295,16.87
X$9394 390 VIA_via2_5
* cell instance $9395 r0 *1 53.295,17.57
X$9395 390 VIA_via1_4
* cell instance $9396 r0 *1 10.355,17.85
X$9396 391 VIA_via2_5
* cell instance $9397 r0 *1 8.835,17.85
X$9397 391 VIA_via2_5
* cell instance $9398 r0 *1 8.835,18.83
X$9398 391 VIA_via1_4
* cell instance $9399 r0 *1 10.355,17.57
X$9399 391 VIA_via1_4
* cell instance $9400 r0 *1 9.405,17.85
X$9400 391 VIA_via1_4
* cell instance $9401 r0 *1 9.405,17.85
X$9401 391 VIA_via2_5
* cell instance $9402 r0 *1 15.105,17.57
X$9402 392 VIA_via2_5
* cell instance $9403 r0 *1 15.105,18.83
X$9403 392 VIA_via1_4
* cell instance $9404 r0 *1 14.345,17.57
X$9404 392 VIA_via1_4
* cell instance $9405 r0 *1 14.345,17.57
X$9405 392 VIA_via2_5
* cell instance $9406 r0 *1 13.965,17.57
X$9406 392 VIA_via1_4
* cell instance $9407 r0 *1 13.965,17.57
X$9407 392 VIA_via2_5
* cell instance $9408 r0 *1 19.665,21.77
X$9408 393 VIA_via1_7
* cell instance $9409 r0 *1 32.775,21.77
X$9409 393 VIA_via1_7
* cell instance $9410 r0 *1 37.525,23.03
X$9410 393 VIA_via1_7
* cell instance $9411 r0 *1 46.835,21.07
X$9411 393 VIA_via2_5
* cell instance $9412 r0 *1 32.775,22.05
X$9412 393 VIA_via2_5
* cell instance $9413 r0 *1 25.555,22.19
X$9413 393 VIA_via2_5
* cell instance $9414 r0 *1 42.655,21.07
X$9414 393 VIA_via2_5
* cell instance $9415 r0 *1 37.525,21.07
X$9415 393 VIA_via2_5
* cell instance $9416 r0 *1 37.525,22.05
X$9416 393 VIA_via2_5
* cell instance $9417 r0 *1 15.865,24.01
X$9417 393 VIA_via2_5
* cell instance $9418 r0 *1 15.865,22.19
X$9418 393 VIA_via2_5
* cell instance $9419 r0 *1 15.485,18.69
X$9419 393 VIA_via2_5
* cell instance $9420 r0 *1 12.635,24.01
X$9420 393 VIA_via2_5
* cell instance $9421 r0 *1 14.155,18.41
X$9421 393 VIA_via2_5
* cell instance $9422 r0 *1 19.665,22.19
X$9422 393 VIA_via2_5
* cell instance $9423 r0 *1 12.445,24.43
X$9423 393 VIA_via1_4
* cell instance $9424 r0 *1 42.655,20.37
X$9424 393 VIA_via1_4
* cell instance $9425 r0 *1 46.835,24.15
X$9425 393 VIA_via1_4
* cell instance $9426 r0 *1 46.835,18.83
X$9426 393 VIA_via1_4
* cell instance $9427 r0 *1 25.555,23.17
X$9427 393 VIA_via1_4
* cell instance $9428 r0 *1 15.865,23.17
X$9428 393 VIA_via1_4
* cell instance $9429 r0 *1 16.245,18.83
X$9429 393 VIA_via1_4
* cell instance $9430 r0 *1 16.245,18.69
X$9430 393 VIA_via2_5
* cell instance $9431 r0 *1 14.155,17.57
X$9431 393 VIA_via1_4
* cell instance $9432 r0 *1 17.385,18.41
X$9432 394 VIA_via1_7
* cell instance $9433 r0 *1 17.195,17.57
X$9433 394 VIA_via1_4
* cell instance $9434 r0 *1 19.665,18.41
X$9434 395 VIA_via1_7
* cell instance $9435 r0 *1 20.045,17.57
X$9435 395 VIA_via1_4
* cell instance $9436 r0 *1 22.135,15.19
X$9436 396 VIA_via1_7
* cell instance $9437 r0 *1 21.755,17.57
X$9437 396 VIA_via1_4
* cell instance $9438 r0 *1 25.555,34.65
X$9438 397 VIA_via2_5
* cell instance $9439 r0 *1 26.885,34.51
X$9439 397 VIA_via2_5
* cell instance $9440 r0 *1 25.555,17.57
X$9440 397 VIA_via1_4
* cell instance $9441 r0 *1 25.745,49.63
X$9441 397 VIA_via1_4
* cell instance $9442 r0 *1 26.315,46.83
X$9442 397 VIA_via1_4
* cell instance $9443 r0 *1 43.415,24.01
X$9443 398 VIA_via1_7
* cell instance $9444 r0 *1 43.415,24.99
X$9444 398 VIA_via1_7
* cell instance $9445 r0 *1 44.365,40.11
X$9445 398 VIA_via2_5
* cell instance $9446 r0 *1 43.415,20.09
X$9446 398 VIA_via2_5
* cell instance $9447 r0 *1 42.845,40.11
X$9447 398 VIA_via2_5
* cell instance $9448 r0 *1 45.695,17.57
X$9448 398 VIA_via2_5
* cell instance $9449 r0 *1 42.655,35.49
X$9449 398 VIA_via2_5
* cell instance $9450 r0 *1 42.655,28.77
X$9450 398 VIA_via2_5
* cell instance $9451 r0 *1 44.175,20.09
X$9451 398 VIA_via2_5
* cell instance $9452 r0 *1 45.885,20.65
X$9452 398 VIA_via2_5
* cell instance $9453 r0 *1 43.415,20.65
X$9453 398 VIA_via2_5
* cell instance $9454 r0 *1 45.695,14.77
X$9454 398 VIA_via1_4
* cell instance $9455 r0 *1 44.365,17.57
X$9455 398 VIA_via1_4
* cell instance $9456 r0 *1 44.365,17.57
X$9456 398 VIA_via2_5
* cell instance $9457 r0 *1 43.415,20.37
X$9457 398 VIA_via1_4
* cell instance $9458 r0 *1 45.885,21.63
X$9458 398 VIA_via1_4
* cell instance $9459 r0 *1 42.845,41.23
X$9459 398 VIA_via1_4
* cell instance $9460 r0 *1 42.845,41.37
X$9460 398 VIA_via2_5
* cell instance $9461 r0 *1 40.375,41.23
X$9461 398 VIA_via1_4
* cell instance $9462 r0 *1 40.375,41.37
X$9462 398 VIA_via2_5
* cell instance $9463 r0 *1 44.365,38.43
X$9463 398 VIA_via1_4
* cell instance $9464 r0 *1 40.945,35.63
X$9464 398 VIA_via1_4
* cell instance $9465 r0 *1 40.945,35.49
X$9465 398 VIA_via2_5
* cell instance $9466 r0 *1 43.605,28.77
X$9466 398 VIA_via1_4
* cell instance $9467 r0 *1 43.605,28.77
X$9467 398 VIA_via2_5
* cell instance $9468 r0 *1 42.655,32.83
X$9468 398 VIA_via1_4
* cell instance $9469 r0 *1 45.125,17.99
X$9469 399 VIA_via1_7
* cell instance $9470 r0 *1 44.745,18.83
X$9470 399 VIA_via1_4
* cell instance $9471 r0 *1 46.075,16.31
X$9471 400 VIA_via1_4
* cell instance $9472 r0 *1 45.505,18.83
X$9472 400 VIA_via1_4
* cell instance $9473 r0 *1 47.975,18.41
X$9473 401 VIA_via1_7
* cell instance $9474 r0 *1 47.595,17.57
X$9474 401 VIA_via1_4
* cell instance $9475 r0 *1 47.025,18.83
X$9475 402 VIA_via1_4
* cell instance $9476 r0 *1 47.025,18.69
X$9476 402 VIA_via2_5
* cell instance $9477 r0 *1 49.875,17.85
X$9477 402 VIA_via1_4
* cell instance $9478 r0 *1 49.685,18.83
X$9478 402 VIA_via1_4
* cell instance $9479 r0 *1 49.685,18.69
X$9479 402 VIA_via2_5
* cell instance $9480 r0 *1 52.535,17.85
X$9480 403 VIA_via2_5
* cell instance $9481 r0 *1 51.205,17.85
X$9481 403 VIA_via2_5
* cell instance $9482 r0 *1 58.425,57.61
X$9482 403 VIA_via2_5
* cell instance $9483 r0 *1 43.415,57.19
X$9483 403 VIA_via2_5
* cell instance $9484 r0 *1 35.815,53.97
X$9484 403 VIA_via2_5
* cell instance $9485 r0 *1 35.815,57.19
X$9485 403 VIA_via2_5
* cell instance $9486 r0 *1 45.885,17.57
X$9486 403 VIA_via1_4
* cell instance $9487 r0 *1 45.885,17.43
X$9487 403 VIA_via2_5
* cell instance $9488 r0 *1 43.415,58.03
X$9488 403 VIA_via1_4
* cell instance $9489 r0 *1 35.815,59.57
X$9489 403 VIA_via1_4
* cell instance $9490 r0 *1 35.815,59.57
X$9490 403 VIA_via2_5
* cell instance $9491 r0 *1 34.105,59.57
X$9491 403 VIA_via1_4
* cell instance $9492 r0 *1 34.105,59.57
X$9492 403 VIA_via2_5
* cell instance $9493 r0 *1 34.675,53.97
X$9493 403 VIA_via1_4
* cell instance $9494 r0 *1 34.675,53.97
X$9494 403 VIA_via2_5
* cell instance $9495 r0 *1 52.535,20.37
X$9495 403 VIA_via1_4
* cell instance $9496 r0 *1 52.535,20.37
X$9496 403 VIA_via2_5
* cell instance $9497 r0 *1 51.205,17.57
X$9497 403 VIA_via1_4
* cell instance $9498 r0 *1 51.205,17.43
X$9498 403 VIA_via2_5
* cell instance $9499 r0 *1 35.815,56.77
X$9499 403 VIA_via1_4
* cell instance $9500 r0 *1 33.155,59.57
X$9500 403 VIA_via1_4
* cell instance $9501 r0 *1 33.155,59.57
X$9501 403 VIA_via2_5
* cell instance $9502 r0 *1 58.805,57.75
X$9502 403 VIA_via1_4
* cell instance $9503 r0 *1 58.805,57.61
X$9503 403 VIA_via2_5
* cell instance $9504 r0 *1 58.425,59.57
X$9504 403 VIA_via1_4
* cell instance $9505 r0 *1 52.735,20.37
X$9505 403 VIA_via3_2
* cell instance $9506 r0 *1 52.735,57.19
X$9506 403 VIA_via3_2
* cell instance $9507 r0 *1 52.155,18.41
X$9507 404 VIA_via1_7
* cell instance $9508 r0 *1 52.345,17.57
X$9508 404 VIA_via1_4
* cell instance $9509 r0 *1 54.245,10.99
X$9509 405 VIA_via1_7
* cell instance $9510 r0 *1 54.625,17.57
X$9510 405 VIA_via1_4
* cell instance $9511 r0 *1 66.025,17.99
X$9511 406 VIA_via1_7
* cell instance $9512 r0 *1 66.025,20.37
X$9512 406 VIA_via1_4
* cell instance $9513 r0 *1 70.775,17.99
X$9513 407 VIA_via1_7
* cell instance $9514 r0 *1 70.775,20.37
X$9514 407 VIA_via1_4
* cell instance $9515 r0 *1 73.055,18.97
X$9515 408 VIA_via2_5
* cell instance $9516 r0 *1 73.815,18.97
X$9516 408 VIA_via1_4
* cell instance $9517 r0 *1 73.815,18.97
X$9517 408 VIA_via2_5
* cell instance $9518 r0 *1 72.865,17.57
X$9518 408 VIA_via1_4
* cell instance $9519 r0 *1 83.505,16.59
X$9519 409 VIA_via1_7
* cell instance $9520 r0 *1 82.935,17.57
X$9520 409 VIA_via1_4
* cell instance $9521 r0 *1 94.145,17.99
X$9521 410 VIA_via1_7
* cell instance $9522 r0 *1 92.245,21.07
X$9522 410 VIA_via2_5
* cell instance $9523 r0 *1 93.955,21.07
X$9523 410 VIA_via2_5
* cell instance $9524 r0 *1 92.245,21.63
X$9524 410 VIA_via1_4
* cell instance $9525 r0 *1 8.455,17.57
X$9525 411 VIA_via2_5
* cell instance $9526 r0 *1 8.455,18.55
X$9526 411 VIA_via1_4
* cell instance $9527 r0 *1 8.835,20.37
X$9527 411 VIA_via1_4
* cell instance $9528 r0 *1 9.785,17.57
X$9528 411 VIA_via1_4
* cell instance $9529 r0 *1 9.785,17.57
X$9529 411 VIA_via2_5
* cell instance $9530 r0 *1 4.465,88.97
X$9530 412 VIA_via1_7
* cell instance $9531 r0 *1 5.985,23.03
X$9531 412 VIA_via1_7
* cell instance $9532 r0 *1 5.985,23.03
X$9532 412 VIA_via2_5
* cell instance $9533 r0 *1 5.225,20.23
X$9533 412 VIA_via1_7
* cell instance $9534 r0 *1 5.225,20.23
X$9534 412 VIA_via2_5
* cell instance $9535 r0 *1 5.415,16.17
X$9535 412 VIA_via1_7
* cell instance $9536 r0 *1 6.745,53.83
X$9536 412 VIA_via1_7
* cell instance $9537 r0 *1 6.745,53.69
X$9537 412 VIA_via2_5
* cell instance $9538 r0 *1 9.595,17.43
X$9538 412 VIA_via1_7
* cell instance $9539 r0 *1 9.595,17.43
X$9539 412 VIA_via2_5
* cell instance $9540 r0 *1 9.615,17.43
X$9540 412 VIA_via3_2
* cell instance $9541 r0 *1 26.695,88.27
X$9541 412 VIA_via2_5
* cell instance $9542 r0 *1 9.215,56.35
X$9542 412 VIA_via2_5
* cell instance $9543 r0 *1 8.455,56.35
X$9543 412 VIA_via2_5
* cell instance $9544 r0 *1 4.275,83.93
X$9544 412 VIA_via2_5
* cell instance $9545 r0 *1 5.035,83.93
X$9545 412 VIA_via2_5
* cell instance $9546 r0 *1 4.465,89.67
X$9546 412 VIA_via2_5
* cell instance $9547 r0 *1 5.035,71.05
X$9547 412 VIA_via2_5
* cell instance $9548 r0 *1 5.795,71.05
X$9548 412 VIA_via2_5
* cell instance $9549 r0 *1 9.025,71.05
X$9549 412 VIA_via2_5
* cell instance $9550 r0 *1 15.485,88.27
X$9550 412 VIA_via2_5
* cell instance $9551 r0 *1 15.485,89.67
X$9551 412 VIA_via2_5
* cell instance $9552 r0 *1 8.455,52.85
X$9552 412 VIA_via2_5
* cell instance $9553 r0 *1 8.455,53.69
X$9553 412 VIA_via2_5
* cell instance $9554 r0 *1 5.795,20.23
X$9554 412 VIA_via2_5
* cell instance $9555 r0 *1 15.485,88.83
X$9555 412 VIA_via1_4
* cell instance $9556 r0 *1 26.695,87.57
X$9556 412 VIA_via1_4
* cell instance $9557 r0 *1 9.025,69.23
X$9557 412 VIA_via1_4
* cell instance $9558 r0 *1 5.795,70.77
X$9558 412 VIA_via1_4
* cell instance $9559 r0 *1 26.505,27.51
X$9559 412 VIA_via1_4
* cell instance $9560 r0 *1 26.505,27.51
X$9560 412 VIA_via2_5
* cell instance $9561 r0 *1 9.615,27.51
X$9561 412 VIA_via3_2
* cell instance $9562 r0 *1 9.615,52.85
X$9562 412 VIA_via3_2
* cell instance $9563 r0 *1 9.615,23.03
X$9563 412 VIA_via3_2
* cell instance $9564 r0 *1 11.685,17.57
X$9564 413 VIA_via1_4
* cell instance $9565 r0 *1 11.685,17.71
X$9565 413 VIA_via2_5
* cell instance $9566 r0 *1 15.295,17.71
X$9566 413 VIA_via1_4
* cell instance $9567 r0 *1 15.295,17.71
X$9567 413 VIA_via2_5
* cell instance $9568 r0 *1 82.365,42.63
X$9568 414 VIA_via1_7
* cell instance $9569 r0 *1 48.735,74.97
X$9569 414 VIA_via1_7
* cell instance $9570 r0 *1 48.735,74.97
X$9570 414 VIA_via2_5
* cell instance $9571 r0 *1 68.685,72.17
X$9571 414 VIA_via1_7
* cell instance $9572 r0 *1 81.985,21.77
X$9572 414 VIA_via1_7
* cell instance $9573 r0 *1 54.415,61.11
X$9573 414 VIA_via5_0
* cell instance $9574 r0 *1 54.415,62.23
X$9574 414 VIA_via5_0
* cell instance $9575 r0 *1 80.085,17.99
X$9575 414 VIA_via2_5
* cell instance $9576 r0 *1 81.985,17.99
X$9576 414 VIA_via2_5
* cell instance $9577 r0 *1 52.345,59.43
X$9577 414 VIA_via2_5
* cell instance $9578 r0 *1 53.485,59.43
X$9578 414 VIA_via2_5
* cell instance $9579 r0 *1 52.535,61.11
X$9579 414 VIA_via2_5
* cell instance $9580 r0 *1 57.475,75.11
X$9580 414 VIA_via2_5
* cell instance $9581 r0 *1 68.685,74.83
X$9581 414 VIA_via2_5
* cell instance $9582 r0 *1 79.135,62.51
X$9582 414 VIA_via2_5
* cell instance $9583 r0 *1 48.545,48.93
X$9583 414 VIA_via2_5
* cell instance $9584 r0 *1 70.965,41.37
X$9584 414 VIA_via2_5
* cell instance $9585 r0 *1 70.935,41.37
X$9585 414 VIA_via3_2
* cell instance $9586 r0 *1 70.965,41.37
X$9586 414 VIA_via1_7
* cell instance $9587 r0 *1 53.675,48.93
X$9587 414 VIA_via2_5
* cell instance $9588 r0 *1 81.985,41.37
X$9588 414 VIA_via2_5
* cell instance $9589 r0 *1 57.475,74.83
X$9589 414 VIA_via1_4
* cell instance $9590 r0 *1 57.475,74.83
X$9590 414 VIA_via2_5
* cell instance $9591 r0 *1 80.085,17.57
X$9591 414 VIA_via1_4
* cell instance $9592 r0 *1 48.545,49.35
X$9592 414 VIA_via1_4
* cell instance $9593 r0 *1 82.365,72.03
X$9593 414 VIA_via1_4
* cell instance $9594 r0 *1 82.365,72.03
X$9594 414 VIA_via2_5
* cell instance $9595 r0 *1 52.345,60.83
X$9595 414 VIA_via1_4
* cell instance $9596 r0 *1 54.415,75.11
X$9596 414 VIA_via4_0
* cell instance $9597 r0 *1 54.415,75.11
X$9597 414 VIA_via3_2
* cell instance $9598 r0 *1 54.415,75.11
X$9598 414 VIA_via5_0
* cell instance $9599 r0 *1 70.935,45.15
X$9599 414 VIA_via4_0
* cell instance $9600 r0 *1 56.655,45.15
X$9600 414 VIA_via4_0
* cell instance $9601 r0 *1 56.655,48.93
X$9601 414 VIA_via3_2
* cell instance $9602 r0 *1 82.135,72.03
X$9602 414 VIA_via3_2
* cell instance $9603 r0 *1 53.575,61.11
X$9603 414 VIA_via3_2
* cell instance $9604 r0 *1 53.575,61.11
X$9604 414 VIA_via4_0
* cell instance $9605 r0 *1 79.055,62.23
X$9605 414 VIA_via3_2
* cell instance $9606 r0 *1 79.055,62.23
X$9606 414 VIA_via4_0
* cell instance $9607 r0 *1 79.135,62.23
X$9607 414 VIA_via2_5
* cell instance $9608 r0 *1 79.135,62.23
X$9608 414 VIA_via1_7
* cell instance $9609 r0 *1 82.135,62.51
X$9609 414 VIA_via3_2
* cell instance $9610 r0 *1 81.225,17.57
X$9610 415 VIA_via1_4
* cell instance $9611 r0 *1 81.225,17.57
X$9611 415 VIA_via2_5
* cell instance $9612 r0 *1 79.515,17.57
X$9612 415 VIA_via1_4
* cell instance $9613 r0 *1 79.515,17.57
X$9613 415 VIA_via2_5
* cell instance $9614 r0 *1 10.735,17.43
X$9614 416 VIA_via1_4
* cell instance $9615 r0 *1 10.735,17.43
X$9615 416 VIA_via2_5
* cell instance $9616 r0 *1 15.865,17.57
X$9616 416 VIA_via1_4
* cell instance $9617 r0 *1 15.865,17.43
X$9617 416 VIA_via2_5
* cell instance $9618 r0 *1 21.565,17.57
X$9618 417 VIA_via1_4
* cell instance $9619 r0 *1 21.565,14.63
X$9619 417 VIA_via1_4
* cell instance $9620 r0 *1 25.365,17.85
X$9620 418 VIA_via2_5
* cell instance $9621 r0 *1 26.885,17.85
X$9621 418 VIA_via1_4
* cell instance $9622 r0 *1 26.885,17.85
X$9622 418 VIA_via2_5
* cell instance $9623 r0 *1 25.365,17.57
X$9623 418 VIA_via1_4
* cell instance $9624 r0 *1 70.015,17.99
X$9624 419 VIA_via1_7
* cell instance $9625 r0 *1 70.015,17.99
X$9625 419 VIA_via2_5
* cell instance $9626 r0 *1 71.155,17.99
X$9626 419 VIA_via2_5
* cell instance $9627 r0 *1 70.965,20.37
X$9627 419 VIA_via1_4
* cell instance $9628 r0 *1 69.825,16.59
X$9628 420 VIA_via1_7
* cell instance $9629 r0 *1 69.825,17.57
X$9629 420 VIA_via1_4
* cell instance $9630 r0 *1 29.355,25.41
X$9630 421 VIA_via1_7
* cell instance $9631 r0 *1 29.355,25.41
X$9631 421 VIA_via2_5
* cell instance $9632 r0 *1 28.975,17.57
X$9632 421 VIA_via2_5
* cell instance $9633 r0 *1 28.025,25.41
X$9633 421 VIA_via2_5
* cell instance $9634 r0 *1 28.595,23.31
X$9634 421 VIA_via2_5
* cell instance $9635 r0 *1 29.355,23.31
X$9635 421 VIA_via2_5
* cell instance $9636 r0 *1 28.595,33.95
X$9636 421 VIA_via2_5
* cell instance $9637 r0 *1 26.505,33.95
X$9637 421 VIA_via2_5
* cell instance $9638 r0 *1 27.455,33.95
X$9638 421 VIA_via2_5
* cell instance $9639 r0 *1 26.315,23.17
X$9639 421 VIA_via1_4
* cell instance $9640 r0 *1 26.315,23.31
X$9640 421 VIA_via2_5
* cell instance $9641 r0 *1 28.975,16.03
X$9641 421 VIA_via1_4
* cell instance $9642 r0 *1 28.975,18.83
X$9642 421 VIA_via1_4
* cell instance $9643 r0 *1 30.875,17.57
X$9643 421 VIA_via1_4
* cell instance $9644 r0 *1 30.875,17.57
X$9644 421 VIA_via2_5
* cell instance $9645 r0 *1 26.505,34.37
X$9645 421 VIA_via1_4
* cell instance $9646 r0 *1 28.025,31.57
X$9646 421 VIA_via1_4
* cell instance $9647 r0 *1 28.595,42.77
X$9647 421 VIA_via1_4
* cell instance $9648 r0 *1 28.595,42.77
X$9648 421 VIA_via2_5
* cell instance $9649 r0 *1 30.115,42.77
X$9649 421 VIA_via1_4
* cell instance $9650 r0 *1 30.115,42.77
X$9650 421 VIA_via2_5
* cell instance $9651 r0 *1 28.215,37.17
X$9651 421 VIA_via1_4
* cell instance $9652 r0 *1 28.025,38.43
X$9652 421 VIA_via1_4
* cell instance $9653 r0 *1 33.155,48.51
X$9653 422 VIA_via2_5
* cell instance $9654 r0 *1 32.015,17.71
X$9654 422 VIA_via1_4
* cell instance $9655 r0 *1 32.015,17.71
X$9655 422 VIA_via2_5
* cell instance $9656 r0 *1 33.155,49.63
X$9656 422 VIA_via1_4
* cell instance $9657 r0 *1 32.205,48.37
X$9657 422 VIA_via1_4
* cell instance $9658 r0 *1 32.205,48.37
X$9658 422 VIA_via2_5
* cell instance $9659 r0 *1 31.735,17.71
X$9659 422 VIA_via3_2
* cell instance $9660 r0 *1 31.735,48.37
X$9660 422 VIA_via3_2
* cell instance $9661 r0 *1 35.245,18.55
X$9661 423 VIA_via1_4
* cell instance $9662 r0 *1 35.815,49.56
X$9662 423 VIA_via1_4
* cell instance $9663 r0 *1 36.005,48.37
X$9663 423 VIA_via1_4
* cell instance $9664 r0 *1 36.005,48.37
X$9664 423 VIA_via2_5
* cell instance $9665 r0 *1 35.375,48.23
X$9665 423 VIA_via3_2
* cell instance $9666 r0 *1 35.375,18.27
X$9666 423 VIA_via3_2
* cell instance $9667 r0 *1 35.245,18.27
X$9667 423 VIA_via2_5
* cell instance $9668 r0 *1 58.425,16.59
X$9668 424 VIA_via1_7
* cell instance $9669 r0 *1 58.425,17.57
X$9669 424 VIA_via1_4
* cell instance $9670 r0 *1 40.565,17.57
X$9670 425 VIA_via1_4
* cell instance $9671 r0 *1 40.565,16.31
X$9671 425 VIA_via1_4
* cell instance $9672 r0 *1 56.335,51.31
X$9672 426 VIA_via2_5
* cell instance $9673 r0 *1 53.295,17.85
X$9673 426 VIA_via1_4
* cell instance $9674 r0 *1 53.295,17.85
X$9674 426 VIA_via2_5
* cell instance $9675 r0 *1 54.055,51.17
X$9675 426 VIA_via1_4
* cell instance $9676 r0 *1 54.055,51.17
X$9676 426 VIA_via2_5
* cell instance $9677 r0 *1 56.335,52.43
X$9677 426 VIA_via1_4
* cell instance $9678 r0 *1 53.855,17.85
X$9678 426 VIA_via3_2
* cell instance $9679 r0 *1 53.855,51.17
X$9679 426 VIA_via3_2
* cell instance $9680 r0 *1 54.815,17.57
X$9680 427 VIA_via1_4
* cell instance $9681 r0 *1 54.815,17.57
X$9681 427 VIA_via2_5
* cell instance $9682 r0 *1 53.105,17.57
X$9682 427 VIA_via1_4
* cell instance $9683 r0 *1 53.105,17.57
X$9683 427 VIA_via2_5
* cell instance $9684 r0 *1 40.755,17.71
X$9684 428 VIA_via1_4
* cell instance $9685 r0 *1 40.755,17.71
X$9685 428 VIA_via2_5
* cell instance $9686 r0 *1 40.695,17.71
X$9686 428 VIA_via3_2
* cell instance $9687 r0 *1 39.235,51.17
X$9687 428 VIA_via1_4
* cell instance $9688 r0 *1 39.235,51.17
X$9688 428 VIA_via2_5
* cell instance $9689 r0 *1 40.755,53.97
X$9689 428 VIA_via1_4
* cell instance $9690 r0 *1 40.755,53.83
X$9690 428 VIA_via2_5
* cell instance $9691 r0 *1 40.135,53.83
X$9691 428 VIA_via3_2
* cell instance $9692 r0 *1 39.855,51.17
X$9692 428 VIA_via3_2
* cell instance $9693 r0 *1 41.325,17.57
X$9693 429 VIA_via1_4
* cell instance $9694 r0 *1 41.325,14.63
X$9694 429 VIA_via1_4
* cell instance $9695 r0 *1 44.555,13.79
X$9695 430 VIA_via1_7
* cell instance $9696 r0 *1 45.315,17.85
X$9696 430 VIA_via2_5
* cell instance $9697 r0 *1 44.555,17.85
X$9697 430 VIA_via2_5
* cell instance $9698 r0 *1 45.315,18.83
X$9698 430 VIA_via1_4
* cell instance $9699 r0 *1 13.205,16.59
X$9699 431 VIA_via1_7
* cell instance $9700 r0 *1 13.585,23.17
X$9700 431 VIA_via1_4
* cell instance $9701 r0 *1 19.475,18.83
X$9701 432 VIA_via2_5
* cell instance $9702 r0 *1 18.715,18.83
X$9702 432 VIA_via1_4
* cell instance $9703 r0 *1 18.715,18.83
X$9703 432 VIA_via2_5
* cell instance $9704 r0 *1 19.475,17.85
X$9704 432 VIA_via1_4
* cell instance $9705 r0 *1 16.435,18.83
X$9705 432 VIA_via1_4
* cell instance $9706 r0 *1 16.435,18.83
X$9706 432 VIA_via2_5
* cell instance $9707 r0 *1 21.565,50.75
X$9707 433 VIA_via2_5
* cell instance $9708 r0 *1 22.515,50.75
X$9708 433 VIA_via2_5
* cell instance $9709 r0 *1 20.045,51.45
X$9709 433 VIA_via2_5
* cell instance $9710 r0 *1 21.565,51.17
X$9710 433 VIA_via1_4
* cell instance $9711 r0 *1 21.565,51.31
X$9711 433 VIA_via2_5
* cell instance $9712 r0 *1 20.045,51.17
X$9712 433 VIA_via1_4
* cell instance $9713 r0 *1 21.185,17.71
X$9713 433 VIA_via1_4
* cell instance $9714 r0 *1 48.535,50.47
X$9714 434 VIA_via6_0
* cell instance $9715 r0 *1 25.015,49.63
X$9715 434 VIA_via5_0
* cell instance $9716 r0 *1 25.015,49.67
X$9716 434 VIA_via6_0
* cell instance $9717 r0 *1 25.015,49.63
X$9717 434 VIA_via4_0
* cell instance $9718 r0 *1 23.275,67.97
X$9718 434 VIA_via2_5
* cell instance $9719 r0 *1 75.525,50.33
X$9719 434 VIA_via2_5
* cell instance $9720 r0 *1 26.125,32.83
X$9720 434 VIA_via2_5
* cell instance $9721 r0 *1 24.795,67.97
X$9721 434 VIA_via2_5
* cell instance $9722 r0 *1 73.435,80.43
X$9722 434 VIA_via1_4
* cell instance $9723 r0 *1 73.435,80.43
X$9723 434 VIA_via2_5
* cell instance $9724 r0 *1 74.005,31.57
X$9724 434 VIA_via1_4
* cell instance $9725 r0 *1 74.015,31.57
X$9725 434 VIA_via3_2
* cell instance $9726 r0 *1 74.005,31.57
X$9726 434 VIA_via2_5
* cell instance $9727 r0 *1 74.005,18.83
X$9727 434 VIA_via1_4
* cell instance $9728 r0 *1 74.015,18.83
X$9728 434 VIA_via3_2
* cell instance $9729 r0 *1 74.005,18.83
X$9729 434 VIA_via2_5
* cell instance $9730 r0 *1 25.745,18.83
X$9730 434 VIA_via1_4
* cell instance $9731 r0 *1 24.985,77.63
X$9731 434 VIA_via1_4
* cell instance $9732 r0 *1 23.085,67.97
X$9732 434 VIA_via1_4
* cell instance $9733 r0 *1 75.145,66.43
X$9733 434 VIA_via1_4
* cell instance $9734 r0 *1 75.145,66.43
X$9734 434 VIA_via2_5
* cell instance $9735 r0 *1 50.065,50.05
X$9735 434 VIA_via1_4
* cell instance $9736 r0 *1 50.065,50.19
X$9736 434 VIA_via2_5
* cell instance $9737 r0 *1 24.985,32.83
X$9737 434 VIA_via1_4
* cell instance $9738 r0 *1 25.015,32.83
X$9738 434 VIA_via3_2
* cell instance $9739 r0 *1 24.985,32.83
X$9739 434 VIA_via2_5
* cell instance $9740 r0 *1 48.535,50.19
X$9740 434 VIA_via4_0
* cell instance $9741 r0 *1 48.535,50.19
X$9741 434 VIA_via3_2
* cell instance $9742 r0 *1 48.535,50.19
X$9742 434 VIA_via5_0
* cell instance $9743 r0 *1 73.735,49.35
X$9743 434 VIA_via4_0
* cell instance $9744 r0 *1 50.215,49.35
X$9744 434 VIA_via4_0
* cell instance $9745 r0 *1 75.415,66.43
X$9745 434 VIA_via3_2
* cell instance $9746 r0 *1 73.735,50.33
X$9746 434 VIA_via3_2
* cell instance $9747 r0 *1 50.215,50.19
X$9747 434 VIA_via3_2
* cell instance $9748 r0 *1 75.415,80.43
X$9748 434 VIA_via3_2
* cell instance $9749 r0 *1 25.015,67.97
X$9749 434 VIA_via3_2
* cell instance $9750 r0 *1 37.145,19.81
X$9750 435 VIA_via1_7
* cell instance $9751 r0 *1 35.625,18.55
X$9751 435 VIA_via2_5
* cell instance $9752 r0 *1 37.145,18.55
X$9752 435 VIA_via2_5
* cell instance $9753 r0 *1 35.435,18.76
X$9753 435 VIA_via1_4
* cell instance $9754 r0 *1 41.515,20.09
X$9754 436 VIA_via1_4
* cell instance $9755 r0 *1 40.375,17.57
X$9755 436 VIA_via1_4
* cell instance $9756 r0 *1 11.305,23.03
X$9756 437 VIA_via1_7
* cell instance $9757 r0 *1 34.295,21.77
X$9757 437 VIA_via1_7
* cell instance $9758 r0 *1 34.295,21.77
X$9758 437 VIA_via2_5
* cell instance $9759 r0 *1 48.165,18.97
X$9759 437 VIA_via1_7
* cell instance $9760 r0 *1 45.125,21.77
X$9760 437 VIA_via1_7
* cell instance $9761 r0 *1 45.125,21.77
X$9761 437 VIA_via2_5
* cell instance $9762 r0 *1 48.355,21.77
X$9762 437 VIA_via2_5
* cell instance $9763 r0 *1 28.215,21.77
X$9763 437 VIA_via2_5
* cell instance $9764 r0 *1 38.855,21.77
X$9764 437 VIA_via2_5
* cell instance $9765 r0 *1 12.825,20.79
X$9765 437 VIA_via2_5
* cell instance $9766 r0 *1 12.825,20.09
X$9766 437 VIA_via2_5
* cell instance $9767 r0 *1 19.095,20.79
X$9767 437 VIA_via2_5
* cell instance $9768 r0 *1 23.655,21.77
X$9768 437 VIA_via2_5
* cell instance $9769 r0 *1 19.095,21.77
X$9769 437 VIA_via2_5
* cell instance $9770 r0 *1 11.115,20.09
X$9770 437 VIA_via2_5
* cell instance $9771 r0 *1 17.385,20.79
X$9771 437 VIA_via2_5
* cell instance $9772 r0 *1 38.855,23.17
X$9772 437 VIA_via1_4
* cell instance $9773 r0 *1 48.355,22.75
X$9773 437 VIA_via1_4
* cell instance $9774 r0 *1 28.215,18.83
X$9774 437 VIA_via1_4
* cell instance $9775 r0 *1 17.385,21.63
X$9775 437 VIA_via1_4
* cell instance $9776 r0 *1 12.825,18.83
X$9776 437 VIA_via1_4
* cell instance $9777 r0 *1 19.095,20.37
X$9777 437 VIA_via1_4
* cell instance $9778 r0 *1 23.655,23.17
X$9778 437 VIA_via1_4
* cell instance $9779 r0 *1 75.335,18.97
X$9779 438 VIA_via1_7
* cell instance $9780 r0 *1 82.555,30.17
X$9780 438 VIA_via1_7
* cell instance $9781 r0 *1 77.425,23.03
X$9781 438 VIA_via1_7
* cell instance $9782 r0 *1 71.155,37.03
X$9782 438 VIA_via1_7
* cell instance $9783 r0 *1 71.155,37.03
X$9783 438 VIA_via2_5
* cell instance $9784 r0 *1 77.615,20.93
X$9784 438 VIA_via2_5
* cell instance $9785 r0 *1 75.145,19.53
X$9785 438 VIA_via2_5
* cell instance $9786 r0 *1 75.145,20.93
X$9786 438 VIA_via2_5
* cell instance $9787 r0 *1 69.065,19.53
X$9787 438 VIA_via2_5
* cell instance $9788 r0 *1 69.065,20.93
X$9788 438 VIA_via2_5
* cell instance $9789 r0 *1 71.155,35.77
X$9789 438 VIA_via2_5
* cell instance $9790 r0 *1 61.845,20.93
X$9790 438 VIA_via2_5
* cell instance $9791 r0 *1 62.415,20.93
X$9791 438 VIA_via2_5
* cell instance $9792 r0 *1 82.175,35.77
X$9792 438 VIA_via2_5
* cell instance $9793 r0 *1 66.215,43.61
X$9793 438 VIA_via2_5
* cell instance $9794 r0 *1 65.835,37.45
X$9794 438 VIA_via2_5
* cell instance $9795 r0 *1 65.835,37.03
X$9795 438 VIA_via2_5
* cell instance $9796 r0 *1 75.335,43.61
X$9796 438 VIA_via2_5
* cell instance $9797 r0 *1 61.845,23.45
X$9797 438 VIA_via2_5
* cell instance $9798 r0 *1 62.225,23.45
X$9798 438 VIA_via2_5
* cell instance $9799 r0 *1 82.175,31.57
X$9799 438 VIA_via1_4
* cell instance $9800 r0 *1 75.335,44.03
X$9800 438 VIA_via1_4
* cell instance $9801 r0 *1 62.035,36.75
X$9801 438 VIA_via1_4
* cell instance $9802 r0 *1 62.415,37.45
X$9802 438 VIA_via1_4
* cell instance $9803 r0 *1 62.415,37.45
X$9803 438 VIA_via2_5
* cell instance $9804 r0 *1 66.215,44.03
X$9804 438 VIA_via1_4
* cell instance $9805 r0 *1 61.845,27.23
X$9805 438 VIA_via1_4
* cell instance $9806 r0 *1 69.065,18.83
X$9806 438 VIA_via1_4
* cell instance $9807 r0 *1 61.845,18.83
X$9807 438 VIA_via1_4
* cell instance $9808 r0 *1 62.225,17.85
X$9808 439 VIA_via1_4
* cell instance $9809 r0 *1 60.705,18.83
X$9809 439 VIA_via1_4
* cell instance $9810 r0 *1 60.705,18.83
X$9810 439 VIA_via2_5
* cell instance $9811 r0 *1 62.035,18.83
X$9811 439 VIA_via1_4
* cell instance $9812 r0 *1 62.035,18.83
X$9812 439 VIA_via2_5
* cell instance $9813 r0 *1 64.885,19.39
X$9813 440 VIA_via1_7
* cell instance $9814 r0 *1 65.075,20.37
X$9814 440 VIA_via1_4
* cell instance $9815 r0 *1 68.495,28.63
X$9815 441 VIA_via1_7
* cell instance $9816 r0 *1 75.145,24.57
X$9816 441 VIA_via1_7
* cell instance $9817 r0 *1 75.525,73.43
X$9817 441 VIA_via1_7
* cell instance $9818 r0 *1 73.245,62.23
X$9818 441 VIA_via1_7
* cell instance $9819 r0 *1 73.245,62.09
X$9819 441 VIA_via2_5
* cell instance $9820 r0 *1 60.515,18.97
X$9820 441 VIA_via1_7
* cell instance $9821 r0 *1 63.175,70.63
X$9821 441 VIA_via1_7
* cell instance $9822 r0 *1 63.175,70.63
X$9822 441 VIA_via2_5
* cell instance $9823 r0 *1 60.515,19.25
X$9823 441 VIA_via2_5
* cell instance $9824 r0 *1 73.435,69.93
X$9824 441 VIA_via2_5
* cell instance $9825 r0 *1 73.435,71.19
X$9825 441 VIA_via2_5
* cell instance $9826 r0 *1 63.745,54.25
X$9826 441 VIA_via2_5
* cell instance $9827 r0 *1 64.505,54.25
X$9827 441 VIA_via2_5
* cell instance $9828 r0 *1 64.125,71.05
X$9828 441 VIA_via2_5
* cell instance $9829 r0 *1 64.125,70.63
X$9829 441 VIA_via2_5
* cell instance $9830 r0 *1 64.315,62.09
X$9830 441 VIA_via2_5
* cell instance $9831 r0 *1 69.635,69.93
X$9831 441 VIA_via2_5
* cell instance $9832 r0 *1 69.635,71.05
X$9832 441 VIA_via2_5
* cell instance $9833 r0 *1 76.095,71.19
X$9833 441 VIA_via2_5
* cell instance $9834 r0 *1 67.735,19.25
X$9834 441 VIA_via2_5
* cell instance $9835 r0 *1 72.675,18.55
X$9835 441 VIA_via2_5
* cell instance $9836 r0 *1 68.495,25.13
X$9836 441 VIA_via2_5
* cell instance $9837 r0 *1 67.925,25.13
X$9837 441 VIA_via2_5
* cell instance $9838 r0 *1 75.145,24.99
X$9838 441 VIA_via2_5
* cell instance $9839 r0 *1 63.745,43.33
X$9839 441 VIA_via2_5
* cell instance $9840 r0 *1 73.625,43.33
X$9840 441 VIA_via2_5
* cell instance $9841 r0 *1 67.735,18.55
X$9841 441 VIA_via2_5
* cell instance $9842 r0 *1 67.925,43.33
X$9842 441 VIA_via2_5
* cell instance $9843 r0 *1 63.745,42.77
X$9843 441 VIA_via1_4
* cell instance $9844 r0 *1 74.005,44.03
X$9844 441 VIA_via1_4
* cell instance $9845 r0 *1 67.735,18.83
X$9845 441 VIA_via1_4
* cell instance $9846 r0 *1 72.675,18.83
X$9846 441 VIA_via1_4
* cell instance $9847 r0 *1 61.655,54.25
X$9847 441 VIA_via1_4
* cell instance $9848 r0 *1 61.655,54.25
X$9848 441 VIA_via2_5
* cell instance $9849 r0 *1 70.015,20.37
X$9849 442 VIA_via1_4
* cell instance $9850 r0 *1 70.585,19.11
X$9850 442 VIA_via1_4
* cell instance $9851 r0 *1 77.995,19.11
X$9851 443 VIA_via1_4
* cell instance $9852 r0 *1 77.615,20.37
X$9852 443 VIA_via1_4
* cell instance $9853 r0 *1 81.225,20.37
X$9853 444 VIA_via2_5
* cell instance $9854 r0 *1 81.415,18.55
X$9854 444 VIA_via1_4
* cell instance $9855 r0 *1 79.895,20.37
X$9855 444 VIA_via1_4
* cell instance $9856 r0 *1 79.895,20.37
X$9856 444 VIA_via2_5
* cell instance $9857 r0 *1 78.755,20.37
X$9857 444 VIA_via1_4
* cell instance $9858 r0 *1 78.755,20.37
X$9858 444 VIA_via2_5
* cell instance $9859 r0 *1 77.995,23.03
X$9859 445 VIA_via2_5
* cell instance $9860 r0 *1 81.415,18.83
X$9860 445 VIA_via2_5
* cell instance $9861 r0 *1 83.695,18.83
X$9861 445 VIA_via2_5
* cell instance $9862 r0 *1 84.835,21.63
X$9862 445 VIA_via2_5
* cell instance $9863 r0 *1 77.995,25.97
X$9863 445 VIA_via2_5
* cell instance $9864 r0 *1 84.835,23.17
X$9864 445 VIA_via1_4
* cell instance $9865 r0 *1 84.835,23.03
X$9865 445 VIA_via2_5
* cell instance $9866 r0 *1 81.415,23.17
X$9866 445 VIA_via1_4
* cell instance $9867 r0 *1 81.415,23.03
X$9867 445 VIA_via2_5
* cell instance $9868 r0 *1 85.025,20.37
X$9868 445 VIA_via1_4
* cell instance $9869 r0 *1 79.895,18.83
X$9869 445 VIA_via1_4
* cell instance $9870 r0 *1 79.895,18.83
X$9870 445 VIA_via2_5
* cell instance $9871 r0 *1 77.995,21.63
X$9871 445 VIA_via1_4
* cell instance $9872 r0 *1 77.995,24.43
X$9872 445 VIA_via1_4
* cell instance $9873 r0 *1 83.695,17.57
X$9873 445 VIA_via1_4
* cell instance $9874 r0 *1 72.865,25.97
X$9874 445 VIA_via1_4
* cell instance $9875 r0 *1 72.865,25.97
X$9875 445 VIA_via2_5
* cell instance $9876 r0 *1 87.305,21.63
X$9876 445 VIA_via1_4
* cell instance $9877 r0 *1 87.305,21.63
X$9877 445 VIA_via2_5
* cell instance $9878 r0 *1 6.175,21.21
X$9878 446 VIA_via1_7
* cell instance $9879 r0 *1 2.945,19.11
X$9879 446 VIA_via2_5
* cell instance $9880 r0 *1 6.175,19.11
X$9880 446 VIA_via2_5
* cell instance $9881 r0 *1 2.945,18.83
X$9881 446 VIA_via1_4
* cell instance $9882 r0 *1 4.085,20.79
X$9882 447 VIA_via2_5
* cell instance $9883 r0 *1 7.505,20.79
X$9883 447 VIA_via2_5
* cell instance $9884 r0 *1 4.465,18.97
X$9884 447 VIA_via2_5
* cell instance $9885 r0 *1 3.705,20.79
X$9885 447 VIA_via2_5
* cell instance $9886 r0 *1 9.595,20.79
X$9886 447 VIA_via2_5
* cell instance $9887 r0 *1 7.885,18.97
X$9887 447 VIA_via2_5
* cell instance $9888 r0 *1 9.595,23.17
X$9888 447 VIA_via1_4
* cell instance $9889 r0 *1 6.935,19.95
X$9889 447 VIA_via1_4
* cell instance $9890 r0 *1 7.315,20.79
X$9890 447 VIA_via1_7
* cell instance $9891 r0 *1 7.315,20.79
X$9891 447 VIA_via2_5
* cell instance $9892 r0 *1 7.505,20.37
X$9892 447 VIA_via1_4
* cell instance $9893 r0 *1 6.935,18.83
X$9893 447 VIA_via1_4
* cell instance $9894 r0 *1 6.935,18.97
X$9894 447 VIA_via2_5
* cell instance $9895 r0 *1 3.705,18.83
X$9895 447 VIA_via1_4
* cell instance $9896 r0 *1 3.705,18.97
X$9896 447 VIA_via2_5
* cell instance $9897 r0 *1 3.895,23.17
X$9897 447 VIA_via1_4
* cell instance $9898 r0 *1 3.515,20.37
X$9898 447 VIA_via1_4
* cell instance $9899 r0 *1 7.885,17.57
X$9899 447 VIA_via1_4
* cell instance $9900 r0 *1 4.465,14.77
X$9900 447 VIA_via1_4
* cell instance $9901 r0 *1 5.985,19.25
X$9901 448 VIA_via2_5
* cell instance $9902 r0 *1 5.985,20.37
X$9902 448 VIA_via1_4
* cell instance $9903 r0 *1 5.225,19.25
X$9903 448 VIA_via1_4
* cell instance $9904 r0 *1 5.225,19.25
X$9904 448 VIA_via2_5
* cell instance $9905 r0 *1 5.225,21.63
X$9905 448 VIA_via1_4
* cell instance $9906 r0 *1 7.125,19.11
X$9906 449 VIA_via2_5
* cell instance $9907 r0 *1 9.785,19.11
X$9907 449 VIA_via1_4
* cell instance $9908 r0 *1 9.785,19.11
X$9908 449 VIA_via2_5
* cell instance $9909 r0 *1 7.125,17.57
X$9909 449 VIA_via1_4
* cell instance $9910 r0 *1 9.785,19.81
X$9910 450 VIA_via1_7
* cell instance $9911 r0 *1 9.595,18.83
X$9911 450 VIA_via2_5
* cell instance $9912 r0 *1 6.175,18.83
X$9912 450 VIA_via1_4
* cell instance $9913 r0 *1 6.175,18.83
X$9913 450 VIA_via2_5
* cell instance $9914 r0 *1 15.675,18.83
X$9914 451 VIA_via1_4
* cell instance $9915 r0 *1 15.675,18.83
X$9915 451 VIA_via2_5
* cell instance $9916 r0 *1 15.675,19.95
X$9916 451 VIA_via1_4
* cell instance $9917 r0 *1 13.015,18.83
X$9917 451 VIA_via1_4
* cell instance $9918 r0 *1 13.015,18.83
X$9918 451 VIA_via2_5
* cell instance $9919 r0 *1 76.475,18.83
X$9919 452 VIA_via1_4
* cell instance $9920 r0 *1 76.665,18.83
X$9920 452 VIA_via1_4
* cell instance $9921 r0 *1 18.145,25.41
X$9921 453 VIA_via1_7
* cell instance $9922 r0 *1 18.145,25.27
X$9922 453 VIA_via2_5
* cell instance $9923 r0 *1 10.925,41.09
X$9923 453 VIA_via2_5
* cell instance $9924 r0 *1 9.215,40.11
X$9924 453 VIA_via2_5
* cell instance $9925 r0 *1 8.645,40.11
X$9925 453 VIA_via2_5
* cell instance $9926 r0 *1 9.405,25.27
X$9926 453 VIA_via2_5
* cell instance $9927 r0 *1 9.405,32.69
X$9927 453 VIA_via2_5
* cell instance $9928 r0 *1 19.665,40.95
X$9928 453 VIA_via2_5
* cell instance $9929 r0 *1 20.425,40.25
X$9929 453 VIA_via2_5
* cell instance $9930 r0 *1 19.665,40.25
X$9930 453 VIA_via2_5
* cell instance $9931 r0 *1 20.045,25.27
X$9931 453 VIA_via2_5
* cell instance $9932 r0 *1 19.855,18.69
X$9932 453 VIA_via2_5
* cell instance $9933 r0 *1 18.715,25.27
X$9933 453 VIA_via2_5
* cell instance $9934 r0 *1 9.405,18.83
X$9934 453 VIA_via1_4
* cell instance $9935 r0 *1 9.405,20.37
X$9935 453 VIA_via1_4
* cell instance $9936 r0 *1 9.025,32.83
X$9936 453 VIA_via1_4
* cell instance $9937 r0 *1 9.025,32.69
X$9937 453 VIA_via2_5
* cell instance $9938 r0 *1 10.925,39.97
X$9938 453 VIA_via1_4
* cell instance $9939 r0 *1 10.925,40.11
X$9939 453 VIA_via2_5
* cell instance $9940 r0 *1 8.645,41.23
X$9940 453 VIA_via1_4
* cell instance $9941 r0 *1 20.425,39.97
X$9941 453 VIA_via1_4
* cell instance $9942 r0 *1 17.005,18.83
X$9942 453 VIA_via1_4
* cell instance $9943 r0 *1 17.005,18.69
X$9943 453 VIA_via2_5
* cell instance $9944 r0 *1 19.855,20.37
X$9944 453 VIA_via1_4
* cell instance $9945 r0 *1 18.715,25.97
X$9945 453 VIA_via1_4
* cell instance $9946 r0 *1 17.575,41.23
X$9946 453 VIA_via1_4
* cell instance $9947 r0 *1 17.575,41.09
X$9947 453 VIA_via2_5
* cell instance $9948 r0 *1 75.145,18.41
X$9948 454 VIA_via2_5
* cell instance $9949 r0 *1 75.525,18.41
X$9949 454 VIA_via2_5
* cell instance $9950 r0 *1 72.865,18.41
X$9950 454 VIA_via2_5
* cell instance $9951 r0 *1 75.525,18.83
X$9951 454 VIA_via1_4
* cell instance $9952 r0 *1 75.145,17.85
X$9952 454 VIA_via1_4
* cell instance $9953 r0 *1 72.865,18.83
X$9953 454 VIA_via1_4
* cell instance $9954 r0 *1 25.175,18.41
X$9954 455 VIA_via1_7
* cell instance $9955 r0 *1 25.175,17.57
X$9955 455 VIA_via1_4
* cell instance $9956 r0 *1 70.395,18.83
X$9956 456 VIA_via1_4
* cell instance $9957 r0 *1 70.205,18.83
X$9957 456 VIA_via1_4
* cell instance $9958 r0 *1 69.255,18.83
X$9958 457 VIA_via1_4
* cell instance $9959 r0 *1 69.255,18.97
X$9959 457 VIA_via2_5
* cell instance $9960 r0 *1 67.925,18.83
X$9960 457 VIA_via1_4
* cell instance $9961 r0 *1 67.925,18.97
X$9961 457 VIA_via2_5
* cell instance $9962 r0 *1 69.255,19.95
X$9962 457 VIA_via1_4
* cell instance $9963 r0 *1 32.585,19.81
X$9963 458 VIA_via1_7
* cell instance $9964 r0 *1 32.585,18.69
X$9964 458 VIA_via2_5
* cell instance $9965 r0 *1 34.485,18.83
X$9965 458 VIA_via1_4
* cell instance $9966 r0 *1 34.485,18.69
X$9966 458 VIA_via2_5
* cell instance $9967 r0 *1 35.625,18.97
X$9967 459 VIA_via1_4
* cell instance $9968 r0 *1 35.625,18.97
X$9968 459 VIA_via2_5
* cell instance $9969 r0 *1 34.295,18.83
X$9969 459 VIA_via1_4
* cell instance $9970 r0 *1 34.295,18.97
X$9970 459 VIA_via2_5
* cell instance $9971 r0 *1 43.605,48.65
X$9971 460 VIA_via2_5
* cell instance $9972 r0 *1 44.745,48.65
X$9972 460 VIA_via2_5
* cell instance $9973 r0 *1 45.505,18.55
X$9973 460 VIA_via1_4
* cell instance $9974 r0 *1 45.505,18.55
X$9974 460 VIA_via2_5
* cell instance $9975 r0 *1 45.455,18.55
X$9975 460 VIA_via3_2
* cell instance $9976 r0 *1 43.605,49.63
X$9976 460 VIA_via1_4
* cell instance $9977 r0 *1 44.745,48.37
X$9977 460 VIA_via1_4
* cell instance $9978 r0 *1 45.455,48.65
X$9978 460 VIA_via3_2
* cell instance $9979 r0 *1 64.505,18.83
X$9979 461 VIA_via1_4
* cell instance $9980 r0 *1 64.505,18.97
X$9980 461 VIA_via2_5
* cell instance $9981 r0 *1 62.985,18.97
X$9981 461 VIA_via1_4
* cell instance $9982 r0 *1 62.985,18.97
X$9982 461 VIA_via2_5
* cell instance $9983 r0 *1 61.655,18.41
X$9983 462 VIA_via1_7
* cell instance $9984 r0 *1 61.655,18.41
X$9984 462 VIA_via2_5
* cell instance $9985 r0 *1 59.945,18.41
X$9985 462 VIA_via2_5
* cell instance $9986 r0 *1 59.945,17.57
X$9986 462 VIA_via1_4
* cell instance $9987 r0 *1 48.355,18.83
X$9987 463 VIA_via1_4
* cell instance $9988 r0 *1 48.355,18.83
X$9988 463 VIA_via2_5
* cell instance $9989 r0 *1 50.255,18.83
X$9989 463 VIA_via1_4
* cell instance $9990 r0 *1 50.255,18.83
X$9990 463 VIA_via2_5
* cell instance $9991 r0 *1 50.255,16.45
X$9991 463 VIA_via1_4
* cell instance $9992 r0 *1 50.635,18.83
X$9992 464 VIA_via1_4
* cell instance $9993 r0 *1 51.965,18.83
X$9993 464 VIA_via1_4
* cell instance $9994 r0 *1 3.895,20.65
X$9994 465 VIA_via2_5
* cell instance $9995 r0 *1 5.035,20.65
X$9995 465 VIA_via1_4
* cell instance $9996 r0 *1 5.035,20.65
X$9996 465 VIA_via2_5
* cell instance $9997 r0 *1 3.895,21.63
X$9997 465 VIA_via1_4
* cell instance $9998 r0 *1 5.415,20.37
X$9998 465 VIA_via1_4
* cell instance $9999 r0 *1 19.285,18.83
X$9999 466 VIA_via1_4
* cell instance $10000 r0 *1 19.285,20.37
X$10000 466 VIA_via1_4
* cell instance $10001 r0 *1 19.285,20.23
X$10001 466 VIA_via2_5
* cell instance $10002 r0 *1 23.465,20.23
X$10002 466 VIA_via1_4
* cell instance $10003 r0 *1 23.465,20.23
X$10003 466 VIA_via2_5
* cell instance $10004 r0 *1 25.365,21.21
X$10004 467 VIA_via1_7
* cell instance $10005 r0 *1 24.985,18.83
X$10005 467 VIA_via1_4
* cell instance $10006 r0 *1 30.115,19.95
X$10006 468 VIA_via2_5
* cell instance $10007 r0 *1 28.405,19.95
X$10007 468 VIA_via2_5
* cell instance $10008 r0 *1 30.115,20.37
X$10008 468 VIA_via1_4
* cell instance $10009 r0 *1 29.165,19.95
X$10009 468 VIA_via1_4
* cell instance $10010 r0 *1 29.165,19.95
X$10010 468 VIA_via2_5
* cell instance $10011 r0 *1 28.405,18.83
X$10011 468 VIA_via1_4
* cell instance $10012 r0 *1 31.255,19.81
X$10012 469 VIA_via1_7
* cell instance $10013 r0 *1 31.635,17.57
X$10013 469 VIA_via1_4
* cell instance $10014 r0 *1 36.195,21.07
X$10014 470 VIA_via2_5
* cell instance $10015 r0 *1 32.965,21.07
X$10015 470 VIA_via2_5
* cell instance $10016 r0 *1 36.195,20.37
X$10016 470 VIA_via1_4
* cell instance $10017 r0 *1 32.965,21.63
X$10017 470 VIA_via1_4
* cell instance $10018 r0 *1 35.815,19.95
X$10018 470 VIA_via1_4
* cell instance $10019 r0 *1 45.505,20.09
X$10019 471 VIA_via1_4
* cell instance $10020 r0 *1 44.555,18.83
X$10020 471 VIA_via1_4
* cell instance $10021 r0 *1 18.525,18.97
X$10021 472 VIA_via1_7
* cell instance $10022 r0 *1 49.495,20.37
X$10022 472 VIA_via2_5
* cell instance $10023 r0 *1 51.015,20.37
X$10023 472 VIA_via2_5
* cell instance $10024 r0 *1 36.005,20.93
X$10024 472 VIA_via2_5
* cell instance $10025 r0 *1 29.355,20.93
X$10025 472 VIA_via2_5
* cell instance $10026 r0 *1 47.405,20.37
X$10026 472 VIA_via2_5
* cell instance $10027 r0 *1 47.405,20.93
X$10027 472 VIA_via2_5
* cell instance $10028 r0 *1 43.985,20.93
X$10028 472 VIA_via2_5
* cell instance $10029 r0 *1 40.185,20.93
X$10029 472 VIA_via2_5
* cell instance $10030 r0 *1 24.225,20.93
X$10030 472 VIA_via2_5
* cell instance $10031 r0 *1 14.915,20.93
X$10031 472 VIA_via2_5
* cell instance $10032 r0 *1 16.055,20.93
X$10032 472 VIA_via2_5
* cell instance $10033 r0 *1 18.525,20.93
X$10033 472 VIA_via2_5
* cell instance $10034 r0 *1 40.185,23.17
X$10034 472 VIA_via1_4
* cell instance $10035 r0 *1 47.405,23.17
X$10035 472 VIA_via1_4
* cell instance $10036 r0 *1 43.985,20.37
X$10036 472 VIA_via1_4
* cell instance $10037 r0 *1 29.355,20.37
X$10037 472 VIA_via1_4
* cell instance $10038 r0 *1 36.005,20.37
X$10038 472 VIA_via1_4
* cell instance $10039 r0 *1 51.015,21.63
X$10039 472 VIA_via1_4
* cell instance $10040 r0 *1 49.495,18.83
X$10040 472 VIA_via1_4
* cell instance $10041 r0 *1 16.055,21.63
X$10041 472 VIA_via1_4
* cell instance $10042 r0 *1 14.915,18.83
X$10042 472 VIA_via1_4
* cell instance $10043 r0 *1 24.225,21.63
X$10043 472 VIA_via1_4
* cell instance $10044 r0 *1 61.465,10.99
X$10044 473 VIA_via1_7
* cell instance $10045 r0 *1 61.465,23.17
X$10045 473 VIA_via2_5
* cell instance $10046 r0 *1 60.515,23.17
X$10046 473 VIA_via1_4
* cell instance $10047 r0 *1 60.515,23.17
X$10047 473 VIA_via2_5
* cell instance $10048 r0 *1 85.025,48.37
X$10048 474 VIA_via2_5
* cell instance $10049 r0 *1 66.025,37.31
X$10049 474 VIA_via2_5
* cell instance $10050 r0 *1 77.235,37.45
X$10050 474 VIA_via2_5
* cell instance $10051 r0 *1 77.615,48.37
X$10051 474 VIA_via2_5
* cell instance $10052 r0 *1 85.215,48.37
X$10052 474 VIA_via1_4
* cell instance $10053 r0 *1 85.215,48.37
X$10053 474 VIA_via2_5
* cell instance $10054 r0 *1 66.025,20.65
X$10054 474 VIA_via1_4
* cell instance $10055 r0 *1 85.025,51.17
X$10055 474 VIA_via1_4
* cell instance $10056 r0 *1 68.115,52.29
X$10056 475 VIA_via1_7
* cell instance $10057 r0 *1 68.115,52.29
X$10057 475 VIA_via2_5
* cell instance $10058 r0 *1 68.135,52.29
X$10058 475 VIA_via3_2
* cell instance $10059 r0 *1 76.285,23.45
X$10059 475 VIA_via2_5
* cell instance $10060 r0 *1 76.475,23.45
X$10060 475 VIA_via2_5
* cell instance $10061 r0 *1 76.475,20.09
X$10061 475 VIA_via2_5
* cell instance $10062 r0 *1 78.755,23.45
X$10062 475 VIA_via2_5
* cell instance $10063 r0 *1 69.255,52.29
X$10063 475 VIA_via2_5
* cell instance $10064 r0 *1 77.805,67.27
X$10064 475 VIA_via2_5
* cell instance $10065 r0 *1 77.235,67.27
X$10065 475 VIA_via2_5
* cell instance $10066 r0 *1 74.195,35.49
X$10066 475 VIA_via2_5
* cell instance $10067 r0 *1 76.095,35.49
X$10067 475 VIA_via2_5
* cell instance $10068 r0 *1 69.445,46.83
X$10068 475 VIA_via2_5
* cell instance $10069 r0 *1 69.825,20.09
X$10069 475 VIA_via2_5
* cell instance $10070 r0 *1 74.575,46.97
X$10070 475 VIA_via2_5
* cell instance $10071 r0 *1 65.835,69.23
X$10071 475 VIA_via1_4
* cell instance $10072 r0 *1 65.835,69.23
X$10072 475 VIA_via2_5
* cell instance $10073 r0 *1 65.895,69.23
X$10073 475 VIA_via3_2
* cell instance $10074 r0 *1 74.005,35.63
X$10074 475 VIA_via1_4
* cell instance $10075 r0 *1 78.565,46.83
X$10075 475 VIA_via1_4
* cell instance $10076 r0 *1 78.565,46.97
X$10076 475 VIA_via2_5
* cell instance $10077 r0 *1 70.205,46.83
X$10077 475 VIA_via1_4
* cell instance $10078 r0 *1 70.205,46.83
X$10078 475 VIA_via2_5
* cell instance $10079 r0 *1 78.755,23.17
X$10079 475 VIA_via1_4
* cell instance $10080 r0 *1 76.665,20.37
X$10080 475 VIA_via1_4
* cell instance $10081 r0 *1 69.825,20.37
X$10081 475 VIA_via1_4
* cell instance $10082 r0 *1 64.885,20.37
X$10082 475 VIA_via1_4
* cell instance $10083 r0 *1 64.885,20.23
X$10083 475 VIA_via2_5
* cell instance $10084 r0 *1 77.235,69.23
X$10084 475 VIA_via1_4
* cell instance $10085 r0 *1 77.805,62.37
X$10085 475 VIA_via1_4
* cell instance $10086 r0 *1 65.895,68.95
X$10086 475 VIA_via4_0
* cell instance $10087 r0 *1 68.135,68.95
X$10087 475 VIA_via4_0
* cell instance $10088 r0 *1 77.095,68.95
X$10088 475 VIA_via4_0
* cell instance $10089 r0 *1 77.095,68.95
X$10089 475 VIA_via3_2
* cell instance $10090 r0 *1 77.235,68.95
X$10090 475 VIA_via2_5
* cell instance $10091 r0 *1 56.905,60.69
X$10091 476 VIA_via2_5
* cell instance $10092 r0 *1 78.375,62.37
X$10092 476 VIA_via2_5
* cell instance $10093 r0 *1 56.905,47.39
X$10093 476 VIA_via2_5
* cell instance $10094 r0 *1 78.755,47.11
X$10094 476 VIA_via2_5
* cell instance $10095 r0 *1 79.325,47.11
X$10095 476 VIA_via2_5
* cell instance $10096 r0 *1 66.595,69.23
X$10096 476 VIA_via1_4
* cell instance $10097 r0 *1 66.595,69.23
X$10097 476 VIA_via2_5
* cell instance $10098 r0 *1 70.965,46.83
X$10098 476 VIA_via1_4
* cell instance $10099 r0 *1 70.965,46.83
X$10099 476 VIA_via2_5
* cell instance $10100 r0 *1 79.515,23.17
X$10100 476 VIA_via1_4
* cell instance $10101 r0 *1 79.515,23.31
X$10101 476 VIA_via2_5
* cell instance $10102 r0 *1 77.425,20.37
X$10102 476 VIA_via1_4
* cell instance $10103 r0 *1 77.425,20.51
X$10103 476 VIA_via2_5
* cell instance $10104 r0 *1 57.665,43.05
X$10104 476 VIA_via1_4
* cell instance $10105 r0 *1 57.665,43.05
X$10105 476 VIA_via2_5
* cell instance $10106 r0 *1 70.585,20.37
X$10106 476 VIA_via1_4
* cell instance $10107 r0 *1 70.585,20.51
X$10107 476 VIA_via2_5
* cell instance $10108 r0 *1 65.645,20.37
X$10108 476 VIA_via1_4
* cell instance $10109 r0 *1 65.645,20.51
X$10109 476 VIA_via2_5
* cell instance $10110 r0 *1 54.625,60.83
X$10110 476 VIA_via1_4
* cell instance $10111 r0 *1 54.625,60.69
X$10111 476 VIA_via2_5
* cell instance $10112 r0 *1 78.565,62.37
X$10112 476 VIA_via1_4
* cell instance $10113 r0 *1 71.215,46.83
X$10113 476 VIA_via4_0
* cell instance $10114 r0 *1 71.215,46.83
X$10114 476 VIA_via3_2
* cell instance $10115 r0 *1 57.215,46.83
X$10115 476 VIA_via4_0
* cell instance $10116 r0 *1 77.935,69.09
X$10116 476 VIA_via3_2
* cell instance $10117 r0 *1 77.935,69.23
X$10117 476 VIA_via4_0
* cell instance $10118 r0 *1 77.995,69.09
X$10118 476 VIA_via2_5
* cell instance $10119 r0 *1 77.995,69.23
X$10119 476 VIA_via1_4
* cell instance $10120 r0 *1 57.215,43.05
X$10120 476 VIA_via3_2
* cell instance $10121 r0 *1 57.215,47.39
X$10121 476 VIA_via3_2
* cell instance $10122 r0 *1 79.335,23.31
X$10122 476 VIA_via3_2
* cell instance $10123 r0 *1 79.335,20.51
X$10123 476 VIA_via3_2
* cell instance $10124 r0 *1 67.015,69.23
X$10124 476 VIA_via3_2
* cell instance $10125 r0 *1 67.015,69.23
X$10125 476 VIA_via4_0
* cell instance $10126 r0 *1 77.935,62.37
X$10126 476 VIA_via3_2
* cell instance $10127 r0 *1 79.335,46.69
X$10127 476 VIA_via3_2
* cell instance $10128 r0 *1 79.325,46.69
X$10128 476 VIA_via2_5
* cell instance $10129 r0 *1 79.335,46.83
X$10129 476 VIA_via4_0
* cell instance $10130 r0 *1 79.325,46.83
X$10130 476 VIA_via1_4
* cell instance $10131 r0 *1 74.385,23.17
X$10131 477 VIA_via1_4
* cell instance $10132 r0 *1 74.385,20.65
X$10132 477 VIA_via1_4
* cell instance $10133 r0 *1 74.575,21.63
X$10133 477 VIA_via1_4
* cell instance $10134 r0 *1 74.765,22.61
X$10134 478 VIA_via1_7
* cell instance $10135 r0 *1 75.525,20.37
X$10135 478 VIA_via1_4
* cell instance $10136 r0 *1 82.935,20.37
X$10136 479 VIA_via1_4
* cell instance $10137 r0 *1 82.935,20.51
X$10137 479 VIA_via2_5
* cell instance $10138 r0 *1 82.745,21.63
X$10138 479 VIA_via1_4
* cell instance $10139 r0 *1 86.545,20.51
X$10139 479 VIA_via1_4
* cell instance $10140 r0 *1 86.545,20.51
X$10140 479 VIA_via2_5
* cell instance $10141 r0 *1 94.335,20.65
X$10141 480 VIA_via2_5
* cell instance $10142 r0 *1 94.335,23.17
X$10142 480 VIA_via1_4
* cell instance $10143 r0 *1 94.335,18.83
X$10143 480 VIA_via1_4
* cell instance $10144 r0 *1 96.425,20.65
X$10144 480 VIA_via1_4
* cell instance $10145 r0 *1 96.425,20.65
X$10145 480 VIA_via2_5
* cell instance $10146 r0 *1 94.715,19.39
X$10146 481 VIA_via1_7
* cell instance $10147 r0 *1 94.715,19.39
X$10147 481 VIA_via2_5
* cell instance $10148 r0 *1 94.145,19.39
X$10148 481 VIA_via2_5
* cell instance $10149 r0 *1 94.145,20.37
X$10149 481 VIA_via1_4
* cell instance $10150 r0 *1 90.155,21.21
X$10150 482 VIA_via1_7
* cell instance $10151 r0 *1 90.155,20.37
X$10151 482 VIA_via2_5
* cell instance $10152 r0 *1 89.015,20.37
X$10152 482 VIA_via1_4
* cell instance $10153 r0 *1 89.015,20.37
X$10153 482 VIA_via2_5
* cell instance $10154 r0 *1 70.395,20.23
X$10154 483 VIA_via1_4
* cell instance $10155 r0 *1 70.395,20.23
X$10155 483 VIA_via2_5
* cell instance $10156 r0 *1 89.775,51.17
X$10156 483 VIA_via1_4
* cell instance $10157 r0 *1 89.775,49.63
X$10157 483 VIA_via1_4
* cell instance $10158 r0 *1 89.775,49.63
X$10158 483 VIA_via2_5
* cell instance $10159 r0 *1 89.695,49.63
X$10159 483 VIA_via3_2
* cell instance $10160 r0 *1 85.215,44.17
X$10160 483 VIA_via3_2
* cell instance $10161 r0 *1 85.215,20.23
X$10161 483 VIA_via3_2
* cell instance $10162 r0 *1 89.695,44.17
X$10162 483 VIA_via3_2
* cell instance $10163 r0 *1 84.265,20.37
X$10163 484 VIA_via1_4
* cell instance $10164 r0 *1 84.265,20.37
X$10164 484 VIA_via2_5
* cell instance $10165 r0 *1 83.315,20.37
X$10165 484 VIA_via1_4
* cell instance $10166 r0 *1 83.315,20.37
X$10166 484 VIA_via2_5
* cell instance $10167 r0 *1 9.975,20.37
X$10167 485 VIA_via1_4
* cell instance $10168 r0 *1 9.975,20.51
X$10168 485 VIA_via2_5
* cell instance $10169 r0 *1 6.365,20.51
X$10169 485 VIA_via1_4
* cell instance $10170 r0 *1 6.365,20.51
X$10170 485 VIA_via2_5
* cell instance $10171 r0 *1 79.705,17.99
X$10171 486 VIA_via1_7
* cell instance $10172 r0 *1 77.805,19.67
X$10172 486 VIA_via2_5
* cell instance $10173 r0 *1 79.705,19.67
X$10173 486 VIA_via2_5
* cell instance $10174 r0 *1 77.805,20.37
X$10174 486 VIA_via1_4
* cell instance $10175 r0 *1 79.135,19.81
X$10175 487 VIA_via1_7
* cell instance $10176 r0 *1 79.135,18.83
X$10176 487 VIA_via1_4
* cell instance $10177 r0 *1 13.965,19.39
X$10177 488 VIA_via1_7
* cell instance $10178 r0 *1 13.965,19.39
X$10178 488 VIA_via2_5
* cell instance $10179 r0 *1 13.395,19.39
X$10179 488 VIA_via2_5
* cell instance $10180 r0 *1 13.395,20.37
X$10180 488 VIA_via1_4
* cell instance $10181 r0 *1 77.045,19.95
X$10181 489 VIA_via2_5
* cell instance $10182 r0 *1 75.905,19.95
X$10182 489 VIA_via1_4
* cell instance $10183 r0 *1 75.905,19.95
X$10183 489 VIA_via2_5
* cell instance $10184 r0 *1 77.045,20.37
X$10184 489 VIA_via1_4
* cell instance $10185 r0 *1 10.355,19.81
X$10185 490 VIA_via1_7
* cell instance $10186 r0 *1 10.355,19.81
X$10186 490 VIA_via2_5
* cell instance $10187 r0 *1 16.245,19.81
X$10187 490 VIA_via2_5
* cell instance $10188 r0 *1 16.245,20.37
X$10188 490 VIA_via1_4
* cell instance $10189 r0 *1 76.855,20.37
X$10189 491 VIA_via1_4
* cell instance $10190 r0 *1 76.855,19.11
X$10190 491 VIA_via1_4
* cell instance $10191 r0 *1 16.055,20.37
X$10191 492 VIA_via1_4
* cell instance $10192 r0 *1 16.055,20.37
X$10192 492 VIA_via2_5
* cell instance $10193 r0 *1 17.385,20.37
X$10193 492 VIA_via1_4
* cell instance $10194 r0 *1 17.385,20.37
X$10194 492 VIA_via2_5
* cell instance $10195 r0 *1 20.235,20.37
X$10195 493 VIA_via1_4
* cell instance $10196 r0 *1 20.235,20.37
X$10196 493 VIA_via2_5
* cell instance $10197 r0 *1 21.185,20.37
X$10197 493 VIA_via1_4
* cell instance $10198 r0 *1 21.185,20.37
X$10198 493 VIA_via2_5
* cell instance $10199 r0 *1 68.875,19.39
X$10199 494 VIA_via1_7
* cell instance $10200 r0 *1 68.875,19.39
X$10200 494 VIA_via2_5
* cell instance $10201 r0 *1 66.975,19.39
X$10201 494 VIA_via2_5
* cell instance $10202 r0 *1 66.975,20.37
X$10202 494 VIA_via1_4
* cell instance $10203 r0 *1 29.355,19.39
X$10203 495 VIA_via1_7
* cell instance $10204 r0 *1 29.355,19.39
X$10204 495 VIA_via2_5
* cell instance $10205 r0 *1 26.885,19.39
X$10205 495 VIA_via2_5
* cell instance $10206 r0 *1 26.885,20.37
X$10206 495 VIA_via1_4
* cell instance $10207 r0 *1 65.835,20.37
X$10207 496 VIA_via1_4
* cell instance $10208 r0 *1 65.835,19.11
X$10208 496 VIA_via1_4
* cell instance $10209 r0 *1 30.495,20.37
X$10209 497 VIA_via1_4
* cell instance $10210 r0 *1 30.875,20.37
X$10210 497 VIA_via1_4
* cell instance $10211 r0 *1 63.935,21.21
X$10211 498 VIA_via1_7
* cell instance $10212 r0 *1 63.935,20.37
X$10212 498 VIA_via2_5
* cell instance $10213 r0 *1 60.705,20.37
X$10213 498 VIA_via1_4
* cell instance $10214 r0 *1 60.705,20.37
X$10214 498 VIA_via2_5
* cell instance $10215 r0 *1 55.575,22.61
X$10215 499 VIA_via1_7
* cell instance $10216 r0 *1 55.575,20.37
X$10216 499 VIA_via2_5
* cell instance $10217 r0 *1 54.625,20.37
X$10217 499 VIA_via1_4
* cell instance $10218 r0 *1 54.625,20.37
X$10218 499 VIA_via2_5
* cell instance $10219 r0 *1 45.315,20.37
X$10219 500 VIA_via1_4
* cell instance $10220 r0 *1 45.125,20.37
X$10220 500 VIA_via1_4
* cell instance $10221 r0 *1 42.845,20.37
X$10221 501 VIA_via1_4
* cell instance $10222 r0 *1 42.845,20.37
X$10222 501 VIA_via2_5
* cell instance $10223 r0 *1 44.365,21.35
X$10223 501 VIA_via1_4
* cell instance $10224 r0 *1 44.175,20.37
X$10224 501 VIA_via1_4
* cell instance $10225 r0 *1 44.175,20.37
X$10225 501 VIA_via2_5
* cell instance $10226 r0 *1 5.795,26.81
X$10226 502 VIA_via1_7
* cell instance $10227 r0 *1 5.795,26.81
X$10227 502 VIA_via2_5
* cell instance $10228 r0 *1 5.985,27.23
X$10228 502 VIA_via1_4
* cell instance $10229 r0 *1 5.795,32.97
X$10229 502 VIA_via2_5
* cell instance $10230 r0 *1 14.535,44.17
X$10230 502 VIA_via2_5
* cell instance $10231 r0 *1 7.315,43.75
X$10231 502 VIA_via2_5
* cell instance $10232 r0 *1 8.265,43.75
X$10232 502 VIA_via2_5
* cell instance $10233 r0 *1 18.145,23.31
X$10233 502 VIA_via2_5
* cell instance $10234 r0 *1 16.625,26.81
X$10234 502 VIA_via2_5
* cell instance $10235 r0 *1 4.465,21.63
X$10235 502 VIA_via1_4
* cell instance $10236 r0 *1 5.795,21.63
X$10236 502 VIA_via1_4
* cell instance $10237 r0 *1 8.265,42.77
X$10237 502 VIA_via1_4
* cell instance $10238 r0 *1 8.265,42.63
X$10238 502 VIA_via2_5
* cell instance $10239 r0 *1 8.215,42.63
X$10239 502 VIA_via3_2
* cell instance $10240 r0 *1 3.895,32.83
X$10240 502 VIA_via1_4
* cell instance $10241 r0 *1 3.895,32.97
X$10241 502 VIA_via2_5
* cell instance $10242 r0 *1 7.315,44.03
X$10242 502 VIA_via1_4
* cell instance $10243 r0 *1 16.625,23.17
X$10243 502 VIA_via1_4
* cell instance $10244 r0 *1 16.625,23.31
X$10244 502 VIA_via2_5
* cell instance $10245 r0 *1 18.145,21.63
X$10245 502 VIA_via1_4
* cell instance $10246 r0 *1 16.625,34.37
X$10246 502 VIA_via1_4
* cell instance $10247 r0 *1 15.675,44.03
X$10247 502 VIA_via1_4
* cell instance $10248 r0 *1 15.675,44.17
X$10248 502 VIA_via2_5
* cell instance $10249 r0 *1 14.535,45.57
X$10249 502 VIA_via1_4
* cell instance $10250 r0 *1 8.215,32.97
X$10250 502 VIA_via3_2
* cell instance $10251 r0 *1 12.445,21.07
X$10251 503 VIA_via2_5
* cell instance $10252 r0 *1 14.725,21.07
X$10252 503 VIA_via2_5
* cell instance $10253 r0 *1 15.485,24.43
X$10253 503 VIA_via2_5
* cell instance $10254 r0 *1 17.955,24.43
X$10254 503 VIA_via2_5
* cell instance $10255 r0 *1 19.475,24.43
X$10255 503 VIA_via2_5
* cell instance $10256 r0 *1 14.155,21.07
X$10256 503 VIA_via2_5
* cell instance $10257 r0 *1 10.735,24.43
X$10257 503 VIA_via1_4
* cell instance $10258 r0 *1 10.735,24.43
X$10258 503 VIA_via2_5
* cell instance $10259 r0 *1 12.445,17.57
X$10259 503 VIA_via1_4
* cell instance $10260 r0 *1 14.725,21.63
X$10260 503 VIA_via1_4
* cell instance $10261 r0 *1 17.005,24.43
X$10261 503 VIA_via1_4
* cell instance $10262 r0 *1 17.005,24.43
X$10262 503 VIA_via2_5
* cell instance $10263 r0 *1 15.485,22.05
X$10263 503 VIA_via1_4
* cell instance $10264 r0 *1 14.155,20.37
X$10264 503 VIA_via1_4
* cell instance $10265 r0 *1 19.475,23.17
X$10265 503 VIA_via1_4
* cell instance $10266 r0 *1 17.955,17.57
X$10266 503 VIA_via1_4
* cell instance $10267 r0 *1 17.575,23.17
X$10267 504 VIA_via2_5
* cell instance $10268 r0 *1 16.815,21.63
X$10268 504 VIA_via1_4
* cell instance $10269 r0 *1 17.575,21.63
X$10269 504 VIA_via1_4
* cell instance $10270 r0 *1 20.995,23.17
X$10270 504 VIA_via1_4
* cell instance $10271 r0 *1 20.995,23.17
X$10271 504 VIA_via2_5
* cell instance $10272 r0 *1 24.035,21.49
X$10272 505 VIA_via1_4
* cell instance $10273 r0 *1 24.035,21.49
X$10273 505 VIA_via2_5
* cell instance $10274 r0 *1 19.855,21.63
X$10274 505 VIA_via1_4
* cell instance $10275 r0 *1 19.855,21.49
X$10275 505 VIA_via2_5
* cell instance $10276 r0 *1 24.415,21.63
X$10276 505 VIA_via1_4
* cell instance $10277 r0 *1 24.415,21.49
X$10277 505 VIA_via2_5
* cell instance $10278 r0 *1 26.695,22.61
X$10278 506 VIA_via1_7
* cell instance $10279 r0 *1 26.505,21.63
X$10279 506 VIA_via1_4
* cell instance $10280 r0 *1 25.745,22.05
X$10280 507 VIA_via2_5
* cell instance $10281 r0 *1 29.545,22.05
X$10281 507 VIA_via2_5
* cell instance $10282 r0 *1 29.545,20.37
X$10282 507 VIA_via1_4
* cell instance $10283 r0 *1 25.745,23.17
X$10283 507 VIA_via1_4
* cell instance $10284 r0 *1 28.785,22.05
X$10284 507 VIA_via1_4
* cell instance $10285 r0 *1 28.785,22.05
X$10285 507 VIA_via2_5
* cell instance $10286 r0 *1 30.685,23.17
X$10286 508 VIA_via2_5
* cell instance $10287 r0 *1 28.785,23.17
X$10287 508 VIA_via1_4
* cell instance $10288 r0 *1 28.785,23.17
X$10288 508 VIA_via2_5
* cell instance $10289 r0 *1 30.875,21.77
X$10289 508 VIA_via1_4
* cell instance $10290 r0 *1 32.015,24.15
X$10290 509 VIA_via2_5
* cell instance $10291 r0 *1 34.865,24.15
X$10291 509 VIA_via1_4
* cell instance $10292 r0 *1 34.865,24.15
X$10292 509 VIA_via2_5
* cell instance $10293 r0 *1 32.015,23.17
X$10293 509 VIA_via1_4
* cell instance $10294 r0 *1 31.825,21.63
X$10294 509 VIA_via1_4
* cell instance $10295 r0 *1 33.345,29.61
X$10295 510 VIA_via1_7
* cell instance $10296 r0 *1 33.345,30.59
X$10296 510 VIA_via1_7
* cell instance $10297 r0 *1 32.395,28.91
X$10297 510 VIA_via2_5
* cell instance $10298 r0 *1 33.345,28.91
X$10298 510 VIA_via2_5
* cell instance $10299 r0 *1 32.585,21.63
X$10299 510 VIA_via2_5
* cell instance $10300 r0 *1 33.345,38.15
X$10300 510 VIA_via2_5
* cell instance $10301 r0 *1 32.015,38.15
X$10301 510 VIA_via2_5
* cell instance $10302 r0 *1 32.585,38.15
X$10302 510 VIA_via2_5
* cell instance $10303 r0 *1 32.585,23.17
X$10303 510 VIA_via1_4
* cell instance $10304 r0 *1 35.055,21.63
X$10304 510 VIA_via1_4
* cell instance $10305 r0 *1 35.055,21.63
X$10305 510 VIA_via2_5
* cell instance $10306 r0 *1 30.495,21.63
X$10306 510 VIA_via1_4
* cell instance $10307 r0 *1 30.495,21.63
X$10307 510 VIA_via2_5
* cell instance $10308 r0 *1 33.535,21.63
X$10308 510 VIA_via1_4
* cell instance $10309 r0 *1 33.535,21.63
X$10309 510 VIA_via2_5
* cell instance $10310 r0 *1 31.255,28.77
X$10310 510 VIA_via1_4
* cell instance $10311 r0 *1 31.255,28.91
X$10311 510 VIA_via2_5
* cell instance $10312 r0 *1 36.385,38.43
X$10312 510 VIA_via1_4
* cell instance $10313 r0 *1 36.385,38.43
X$10313 510 VIA_via2_5
* cell instance $10314 r0 *1 33.345,38.43
X$10314 510 VIA_via1_4
* cell instance $10315 r0 *1 32.015,38.43
X$10315 510 VIA_via1_4
* cell instance $10316 r0 *1 35.055,38.43
X$10316 510 VIA_via1_4
* cell instance $10317 r0 *1 35.055,38.29
X$10317 510 VIA_via2_5
* cell instance $10318 r0 *1 32.585,34.37
X$10318 510 VIA_via1_4
* cell instance $10319 r0 *1 33.915,21.21
X$10319 511 VIA_via1_7
* cell instance $10320 r0 *1 33.535,20.37
X$10320 511 VIA_via1_4
* cell instance $10321 r0 *1 45.885,22.75
X$10321 512 VIA_via1_4
* cell instance $10322 r0 *1 45.315,21.63
X$10322 512 VIA_via1_4
* cell instance $10323 r0 *1 44.745,20.37
X$10323 512 VIA_via1_4
* cell instance $10324 r0 *1 50.825,23.17
X$10324 513 VIA_via2_5
* cell instance $10325 r0 *1 51.205,21.63
X$10325 513 VIA_via1_4
* cell instance $10326 r0 *1 50.825,22.05
X$10326 513 VIA_via1_4
* cell instance $10327 r0 *1 50.445,23.17
X$10327 513 VIA_via1_4
* cell instance $10328 r0 *1 50.445,23.17
X$10328 513 VIA_via2_5
* cell instance $10329 r0 *1 54.625,23.45
X$10329 514 VIA_via2_5
* cell instance $10330 r0 *1 56.715,23.45
X$10330 514 VIA_via2_5
* cell instance $10331 r0 *1 56.715,23.17
X$10331 514 VIA_via1_4
* cell instance $10332 r0 *1 56.905,20.65
X$10332 514 VIA_via1_4
* cell instance $10333 r0 *1 54.625,23.17
X$10333 514 VIA_via1_4
* cell instance $10334 r0 *1 69.445,52.01
X$10334 515 VIA_via1_7
* cell instance $10335 r0 *1 69.445,52.01
X$10335 515 VIA_via2_5
* cell instance $10336 r0 *1 58.045,21.35
X$10336 515 VIA_via2_5
* cell instance $10337 r0 *1 52.535,21.35
X$10337 515 VIA_via2_5
* cell instance $10338 r0 *1 58.045,22.89
X$10338 515 VIA_via2_5
* cell instance $10339 r0 *1 62.035,52.57
X$10339 515 VIA_via2_5
* cell instance $10340 r0 *1 62.035,51.87
X$10340 515 VIA_via2_5
* cell instance $10341 r0 *1 52.915,52.57
X$10341 515 VIA_via2_5
* cell instance $10342 r0 *1 67.925,49.35
X$10342 515 VIA_via2_5
* cell instance $10343 r0 *1 67.925,52.01
X$10343 515 VIA_via2_5
* cell instance $10344 r0 *1 65.455,49.35
X$10344 515 VIA_via2_5
* cell instance $10345 r0 *1 65.645,24.57
X$10345 515 VIA_via2_5
* cell instance $10346 r0 *1 62.225,23.87
X$10346 515 VIA_via2_5
* cell instance $10347 r0 *1 62.795,22.89
X$10347 515 VIA_via2_5
* cell instance $10348 r0 *1 62.795,23.87
X$10348 515 VIA_via2_5
* cell instance $10349 r0 *1 58.045,21.63
X$10349 515 VIA_via1_4
* cell instance $10350 r0 *1 52.535,21.63
X$10350 515 VIA_via1_4
* cell instance $10351 r0 *1 62.225,24.43
X$10351 515 VIA_via1_4
* cell instance $10352 r0 *1 62.225,24.57
X$10352 515 VIA_via2_5
* cell instance $10353 r0 *1 68.115,49.63
X$10353 515 VIA_via1_4
* cell instance $10354 r0 *1 52.915,53.97
X$10354 515 VIA_via1_4
* cell instance $10355 r0 *1 58.045,20.79
X$10355 516 VIA_via1_7
* cell instance $10356 r0 *1 58.425,21.63
X$10356 516 VIA_via1_4
* cell instance $10357 r0 *1 58.615,17.99
X$10357 517 VIA_via1_7
* cell instance $10358 r0 *1 58.995,21.63
X$10358 517 VIA_via1_4
* cell instance $10359 r0 *1 58.995,20.79
X$10359 518 VIA_via1_7
* cell instance $10360 r0 *1 59.185,21.63
X$10360 518 VIA_via1_4
* cell instance $10361 r0 *1 63.175,23.17
X$10361 519 VIA_via1_4
* cell instance $10362 r0 *1 62.985,21.63
X$10362 519 VIA_via1_4
* cell instance $10363 r0 *1 62.985,20.65
X$10363 519 VIA_via1_4
* cell instance $10364 r0 *1 66.595,21.77
X$10364 520 VIA_via1_7
* cell instance $10365 r0 *1 66.595,21.77
X$10365 520 VIA_via2_5
* cell instance $10366 r0 *1 72.485,60.97
X$10366 520 VIA_via1_7
* cell instance $10367 r0 *1 62.795,21.77
X$10367 520 VIA_via1_7
* cell instance $10368 r0 *1 62.795,21.77
X$10368 520 VIA_via2_5
* cell instance $10369 r0 *1 73.625,30.17
X$10369 520 VIA_via1_7
* cell instance $10370 r0 *1 73.625,30.17
X$10370 520 VIA_via2_5
* cell instance $10371 r0 *1 75.145,48.23
X$10371 520 VIA_via1_7
* cell instance $10372 r0 *1 75.145,48.09
X$10372 520 VIA_via2_5
* cell instance $10373 r0 *1 74.385,21.77
X$10373 520 VIA_via1_7
* cell instance $10374 r0 *1 74.385,21.77
X$10374 520 VIA_via2_5
* cell instance $10375 r0 *1 74.295,21.77
X$10375 520 VIA_via3_2
* cell instance $10376 r0 *1 72.485,65.17
X$10376 520 VIA_via2_5
* cell instance $10377 r0 *1 63.555,52.57
X$10377 520 VIA_via2_5
* cell instance $10378 r0 *1 63.175,53.83
X$10378 520 VIA_via2_5
* cell instance $10379 r0 *1 63.555,53.83
X$10379 520 VIA_via2_5
* cell instance $10380 r0 *1 63.555,52.99
X$10380 520 VIA_via2_5
* cell instance $10381 r0 *1 65.455,52.99
X$10381 520 VIA_via2_5
* cell instance $10382 r0 *1 73.815,65.17
X$10382 520 VIA_via2_5
* cell instance $10383 r0 *1 66.215,30.31
X$10383 520 VIA_via2_5
* cell instance $10384 r0 *1 65.835,30.31
X$10384 520 VIA_via2_5
* cell instance $10385 r0 *1 66.785,48.09
X$10385 520 VIA_via2_5
* cell instance $10386 r0 *1 73.625,26.11
X$10386 520 VIA_via2_5
* cell instance $10387 r0 *1 65.835,21.77
X$10387 520 VIA_via2_5
* cell instance $10388 r0 *1 65.645,48.09
X$10388 520 VIA_via2_5
* cell instance $10389 r0 *1 63.365,65.17
X$10389 520 VIA_via1_4
* cell instance $10390 r0 *1 63.365,65.17
X$10390 520 VIA_via2_5
* cell instance $10391 r0 *1 74.575,25.97
X$10391 520 VIA_via1_4
* cell instance $10392 r0 *1 74.575,26.11
X$10392 520 VIA_via2_5
* cell instance $10393 r0 *1 66.405,38.43
X$10393 520 VIA_via1_4
* cell instance $10394 r0 *1 73.815,66.43
X$10394 520 VIA_via1_4
* cell instance $10395 r0 *1 62.795,52.57
X$10395 520 VIA_via1_4
* cell instance $10396 r0 *1 62.795,52.57
X$10396 520 VIA_via2_5
* cell instance $10397 r0 *1 74.295,26.11
X$10397 520 VIA_via3_2
* cell instance $10398 r0 *1 70.015,21.21
X$10398 521 VIA_via1_7
* cell instance $10399 r0 *1 70.205,20.37
X$10399 521 VIA_via1_4
* cell instance $10400 r0 *1 83.315,52.15
X$10400 522 VIA_via2_5
* cell instance $10401 r0 *1 71.725,21.35
X$10401 522 VIA_via2_5
* cell instance $10402 r0 *1 71.535,27.23
X$10402 522 VIA_via2_5
* cell instance $10403 r0 *1 59.185,21.35
X$10403 522 VIA_via1_4
* cell instance $10404 r0 *1 59.185,21.35
X$10404 522 VIA_via2_5
* cell instance $10405 r0 *1 79.895,52.43
X$10405 522 VIA_via1_4
* cell instance $10406 r0 *1 79.895,52.43
X$10406 522 VIA_via3_2
* cell instance $10407 r0 *1 79.895,52.43
X$10407 522 VIA_via2_5
* cell instance $10408 r0 *1 83.315,52.43
X$10408 522 VIA_via1_4
* cell instance $10409 r0 *1 79.895,27.23
X$10409 522 VIA_via3_2
* cell instance $10410 r0 *1 77.045,22.61
X$10410 523 VIA_via1_7
* cell instance $10411 r0 *1 77.235,21.63
X$10411 523 VIA_via1_4
* cell instance $10412 r0 *1 89.775,23.03
X$10412 524 VIA_via2_5
* cell instance $10413 r0 *1 85.405,23.03
X$10413 524 VIA_via2_5
* cell instance $10414 r0 *1 76.665,21.77
X$10414 524 VIA_via2_5
* cell instance $10415 r0 *1 78.185,21.77
X$10415 524 VIA_via2_5
* cell instance $10416 r0 *1 76.665,24.15
X$10416 524 VIA_via2_5
* cell instance $10417 r0 *1 82.175,21.91
X$10417 524 VIA_via2_5
* cell instance $10418 r0 *1 75.905,24.15
X$10418 524 VIA_via2_5
* cell instance $10419 r0 *1 83.885,21.91
X$10419 524 VIA_via2_5
* cell instance $10420 r0 *1 73.055,24.15
X$10420 524 VIA_via2_5
* cell instance $10421 r0 *1 75.905,25.13
X$10421 524 VIA_via2_5
* cell instance $10422 r0 *1 75.335,25.13
X$10422 524 VIA_via2_5
* cell instance $10423 r0 *1 82.175,23.17
X$10423 524 VIA_via1_4
* cell instance $10424 r0 *1 85.405,22.05
X$10424 524 VIA_via1_4
* cell instance $10425 r0 *1 85.405,21.91
X$10425 524 VIA_via2_5
* cell instance $10426 r0 *1 87.495,25.97
X$10426 524 VIA_via1_4
* cell instance $10427 r0 *1 84.265,25.97
X$10427 524 VIA_via1_4
* cell instance $10428 r0 *1 75.335,25.97
X$10428 524 VIA_via1_4
* cell instance $10429 r0 *1 75.905,24.43
X$10429 524 VIA_via1_4
* cell instance $10430 r0 *1 76.665,23.17
X$10430 524 VIA_via1_4
* cell instance $10431 r0 *1 78.185,20.37
X$10431 524 VIA_via1_4
* cell instance $10432 r0 *1 73.055,24.43
X$10432 524 VIA_via1_4
* cell instance $10433 r0 *1 87.305,23.17
X$10433 524 VIA_via1_4
* cell instance $10434 r0 *1 87.305,23.03
X$10434 524 VIA_via2_5
* cell instance $10435 r0 *1 89.775,21.63
X$10435 524 VIA_via1_4
* cell instance $10436 r0 *1 82.365,23.17
X$10436 525 VIA_via2_5
* cell instance $10437 r0 *1 82.175,21.63
X$10437 525 VIA_via1_4
* cell instance $10438 r0 *1 82.745,23.17
X$10438 525 VIA_via1_4
* cell instance $10439 r0 *1 82.745,23.17
X$10439 525 VIA_via2_5
* cell instance $10440 r0 *1 86.355,23.17
X$10440 525 VIA_via1_4
* cell instance $10441 r0 *1 86.355,23.17
X$10441 525 VIA_via2_5
* cell instance $10442 r0 *1 4.845,21.21
X$10442 526 VIA_via1_7
* cell instance $10443 r0 *1 4.845,21.21
X$10443 526 VIA_via2_5
* cell instance $10444 r0 *1 2.755,21.21
X$10444 526 VIA_via2_5
* cell instance $10445 r0 *1 2.755,20.37
X$10445 526 VIA_via1_4
* cell instance $10446 r0 *1 96.045,22.61
X$10446 527 VIA_via1_7
* cell instance $10447 r0 *1 96.045,21.63
X$10447 527 VIA_via2_5
* cell instance $10448 r0 *1 93.955,21.63
X$10448 527 VIA_via1_4
* cell instance $10449 r0 *1 93.955,21.63
X$10449 527 VIA_via2_5
* cell instance $10450 r0 *1 7.125,22.61
X$10450 528 VIA_via1_7
* cell instance $10451 r0 *1 7.125,21.63
X$10451 528 VIA_via2_5
* cell instance $10452 r0 *1 10.925,21.63
X$10452 528 VIA_via1_4
* cell instance $10453 r0 *1 10.925,21.63
X$10453 528 VIA_via2_5
* cell instance $10454 r0 *1 89.965,21.63
X$10454 529 VIA_via2_5
* cell instance $10455 r0 *1 91.295,21.63
X$10455 529 VIA_via2_5
* cell instance $10456 r0 *1 89.205,21.63
X$10456 529 VIA_via1_4
* cell instance $10457 r0 *1 89.205,21.63
X$10457 529 VIA_via2_5
* cell instance $10458 r0 *1 89.965,23.17
X$10458 529 VIA_via1_4
* cell instance $10459 r0 *1 91.295,20.65
X$10459 529 VIA_via1_4
* cell instance $10460 r0 *1 17.195,21.21
X$10460 530 VIA_via1_7
* cell instance $10461 r0 *1 17.195,20.37
X$10461 530 VIA_via1_4
* cell instance $10462 r0 *1 18.905,45.57
X$10462 531 VIA_via2_5
* cell instance $10463 r0 *1 16.435,21.07
X$10463 531 VIA_via2_5
* cell instance $10464 r0 *1 16.435,20.51
X$10464 531 VIA_via1_4
* cell instance $10465 r0 *1 18.905,46.83
X$10465 531 VIA_via1_4
* cell instance $10466 r0 *1 19.665,45.57
X$10466 531 VIA_via1_4
* cell instance $10467 r0 *1 19.695,45.57
X$10467 531 VIA_via3_2
* cell instance $10468 r0 *1 19.665,45.57
X$10468 531 VIA_via2_5
* cell instance $10469 r0 *1 19.695,21.07
X$10469 531 VIA_via3_2
* cell instance $10470 r0 *1 80.845,20.79
X$10470 532 VIA_via1_7
* cell instance $10471 r0 *1 80.845,21.63
X$10471 532 VIA_via2_5
* cell instance $10472 r0 *1 79.705,21.63
X$10472 532 VIA_via1_4
* cell instance $10473 r0 *1 79.705,21.63
X$10473 532 VIA_via2_5
* cell instance $10474 r0 *1 20.805,21.63
X$10474 533 VIA_via1_4
* cell instance $10475 r0 *1 20.805,21.63
X$10475 533 VIA_via2_5
* cell instance $10476 r0 *1 21.755,21.63
X$10476 533 VIA_via1_4
* cell instance $10477 r0 *1 21.755,21.63
X$10477 533 VIA_via2_5
* cell instance $10478 r0 *1 87.685,49.35
X$10478 534 VIA_via2_5
* cell instance $10479 r0 *1 87.685,52.43
X$10479 534 VIA_via2_5
* cell instance $10480 r0 *1 77.615,20.65
X$10480 534 VIA_via2_5
* cell instance $10481 r0 *1 77.805,20.65
X$10481 534 VIA_via1_4
* cell instance $10482 r0 *1 90.725,52.5
X$10482 534 VIA_via1_4
* cell instance $10483 r0 *1 90.725,52.57
X$10483 534 VIA_via2_5
* cell instance $10484 r0 *1 89.775,52.43
X$10484 534 VIA_via1_4
* cell instance $10485 r0 *1 89.775,52.43
X$10485 534 VIA_via2_5
* cell instance $10486 r0 *1 77.375,20.65
X$10486 534 VIA_via3_2
* cell instance $10487 r0 *1 77.375,49.35
X$10487 534 VIA_via3_2
* cell instance $10488 r0 *1 75.525,21.21
X$10488 535 VIA_via1_7
* cell instance $10489 r0 *1 75.525,21.21
X$10489 535 VIA_via2_5
* cell instance $10490 r0 *1 72.105,21.21
X$10490 535 VIA_via2_5
* cell instance $10491 r0 *1 72.105,20.37
X$10491 535 VIA_via1_4
* cell instance $10492 r0 *1 32.205,21.21
X$10492 536 VIA_via1_7
* cell instance $10493 r0 *1 32.205,20.37
X$10493 536 VIA_via1_4
* cell instance $10494 r0 *1 73.435,22.61
X$10494 537 VIA_via1_7
* cell instance $10495 r0 *1 73.435,21.63
X$10495 537 VIA_via2_5
* cell instance $10496 r0 *1 71.535,21.63
X$10496 537 VIA_via1_4
* cell instance $10497 r0 *1 71.535,21.63
X$10497 537 VIA_via2_5
* cell instance $10498 r0 *1 68.875,22.75
X$10498 538 VIA_via1_4
* cell instance $10499 r0 *1 69.255,21.63
X$10499 538 VIA_via1_4
* cell instance $10500 r0 *1 69.255,21.63
X$10500 538 VIA_via2_5
* cell instance $10501 r0 *1 66.785,21.63
X$10501 538 VIA_via1_4
* cell instance $10502 r0 *1 66.785,21.63
X$10502 538 VIA_via2_5
* cell instance $10503 r0 *1 69.635,21.63
X$10503 539 VIA_via1_4
* cell instance $10504 r0 *1 69.825,21.63
X$10504 539 VIA_via1_4
* cell instance $10505 r0 *1 36.765,21.49
X$10505 540 VIA_via2_5
* cell instance $10506 r0 *1 36.765,22.75
X$10506 540 VIA_via2_5
* cell instance $10507 r0 *1 34.485,21.63
X$10507 540 VIA_via1_4
* cell instance $10508 r0 *1 34.485,21.49
X$10508 540 VIA_via2_5
* cell instance $10509 r0 *1 37.335,22.75
X$10509 540 VIA_via1_4
* cell instance $10510 r0 *1 37.335,22.75
X$10510 540 VIA_via2_5
* cell instance $10511 r0 *1 36.765,20.37
X$10511 540 VIA_via1_4
* cell instance $10512 r0 *1 47.975,60.97
X$10512 541 VIA_via1_7
* cell instance $10513 r0 *1 47.975,60.97
X$10513 541 VIA_via2_5
* cell instance $10514 r0 *1 68.495,21.77
X$10514 541 VIA_via1_7
* cell instance $10515 r0 *1 68.495,21.77
X$10515 541 VIA_via2_5
* cell instance $10516 r0 *1 49.495,61.81
X$10516 541 VIA_via2_5
* cell instance $10517 r0 *1 50.825,61.81
X$10517 541 VIA_via2_5
* cell instance $10518 r0 *1 73.625,23.45
X$10518 541 VIA_via2_5
* cell instance $10519 r0 *1 49.495,60.97
X$10519 541 VIA_via2_5
* cell instance $10520 r0 *1 74.195,67.13
X$10520 541 VIA_via2_5
* cell instance $10521 r0 *1 65.645,40.25
X$10521 541 VIA_via2_5
* cell instance $10522 r0 *1 66.025,40.25
X$10522 541 VIA_via2_5
* cell instance $10523 r0 *1 65.645,43.05
X$10523 541 VIA_via2_5
* cell instance $10524 r0 *1 51.015,66.43
X$10524 541 VIA_via1_4
* cell instance $10525 r0 *1 51.015,66.29
X$10525 541 VIA_via2_5
* cell instance $10526 r0 *1 63.175,66.43
X$10526 541 VIA_via1_4
* cell instance $10527 r0 *1 63.175,66.29
X$10527 541 VIA_via2_5
* cell instance $10528 r0 *1 73.815,48.37
X$10528 541 VIA_via1_4
* cell instance $10529 r0 *1 73.815,48.37
X$10529 541 VIA_via2_5
* cell instance $10530 r0 *1 49.115,51.45
X$10530 541 VIA_via1_4
* cell instance $10531 r0 *1 49.115,51.45
X$10531 541 VIA_via2_5
* cell instance $10532 r0 *1 66.025,39.97
X$10532 541 VIA_via1_4
* cell instance $10533 r0 *1 73.625,23.17
X$10533 541 VIA_via1_4
* cell instance $10534 r0 *1 73.625,24.43
X$10534 541 VIA_via1_4
* cell instance $10535 r0 *1 74.195,69.23
X$10535 541 VIA_via1_4
* cell instance $10536 r0 *1 73.815,60.83
X$10536 541 VIA_via1_4
* cell instance $10537 r0 *1 73.815,60.83
X$10537 541 VIA_via2_5
* cell instance $10538 r0 *1 73.735,67.13
X$10538 541 VIA_via3_2
* cell instance $10539 r0 *1 68.135,40.25
X$10539 541 VIA_via3_2
* cell instance $10540 r0 *1 73.735,66.29
X$10540 541 VIA_via3_2
* cell instance $10541 r0 *1 74.015,60.83
X$10541 541 VIA_via3_2
* cell instance $10542 r0 *1 68.135,21.77
X$10542 541 VIA_via3_2
* cell instance $10543 r0 *1 68.135,23.45
X$10543 541 VIA_via3_2
* cell instance $10544 r0 *1 74.015,48.37
X$10544 541 VIA_via3_2
* cell instance $10545 r0 *1 49.375,51.45
X$10545 541 VIA_via3_2
* cell instance $10546 r0 *1 49.375,43.19
X$10546 541 VIA_via3_2
* cell instance $10547 r0 *1 39.995,22.61
X$10547 542 VIA_via1_7
* cell instance $10548 r0 *1 39.995,21.63
X$10548 542 VIA_via2_5
* cell instance $10549 r0 *1 38.665,21.63
X$10549 542 VIA_via1_4
* cell instance $10550 r0 *1 38.665,21.63
X$10550 542 VIA_via2_5
* cell instance $10551 r0 *1 66.785,25.97
X$10551 543 VIA_via2_5
* cell instance $10552 r0 *1 70.205,25.27
X$10552 543 VIA_via2_5
* cell instance $10553 r0 *1 67.355,25.27
X$10553 543 VIA_via2_5
* cell instance $10554 r0 *1 63.745,25.97
X$10554 543 VIA_via2_5
* cell instance $10555 r0 *1 63.745,27.23
X$10555 543 VIA_via2_5
* cell instance $10556 r0 *1 62.225,27.23
X$10556 543 VIA_via2_5
* cell instance $10557 r0 *1 61.465,21.63
X$10557 543 VIA_via2_5
* cell instance $10558 r0 *1 63.745,21.63
X$10558 543 VIA_via2_5
* cell instance $10559 r0 *1 70.205,24.43
X$10559 543 VIA_via1_4
* cell instance $10560 r0 *1 64.885,24.43
X$10560 543 VIA_via1_4
* cell instance $10561 r0 *1 66.975,25.97
X$10561 543 VIA_via1_4
* cell instance $10562 r0 *1 66.975,25.97
X$10562 543 VIA_via2_5
* cell instance $10563 r0 *1 67.355,25.55
X$10563 543 VIA_via1_4
* cell instance $10564 r0 *1 64.885,25.97
X$10564 543 VIA_via1_4
* cell instance $10565 r0 *1 64.885,25.97
X$10565 543 VIA_via2_5
* cell instance $10566 r0 *1 66.785,28.77
X$10566 543 VIA_via1_4
* cell instance $10567 r0 *1 61.085,21.63
X$10567 543 VIA_via1_4
* cell instance $10568 r0 *1 61.085,21.63
X$10568 543 VIA_via2_5
* cell instance $10569 r0 *1 67.355,23.17
X$10569 543 VIA_via1_4
* cell instance $10570 r0 *1 61.465,20.37
X$10570 543 VIA_via1_4
* cell instance $10571 r0 *1 62.035,28.77
X$10571 543 VIA_via1_4
* cell instance $10572 r0 *1 43.795,20.79
X$10572 544 VIA_via1_7
* cell instance $10573 r0 *1 43.795,20.79
X$10573 544 VIA_via2_5
* cell instance $10574 r0 *1 42.085,20.79
X$10574 544 VIA_via2_5
* cell instance $10575 r0 *1 42.085,21.63
X$10575 544 VIA_via1_4
* cell instance $10576 r0 *1 51.395,22.61
X$10576 545 VIA_via1_7
* cell instance $10577 r0 *1 51.395,21.63
X$10577 545 VIA_via2_5
* cell instance $10578 r0 *1 48.545,21.63
X$10578 545 VIA_via1_4
* cell instance $10579 r0 *1 48.545,21.63
X$10579 545 VIA_via2_5
* cell instance $10580 r0 *1 56.715,21.63
X$10580 546 VIA_via1_4
* cell instance $10581 r0 *1 56.715,21.77
X$10581 546 VIA_via2_5
* cell instance $10582 r0 *1 52.155,21.77
X$10582 546 VIA_via1_4
* cell instance $10583 r0 *1 52.155,21.77
X$10583 546 VIA_via2_5
* cell instance $10584 r0 *1 11.305,22.19
X$10584 547 VIA_via1_7
* cell instance $10585 r0 *1 11.685,23.31
X$10585 547 VIA_via2_5
* cell instance $10586 r0 *1 13.015,23.17
X$10586 547 VIA_via1_4
* cell instance $10587 r0 *1 13.015,23.31
X$10587 547 VIA_via2_5
* cell instance $10588 r0 *1 12.825,90.93
X$10588 548 VIA_via2_5
* cell instance $10589 r0 *1 11.115,29.33
X$10589 548 VIA_via2_5
* cell instance $10590 r0 *1 55.765,86.03
X$10590 548 VIA_via1_4
* cell instance $10591 r0 *1 55.765,86.03
X$10591 548 VIA_via2_5
* cell instance $10592 r0 *1 51.205,91.63
X$10592 548 VIA_via1_4
* cell instance $10593 r0 *1 12.825,90.37
X$10593 548 VIA_via1_4
* cell instance $10594 r0 *1 41.135,90.37
X$10594 548 VIA_via1_4
* cell instance $10595 r0 *1 33.155,88.83
X$10595 548 VIA_via1_4
* cell instance $10596 r0 *1 33.155,88.83
X$10596 548 VIA_via2_5
* cell instance $10597 r0 *1 33.135,88.83
X$10597 548 VIA_via3_2
* cell instance $10598 r0 *1 56.905,24.15
X$10598 548 VIA_via1_4
* cell instance $10599 r0 *1 12.255,55.23
X$10599 548 VIA_via1_4
* cell instance $10600 r0 *1 12.255,55.37
X$10600 548 VIA_via2_5
* cell instance $10601 r0 *1 12.135,55.37
X$10601 548 VIA_via3_2
* cell instance $10602 r0 *1 11.875,65.17
X$10602 548 VIA_via1_4
* cell instance $10603 r0 *1 11.875,65.17
X$10603 548 VIA_via2_5
* cell instance $10604 r0 *1 12.635,74.83
X$10604 548 VIA_via1_4
* cell instance $10605 r0 *1 12.635,74.83
X$10605 548 VIA_via2_5
* cell instance $10606 r0 *1 13.395,23.17
X$10606 548 VIA_via1_4
* cell instance $10607 r0 *1 13.395,23.17
X$10607 548 VIA_via2_5
* cell instance $10608 r0 *1 13.255,23.17
X$10608 548 VIA_via3_2
* cell instance $10609 r0 *1 13.255,23.31
X$10609 548 VIA_via4_0
* cell instance $10610 r0 *1 12.975,90.51
X$10610 548 VIA_via4_0
* cell instance $10611 r0 *1 14.375,90.51
X$10611 548 VIA_via4_0
* cell instance $10612 r0 *1 14.375,65.31
X$10612 548 VIA_via4_0
* cell instance $10613 r0 *1 31.735,90.51
X$10613 548 VIA_via4_0
* cell instance $10614 r0 *1 55.535,91.35
X$10614 548 VIA_via4_0
* cell instance $10615 r0 *1 12.135,65.17
X$10615 548 VIA_via3_2
* cell instance $10616 r0 *1 12.135,65.31
X$10616 548 VIA_via4_0
* cell instance $10617 r0 *1 20.255,90.51
X$10617 548 VIA_via3_2
* cell instance $10618 r0 *1 20.235,90.51
X$10618 548 VIA_via2_5
* cell instance $10619 r0 *1 20.255,90.51
X$10619 548 VIA_via4_0
* cell instance $10620 r0 *1 20.235,90.37
X$10620 548 VIA_via1_4
* cell instance $10621 r0 *1 55.535,86.03
X$10621 548 VIA_via3_2
* cell instance $10622 r0 *1 12.975,90.93
X$10622 548 VIA_via3_2
* cell instance $10623 r0 *1 56.935,23.31
X$10623 548 VIA_via3_2
* cell instance $10624 r0 *1 56.905,23.31
X$10624 548 VIA_via2_5
* cell instance $10625 r0 *1 56.935,23.31
X$10625 548 VIA_via4_0
* cell instance $10626 r0 *1 14.375,74.83
X$10626 548 VIA_via3_2
* cell instance $10627 r0 *1 51.335,91.35
X$10627 548 VIA_via3_2
* cell instance $10628 r0 *1 51.205,91.35
X$10628 548 VIA_via2_5
* cell instance $10629 r0 *1 51.335,91.35
X$10629 548 VIA_via4_0
* cell instance $10630 r0 *1 41.255,90.79
X$10630 548 VIA_via3_2
* cell instance $10631 r0 *1 41.135,90.79
X$10631 548 VIA_via2_5
* cell instance $10632 r0 *1 41.255,90.79
X$10632 548 VIA_via4_0
* cell instance $10633 r0 *1 33.135,90.79
X$10633 548 VIA_via3_2
* cell instance $10634 r0 *1 31.735,90.79
X$10634 548 VIA_via3_2
* cell instance $10635 r0 *1 13.255,29.33
X$10635 548 VIA_via3_2
* cell instance $10636 r0 *1 16.055,24.15
X$10636 549 VIA_via2_5
* cell instance $10637 r0 *1 16.245,21.63
X$10637 549 VIA_via1_4
* cell instance $10638 r0 *1 18.525,24.15
X$10638 549 VIA_via1_4
* cell instance $10639 r0 *1 18.525,24.15
X$10639 549 VIA_via2_5
* cell instance $10640 r0 *1 16.055,23.17
X$10640 549 VIA_via1_4
* cell instance $10641 r0 *1 18.525,22.19
X$10641 550 VIA_via1_7
* cell instance $10642 r0 *1 18.715,23.17
X$10642 550 VIA_via1_4
* cell instance $10643 r0 *1 31.255,22.19
X$10643 551 VIA_via2_5
* cell instance $10644 r0 *1 29.925,22.61
X$10644 551 VIA_via2_5
* cell instance $10645 r0 *1 29.925,21.63
X$10645 551 VIA_via1_4
* cell instance $10646 r0 *1 31.065,22.75
X$10646 551 VIA_via1_4
* cell instance $10647 r0 *1 31.065,22.61
X$10647 551 VIA_via2_5
* cell instance $10648 r0 *1 31.255,21.63
X$10648 551 VIA_via1_4
* cell instance $10649 r0 *1 35.435,22.19
X$10649 552 VIA_via1_7
* cell instance $10650 r0 *1 35.055,23.17
X$10650 552 VIA_via1_4
* cell instance $10651 r0 *1 38.665,22.61
X$10651 553 VIA_via1_7
* cell instance $10652 r0 *1 38.285,20.37
X$10652 553 VIA_via1_4
* cell instance $10653 r0 *1 37.715,23.17
X$10653 554 VIA_via1_4
* cell instance $10654 r0 *1 37.715,23.31
X$10654 554 VIA_via2_5
* cell instance $10655 r0 *1 40.565,20.65
X$10655 554 VIA_via1_4
* cell instance $10656 r0 *1 40.375,23.17
X$10656 554 VIA_via1_4
* cell instance $10657 r0 *1 40.375,23.31
X$10657 554 VIA_via2_5
* cell instance $10658 r0 *1 51.775,24.15
X$10658 555 VIA_via2_5
* cell instance $10659 r0 *1 53.295,24.15
X$10659 555 VIA_via1_4
* cell instance $10660 r0 *1 53.295,24.15
X$10660 555 VIA_via2_5
* cell instance $10661 r0 *1 51.775,21.63
X$10661 555 VIA_via1_4
* cell instance $10662 r0 *1 51.775,23.17
X$10662 555 VIA_via1_4
* cell instance $10663 r0 *1 53.105,48.51
X$10663 556 VIA_via2_5
* cell instance $10664 r0 *1 51.965,48.51
X$10664 556 VIA_via2_5
* cell instance $10665 r0 *1 53.105,45.57
X$10665 556 VIA_via2_5
* cell instance $10666 r0 *1 53.865,45.57
X$10666 556 VIA_via2_5
* cell instance $10667 r0 *1 53.865,24.99
X$10667 556 VIA_via2_5
* cell instance $10668 r0 *1 53.865,37.17
X$10668 556 VIA_via1_4
* cell instance $10669 r0 *1 53.105,46.83
X$10669 556 VIA_via1_4
* cell instance $10670 r0 *1 51.775,48.37
X$10670 556 VIA_via1_4
* cell instance $10671 r0 *1 50.445,48.37
X$10671 556 VIA_via1_4
* cell instance $10672 r0 *1 50.445,48.51
X$10672 556 VIA_via2_5
* cell instance $10673 r0 *1 55.385,45.57
X$10673 556 VIA_via1_4
* cell instance $10674 r0 *1 55.385,45.57
X$10674 556 VIA_via2_5
* cell instance $10675 r0 *1 55.195,24.43
X$10675 556 VIA_via1_4
* cell instance $10676 r0 *1 55.005,24.99
X$10676 556 VIA_via1_7
* cell instance $10677 r0 *1 55.005,24.99
X$10677 556 VIA_via2_5
* cell instance $10678 r0 *1 55.195,23.17
X$10678 556 VIA_via1_4
* cell instance $10679 r0 *1 52.345,23.17
X$10679 556 VIA_via1_4
* cell instance $10680 r0 *1 52.345,23.31
X$10680 556 VIA_via2_5
* cell instance $10681 r0 *1 53.865,23.17
X$10681 556 VIA_via1_4
* cell instance $10682 r0 *1 53.865,23.31
X$10682 556 VIA_via2_5
* cell instance $10683 r0 *1 51.015,23.17
X$10683 556 VIA_via1_4
* cell instance $10684 r0 *1 51.015,23.31
X$10684 556 VIA_via2_5
* cell instance $10685 r0 *1 54.245,34.37
X$10685 556 VIA_via1_4
* cell instance $10686 r0 *1 55.385,23.31
X$10686 557 VIA_via2_5
* cell instance $10687 r0 *1 54.435,23.73
X$10687 557 VIA_via2_5
* cell instance $10688 r0 *1 63.175,52.01
X$10688 557 VIA_via2_5
* cell instance $10689 r0 *1 50.255,52.01
X$10689 557 VIA_via2_5
* cell instance $10690 r0 *1 48.925,23.73
X$10690 557 VIA_via2_5
* cell instance $10691 r0 *1 59.755,26.95
X$10691 557 VIA_via2_5
* cell instance $10692 r0 *1 55.385,24.99
X$10692 557 VIA_via2_5
* cell instance $10693 r0 *1 59.755,24.99
X$10693 557 VIA_via2_5
* cell instance $10694 r0 *1 48.925,23.17
X$10694 557 VIA_via1_4
* cell instance $10695 r0 *1 54.435,23.17
X$10695 557 VIA_via1_4
* cell instance $10696 r0 *1 54.435,23.31
X$10696 557 VIA_via2_5
* cell instance $10697 r0 *1 59.185,27.23
X$10697 557 VIA_via1_4
* cell instance $10698 r0 *1 50.255,52.43
X$10698 557 VIA_via1_4
* cell instance $10699 r0 *1 63.175,53.55
X$10699 557 VIA_via1_4
* cell instance $10700 r0 *1 63.555,54.39
X$10700 557 VIA_via1_7
* cell instance $10701 r0 *1 63.745,55.23
X$10701 557 VIA_via1_4
* cell instance $10702 r0 *1 60.015,26.95
X$10702 557 VIA_via4_0
* cell instance $10703 r0 *1 60.015,26.95
X$10703 557 VIA_via5_0
* cell instance $10704 r0 *1 60.015,26.95
X$10704 557 VIA_via3_2
* cell instance $10705 r0 *1 60.015,51.03
X$10705 557 VIA_via4_0
* cell instance $10706 r0 *1 60.015,51.03
X$10706 557 VIA_via5_0
* cell instance $10707 r0 *1 60.015,52.01
X$10707 557 VIA_via3_2
* cell instance $10708 r0 *1 56.525,23.17
X$10708 558 VIA_via2_5
* cell instance $10709 r0 *1 56.525,22.05
X$10709 558 VIA_via1_4
* cell instance $10710 r0 *1 56.145,23.17
X$10710 558 VIA_via1_4
* cell instance $10711 r0 *1 56.145,23.17
X$10711 558 VIA_via2_5
* cell instance $10712 r0 *1 53.295,23.17
X$10712 558 VIA_via1_4
* cell instance $10713 r0 *1 53.295,23.17
X$10713 558 VIA_via2_5
* cell instance $10714 r0 *1 70.965,31.43
X$10714 559 VIA_via1_7
* cell instance $10715 r0 *1 69.065,23.03
X$10715 559 VIA_via1_7
* cell instance $10716 r0 *1 72.485,46.97
X$10716 559 VIA_via1_7
* cell instance $10717 r0 *1 71.915,67.83
X$10717 559 VIA_via1_7
* cell instance $10718 r0 *1 61.275,67.83
X$10718 559 VIA_via1_7
* cell instance $10719 r0 *1 64.695,52.85
X$10719 559 VIA_via2_5
* cell instance $10720 r0 *1 71.915,67.55
X$10720 559 VIA_via2_5
* cell instance $10721 r0 *1 72.295,23.59
X$10721 559 VIA_via2_5
* cell instance $10722 r0 *1 69.065,23.59
X$10722 559 VIA_via2_5
* cell instance $10723 r0 *1 69.255,40.67
X$10723 559 VIA_via2_5
* cell instance $10724 r0 *1 69.255,40.11
X$10724 559 VIA_via2_5
* cell instance $10725 r0 *1 70.965,23.59
X$10725 559 VIA_via2_5
* cell instance $10726 r0 *1 71.155,40.11
X$10726 559 VIA_via2_5
* cell instance $10727 r0 *1 65.075,40.67
X$10727 559 VIA_via2_5
* cell instance $10728 r0 *1 63.555,40.67
X$10728 559 VIA_via2_5
* cell instance $10729 r0 *1 65.075,47.25
X$10729 559 VIA_via2_5
* cell instance $10730 r0 *1 64.695,47.25
X$10730 559 VIA_via2_5
* cell instance $10731 r0 *1 72.485,47.25
X$10731 559 VIA_via2_5
* cell instance $10732 r0 *1 63.555,39.97
X$10732 559 VIA_via1_4
* cell instance $10733 r0 *1 72.295,24.43
X$10733 559 VIA_via1_4
* cell instance $10734 r0 *1 72.295,23.17
X$10734 559 VIA_via1_4
* cell instance $10735 r0 *1 61.085,23.17
X$10735 559 VIA_via1_4
* cell instance $10736 r0 *1 61.085,23.31
X$10736 559 VIA_via2_5
* cell instance $10737 r0 *1 61.465,52.85
X$10737 559 VIA_via1_4
* cell instance $10738 r0 *1 61.465,52.85
X$10738 559 VIA_via2_5
* cell instance $10739 r0 *1 72.485,59.57
X$10739 559 VIA_via1_4
* cell instance $10740 r0 *1 61.135,67.55
X$10740 559 VIA_via4_0
* cell instance $10741 r0 *1 61.135,67.55
X$10741 559 VIA_via3_2
* cell instance $10742 r0 *1 61.275,67.55
X$10742 559 VIA_via2_5
* cell instance $10743 r0 *1 71.495,67.55
X$10743 559 VIA_via3_2
* cell instance $10744 r0 *1 71.495,67.55
X$10744 559 VIA_via4_0
* cell instance $10745 r0 *1 61.135,52.85
X$10745 559 VIA_via3_2
* cell instance $10746 r0 *1 65.075,22.61
X$10746 560 VIA_via1_7
* cell instance $10747 r0 *1 65.265,20.37
X$10747 560 VIA_via1_4
* cell instance $10748 r0 *1 71.725,23.17
X$10748 561 VIA_via2_5
* cell instance $10749 r0 *1 68.685,23.17
X$10749 561 VIA_via2_5
* cell instance $10750 r0 *1 69.255,23.17
X$10750 561 VIA_via1_4
* cell instance $10751 r0 *1 69.255,23.17
X$10751 561 VIA_via2_5
* cell instance $10752 r0 *1 68.685,21.63
X$10752 561 VIA_via1_4
* cell instance $10753 r0 *1 71.725,24.15
X$10753 561 VIA_via1_4
* cell instance $10754 r0 *1 78.185,22.05
X$10754 562 VIA_via2_5
* cell instance $10755 r0 *1 78.185,23.59
X$10755 562 VIA_via2_5
* cell instance $10756 r0 *1 76.095,23.59
X$10756 562 VIA_via2_5
* cell instance $10757 r0 *1 78.185,23.17
X$10757 562 VIA_via1_4
* cell instance $10758 r0 *1 79.515,22.05
X$10758 562 VIA_via1_4
* cell instance $10759 r0 *1 79.515,22.05
X$10759 562 VIA_via2_5
* cell instance $10760 r0 *1 76.095,23.17
X$10760 562 VIA_via1_4
* cell instance $10761 r0 *1 79.705,23.17
X$10761 563 VIA_via1_4
* cell instance $10762 r0 *1 79.895,21.91
X$10762 563 VIA_via1_4
* cell instance $10763 r0 *1 79.895,23.17
X$10763 564 VIA_via1_4
* cell instance $10764 r0 *1 80.275,22.89
X$10764 564 VIA_via1_4
* cell instance $10765 r0 *1 83.125,22.19
X$10765 565 VIA_via1_7
* cell instance $10766 r0 *1 82.935,23.31
X$10766 565 VIA_via2_5
* cell instance $10767 r0 *1 80.085,23.17
X$10767 565 VIA_via1_4
* cell instance $10768 r0 *1 80.085,23.31
X$10768 565 VIA_via2_5
* cell instance $10769 r0 *1 87.685,22.61
X$10769 566 VIA_via1_7
* cell instance $10770 r0 *1 86.545,21.63
X$10770 566 VIA_via1_4
* cell instance $10771 r0 *1 92.435,21.91
X$10771 567 VIA_via1_4
* cell instance $10772 r0 *1 92.245,24.43
X$10772 567 VIA_via1_4
* cell instance $10773 r0 *1 96.235,23.17
X$10773 568 VIA_via2_5
* cell instance $10774 r0 *1 96.235,22.05
X$10774 568 VIA_via1_4
* cell instance $10775 r0 *1 95.665,23.17
X$10775 568 VIA_via1_4
* cell instance $10776 r0 *1 95.665,23.17
X$10776 568 VIA_via2_5
* cell instance $10777 r0 *1 93.765,23.17
X$10777 568 VIA_via1_4
* cell instance $10778 r0 *1 93.765,23.31
X$10778 568 VIA_via2_5
* cell instance $10779 r0 *1 7.125,24.01
X$10779 569 VIA_via1_7
* cell instance $10780 r0 *1 7.125,23.17
X$10780 569 VIA_via2_5
* cell instance $10781 r0 *1 3.135,23.17
X$10781 569 VIA_via1_4
* cell instance $10782 r0 *1 3.135,23.17
X$10782 569 VIA_via2_5
* cell instance $10783 r0 *1 94.715,23.17
X$10783 570 VIA_via1_4
* cell instance $10784 r0 *1 94.715,23.17
X$10784 570 VIA_via2_5
* cell instance $10785 r0 *1 92.435,23.17
X$10785 570 VIA_via1_4
* cell instance $10786 r0 *1 92.435,23.17
X$10786 570 VIA_via2_5
* cell instance $10787 r0 *1 12.445,23.17
X$10787 571 VIA_via1_4
* cell instance $10788 r0 *1 12.445,23.17
X$10788 571 VIA_via2_5
* cell instance $10789 r0 *1 8.835,23.17
X$10789 571 VIA_via1_4
* cell instance $10790 r0 *1 8.835,23.17
X$10790 571 VIA_via2_5
* cell instance $10791 r0 *1 90.535,23.17
X$10791 572 VIA_via1_4
* cell instance $10792 r0 *1 90.345,23.17
X$10792 572 VIA_via1_4
* cell instance $10793 r0 *1 88.825,23.17
X$10793 573 VIA_via2_5
* cell instance $10794 r0 *1 88.825,22.05
X$10794 573 VIA_via1_4
* cell instance $10795 r0 *1 86.735,23.17
X$10795 573 VIA_via1_4
* cell instance $10796 r0 *1 86.735,23.17
X$10796 573 VIA_via2_5
* cell instance $10797 r0 *1 89.395,23.17
X$10797 573 VIA_via1_4
* cell instance $10798 r0 *1 89.395,23.17
X$10798 573 VIA_via2_5
* cell instance $10799 r0 *1 16.245,23.03
X$10799 574 VIA_via2_5
* cell instance $10800 r0 *1 16.245,24.43
X$10800 574 VIA_via1_4
* cell instance $10801 r0 *1 17.005,23.03
X$10801 574 VIA_via1_4
* cell instance $10802 r0 *1 17.005,23.03
X$10802 574 VIA_via2_5
* cell instance $10803 r0 *1 84.075,22.89
X$10803 575 VIA_via2_5
* cell instance $10804 r0 *1 84.075,23.17
X$10804 575 VIA_via1_4
* cell instance $10805 r0 *1 83.125,22.89
X$10805 575 VIA_via1_4
* cell instance $10806 r0 *1 83.125,22.89
X$10806 575 VIA_via2_5
* cell instance $10807 r0 *1 24.985,23.17
X$10807 576 VIA_via2_5
* cell instance $10808 r0 *1 25.365,23.17
X$10808 576 VIA_via2_5
* cell instance $10809 r0 *1 24.985,21.63
X$10809 576 VIA_via1_4
* cell instance $10810 r0 *1 25.365,24.15
X$10810 576 VIA_via1_4
* cell instance $10811 r0 *1 23.845,23.17
X$10811 576 VIA_via1_4
* cell instance $10812 r0 *1 23.845,23.17
X$10812 576 VIA_via2_5
* cell instance $10813 r0 *1 75.335,23.17
X$10813 577 VIA_via1_4
* cell instance $10814 r0 *1 75.335,23.17
X$10814 577 VIA_via2_5
* cell instance $10815 r0 *1 79.135,23.17
X$10815 577 VIA_via1_4
* cell instance $10816 r0 *1 79.135,23.17
X$10816 577 VIA_via2_5
* cell instance $10817 r0 *1 40.945,22.05
X$10817 578 VIA_via1_4
* cell instance $10818 r0 *1 39.045,23.17
X$10818 578 VIA_via1_4
* cell instance $10819 r0 *1 39.045,23.17
X$10819 578 VIA_via2_5
* cell instance $10820 r0 *1 40.945,23.17
X$10820 578 VIA_via1_4
* cell instance $10821 r0 *1 40.945,23.17
X$10821 578 VIA_via2_5
* cell instance $10822 r0 *1 41.325,22.61
X$10822 579 VIA_via1_7
* cell instance $10823 r0 *1 41.325,20.37
X$10823 579 VIA_via1_4
* cell instance $10824 r0 *1 73.815,22.05
X$10824 580 VIA_via1_4
* cell instance $10825 r0 *1 73.815,23.17
X$10825 580 VIA_via1_4
* cell instance $10826 r0 *1 73.815,23.17
X$10826 580 VIA_via2_5
* cell instance $10827 r0 *1 72.485,23.17
X$10827 580 VIA_via1_4
* cell instance $10828 r0 *1 72.485,23.17
X$10828 580 VIA_via2_5
* cell instance $10829 r0 *1 46.265,22.19
X$10829 581 VIA_via1_7
* cell instance $10830 r0 *1 46.265,23.17
X$10830 581 VIA_via2_5
* cell instance $10831 r0 *1 43.605,23.17
X$10831 581 VIA_via1_4
* cell instance $10832 r0 *1 43.605,23.17
X$10832 581 VIA_via2_5
* cell instance $10833 r0 *1 67.735,22.19
X$10833 582 VIA_via1_7
* cell instance $10834 r0 *1 67.735,23.17
X$10834 582 VIA_via2_5
* cell instance $10835 r0 *1 66.595,23.17
X$10835 582 VIA_via1_4
* cell instance $10836 r0 *1 66.595,23.17
X$10836 582 VIA_via2_5
* cell instance $10837 r0 *1 64.695,23.17
X$10837 583 VIA_via1_4
* cell instance $10838 r0 *1 64.695,23.17
X$10838 583 VIA_via2_5
* cell instance $10839 r0 *1 63.555,23.17
X$10839 583 VIA_via1_4
* cell instance $10840 r0 *1 63.555,23.17
X$10840 583 VIA_via2_5
* cell instance $10841 r0 *1 62.225,22.61
X$10841 584 VIA_via1_7
* cell instance $10842 r0 *1 62.225,22.61
X$10842 584 VIA_via2_5
* cell instance $10843 r0 *1 60.325,22.61
X$10843 584 VIA_via2_5
* cell instance $10844 r0 *1 60.325,21.63
X$10844 584 VIA_via1_4
* cell instance $10845 r0 *1 61.275,23.17
X$10845 585 VIA_via1_4
* cell instance $10846 r0 *1 61.275,23.03
X$10846 585 VIA_via2_5
* cell instance $10847 r0 *1 62.605,22.05
X$10847 585 VIA_via1_4
* cell instance $10848 r0 *1 62.605,23.17
X$10848 585 VIA_via1_4
* cell instance $10849 r0 *1 62.605,23.03
X$10849 585 VIA_via2_5
* cell instance $10850 r0 *1 54.245,22.61
X$10850 586 VIA_via1_7
* cell instance $10851 r0 *1 54.245,21.63
X$10851 586 VIA_via1_4
* cell instance $10852 r0 *1 58.235,22.05
X$10852 587 VIA_via2_5
* cell instance $10853 r0 *1 57.095,22.05
X$10853 587 VIA_via1_4
* cell instance $10854 r0 *1 57.095,22.05
X$10854 587 VIA_via2_5
* cell instance $10855 r0 *1 58.235,21.63
X$10855 587 VIA_via1_4
* cell instance $10856 r0 *1 57.095,22.61
X$10856 588 VIA_via1_7
* cell instance $10857 r0 *1 57.095,22.61
X$10857 588 VIA_via2_5
* cell instance $10858 r0 *1 57.855,22.61
X$10858 588 VIA_via2_5
* cell instance $10859 r0 *1 57.855,20.37
X$10859 588 VIA_via1_4
* cell instance $10860 r0 *1 5.225,24.99
X$10860 589 VIA_via1_7
* cell instance $10861 r0 *1 4.275,25.97
X$10861 589 VIA_via1_4
* cell instance $10862 r0 *1 6.365,25.27
X$10862 590 VIA_via2_5
* cell instance $10863 r0 *1 4.275,25.27
X$10863 590 VIA_via2_5
* cell instance $10864 r0 *1 6.175,23.17
X$10864 590 VIA_via1_4
* cell instance $10865 r0 *1 4.275,24.43
X$10865 590 VIA_via1_4
* cell instance $10866 r0 *1 6.555,25.55
X$10866 590 VIA_via1_4
* cell instance $10867 r0 *1 7.885,26.81
X$10867 591 VIA_via1_7
* cell instance $10868 r0 *1 7.885,27.79
X$10868 591 VIA_via1_7
* cell instance $10869 r0 *1 7.885,35.49
X$10869 591 VIA_via2_5
* cell instance $10870 r0 *1 12.065,24.57
X$10870 591 VIA_via2_5
* cell instance $10871 r0 *1 4.275,46.83
X$10871 591 VIA_via2_5
* cell instance $10872 r0 *1 7.885,24.71
X$10872 591 VIA_via2_5
* cell instance $10873 r0 *1 6.745,24.71
X$10873 591 VIA_via2_5
* cell instance $10874 r0 *1 4.845,24.71
X$10874 591 VIA_via2_5
* cell instance $10875 r0 *1 13.015,46.55
X$10875 591 VIA_via2_5
* cell instance $10876 r0 *1 14.155,46.55
X$10876 591 VIA_via2_5
* cell instance $10877 r0 *1 6.745,24.43
X$10877 591 VIA_via1_4
* cell instance $10878 r0 *1 12.065,23.17
X$10878 591 VIA_via1_4
* cell instance $10879 r0 *1 4.845,24.43
X$10879 591 VIA_via1_4
* cell instance $10880 r0 *1 4.275,35.63
X$10880 591 VIA_via1_4
* cell instance $10881 r0 *1 4.275,35.63
X$10881 591 VIA_via2_5
* cell instance $10882 r0 *1 5.795,46.83
X$10882 591 VIA_via1_4
* cell instance $10883 r0 *1 5.795,46.83
X$10883 591 VIA_via2_5
* cell instance $10884 r0 *1 4.275,45.57
X$10884 591 VIA_via1_4
* cell instance $10885 r0 *1 13.205,24.43
X$10885 591 VIA_via1_4
* cell instance $10886 r0 *1 13.205,24.57
X$10886 591 VIA_via2_5
* cell instance $10887 r0 *1 14.345,35.63
X$10887 591 VIA_via1_4
* cell instance $10888 r0 *1 14.345,35.49
X$10888 591 VIA_via2_5
* cell instance $10889 r0 *1 14.155,46.83
X$10889 591 VIA_via1_4
* cell instance $10890 r0 *1 13.395,48.37
X$10890 591 VIA_via1_4
* cell instance $10891 r0 *1 11.495,25.13
X$10891 592 VIA_via2_5
* cell instance $10892 r0 *1 12.635,25.13
X$10892 592 VIA_via2_5
* cell instance $10893 r0 *1 11.495,23.17
X$10893 592 VIA_via1_4
* cell instance $10894 r0 *1 11.115,23.45
X$10894 592 VIA_via1_4
* cell instance $10895 r0 *1 12.635,25.97
X$10895 592 VIA_via1_4
* cell instance $10896 r0 *1 12.255,24.85
X$10896 593 VIA_via1_4
* cell instance $10897 r0 *1 12.065,25.97
X$10897 593 VIA_via1_4
* cell instance $10898 r0 *1 12.635,24.43
X$10898 593 VIA_via1_4
* cell instance $10899 r0 *1 13.965,24.01
X$10899 594 VIA_via1_7
* cell instance $10900 r0 *1 12.825,23.17
X$10900 594 VIA_via1_4
* cell instance $10901 r0 *1 13.015,25.41
X$10901 595 VIA_via1_7
* cell instance $10902 r0 *1 13.775,24.43
X$10902 595 VIA_via1_4
* cell instance $10903 r0 *1 32.965,23.59
X$10903 596 VIA_via1_7
* cell instance $10904 r0 *1 32.585,24.43
X$10904 596 VIA_via1_4
* cell instance $10905 r0 *1 58.235,25.83
X$10905 597 VIA_via1_7
* cell instance $10906 r0 *1 58.235,23.59
X$10906 597 VIA_via2_5
* cell instance $10907 r0 *1 53.105,23.45
X$10907 597 VIA_via2_5
* cell instance $10908 r0 *1 48.735,23.45
X$10908 597 VIA_via2_5
* cell instance $10909 r0 *1 48.355,24.43
X$10909 597 VIA_via1_4
* cell instance $10910 r0 *1 48.925,52.43
X$10910 597 VIA_via1_4
* cell instance $10911 r0 *1 48.925,52.43
X$10911 597 VIA_via2_5
* cell instance $10912 r0 *1 53.105,23.17
X$10912 597 VIA_via1_4
* cell instance $10913 r0 *1 65.455,53.55
X$10913 597 VIA_via1_4
* cell instance $10914 r0 *1 65.455,53.55
X$10914 597 VIA_via2_5
* cell instance $10915 r0 *1 65.645,53.97
X$10915 597 VIA_via1_4
* cell instance $10916 r0 *1 49.095,52.15
X$10916 597 VIA_via4_0
* cell instance $10917 r0 *1 65.615,52.43
X$10917 597 VIA_via4_0
* cell instance $10918 r0 *1 65.615,53.55
X$10918 597 VIA_via3_2
* cell instance $10919 r0 *1 49.095,52.43
X$10919 597 VIA_via3_2
* cell instance $10920 r0 *1 60.515,27.37
X$10920 598 VIA_via1_7
* cell instance $10921 r0 *1 60.515,27.37
X$10921 598 VIA_via2_5
* cell instance $10922 r0 *1 60.575,27.37
X$10922 598 VIA_via3_2
* cell instance $10923 r0 *1 60.325,53.83
X$10923 598 VIA_via2_5
* cell instance $10924 r0 *1 46.455,23.31
X$10924 598 VIA_via2_5
* cell instance $10925 r0 *1 50.445,27.23
X$10925 598 VIA_via2_5
* cell instance $10926 r0 *1 46.455,24.43
X$10926 598 VIA_via1_4
* cell instance $10927 r0 *1 61.275,41.23
X$10927 598 VIA_via1_4
* cell instance $10928 r0 *1 61.275,41.23
X$10928 598 VIA_via2_5
* cell instance $10929 r0 *1 46.645,53.97
X$10929 598 VIA_via1_4
* cell instance $10930 r0 *1 46.645,53.83
X$10930 598 VIA_via2_5
* cell instance $10931 r0 *1 50.255,23.17
X$10931 598 VIA_via1_4
* cell instance $10932 r0 *1 50.255,23.31
X$10932 598 VIA_via2_5
* cell instance $10933 r0 *1 60.325,53.55
X$10933 598 VIA_via1_4
* cell instance $10934 r0 *1 60.575,41.23
X$10934 598 VIA_via3_2
* cell instance $10935 r0 *1 60.575,53.83
X$10935 598 VIA_via3_2
* cell instance $10936 r0 *1 63.365,54.81
X$10936 599 VIA_via1_7
* cell instance $10937 r0 *1 62.035,25.83
X$10937 599 VIA_via1_7
* cell instance $10938 r0 *1 51.585,23.59
X$10938 599 VIA_via2_5
* cell instance $10939 r0 *1 63.175,51.03
X$10939 599 VIA_via2_5
* cell instance $10940 r0 *1 63.365,51.03
X$10940 599 VIA_via2_5
* cell instance $10941 r0 *1 47.975,23.59
X$10941 599 VIA_via2_5
* cell instance $10942 r0 *1 51.585,25.13
X$10942 599 VIA_via2_5
* cell instance $10943 r0 *1 62.035,26.39
X$10943 599 VIA_via2_5
* cell instance $10944 r0 *1 62.035,25.13
X$10944 599 VIA_via2_5
* cell instance $10945 r0 *1 63.175,26.39
X$10945 599 VIA_via2_5
* cell instance $10946 r0 *1 47.975,23.17
X$10946 599 VIA_via1_4
* cell instance $10947 r0 *1 62.985,37.17
X$10947 599 VIA_via1_4
* cell instance $10948 r0 *1 46.835,51.17
X$10948 599 VIA_via1_4
* cell instance $10949 r0 *1 46.835,51.03
X$10949 599 VIA_via2_5
* cell instance $10950 r0 *1 51.585,23.17
X$10950 599 VIA_via1_4
* cell instance $10951 r0 *1 57.665,24.29
X$10951 600 VIA_via2_5
* cell instance $10952 r0 *1 69.635,46.69
X$10952 600 VIA_via2_5
* cell instance $10953 r0 *1 78.375,35.63
X$10953 600 VIA_via1_4
* cell instance $10954 r0 *1 78.375,35.63
X$10954 600 VIA_via2_5
* cell instance $10955 r0 *1 60.325,46.83
X$10955 600 VIA_via1_4
* cell instance $10956 r0 *1 60.325,46.69
X$10956 600 VIA_via2_5
* cell instance $10957 r0 *1 55.955,24.43
X$10957 600 VIA_via1_4
* cell instance $10958 r0 *1 55.955,24.29
X$10958 600 VIA_via2_5
* cell instance $10959 r0 *1 57.665,23.17
X$10959 600 VIA_via1_4
* cell instance $10960 r0 *1 62.985,24.43
X$10960 600 VIA_via1_4
* cell instance $10961 r0 *1 62.985,24.43
X$10961 600 VIA_via2_5
* cell instance $10962 r0 *1 69.635,49.91
X$10962 600 VIA_via1_4
* cell instance $10963 r0 *1 77.935,46.69
X$10963 600 VIA_via3_2
* cell instance $10964 r0 *1 62.815,24.43
X$10964 600 VIA_via3_2
* cell instance $10965 r0 *1 77.935,35.63
X$10965 600 VIA_via3_2
* cell instance $10966 r0 *1 62.815,46.69
X$10966 600 VIA_via3_2
* cell instance $10967 r0 *1 62.415,24.43
X$10967 601 VIA_via1_4
* cell instance $10968 r0 *1 62.035,24.85
X$10968 601 VIA_via1_4
* cell instance $10969 r0 *1 55.385,34.23
X$10969 602 VIA_via1_7
* cell instance $10970 r0 *1 55.385,34.23
X$10970 602 VIA_via2_5
* cell instance $10971 r0 *1 61.275,34.23
X$10971 602 VIA_via1_7
* cell instance $10972 r0 *1 61.275,34.23
X$10972 602 VIA_via2_5
* cell instance $10973 r0 *1 34.485,28.63
X$10973 602 VIA_via1_7
* cell instance $10974 r0 *1 34.485,28.49
X$10974 602 VIA_via2_5
* cell instance $10975 r0 *1 29.355,31.43
X$10975 602 VIA_via1_7
* cell instance $10976 r0 *1 37.715,31.43
X$10976 602 VIA_via1_7
* cell instance $10977 r0 *1 45.315,28.63
X$10977 602 VIA_via1_7
* cell instance $10978 r0 *1 45.315,28.49
X$10978 602 VIA_via2_5
* cell instance $10979 r0 *1 51.205,28.49
X$10979 602 VIA_via2_5
* cell instance $10980 r0 *1 62.795,34.23
X$10980 602 VIA_via2_5
* cell instance $10981 r0 *1 24.795,29.05
X$10981 602 VIA_via2_5
* cell instance $10982 r0 *1 29.735,29.05
X$10982 602 VIA_via2_5
* cell instance $10983 r0 *1 34.485,29.05
X$10983 602 VIA_via2_5
* cell instance $10984 r0 *1 42.275,28.49
X$10984 602 VIA_via2_5
* cell instance $10985 r0 *1 37.905,28.49
X$10985 602 VIA_via2_5
* cell instance $10986 r0 *1 55.385,28.91
X$10986 602 VIA_via2_5
* cell instance $10987 r0 *1 20.235,29.05
X$10987 602 VIA_via2_5
* cell instance $10988 r0 *1 62.415,23.17
X$10988 602 VIA_via1_4
* cell instance $10989 r0 *1 51.205,28.77
X$10989 602 VIA_via1_4
* cell instance $10990 r0 *1 51.205,28.91
X$10990 602 VIA_via2_5
* cell instance $10991 r0 *1 20.235,30.03
X$10991 602 VIA_via1_4
* cell instance $10992 r0 *1 24.795,28.77
X$10992 602 VIA_via1_4
* cell instance $10993 r0 *1 42.275,24.85
X$10993 602 VIA_via1_4
* cell instance $10994 r0 *1 63.365,20.79
X$10994 603 VIA_via1_7
* cell instance $10995 r0 *1 63.365,24.43
X$10995 603 VIA_via1_4
* cell instance $10996 r0 *1 70.205,23.59
X$10996 604 VIA_via1_7
* cell instance $10997 r0 *1 69.445,24.43
X$10997 604 VIA_via1_4
* cell instance $10998 r0 *1 73.435,24.99
X$10998 605 VIA_via1_7
* cell instance $10999 r0 *1 72.105,25.97
X$10999 605 VIA_via1_4
* cell instance $11000 r0 *1 72.485,24.71
X$11000 606 VIA_via2_5
* cell instance $11001 r0 *1 74.385,24.71
X$11001 606 VIA_via2_5
* cell instance $11002 r0 *1 73.815,24.71
X$11002 606 VIA_via2_5
* cell instance $11003 r0 *1 74.385,25.55
X$11003 606 VIA_via1_4
* cell instance $11004 r0 *1 73.815,24.43
X$11004 606 VIA_via1_4
* cell instance $11005 r0 *1 72.485,24.43
X$11005 606 VIA_via1_4
* cell instance $11006 r0 *1 74.765,24.01
X$11006 607 VIA_via1_7
* cell instance $11007 r0 *1 75.145,23.17
X$11007 607 VIA_via1_4
* cell instance $11008 r0 *1 92.245,48.51
X$11008 608 VIA_via2_5
* cell instance $11009 r0 *1 92.245,24.71
X$11009 608 VIA_via2_5
* cell instance $11010 r0 *1 91.675,48.37
X$11010 608 VIA_via1_4
* cell instance $11011 r0 *1 91.675,48.51
X$11011 608 VIA_via2_5
* cell instance $11012 r0 *1 91.865,24.29
X$11012 608 VIA_via1_4
* cell instance $11013 r0 *1 91.865,24.29
X$11013 608 VIA_via2_5
* cell instance $11014 r0 *1 92.245,51.17
X$11014 608 VIA_via1_4
* cell instance $11015 r0 *1 92.625,23.59
X$11015 609 VIA_via1_7
* cell instance $11016 r0 *1 92.435,24.43
X$11016 609 VIA_via1_4
* cell instance $11017 r0 *1 5.415,24.43
X$11017 610 VIA_via2_5
* cell instance $11018 r0 *1 6.745,23.17
X$11018 610 VIA_via1_4
* cell instance $11019 r0 *1 6.745,23.31
X$11019 610 VIA_via2_5
* cell instance $11020 r0 *1 5.415,23.31
X$11020 610 VIA_via1_4
* cell instance $11021 r0 *1 5.415,23.31
X$11021 610 VIA_via2_5
* cell instance $11022 r0 *1 6.175,24.43
X$11022 610 VIA_via1_4
* cell instance $11023 r0 *1 6.175,24.43
X$11023 610 VIA_via2_5
* cell instance $11024 r0 *1 9.975,24.43
X$11024 611 VIA_via1_4
* cell instance $11025 r0 *1 9.975,24.29
X$11025 611 VIA_via2_5
* cell instance $11026 r0 *1 13.585,24.29
X$11026 611 VIA_via1_4
* cell instance $11027 r0 *1 13.585,24.29
X$11027 611 VIA_via2_5
* cell instance $11028 r0 *1 90.725,23.59
X$11028 612 VIA_via1_7
* cell instance $11029 r0 *1 91.485,23.87
X$11029 612 VIA_via2_5
* cell instance $11030 r0 *1 90.725,23.87
X$11030 612 VIA_via2_5
* cell instance $11031 r0 *1 91.485,24.43
X$11031 612 VIA_via1_4
* cell instance $11032 r0 *1 91.675,24.43
X$11032 613 VIA_via1_4
* cell instance $11033 r0 *1 91.675,24.43
X$11033 613 VIA_via2_5
* cell instance $11034 r0 *1 86.735,24.43
X$11034 613 VIA_via1_4
* cell instance $11035 r0 *1 86.735,24.43
X$11035 613 VIA_via2_5
* cell instance $11036 r0 *1 20.045,48.65
X$11036 614 VIA_via2_5
* cell instance $11037 r0 *1 13.775,23.45
X$11037 614 VIA_via1_4
* cell instance $11038 r0 *1 13.775,23.45
X$11038 614 VIA_via2_5
* cell instance $11039 r0 *1 18.335,48.37
X$11039 614 VIA_via1_4
* cell instance $11040 r0 *1 18.335,48.51
X$11040 614 VIA_via2_5
* cell instance $11041 r0 *1 20.045,48.37
X$11041 614 VIA_via1_4
* cell instance $11042 r0 *1 16.055,23.45
X$11042 614 VIA_via3_2
* cell instance $11043 r0 *1 16.055,48.51
X$11043 614 VIA_via3_2
* cell instance $11044 r0 *1 24.795,23.59
X$11044 615 VIA_via1_7
* cell instance $11045 r0 *1 24.795,24.43
X$11045 615 VIA_via2_5
* cell instance $11046 r0 *1 23.085,24.43
X$11046 615 VIA_via1_4
* cell instance $11047 r0 *1 23.085,24.43
X$11047 615 VIA_via2_5
* cell instance $11048 r0 *1 77.615,24.15
X$11048 616 VIA_via2_5
* cell instance $11049 r0 *1 77.615,24.43
X$11049 616 VIA_via2_5
* cell instance $11050 r0 *1 75.335,24.43
X$11050 616 VIA_via1_4
* cell instance $11051 r0 *1 75.335,24.43
X$11051 616 VIA_via2_5
* cell instance $11052 r0 *1 79.515,24.15
X$11052 616 VIA_via1_4
* cell instance $11053 r0 *1 79.515,24.15
X$11053 616 VIA_via2_5
* cell instance $11054 r0 *1 77.615,23.17
X$11054 616 VIA_via1_4
* cell instance $11055 r0 *1 79.895,24.01
X$11055 617 VIA_via1_7
* cell instance $11056 r0 *1 79.895,24.01
X$11056 617 VIA_via2_5
* cell instance $11057 r0 *1 78.945,24.01
X$11057 617 VIA_via2_5
* cell instance $11058 r0 *1 78.945,23.17
X$11058 617 VIA_via1_4
* cell instance $11059 r0 *1 78.565,23.59
X$11059 618 VIA_via1_7
* cell instance $11060 r0 *1 78.565,23.59
X$11060 618 VIA_via2_5
* cell instance $11061 r0 *1 79.705,23.59
X$11061 618 VIA_via2_5
* cell instance $11062 r0 *1 79.705,24.43
X$11062 618 VIA_via1_4
* cell instance $11063 r0 *1 76.285,24.43
X$11063 619 VIA_via1_4
* cell instance $11064 r0 *1 77.235,24.43
X$11064 619 VIA_via1_4
* cell instance $11065 r0 *1 52.725,50.89
X$11065 620 VIA_via2_5
* cell instance $11066 r0 *1 47.975,42.21
X$11066 620 VIA_via2_5
* cell instance $11067 r0 *1 47.215,42.21
X$11067 620 VIA_via2_5
* cell instance $11068 r0 *1 47.405,23.45
X$11068 620 VIA_via2_5
* cell instance $11069 r0 *1 47.405,24.43
X$11069 620 VIA_via2_5
* cell instance $11070 r0 *1 47.025,23.45
X$11070 620 VIA_via2_5
* cell instance $11071 r0 *1 48.165,50.89
X$11071 620 VIA_via2_5
* cell instance $11072 r0 *1 42.655,52.85
X$11072 620 VIA_via2_5
* cell instance $11073 r0 *1 39.615,54.25
X$11073 620 VIA_via2_5
* cell instance $11074 r0 *1 38.665,54.25
X$11074 620 VIA_via2_5
* cell instance $11075 r0 *1 39.615,52.85
X$11075 620 VIA_via2_5
* cell instance $11076 r0 *1 58.995,42.21
X$11076 620 VIA_via2_5
* cell instance $11077 r0 *1 61.465,42.21
X$11077 620 VIA_via2_5
* cell instance $11078 r0 *1 58.995,42.77
X$11078 620 VIA_via1_4
* cell instance $11079 r0 *1 41.705,24.43
X$11079 620 VIA_via1_4
* cell instance $11080 r0 *1 41.705,24.43
X$11080 620 VIA_via2_5
* cell instance $11081 r0 *1 47.025,23.17
X$11081 620 VIA_via1_4
* cell instance $11082 r0 *1 61.465,37.17
X$11082 620 VIA_via1_4
* cell instance $11083 r0 *1 38.665,55.23
X$11083 620 VIA_via1_4
* cell instance $11084 r0 *1 42.655,51.17
X$11084 620 VIA_via1_4
* cell instance $11085 r0 *1 42.655,51.03
X$11085 620 VIA_via2_5
* cell instance $11086 r0 *1 45.885,51.03
X$11086 620 VIA_via1_4
* cell instance $11087 r0 *1 45.885,51.03
X$11087 620 VIA_via2_5
* cell instance $11088 r0 *1 48.165,51.17
X$11088 620 VIA_via1_4
* cell instance $11089 r0 *1 39.805,48.37
X$11089 620 VIA_via1_4
* cell instance $11090 r0 *1 52.725,52.43
X$11090 620 VIA_via1_4
* cell instance $11091 r0 *1 47.405,25.97
X$11091 620 VIA_via1_4
* cell instance $11092 r0 *1 52.725,24.43
X$11092 621 VIA_via2_5
* cell instance $11093 r0 *1 51.015,24.43
X$11093 621 VIA_via1_4
* cell instance $11094 r0 *1 51.015,24.43
X$11094 621 VIA_via2_5
* cell instance $11095 r0 *1 52.725,23.03
X$11095 621 VIA_via1_4
* cell instance $11096 r0 *1 59.755,24.43
X$11096 622 VIA_via1_4
* cell instance $11097 r0 *1 59.755,24.43
X$11097 622 VIA_via2_5
* cell instance $11098 r0 *1 62.605,24.43
X$11098 622 VIA_via1_4
* cell instance $11099 r0 *1 62.605,24.43
X$11099 622 VIA_via2_5
* cell instance $11100 r0 *1 60.705,23.59
X$11100 623 VIA_via1_7
* cell instance $11101 r0 *1 60.705,23.59
X$11101 623 VIA_via2_5
* cell instance $11102 r0 *1 63.175,23.59
X$11102 623 VIA_via2_5
* cell instance $11103 r0 *1 63.175,24.43
X$11103 623 VIA_via1_4
* cell instance $11104 r0 *1 64.315,36.89
X$11104 624 VIA_via2_5
* cell instance $11105 r0 *1 64.315,24.15
X$11105 624 VIA_via2_5
* cell instance $11106 r0 *1 63.365,24.15
X$11106 624 VIA_via1_4
* cell instance $11107 r0 *1 63.365,24.15
X$11107 624 VIA_via2_5
* cell instance $11108 r0 *1 83.505,51.17
X$11108 624 VIA_via1_4
* cell instance $11109 r0 *1 83.505,51.03
X$11109 624 VIA_via2_5
* cell instance $11110 r0 *1 82.175,51.17
X$11110 624 VIA_via1_4
* cell instance $11111 r0 *1 82.175,51.17
X$11111 624 VIA_via2_5
* cell instance $11112 r0 *1 82.415,36.61
X$11112 624 VIA_via3_2
* cell instance $11113 r0 *1 82.415,51.17
X$11113 624 VIA_via3_2
* cell instance $11114 r0 *1 1.615,25.27
X$11114 625 VIA_via2_5
* cell instance $11115 r0 *1 1.615,25.97
X$11115 625 VIA_via1_4
* cell instance $11116 r0 *1 0.935,25.27
X$11116 625 VIA_via3_2
* cell instance $11117 r0 *1 0.935,25.27
X$11117 625 VIA_via4_0
* cell instance $11118 r0 *1 2.375,26.39
X$11118 626 VIA_via2_5
* cell instance $11119 r0 *1 2.375,25.97
X$11119 626 VIA_via1_4
* cell instance $11120 r0 *1 1.215,26.39
X$11120 626 VIA_via3_2
* cell instance $11121 r0 *1 1.215,26.39
X$11121 626 VIA_via4_0
* cell instance $11122 r0 *1 20.805,88.97
X$11122 627 VIA_via1_7
* cell instance $11123 r0 *1 30.305,88.97
X$11123 627 VIA_via1_7
* cell instance $11124 r0 *1 14.345,53.83
X$11124 627 VIA_via1_7
* cell instance $11125 r0 *1 14.345,53.69
X$11125 627 VIA_via2_5
* cell instance $11126 r0 *1 30.305,89.25
X$11126 627 VIA_via2_5
* cell instance $11127 r0 *1 30.305,89.81
X$11127 627 VIA_via2_5
* cell instance $11128 r0 *1 47.595,91.07
X$11128 627 VIA_via2_5
* cell instance $11129 r0 *1 48.165,91.07
X$11129 627 VIA_via2_5
* cell instance $11130 r0 *1 11.685,74.13
X$11130 627 VIA_via2_5
* cell instance $11131 r0 *1 11.875,87.99
X$11131 627 VIA_via2_5
* cell instance $11132 r0 *1 11.305,87.99
X$11132 627 VIA_via2_5
* cell instance $11133 r0 *1 12.445,74.13
X$11133 627 VIA_via2_5
* cell instance $11134 r0 *1 20.805,89.25
X$11134 627 VIA_via2_5
* cell instance $11135 r0 *1 20.805,87.99
X$11135 627 VIA_via2_5
* cell instance $11136 r0 *1 36.955,91.07
X$11136 627 VIA_via2_5
* cell instance $11137 r0 *1 36.955,89.25
X$11137 627 VIA_via2_5
* cell instance $11138 r0 *1 36.955,90.37
X$11138 627 VIA_via1_4
* cell instance $11139 r0 *1 47.595,90.37
X$11139 627 VIA_via1_4
* cell instance $11140 r0 *1 48.165,87.57
X$11140 627 VIA_via1_4
* cell instance $11141 r0 *1 12.635,65.17
X$11141 627 VIA_via1_4
* cell instance $11142 r0 *1 12.635,65.17
X$11142 627 VIA_via2_5
* cell instance $11143 r0 *1 12.695,65.17
X$11143 627 VIA_via3_2
* cell instance $11144 r0 *1 11.305,87.57
X$11144 627 VIA_via1_4
* cell instance $11145 r0 *1 11.875,25.97
X$11145 627 VIA_via1_4
* cell instance $11146 r0 *1 11.875,25.97
X$11146 627 VIA_via2_5
* cell instance $11147 r0 *1 11.685,73.57
X$11147 627 VIA_via1_4
* cell instance $11148 r0 *1 47.975,25.83
X$11148 627 VIA_via1_4
* cell instance $11149 r0 *1 47.975,25.83
X$11149 627 VIA_via2_5
* cell instance $11150 r0 *1 12.695,53.69
X$11150 627 VIA_via3_2
* cell instance $11151 r0 *1 12.695,74.13
X$11151 627 VIA_via3_2
* cell instance $11152 r0 *1 12.695,25.97
X$11152 627 VIA_via3_2
* cell instance $11153 r0 *1 16.435,34.23
X$11153 628 VIA_via1_7
* cell instance $11154 r0 *1 16.435,34.23
X$11154 628 VIA_via2_5
* cell instance $11155 r0 *1 27.835,31.43
X$11155 628 VIA_via1_7
* cell instance $11156 r0 *1 31.065,28.63
X$11156 628 VIA_via1_7
* cell instance $11157 r0 *1 31.065,28.63
X$11157 628 VIA_via2_5
* cell instance $11158 r0 *1 50.445,28.91
X$11158 628 VIA_via2_5
* cell instance $11159 r0 *1 27.645,28.63
X$11159 628 VIA_via2_5
* cell instance $11160 r0 *1 31.065,29.19
X$11160 628 VIA_via2_5
* cell instance $11161 r0 *1 36.575,29.19
X$11161 628 VIA_via2_5
* cell instance $11162 r0 *1 21.945,28.63
X$11162 628 VIA_via2_5
* cell instance $11163 r0 *1 18.145,34.23
X$11163 628 VIA_via2_5
* cell instance $11164 r0 *1 18.145,27.37
X$11164 628 VIA_via2_5
* cell instance $11165 r0 *1 21.945,27.37
X$11165 628 VIA_via2_5
* cell instance $11166 r0 *1 14.155,34.23
X$11166 628 VIA_via2_5
* cell instance $11167 r0 *1 49.875,28.77
X$11167 628 VIA_via1_4
* cell instance $11168 r0 *1 49.875,28.91
X$11168 628 VIA_via2_5
* cell instance $11169 r0 *1 12.825,35.63
X$11169 628 VIA_via1_4
* cell instance $11170 r0 *1 12.825,35.63
X$11170 628 VIA_via2_5
* cell instance $11171 r0 *1 14.155,35.63
X$11171 628 VIA_via1_4
* cell instance $11172 r0 *1 14.155,35.63
X$11172 628 VIA_via2_5
* cell instance $11173 r0 *1 50.825,33.95
X$11173 628 VIA_via1_4
* cell instance $11174 r0 *1 18.525,25.97
X$11174 628 VIA_via1_4
* cell instance $11175 r0 *1 21.945,25.97
X$11175 628 VIA_via1_4
* cell instance $11176 r0 *1 36.575,28.77
X$11176 628 VIA_via1_4
* cell instance $11177 r0 *1 36.575,28.91
X$11177 628 VIA_via2_5
* cell instance $11178 r0 *1 43.415,28.77
X$11178 628 VIA_via1_4
* cell instance $11179 r0 *1 43.415,28.91
X$11179 628 VIA_via2_5
* cell instance $11180 r0 *1 20.425,30.03
X$11180 629 VIA_via1_4
* cell instance $11181 r0 *1 20.805,27.23
X$11181 629 VIA_via1_4
* cell instance $11182 r0 *1 19.285,25.97
X$11182 629 VIA_via1_4
* cell instance $11183 r0 *1 22.135,27.23
X$11183 630 VIA_via1_4
* cell instance $11184 r0 *1 23.085,25.69
X$11184 630 VIA_via1_4
* cell instance $11185 r0 *1 24.985,26.95
X$11185 631 VIA_via2_5
* cell instance $11186 r0 *1 22.705,26.95
X$11186 631 VIA_via2_5
* cell instance $11187 r0 *1 24.415,26.95
X$11187 631 VIA_via1_4
* cell instance $11188 r0 *1 24.415,26.95
X$11188 631 VIA_via2_5
* cell instance $11189 r0 *1 22.705,25.97
X$11189 631 VIA_via1_4
* cell instance $11190 r0 *1 24.985,28.77
X$11190 631 VIA_via1_4
* cell instance $11191 r0 *1 52.535,28.63
X$11191 632 VIA_via1_7
* cell instance $11192 r0 *1 20.805,28.63
X$11192 632 VIA_via1_7
* cell instance $11193 r0 *1 27.075,28.63
X$11193 632 VIA_via1_7
* cell instance $11194 r0 *1 52.535,27.09
X$11194 632 VIA_via2_5
* cell instance $11195 r0 *1 27.455,26.95
X$11195 632 VIA_via2_5
* cell instance $11196 r0 *1 40.375,27.09
X$11196 632 VIA_via2_5
* cell instance $11197 r0 *1 20.805,29.47
X$11197 632 VIA_via2_5
* cell instance $11198 r0 *1 20.995,27.09
X$11198 632 VIA_via2_5
* cell instance $11199 r0 *1 15.675,29.47
X$11199 632 VIA_via2_5
* cell instance $11200 r0 *1 13.965,27.23
X$11200 632 VIA_via1_4
* cell instance $11201 r0 *1 15.675,30.03
X$11201 632 VIA_via1_4
* cell instance $11202 r0 *1 15.675,30.03
X$11202 632 VIA_via2_5
* cell instance $11203 r0 *1 14.155,30.03
X$11203 632 VIA_via1_4
* cell instance $11204 r0 *1 14.155,30.03
X$11204 632 VIA_via2_5
* cell instance $11205 r0 *1 24.605,27.23
X$11205 632 VIA_via1_4
* cell instance $11206 r0 *1 24.605,27.09
X$11206 632 VIA_via2_5
* cell instance $11207 r0 *1 52.915,31.57
X$11207 632 VIA_via1_4
* cell instance $11208 r0 *1 34.295,27.23
X$11208 632 VIA_via1_4
* cell instance $11209 r0 *1 34.295,27.09
X$11209 632 VIA_via2_5
* cell instance $11210 r0 *1 42.655,27.23
X$11210 632 VIA_via1_4
* cell instance $11211 r0 *1 42.655,27.09
X$11211 632 VIA_via2_5
* cell instance $11212 r0 *1 40.375,30.03
X$11212 632 VIA_via1_4
* cell instance $11213 r0 *1 35.435,26.81
X$11213 633 VIA_via1_7
* cell instance $11214 r0 *1 34.865,25.97
X$11214 633 VIA_via1_4
* cell instance $11215 r0 *1 40.945,45.85
X$11215 634 VIA_via2_5
* cell instance $11216 r0 *1 44.555,52.85
X$11216 634 VIA_via2_5
* cell instance $11217 r0 *1 43.985,45.29
X$11217 634 VIA_via2_5
* cell instance $11218 r0 *1 42.465,45.29
X$11218 634 VIA_via2_5
* cell instance $11219 r0 *1 41.895,45.29
X$11219 634 VIA_via2_5
* cell instance $11220 r0 *1 41.895,45.85
X$11220 634 VIA_via2_5
* cell instance $11221 r0 *1 47.405,52.85
X$11221 634 VIA_via2_5
* cell instance $11222 r0 *1 44.555,53.97
X$11222 634 VIA_via2_5
* cell instance $11223 r0 *1 43.035,26.81
X$11223 634 VIA_via2_5
* cell instance $11224 r0 *1 25.745,27.09
X$11224 634 VIA_via2_5
* cell instance $11225 r0 *1 32.775,26.81
X$11225 634 VIA_via2_5
* cell instance $11226 r0 *1 32.775,27.09
X$11226 634 VIA_via2_5
* cell instance $11227 r0 *1 40.755,26.81
X$11227 634 VIA_via2_5
* cell instance $11228 r0 *1 47.595,26.81
X$11228 634 VIA_via2_5
* cell instance $11229 r0 *1 40.945,46.83
X$11229 634 VIA_via1_4
* cell instance $11230 r0 *1 31.825,45.57
X$11230 634 VIA_via1_4
* cell instance $11231 r0 *1 31.825,45.57
X$11231 634 VIA_via2_5
* cell instance $11232 r0 *1 44.555,51.45
X$11232 634 VIA_via1_4
* cell instance $11233 r0 *1 47.595,49.63
X$11233 634 VIA_via1_4
* cell instance $11234 r0 *1 43.035,53.97
X$11234 634 VIA_via1_4
* cell instance $11235 r0 *1 43.035,53.97
X$11235 634 VIA_via2_5
* cell instance $11236 r0 *1 25.935,27.23
X$11236 634 VIA_via1_4
* cell instance $11237 r0 *1 32.775,25.97
X$11237 634 VIA_via1_4
* cell instance $11238 r0 *1 24.795,45.57
X$11238 634 VIA_via1_4
* cell instance $11239 r0 *1 24.795,45.57
X$11239 634 VIA_via2_5
* cell instance $11240 r0 *1 47.595,27.23
X$11240 634 VIA_via1_4
* cell instance $11241 r0 *1 40.755,27.23
X$11241 634 VIA_via1_4
* cell instance $11242 r0 *1 43.035,30.03
X$11242 634 VIA_via1_4
* cell instance $11243 r0 *1 43.795,26.81
X$11243 635 VIA_via1_7
* cell instance $11244 r0 *1 43.605,25.97
X$11244 635 VIA_via1_4
* cell instance $11245 r0 *1 44.365,32.83
X$11245 636 VIA_via2_5
* cell instance $11246 r0 *1 41.515,32.83
X$11246 636 VIA_via2_5
* cell instance $11247 r0 *1 41.325,37.17
X$11247 636 VIA_via1_4
* cell instance $11248 r0 *1 40.375,38.43
X$11248 636 VIA_via1_4
* cell instance $11249 r0 *1 45.505,31.57
X$11249 636 VIA_via1_4
* cell instance $11250 r0 *1 44.365,33.95
X$11250 636 VIA_via1_4
* cell instance $11251 r0 *1 44.745,34.79
X$11251 636 VIA_via1_7
* cell instance $11252 r0 *1 44.935,35.63
X$11252 636 VIA_via1_4
* cell instance $11253 r0 *1 45.315,32.83
X$11253 636 VIA_via1_4
* cell instance $11254 r0 *1 45.315,32.83
X$11254 636 VIA_via2_5
* cell instance $11255 r0 *1 42.085,32.83
X$11255 636 VIA_via1_4
* cell instance $11256 r0 *1 42.085,32.83
X$11256 636 VIA_via2_5
* cell instance $11257 r0 *1 44.365,25.97
X$11257 636 VIA_via1_4
* cell instance $11258 r0 *1 45.505,27.23
X$11258 636 VIA_via1_4
* cell instance $11259 r0 *1 46.075,27.23
X$11259 637 VIA_via2_5
* cell instance $11260 r0 *1 45.885,26.25
X$11260 637 VIA_via1_4
* cell instance $11261 r0 *1 46.075,28.77
X$11261 637 VIA_via1_4
* cell instance $11262 r0 *1 43.415,27.23
X$11262 637 VIA_via1_4
* cell instance $11263 r0 *1 43.415,27.23
X$11263 637 VIA_via2_5
* cell instance $11264 r0 *1 58.425,25.97
X$11264 638 VIA_via1_4
* cell instance $11265 r0 *1 58.045,27.23
X$11265 638 VIA_via1_4
* cell instance $11266 r0 *1 58.045,26.25
X$11266 638 VIA_via1_4
* cell instance $11267 r0 *1 58.995,26.81
X$11267 639 VIA_via1_7
* cell instance $11268 r0 *1 59.565,24.43
X$11268 639 VIA_via1_4
* cell instance $11269 r0 *1 60.135,48.09
X$11269 640 VIA_via2_5
* cell instance $11270 r0 *1 58.805,48.09
X$11270 640 VIA_via2_5
* cell instance $11271 r0 *1 61.465,31.71
X$11271 640 VIA_via2_5
* cell instance $11272 r0 *1 60.135,45.29
X$11272 640 VIA_via2_5
* cell instance $11273 r0 *1 60.705,45.29
X$11273 640 VIA_via2_5
* cell instance $11274 r0 *1 58.425,45.29
X$11274 640 VIA_via2_5
* cell instance $11275 r0 *1 60.705,31.71
X$11275 640 VIA_via2_5
* cell instance $11276 r0 *1 61.275,25.83
X$11276 640 VIA_via2_5
* cell instance $11277 r0 *1 60.705,38.15
X$11277 640 VIA_via2_5
* cell instance $11278 r0 *1 59.375,38.15
X$11278 640 VIA_via2_5
* cell instance $11279 r0 *1 59.945,31.57
X$11279 640 VIA_via2_5
* cell instance $11280 r0 *1 59.185,31.57
X$11280 640 VIA_via1_4
* cell instance $11281 r0 *1 59.185,31.57
X$11281 640 VIA_via2_5
* cell instance $11282 r0 *1 59.375,38.43
X$11282 640 VIA_via1_4
* cell instance $11283 r0 *1 61.275,27.23
X$11283 640 VIA_via1_4
* cell instance $11284 r0 *1 61.275,27.23
X$11284 640 VIA_via2_5
* cell instance $11285 r0 *1 58.425,45.57
X$11285 640 VIA_via1_4
* cell instance $11286 r0 *1 60.705,44.03
X$11286 640 VIA_via1_4
* cell instance $11287 r0 *1 60.135,48.37
X$11287 640 VIA_via1_4
* cell instance $11288 r0 *1 58.805,48.37
X$11288 640 VIA_via1_4
* cell instance $11289 r0 *1 58.995,25.97
X$11289 640 VIA_via1_4
* cell instance $11290 r0 *1 58.995,25.83
X$11290 640 VIA_via2_5
* cell instance $11291 r0 *1 59.945,27.23
X$11291 640 VIA_via1_4
* cell instance $11292 r0 *1 59.945,27.23
X$11292 640 VIA_via2_5
* cell instance $11293 r0 *1 61.465,32.83
X$11293 640 VIA_via1_4
* cell instance $11294 r0 *1 62.795,25.97
X$11294 640 VIA_via1_4
* cell instance $11295 r0 *1 62.795,25.83
X$11295 640 VIA_via2_5
* cell instance $11296 r0 *1 62.605,25.97
X$11296 641 VIA_via2_5
* cell instance $11297 r0 *1 62.225,25.97
X$11297 641 VIA_via1_4
* cell instance $11298 r0 *1 62.225,25.97
X$11298 641 VIA_via2_5
* cell instance $11299 r0 *1 62.605,27.23
X$11299 641 VIA_via1_4
* cell instance $11300 r0 *1 66.405,25.83
X$11300 641 VIA_via1_4
* cell instance $11301 r0 *1 66.405,25.83
X$11301 641 VIA_via2_5
* cell instance $11302 r0 *1 75.335,26.95
X$11302 642 VIA_via1_4
* cell instance $11303 r0 *1 74.765,25.97
X$11303 642 VIA_via1_4
* cell instance $11304 r0 *1 74.385,24.43
X$11304 642 VIA_via1_4
* cell instance $11305 r0 *1 84.645,26.39
X$11305 643 VIA_via1_7
* cell instance $11306 r0 *1 84.455,27.23
X$11306 643 VIA_via1_4
* cell instance $11307 r0 *1 90.345,25.97
X$11307 644 VIA_via2_5
* cell instance $11308 r0 *1 90.345,26.95
X$11308 644 VIA_via1_4
* cell instance $11309 r0 *1 86.925,25.97
X$11309 644 VIA_via1_4
* cell instance $11310 r0 *1 86.925,25.97
X$11310 644 VIA_via2_5
* cell instance $11311 r0 *1 86.165,25.97
X$11311 644 VIA_via1_4
* cell instance $11312 r0 *1 86.165,25.97
X$11312 644 VIA_via2_5
* cell instance $11313 r0 *1 87.875,26.39
X$11313 645 VIA_via1_7
* cell instance $11314 r0 *1 88.065,27.23
X$11314 645 VIA_via1_4
* cell instance $11315 r0 *1 94.145,27.23
X$11315 646 VIA_via1_4
* cell instance $11316 r0 *1 94.145,27.23
X$11316 646 VIA_via2_5
* cell instance $11317 r0 *1 96.615,26.25
X$11317 646 VIA_via1_4
* cell instance $11318 r0 *1 96.235,27.23
X$11318 646 VIA_via1_4
* cell instance $11319 r0 *1 96.235,27.23
X$11319 646 VIA_via2_5
* cell instance $11320 r0 *1 92.625,30.03
X$11320 647 VIA_via2_5
* cell instance $11321 r0 *1 93.005,35.63
X$11321 647 VIA_via2_5
* cell instance $11322 r0 *1 93.005,34.37
X$11322 647 VIA_via2_5
* cell instance $11323 r0 *1 93.005,33.67
X$11323 647 VIA_via2_5
* cell instance $11324 r0 *1 88.445,33.67
X$11324 647 VIA_via2_5
* cell instance $11325 r0 *1 91.675,30.03
X$11325 647 VIA_via2_5
* cell instance $11326 r0 *1 91.675,25.97
X$11326 647 VIA_via2_5
* cell instance $11327 r0 *1 88.065,33.67
X$11327 647 VIA_via2_5
* cell instance $11328 r0 *1 91.485,30.03
X$11328 647 VIA_via1_4
* cell instance $11329 r0 *1 95.095,25.97
X$11329 647 VIA_via1_4
* cell instance $11330 r0 *1 95.095,25.97
X$11330 647 VIA_via2_5
* cell instance $11331 r0 *1 88.445,32.83
X$11331 647 VIA_via1_4
* cell instance $11332 r0 *1 91.295,25.97
X$11332 647 VIA_via1_4
* cell instance $11333 r0 *1 91.295,25.97
X$11333 647 VIA_via2_5
* cell instance $11334 r0 *1 95.095,28.77
X$11334 647 VIA_via1_4
* cell instance $11335 r0 *1 94.525,35.63
X$11335 647 VIA_via1_4
* cell instance $11336 r0 *1 94.525,35.63
X$11336 647 VIA_via2_5
* cell instance $11337 r0 *1 88.065,34.37
X$11337 647 VIA_via1_4
* cell instance $11338 r0 *1 92.625,31.57
X$11338 647 VIA_via1_4
* cell instance $11339 r0 *1 93.005,31.99
X$11339 647 VIA_via1_7
* cell instance $11340 r0 *1 92.625,34.37
X$11340 647 VIA_via1_4
* cell instance $11341 r0 *1 92.625,34.37
X$11341 647 VIA_via2_5
* cell instance $11342 r0 *1 92.435,26.81
X$11342 648 VIA_via1_7
* cell instance $11343 r0 *1 92.435,26.81
X$11343 648 VIA_via2_5
* cell instance $11344 r0 *1 90.535,26.81
X$11344 648 VIA_via2_5
* cell instance $11345 r0 *1 90.535,25.97
X$11345 648 VIA_via1_4
* cell instance $11346 r0 *1 91.485,50.89
X$11346 649 VIA_via2_5
* cell instance $11347 r0 *1 92.055,50.89
X$11347 649 VIA_via2_5
* cell instance $11348 r0 *1 79.325,25.41
X$11348 649 VIA_via2_5
* cell instance $11349 r0 *1 79.325,23.31
X$11349 649 VIA_via1_4
* cell instance $11350 r0 *1 91.485,48.37
X$11350 649 VIA_via1_4
* cell instance $11351 r0 *1 91.485,48.37
X$11351 649 VIA_via2_5
* cell instance $11352 r0 *1 92.055,51.17
X$11352 649 VIA_via1_4
* cell instance $11353 r0 *1 89.135,25.41
X$11353 649 VIA_via3_2
* cell instance $11354 r0 *1 89.135,48.37
X$11354 649 VIA_via3_2
* cell instance $11355 r0 *1 86.545,25.41
X$11355 650 VIA_via1_7
* cell instance $11356 r0 *1 86.545,24.43
X$11356 650 VIA_via1_4
* cell instance $11357 r0 *1 85.595,26.95
X$11357 651 VIA_via2_5
* cell instance $11358 r0 *1 86.735,26.95
X$11358 651 VIA_via1_4
* cell instance $11359 r0 *1 86.735,26.95
X$11359 651 VIA_via2_5
* cell instance $11360 r0 *1 83.695,25.97
X$11360 651 VIA_via1_4
* cell instance $11361 r0 *1 83.695,25.97
X$11361 651 VIA_via2_5
* cell instance $11362 r0 *1 85.595,25.97
X$11362 651 VIA_via1_4
* cell instance $11363 r0 *1 85.595,25.97
X$11363 651 VIA_via2_5
* cell instance $11364 r0 *1 19.665,26.39
X$11364 652 VIA_via1_7
* cell instance $11365 r0 *1 19.665,26.39
X$11365 652 VIA_via2_5
* cell instance $11366 r0 *1 18.525,26.39
X$11366 652 VIA_via2_5
* cell instance $11367 r0 *1 18.525,27.23
X$11367 652 VIA_via1_4
* cell instance $11368 r0 *1 22.895,25.97
X$11368 653 VIA_via2_5
* cell instance $11369 r0 *1 22.515,27.23
X$11369 653 VIA_via2_5
* cell instance $11370 r0 *1 23.845,25.97
X$11370 653 VIA_via2_5
* cell instance $11371 r0 *1 16.245,31.57
X$11371 653 VIA_via2_5
* cell instance $11372 r0 *1 19.665,31.57
X$11372 653 VIA_via2_5
* cell instance $11373 r0 *1 23.845,24.43
X$11373 653 VIA_via1_4
* cell instance $11374 r0 *1 17.195,31.57
X$11374 653 VIA_via1_4
* cell instance $11375 r0 *1 17.195,31.57
X$11375 653 VIA_via2_5
* cell instance $11376 r0 *1 16.245,32.83
X$11376 653 VIA_via1_4
* cell instance $11377 r0 *1 19.095,28.77
X$11377 653 VIA_via1_4
* cell instance $11378 r0 *1 19.285,27.23
X$11378 653 VIA_via1_4
* cell instance $11379 r0 *1 19.285,27.23
X$11379 653 VIA_via2_5
* cell instance $11380 r0 *1 19.665,30.03
X$11380 653 VIA_via1_4
* cell instance $11381 r0 *1 22.515,28.35
X$11381 653 VIA_via1_4
* cell instance $11382 r0 *1 22.895,27.23
X$11382 653 VIA_via1_4
* cell instance $11383 r0 *1 22.895,27.23
X$11383 653 VIA_via2_5
* cell instance $11384 r0 *1 15.865,28.77
X$11384 653 VIA_via1_4
* cell instance $11385 r0 *1 24.795,25.97
X$11385 653 VIA_via1_4
* cell instance $11386 r0 *1 24.795,25.97
X$11386 653 VIA_via2_5
* cell instance $11387 r0 *1 75.715,26.39
X$11387 654 VIA_via1_7
* cell instance $11388 r0 *1 75.715,26.39
X$11388 654 VIA_via2_5
* cell instance $11389 r0 *1 73.055,26.39
X$11389 654 VIA_via2_5
* cell instance $11390 r0 *1 73.055,27.23
X$11390 654 VIA_via1_4
* cell instance $11391 r0 *1 38.665,31.71
X$11391 655 VIA_via2_5
* cell instance $11392 r0 *1 39.615,31.71
X$11392 655 VIA_via2_5
* cell instance $11393 r0 *1 32.585,25.97
X$11393 655 VIA_via2_5
* cell instance $11394 r0 *1 33.915,29.75
X$11394 655 VIA_via2_5
* cell instance $11395 r0 *1 33.915,25.97
X$11395 655 VIA_via2_5
* cell instance $11396 r0 *1 34.295,30.03
X$11396 655 VIA_via2_5
* cell instance $11397 r0 *1 39.995,31.71
X$11397 655 VIA_via2_5
* cell instance $11398 r0 *1 30.685,30.03
X$11398 655 VIA_via1_4
* cell instance $11399 r0 *1 30.685,30.03
X$11399 655 VIA_via2_5
* cell instance $11400 r0 *1 39.995,32.83
X$11400 655 VIA_via1_4
* cell instance $11401 r0 *1 32.585,27.23
X$11401 655 VIA_via1_4
* cell instance $11402 r0 *1 35.625,25.97
X$11402 655 VIA_via1_4
* cell instance $11403 r0 *1 35.625,25.97
X$11403 655 VIA_via2_5
* cell instance $11404 r0 *1 34.485,31.57
X$11404 655 VIA_via1_4
* cell instance $11405 r0 *1 34.485,31.71
X$11405 655 VIA_via2_5
* cell instance $11406 r0 *1 36.575,31.71
X$11406 655 VIA_via1_4
* cell instance $11407 r0 *1 36.575,31.71
X$11407 655 VIA_via2_5
* cell instance $11408 r0 *1 38.665,30.03
X$11408 655 VIA_via1_4
* cell instance $11409 r0 *1 37.145,31.57
X$11409 655 VIA_via1_4
* cell instance $11410 r0 *1 37.145,31.71
X$11410 655 VIA_via2_5
* cell instance $11411 r0 *1 37.145,34.37
X$11411 655 VIA_via1_4
* cell instance $11412 r0 *1 39.615,28.77
X$11412 655 VIA_via1_4
* cell instance $11413 r0 *1 62.985,26.81
X$11413 656 VIA_via1_7
* cell instance $11414 r0 *1 62.985,26.81
X$11414 656 VIA_via2_5
* cell instance $11415 r0 *1 61.655,26.81
X$11415 656 VIA_via2_5
* cell instance $11416 r0 *1 61.655,24.43
X$11416 656 VIA_via1_4
* cell instance $11417 r0 *1 63.175,26.11
X$11417 657 VIA_via1_4
* cell instance $11418 r0 *1 63.175,26.11
X$11418 657 VIA_via2_5
* cell instance $11419 r0 *1 64.125,25.97
X$11419 657 VIA_via1_4
* cell instance $11420 r0 *1 64.125,26.11
X$11420 657 VIA_via2_5
* cell instance $11421 r0 *1 55.765,25.97
X$11421 658 VIA_via1_4
* cell instance $11422 r0 *1 55.765,25.97
X$11422 658 VIA_via2_5
* cell instance $11423 r0 *1 59.375,25.97
X$11423 658 VIA_via1_4
* cell instance $11424 r0 *1 59.375,25.97
X$11424 658 VIA_via2_5
* cell instance $11425 r0 *1 4.085,27.37
X$11425 659 VIA_via1_7
* cell instance $11426 r0 *1 4.085,27.37
X$11426 659 VIA_via2_5
* cell instance $11427 r0 *1 49.875,30.17
X$11427 659 VIA_via1_7
* cell instance $11428 r0 *1 49.875,30.17
X$11428 659 VIA_via2_5
* cell instance $11429 r0 *1 33.725,30.17
X$11429 659 VIA_via1_7
* cell instance $11430 r0 *1 33.725,30.31
X$11430 659 VIA_via2_5
* cell instance $11431 r0 *1 44.745,30.17
X$11431 659 VIA_via1_7
* cell instance $11432 r0 *1 44.745,30.17
X$11432 659 VIA_via2_5
* cell instance $11433 r0 *1 9.785,30.45
X$11433 659 VIA_via2_5
* cell instance $11434 r0 *1 51.395,30.17
X$11434 659 VIA_via2_5
* cell instance $11435 r0 *1 28.785,30.17
X$11435 659 VIA_via2_5
* cell instance $11436 r0 *1 39.045,30.31
X$11436 659 VIA_via2_5
* cell instance $11437 r0 *1 21.945,30.45
X$11437 659 VIA_via2_5
* cell instance $11438 r0 *1 8.455,27.23
X$11438 659 VIA_via1_4
* cell instance $11439 r0 *1 8.455,27.37
X$11439 659 VIA_via2_5
* cell instance $11440 r0 *1 9.785,27.23
X$11440 659 VIA_via1_4
* cell instance $11441 r0 *1 9.785,27.37
X$11441 659 VIA_via2_5
* cell instance $11442 r0 *1 3.895,30.03
X$11442 659 VIA_via1_4
* cell instance $11443 r0 *1 21.945,30.03
X$11443 659 VIA_via1_4
* cell instance $11444 r0 *1 21.945,30.03
X$11444 659 VIA_via2_5
* cell instance $11445 r0 *1 51.395,32.55
X$11445 659 VIA_via1_4
* cell instance $11446 r0 *1 28.785,28.77
X$11446 659 VIA_via1_4
* cell instance $11447 r0 *1 39.045,31.57
X$11447 659 VIA_via1_4
* cell instance $11448 r0 *1 6.745,28.77
X$11448 660 VIA_via2_5
* cell instance $11449 r0 *1 10.735,30.03
X$11449 660 VIA_via2_5
* cell instance $11450 r0 *1 5.035,28.77
X$11450 660 VIA_via2_5
* cell instance $11451 r0 *1 13.015,30.03
X$11451 660 VIA_via2_5
* cell instance $11452 r0 *1 10.735,28.77
X$11452 660 VIA_via1_4
* cell instance $11453 r0 *1 6.745,30.03
X$11453 660 VIA_via1_4
* cell instance $11454 r0 *1 6.745,30.03
X$11454 660 VIA_via2_5
* cell instance $11455 r0 *1 8.455,30.03
X$11455 660 VIA_via1_4
* cell instance $11456 r0 *1 8.455,30.03
X$11456 660 VIA_via2_5
* cell instance $11457 r0 *1 9.405,30.03
X$11457 660 VIA_via1_4
* cell instance $11458 r0 *1 9.405,30.03
X$11458 660 VIA_via2_5
* cell instance $11459 r0 *1 7.125,28.77
X$11459 660 VIA_via1_4
* cell instance $11460 r0 *1 7.125,28.77
X$11460 660 VIA_via2_5
* cell instance $11461 r0 *1 11.685,30.03
X$11461 660 VIA_via1_4
* cell instance $11462 r0 *1 11.685,30.03
X$11462 660 VIA_via2_5
* cell instance $11463 r0 *1 3.705,28.77
X$11463 660 VIA_via1_4
* cell instance $11464 r0 *1 3.705,28.77
X$11464 660 VIA_via2_5
* cell instance $11465 r0 *1 5.035,25.97
X$11465 660 VIA_via1_4
* cell instance $11466 r0 *1 13.015,32.83
X$11466 660 VIA_via1_4
* cell instance $11467 r0 *1 13.395,34.37
X$11467 660 VIA_via1_4
* cell instance $11468 r0 *1 11.495,35.63
X$11468 661 VIA_via1_4
* cell instance $11469 r0 *1 10.545,27.23
X$11469 661 VIA_via1_4
* cell instance $11470 r0 *1 12.255,29.05
X$11470 661 VIA_via1_4
* cell instance $11471 r0 *1 28.215,28.21
X$11471 662 VIA_via1_7
* cell instance $11472 r0 *1 28.595,27.23
X$11472 662 VIA_via1_4
* cell instance $11473 r0 *1 32.205,28.21
X$11473 663 VIA_via1_7
* cell instance $11474 r0 *1 31.825,27.23
X$11474 663 VIA_via1_4
* cell instance $11475 r0 *1 44.555,28.21
X$11475 664 VIA_via1_7
* cell instance $11476 r0 *1 44.745,27.23
X$11476 664 VIA_via1_4
* cell instance $11477 r0 *1 47.025,28.77
X$11477 665 VIA_via2_5
* cell instance $11478 r0 *1 45.505,28.77
X$11478 665 VIA_via1_4
* cell instance $11479 r0 *1 45.505,28.77
X$11479 665 VIA_via2_5
* cell instance $11480 r0 *1 47.025,27.65
X$11480 665 VIA_via1_4
* cell instance $11481 r0 *1 44.175,28.77
X$11481 665 VIA_via1_4
* cell instance $11482 r0 *1 44.175,28.77
X$11482 665 VIA_via2_5
* cell instance $11483 r0 *1 50.825,30.03
X$11483 666 VIA_via2_5
* cell instance $11484 r0 *1 55.955,30.03
X$11484 666 VIA_via2_5
* cell instance $11485 r0 *1 55.955,33.11
X$11485 666 VIA_via2_5
* cell instance $11486 r0 *1 59.565,33.11
X$11486 666 VIA_via2_5
* cell instance $11487 r0 *1 61.085,33.11
X$11487 666 VIA_via2_5
* cell instance $11488 r0 *1 61.085,31.57
X$11488 666 VIA_via1_4
* cell instance $11489 r0 *1 55.955,31.57
X$11489 666 VIA_via1_4
* cell instance $11490 r0 *1 50.825,31.57
X$11490 666 VIA_via1_4
* cell instance $11491 r0 *1 53.295,30.03
X$11491 666 VIA_via1_4
* cell instance $11492 r0 *1 53.295,30.03
X$11492 666 VIA_via2_5
* cell instance $11493 r0 *1 50.635,27.23
X$11493 666 VIA_via1_4
* cell instance $11494 r0 *1 56.145,27.23
X$11494 666 VIA_via1_4
* cell instance $11495 r0 *1 55.955,30.45
X$11495 666 VIA_via1_4
* cell instance $11496 r0 *1 56.525,25.97
X$11496 666 VIA_via1_4
* cell instance $11497 r0 *1 59.565,34.37
X$11497 666 VIA_via1_4
* cell instance $11498 r0 *1 52.155,27.65
X$11498 667 VIA_via1_4
* cell instance $11499 r0 *1 51.395,28.77
X$11499 667 VIA_via1_4
* cell instance $11500 r0 *1 51.395,28.77
X$11500 667 VIA_via2_5
* cell instance $11501 r0 *1 50.635,28.77
X$11501 667 VIA_via1_4
* cell instance $11502 r0 *1 50.635,28.77
X$11502 667 VIA_via2_5
* cell instance $11503 r0 *1 54.815,28.77
X$11503 668 VIA_via2_5
* cell instance $11504 r0 *1 53.295,28.77
X$11504 668 VIA_via1_4
* cell instance $11505 r0 *1 53.295,28.77
X$11505 668 VIA_via2_5
* cell instance $11506 r0 *1 54.815,29.75
X$11506 668 VIA_via1_4
* cell instance $11507 r0 *1 51.965,28.77
X$11507 668 VIA_via1_4
* cell instance $11508 r0 *1 51.965,28.77
X$11508 668 VIA_via2_5
* cell instance $11509 r0 *1 58.615,27.23
X$11509 669 VIA_via1_4
* cell instance $11510 r0 *1 58.615,27.23
X$11510 669 VIA_via2_5
* cell instance $11511 r0 *1 59.375,27.23
X$11511 669 VIA_via1_4
* cell instance $11512 r0 *1 59.375,27.23
X$11512 669 VIA_via2_5
* cell instance $11513 r0 *1 57.665,27.23
X$11513 669 VIA_via1_4
* cell instance $11514 r0 *1 57.665,27.23
X$11514 669 VIA_via2_5
* cell instance $11515 r0 *1 61.655,27.79
X$11515 670 VIA_via1_7
* cell instance $11516 r0 *1 61.275,28.77
X$11516 670 VIA_via1_4
* cell instance $11517 r0 *1 63.555,27.09
X$11517 671 VIA_via2_5
* cell instance $11518 r0 *1 60.705,27.23
X$11518 671 VIA_via1_4
* cell instance $11519 r0 *1 60.705,27.09
X$11519 671 VIA_via2_5
* cell instance $11520 r0 *1 62.035,27.23
X$11520 671 VIA_via1_4
* cell instance $11521 r0 *1 62.035,27.09
X$11521 671 VIA_via2_5
* cell instance $11522 r0 *1 63.555,28.35
X$11522 671 VIA_via1_4
* cell instance $11523 r0 *1 79.325,32.41
X$11523 672 VIA_via1_7
* cell instance $11524 r0 *1 79.325,32.41
X$11524 672 VIA_via2_5
* cell instance $11525 r0 *1 69.255,30.17
X$11525 672 VIA_via2_5
* cell instance $11526 r0 *1 71.725,32.27
X$11526 672 VIA_via2_5
* cell instance $11527 r0 *1 70.585,32.27
X$11527 672 VIA_via2_5
* cell instance $11528 r0 *1 69.255,32.27
X$11528 672 VIA_via2_5
* cell instance $11529 r0 *1 79.135,32.41
X$11529 672 VIA_via2_5
* cell instance $11530 r0 *1 77.805,32.13
X$11530 672 VIA_via2_5
* cell instance $11531 r0 *1 74.575,32.27
X$11531 672 VIA_via2_5
* cell instance $11532 r0 *1 75.905,32.27
X$11532 672 VIA_via2_5
* cell instance $11533 r0 *1 80.655,32.41
X$11533 672 VIA_via2_5
* cell instance $11534 r0 *1 80.655,31.57
X$11534 672 VIA_via1_4
* cell instance $11535 r0 *1 75.905,32.83
X$11535 672 VIA_via1_4
* cell instance $11536 r0 *1 79.135,30.03
X$11536 672 VIA_via1_4
* cell instance $11537 r0 *1 77.045,28.77
X$11537 672 VIA_via1_4
* cell instance $11538 r0 *1 74.385,30.03
X$11538 672 VIA_via1_4
* cell instance $11539 r0 *1 77.805,30.03
X$11539 672 VIA_via1_4
* cell instance $11540 r0 *1 67.735,30.03
X$11540 672 VIA_via1_4
* cell instance $11541 r0 *1 67.735,30.17
X$11541 672 VIA_via2_5
* cell instance $11542 r0 *1 69.255,28.77
X$11542 672 VIA_via1_4
* cell instance $11543 r0 *1 71.725,31.57
X$11543 672 VIA_via1_4
* cell instance $11544 r0 *1 70.585,34.37
X$11544 672 VIA_via1_4
* cell instance $11545 r0 *1 88.255,28.77
X$11545 673 VIA_via2_5
* cell instance $11546 r0 *1 88.825,28.77
X$11546 673 VIA_via2_5
* cell instance $11547 r0 *1 85.025,28.77
X$11547 673 VIA_via2_5
* cell instance $11548 r0 *1 85.215,28.77
X$11548 673 VIA_via2_5
* cell instance $11549 r0 *1 81.795,28.77
X$11549 673 VIA_via2_5
* cell instance $11550 r0 *1 81.795,32.83
X$11550 673 VIA_via1_4
* cell instance $11551 r0 *1 85.215,31.57
X$11551 673 VIA_via1_4
* cell instance $11552 r0 *1 88.825,27.23
X$11552 673 VIA_via1_4
* cell instance $11553 r0 *1 88.255,30.03
X$11553 673 VIA_via1_4
* cell instance $11554 r0 *1 79.135,27.23
X$11554 673 VIA_via1_4
* cell instance $11555 r0 *1 85.215,27.23
X$11555 673 VIA_via1_4
* cell instance $11556 r0 *1 79.135,28.77
X$11556 673 VIA_via1_4
* cell instance $11557 r0 *1 79.135,28.77
X$11557 673 VIA_via2_5
* cell instance $11558 r0 *1 83.505,28.77
X$11558 673 VIA_via1_4
* cell instance $11559 r0 *1 83.505,28.77
X$11559 673 VIA_via2_5
* cell instance $11560 r0 *1 85.595,28.77
X$11560 673 VIA_via1_4
* cell instance $11561 r0 *1 85.595,28.77
X$11561 673 VIA_via2_5
* cell instance $11562 r0 *1 91.485,30.31
X$11562 674 VIA_via2_5
* cell instance $11563 r0 *1 92.055,30.17
X$11563 674 VIA_via2_5
* cell instance $11564 r0 *1 91.865,28.35
X$11564 674 VIA_via1_4
* cell instance $11565 r0 *1 91.485,31.57
X$11565 674 VIA_via1_4
* cell instance $11566 r0 *1 70.965,40.53
X$11566 675 VIA_via2_5
* cell instance $11567 r0 *1 70.015,40.53
X$11567 675 VIA_via2_5
* cell instance $11568 r0 *1 96.425,40.25
X$11568 675 VIA_via2_5
* cell instance $11569 r0 *1 95.665,30.03
X$11569 675 VIA_via2_5
* cell instance $11570 r0 *1 96.425,30.03
X$11570 675 VIA_via2_5
* cell instance $11571 r0 *1 84.455,40.25
X$11571 675 VIA_via2_5
* cell instance $11572 r0 *1 84.455,40.53
X$11572 675 VIA_via2_5
* cell instance $11573 r0 *1 84.455,41.23
X$11573 675 VIA_via1_4
* cell instance $11574 r0 *1 94.905,30.03
X$11574 675 VIA_via1_4
* cell instance $11575 r0 *1 94.905,30.03
X$11575 675 VIA_via2_5
* cell instance $11576 r0 *1 93.385,30.03
X$11576 675 VIA_via1_4
* cell instance $11577 r0 *1 93.385,30.03
X$11577 675 VIA_via2_5
* cell instance $11578 r0 *1 91.485,27.23
X$11578 675 VIA_via1_4
* cell instance $11579 r0 *1 91.485,27.09
X$11579 675 VIA_via2_5
* cell instance $11580 r0 *1 95.665,27.23
X$11580 675 VIA_via1_4
* cell instance $11581 r0 *1 95.665,27.09
X$11581 675 VIA_via2_5
* cell instance $11582 r0 *1 96.615,36.05
X$11582 675 VIA_via1_4
* cell instance $11583 r0 *1 69.825,42.77
X$11583 675 VIA_via1_4
* cell instance $11584 r0 *1 70.965,39.97
X$11584 675 VIA_via1_4
* cell instance $11585 r0 *1 94.335,27.37
X$11585 676 VIA_via2_5
* cell instance $11586 r0 *1 96.615,27.37
X$11586 676 VIA_via1_4
* cell instance $11587 r0 *1 96.615,27.37
X$11587 676 VIA_via2_5
* cell instance $11588 r0 *1 94.335,25.97
X$11588 676 VIA_via1_4
* cell instance $11589 r0 *1 5.225,27.79
X$11589 677 VIA_via1_7
* cell instance $11590 r0 *1 5.225,27.79
X$11590 677 VIA_via2_5
* cell instance $11591 r0 *1 2.945,27.79
X$11591 677 VIA_via2_5
* cell instance $11592 r0 *1 2.945,28.77
X$11592 677 VIA_via1_4
* cell instance $11593 r0 *1 94.525,27.79
X$11593 678 VIA_via1_7
* cell instance $11594 r0 *1 94.525,27.79
X$11594 678 VIA_via2_5
* cell instance $11595 r0 *1 91.485,27.79
X$11595 678 VIA_via2_5
* cell instance $11596 r0 *1 91.485,28.77
X$11596 678 VIA_via1_4
* cell instance $11597 r0 *1 9.595,27.79
X$11597 679 VIA_via1_7
* cell instance $11598 r0 *1 9.595,27.79
X$11598 679 VIA_via2_5
* cell instance $11599 r0 *1 6.365,27.79
X$11599 679 VIA_via2_5
* cell instance $11600 r0 *1 6.365,28.77
X$11600 679 VIA_via1_4
* cell instance $11601 r0 *1 92.815,27.23
X$11601 680 VIA_via2_5
* cell instance $11602 r0 *1 93.575,27.23
X$11602 680 VIA_via1_4
* cell instance $11603 r0 *1 93.575,27.23
X$11603 680 VIA_via2_5
* cell instance $11604 r0 *1 92.055,27.23
X$11604 680 VIA_via1_4
* cell instance $11605 r0 *1 92.055,27.23
X$11605 680 VIA_via2_5
* cell instance $11606 r0 *1 92.815,26.25
X$11606 680 VIA_via1_4
* cell instance $11607 r0 *1 10.925,27.79
X$11607 681 VIA_via1_7
* cell instance $11608 r0 *1 10.925,27.79
X$11608 681 VIA_via2_5
* cell instance $11609 r0 *1 9.975,27.79
X$11609 681 VIA_via2_5
* cell instance $11610 r0 *1 9.975,28.77
X$11610 681 VIA_via1_4
* cell instance $11611 r0 *1 79.895,27.65
X$11611 682 VIA_via2_5
* cell instance $11612 r0 *1 79.895,28.91
X$11612 682 VIA_via2_5
* cell instance $11613 r0 *1 76.475,28.77
X$11613 682 VIA_via1_4
* cell instance $11614 r0 *1 76.475,28.91
X$11614 682 VIA_via2_5
* cell instance $11615 r0 *1 79.895,30.03
X$11615 682 VIA_via1_4
* cell instance $11616 r0 *1 80.655,27.65
X$11616 682 VIA_via1_4
* cell instance $11617 r0 *1 80.655,27.65
X$11617 682 VIA_via2_5
* cell instance $11618 r0 *1 77.425,28.21
X$11618 683 VIA_via1_7
* cell instance $11619 r0 *1 77.425,28.21
X$11619 683 VIA_via2_5
* cell instance $11620 r0 *1 78.375,28.21
X$11620 683 VIA_via2_5
* cell instance $11621 r0 *1 78.375,27.23
X$11621 683 VIA_via1_4
* cell instance $11622 r0 *1 24.035,27.37
X$11622 684 VIA_via2_5
* cell instance $11623 r0 *1 24.035,25.97
X$11623 684 VIA_via1_4
* cell instance $11624 r0 *1 25.745,27.37
X$11624 684 VIA_via1_4
* cell instance $11625 r0 *1 25.745,27.37
X$11625 684 VIA_via2_5
* cell instance $11626 r0 *1 25.555,27.23
X$11626 685 VIA_via2_5
* cell instance $11627 r0 *1 26.315,27.23
X$11627 685 VIA_via2_5
* cell instance $11628 r0 *1 25.365,27.23
X$11628 685 VIA_via1_4
* cell instance $11629 r0 *1 25.365,27.23
X$11629 685 VIA_via2_5
* cell instance $11630 r0 *1 26.315,26.25
X$11630 685 VIA_via1_4
* cell instance $11631 r0 *1 25.555,28.77
X$11631 685 VIA_via1_4
* cell instance $11632 r0 *1 30.115,27.65
X$11632 686 VIA_via2_5
* cell instance $11633 r0 *1 27.835,27.65
X$11633 686 VIA_via2_5
* cell instance $11634 r0 *1 27.835,28.77
X$11634 686 VIA_via1_4
* cell instance $11635 r0 *1 30.115,31.57
X$11635 686 VIA_via1_4
* cell instance $11636 r0 *1 30.875,27.65
X$11636 686 VIA_via1_4
* cell instance $11637 r0 *1 30.875,27.65
X$11637 686 VIA_via2_5
* cell instance $11638 r0 *1 55.385,27.23
X$11638 687 VIA_via1_4
* cell instance $11639 r0 *1 55.385,27.09
X$11639 687 VIA_via2_5
* cell instance $11640 r0 *1 60.325,27.09
X$11640 687 VIA_via1_4
* cell instance $11641 r0 *1 60.325,27.09
X$11641 687 VIA_via2_5
* cell instance $11642 r0 *1 35.245,27.23
X$11642 688 VIA_via2_5
* cell instance $11643 r0 *1 37.145,27.23
X$11643 688 VIA_via2_5
* cell instance $11644 r0 *1 35.245,28.77
X$11644 688 VIA_via1_4
* cell instance $11645 r0 *1 35.055,27.23
X$11645 688 VIA_via1_4
* cell instance $11646 r0 *1 35.055,27.23
X$11646 688 VIA_via2_5
* cell instance $11647 r0 *1 37.145,26.25
X$11647 688 VIA_via1_4
* cell instance $11648 r0 *1 51.015,28.21
X$11648 689 VIA_via1_7
* cell instance $11649 r0 *1 51.015,28.21
X$11649 689 VIA_via2_5
* cell instance $11650 r0 *1 49.875,28.21
X$11650 689 VIA_via2_5
* cell instance $11651 r0 *1 49.875,27.23
X$11651 689 VIA_via1_4
* cell instance $11652 r0 *1 38.095,28.63
X$11652 690 VIA_via2_5
* cell instance $11653 r0 *1 41.135,28.63
X$11653 690 VIA_via1_4
* cell instance $11654 r0 *1 41.135,28.63
X$11654 690 VIA_via2_5
* cell instance $11655 r0 *1 37.905,31.57
X$11655 690 VIA_via1_4
* cell instance $11656 r0 *1 37.335,28.77
X$11656 690 VIA_via1_4
* cell instance $11657 r0 *1 37.335,28.63
X$11657 690 VIA_via2_5
* cell instance $11658 r0 *1 7.315,35.91
X$11658 691 VIA_via2_5
* cell instance $11659 r0 *1 5.225,35.91
X$11659 691 VIA_via2_5
* cell instance $11660 r0 *1 7.315,37.17
X$11660 691 VIA_via1_4
* cell instance $11661 r0 *1 5.225,29.05
X$11661 691 VIA_via1_4
* cell instance $11662 r0 *1 4.845,27.23
X$11662 691 VIA_via1_4
* cell instance $11663 r0 *1 8.835,35.63
X$11663 692 VIA_via2_5
* cell instance $11664 r0 *1 9.215,35.63
X$11664 692 VIA_via1_4
* cell instance $11665 r0 *1 9.215,35.63
X$11665 692 VIA_via2_5
* cell instance $11666 r0 *1 8.645,29.05
X$11666 692 VIA_via1_4
* cell instance $11667 r0 *1 9.215,27.23
X$11667 692 VIA_via1_4
* cell instance $11668 r0 *1 9.025,37.17
X$11668 693 VIA_via2_5
* cell instance $11669 r0 *1 26.505,42.91
X$11669 693 VIA_via2_5
* cell instance $11670 r0 *1 9.215,30.17
X$11670 693 VIA_via2_5
* cell instance $11671 r0 *1 45.505,34.37
X$11671 693 VIA_via2_5
* cell instance $11672 r0 *1 43.985,31.57
X$11672 693 VIA_via2_5
* cell instance $11673 r0 *1 25.745,29.47
X$11673 693 VIA_via2_5
* cell instance $11674 r0 *1 21.185,42.91
X$11674 693 VIA_via2_5
* cell instance $11675 r0 *1 8.835,44.03
X$11675 693 VIA_via2_5
* cell instance $11676 r0 *1 36.195,32.55
X$11676 693 VIA_via2_5
* cell instance $11677 r0 *1 26.695,32.55
X$11677 693 VIA_via2_5
* cell instance $11678 r0 *1 25.935,32.55
X$11678 693 VIA_via2_5
* cell instance $11679 r0 *1 21.755,30.17
X$11679 693 VIA_via2_5
* cell instance $11680 r0 *1 21.755,29.47
X$11680 693 VIA_via2_5
* cell instance $11681 r0 *1 22.135,29.47
X$11681 693 VIA_via2_5
* cell instance $11682 r0 *1 46.075,44.03
X$11682 693 VIA_via1_4
* cell instance $11683 r0 *1 7.885,37.17
X$11683 693 VIA_via1_4
* cell instance $11684 r0 *1 7.885,37.17
X$11684 693 VIA_via2_5
* cell instance $11685 r0 *1 9.025,30.03
X$11685 693 VIA_via1_4
* cell instance $11686 r0 *1 8.645,46.83
X$11686 693 VIA_via1_4
* cell instance $11687 r0 *1 22.135,28.77
X$11687 693 VIA_via1_4
* cell instance $11688 r0 *1 26.505,35.63
X$11688 693 VIA_via1_4
* cell instance $11689 r0 *1 25.745,32.55
X$11689 693 VIA_via1_4
* cell instance $11690 r0 *1 25.935,32.83
X$11690 693 VIA_via1_4
* cell instance $11691 r0 *1 43.985,34.37
X$11691 693 VIA_via1_4
* cell instance $11692 r0 *1 43.985,34.37
X$11692 693 VIA_via2_5
* cell instance $11693 r0 *1 36.195,31.57
X$11693 693 VIA_via1_4
* cell instance $11694 r0 *1 36.195,31.57
X$11694 693 VIA_via2_5
* cell instance $11695 r0 *1 32.775,42.77
X$11695 693 VIA_via1_4
* cell instance $11696 r0 *1 32.775,42.91
X$11696 693 VIA_via2_5
* cell instance $11697 r0 *1 21.185,44.03
X$11697 693 VIA_via1_4
* cell instance $11698 r0 *1 21.185,44.03
X$11698 693 VIA_via2_5
* cell instance $11699 r0 *1 14.915,30.31
X$11699 694 VIA_via2_5
* cell instance $11700 r0 *1 15.865,30.31
X$11700 694 VIA_via2_5
* cell instance $11701 r0 *1 14.915,30.03
X$11701 694 VIA_via1_4
* cell instance $11702 r0 *1 13.205,30.31
X$11702 694 VIA_via1_4
* cell instance $11703 r0 *1 13.205,30.31
X$11703 694 VIA_via2_5
* cell instance $11704 r0 *1 15.865,34.37
X$11704 694 VIA_via1_4
* cell instance $11705 r0 *1 14.725,29.05
X$11705 695 VIA_via2_5
* cell instance $11706 r0 *1 16.815,35.07
X$11706 695 VIA_via2_5
* cell instance $11707 r0 *1 15.675,35.07
X$11707 695 VIA_via2_5
* cell instance $11708 r0 *1 15.485,29.05
X$11708 695 VIA_via2_5
* cell instance $11709 r0 *1 16.625,35.63
X$11709 695 VIA_via1_4
* cell instance $11710 r0 *1 14.725,27.23
X$11710 695 VIA_via1_4
* cell instance $11711 r0 *1 17.385,29.05
X$11711 695 VIA_via1_4
* cell instance $11712 r0 *1 17.385,29.05
X$11712 695 VIA_via2_5
* cell instance $11713 r0 *1 21.185,28.77
X$11713 696 VIA_via2_5
* cell instance $11714 r0 *1 21.565,28.77
X$11714 696 VIA_via1_4
* cell instance $11715 r0 *1 21.565,28.77
X$11715 696 VIA_via2_5
* cell instance $11716 r0 *1 20.995,30.03
X$11716 696 VIA_via1_4
* cell instance $11717 r0 *1 20.615,28.77
X$11717 696 VIA_via1_4
* cell instance $11718 r0 *1 20.615,28.77
X$11718 696 VIA_via2_5
* cell instance $11719 r0 *1 22.515,31.85
X$11719 697 VIA_via2_5
* cell instance $11720 r0 *1 22.705,30.03
X$11720 697 VIA_via1_4
* cell instance $11721 r0 *1 25.555,34.37
X$11721 697 VIA_via1_4
* cell instance $11722 r0 *1 24.985,31.85
X$11722 697 VIA_via1_4
* cell instance $11723 r0 *1 24.985,31.85
X$11723 697 VIA_via2_5
* cell instance $11724 r0 *1 25.935,29.19
X$11724 698 VIA_via1_7
* cell instance $11725 r0 *1 25.935,37.17
X$11725 698 VIA_via1_4
* cell instance $11726 r0 *1 34.675,31.85
X$11726 699 VIA_via2_5
* cell instance $11727 r0 *1 36.005,31.85
X$11727 699 VIA_via1_4
* cell instance $11728 r0 *1 36.005,31.85
X$11728 699 VIA_via2_5
* cell instance $11729 r0 *1 34.675,34.37
X$11729 699 VIA_via1_4
* cell instance $11730 r0 *1 34.485,30.03
X$11730 699 VIA_via1_4
* cell instance $11731 r0 *1 35.625,29.19
X$11731 700 VIA_via1_7
* cell instance $11732 r0 *1 35.435,35.63
X$11732 700 VIA_via1_4
* cell instance $11733 r0 *1 46.455,29.19
X$11733 701 VIA_via1_7
* cell instance $11734 r0 *1 46.265,30.03
X$11734 701 VIA_via1_4
* cell instance $11735 r0 *1 52.345,29.19
X$11735 702 VIA_via1_7
* cell instance $11736 r0 *1 52.535,35.63
X$11736 702 VIA_via1_4
* cell instance $11737 r0 *1 68.305,29.75
X$11737 703 VIA_via2_5
* cell instance $11738 r0 *1 69.065,30.03
X$11738 703 VIA_via1_4
* cell instance $11739 r0 *1 69.065,30.03
X$11739 703 VIA_via2_5
* cell instance $11740 r0 *1 68.305,29.05
X$11740 703 VIA_via1_4
* cell instance $11741 r0 *1 67.165,30.03
X$11741 703 VIA_via1_4
* cell instance $11742 r0 *1 67.165,30.03
X$11742 703 VIA_via2_5
* cell instance $11743 r0 *1 72.865,28.77
X$11743 704 VIA_via1_4
* cell instance $11744 r0 *1 72.865,28.77
X$11744 704 VIA_via2_5
* cell instance $11745 r0 *1 68.495,30.03
X$11745 704 VIA_via1_4
* cell instance $11746 r0 *1 68.685,28.77
X$11746 704 VIA_via1_4
* cell instance $11747 r0 *1 68.685,28.77
X$11747 704 VIA_via2_5
* cell instance $11748 r0 *1 71.345,29.47
X$11748 705 VIA_via2_5
* cell instance $11749 r0 *1 70.775,29.47
X$11749 705 VIA_via2_5
* cell instance $11750 r0 *1 71.915,29.47
X$11750 705 VIA_via2_5
* cell instance $11751 r0 *1 65.835,32.83
X$11751 705 VIA_via2_5
* cell instance $11752 r0 *1 70.775,32.83
X$11752 705 VIA_via2_5
* cell instance $11753 r0 *1 70.015,32.83
X$11753 705 VIA_via2_5
* cell instance $11754 r0 *1 73.815,29.47
X$11754 705 VIA_via2_5
* cell instance $11755 r0 *1 73.815,27.23
X$11755 705 VIA_via1_4
* cell instance $11756 r0 *1 71.345,28.77
X$11756 705 VIA_via1_4
* cell instance $11757 r0 *1 71.915,30.03
X$11757 705 VIA_via1_4
* cell instance $11758 r0 *1 65.835,34.37
X$11758 705 VIA_via1_4
* cell instance $11759 r0 *1 65.455,32.83
X$11759 705 VIA_via1_4
* cell instance $11760 r0 *1 65.455,32.83
X$11760 705 VIA_via2_5
* cell instance $11761 r0 *1 70.775,31.57
X$11761 705 VIA_via1_4
* cell instance $11762 r0 *1 71.155,32.83
X$11762 705 VIA_via1_4
* cell instance $11763 r0 *1 71.155,32.83
X$11763 705 VIA_via2_5
* cell instance $11764 r0 *1 69.065,32.83
X$11764 705 VIA_via1_4
* cell instance $11765 r0 *1 69.065,32.83
X$11765 705 VIA_via2_5
* cell instance $11766 r0 *1 70.015,35.63
X$11766 705 VIA_via1_4
* cell instance $11767 r0 *1 74.955,35.63
X$11767 706 VIA_via2_5
* cell instance $11768 r0 *1 75.145,30.31
X$11768 706 VIA_via1_4
* cell instance $11769 r0 *1 72.865,35.63
X$11769 706 VIA_via1_4
* cell instance $11770 r0 *1 72.865,35.63
X$11770 706 VIA_via2_5
* cell instance $11771 r0 *1 83.315,31.01
X$11771 707 VIA_via1_7
* cell instance $11772 r0 *1 83.315,30.31
X$11772 707 VIA_via2_5
* cell instance $11773 r0 *1 74.955,30.03
X$11773 707 VIA_via1_4
* cell instance $11774 r0 *1 74.955,30.03
X$11774 707 VIA_via2_5
* cell instance $11775 r0 *1 79.515,29.61
X$11775 708 VIA_via1_7
* cell instance $11776 r0 *1 78.375,28.77
X$11776 708 VIA_via1_4
* cell instance $11777 r0 *1 78.565,30.03
X$11777 709 VIA_via1_4
* cell instance $11778 r0 *1 78.565,30.03
X$11778 709 VIA_via2_5
* cell instance $11779 r0 *1 80.465,30.03
X$11779 709 VIA_via1_4
* cell instance $11780 r0 *1 80.465,30.03
X$11780 709 VIA_via2_5
* cell instance $11781 r0 *1 80.655,29.05
X$11781 709 VIA_via1_4
* cell instance $11782 r0 *1 87.305,37.17
X$11782 710 VIA_via2_5
* cell instance $11783 r0 *1 83.315,32.83
X$11783 710 VIA_via2_5
* cell instance $11784 r0 *1 84.075,30.31
X$11784 710 VIA_via2_5
* cell instance $11785 r0 *1 85.595,30.31
X$11785 710 VIA_via2_5
* cell instance $11786 r0 *1 75.905,36.89
X$11786 710 VIA_via2_5
* cell instance $11787 r0 *1 79.515,36.89
X$11787 710 VIA_via2_5
* cell instance $11788 r0 *1 79.515,37.45
X$11788 710 VIA_via2_5
* cell instance $11789 r0 *1 83.315,37.17
X$11789 710 VIA_via1_4
* cell instance $11790 r0 *1 83.315,37.17
X$11790 710 VIA_via2_5
* cell instance $11791 r0 *1 80.085,37.17
X$11791 710 VIA_via1_4
* cell instance $11792 r0 *1 80.085,37.31
X$11792 710 VIA_via2_5
* cell instance $11793 r0 *1 75.905,37.17
X$11793 710 VIA_via1_4
* cell instance $11794 r0 *1 83.695,32.83
X$11794 710 VIA_via1_4
* cell instance $11795 r0 *1 83.695,32.83
X$11795 710 VIA_via2_5
* cell instance $11796 r0 *1 78.945,32.83
X$11796 710 VIA_via1_4
* cell instance $11797 r0 *1 84.265,30.03
X$11797 710 VIA_via1_4
* cell instance $11798 r0 *1 85.595,30.03
X$11798 710 VIA_via1_4
* cell instance $11799 r0 *1 88.065,40.95
X$11799 710 VIA_via1_4
* cell instance $11800 r0 *1 87.115,29.75
X$11800 711 VIA_via2_5
* cell instance $11801 r0 *1 87.115,29.05
X$11801 711 VIA_via1_4
* cell instance $11802 r0 *1 82.745,30.03
X$11802 711 VIA_via1_4
* cell instance $11803 r0 *1 82.745,29.89
X$11803 711 VIA_via2_5
* cell instance $11804 r0 *1 84.835,30.03
X$11804 711 VIA_via1_4
* cell instance $11805 r0 *1 84.835,29.89
X$11805 711 VIA_via2_5
* cell instance $11806 r0 *1 89.775,30.03
X$11806 712 VIA_via1_4
* cell instance $11807 r0 *1 89.775,30.03
X$11807 712 VIA_via2_5
* cell instance $11808 r0 *1 86.165,30.03
X$11808 712 VIA_via1_4
* cell instance $11809 r0 *1 86.165,30.03
X$11809 712 VIA_via2_5
* cell instance $11810 r0 *1 83.315,30.03
X$11810 712 VIA_via1_4
* cell instance $11811 r0 *1 83.315,30.03
X$11811 712 VIA_via2_5
* cell instance $11812 r0 *1 93.765,30.45
X$11812 713 VIA_via2_5
* cell instance $11813 r0 *1 93.005,30.45
X$11813 713 VIA_via1_4
* cell instance $11814 r0 *1 93.005,30.45
X$11814 713 VIA_via2_5
* cell instance $11815 r0 *1 93.955,30.03
X$11815 713 VIA_via1_4
* cell instance $11816 r0 *1 93.765,31.57
X$11816 713 VIA_via1_4
* cell instance $11817 r0 *1 95.475,31.57
X$11817 714 VIA_via2_5
* cell instance $11818 r0 *1 95.475,29.05
X$11818 714 VIA_via2_5
* cell instance $11819 r0 *1 95.475,30.03
X$11819 714 VIA_via1_4
* cell instance $11820 r0 *1 96.615,29.05
X$11820 714 VIA_via1_4
* cell instance $11821 r0 *1 96.615,29.05
X$11821 714 VIA_via2_5
* cell instance $11822 r0 *1 94.335,31.57
X$11822 714 VIA_via1_4
* cell instance $11823 r0 *1 94.335,31.57
X$11823 714 VIA_via2_5
* cell instance $11824 r0 *1 5.985,30.03
X$11824 715 VIA_via1_4
* cell instance $11825 r0 *1 5.985,30.03
X$11825 715 VIA_via2_5
* cell instance $11826 r0 *1 5.035,30.03
X$11826 715 VIA_via1_4
* cell instance $11827 r0 *1 5.035,30.03
X$11827 715 VIA_via2_5
* cell instance $11828 r0 *1 95.855,29.61
X$11828 716 VIA_via1_7
* cell instance $11829 r0 *1 95.855,29.61
X$11829 716 VIA_via2_5
* cell instance $11830 r0 *1 94.335,29.61
X$11830 716 VIA_via2_5
* cell instance $11831 r0 *1 94.335,28.77
X$11831 716 VIA_via1_4
* cell instance $11832 r0 *1 94.335,29.89
X$11832 717 VIA_via1_4
* cell instance $11833 r0 *1 94.335,29.89
X$11833 717 VIA_via2_5
* cell instance $11834 r0 *1 90.725,30.03
X$11834 717 VIA_via1_4
* cell instance $11835 r0 *1 90.725,29.89
X$11835 717 VIA_via2_5
* cell instance $11836 r0 *1 10.925,30.03
X$11836 718 VIA_via1_4
* cell instance $11837 r0 *1 10.925,29.89
X$11837 718 VIA_via2_5
* cell instance $11838 r0 *1 15.295,29.89
X$11838 718 VIA_via1_4
* cell instance $11839 r0 *1 15.295,29.89
X$11839 718 VIA_via2_5
* cell instance $11840 r0 *1 15.105,27.79
X$11840 719 VIA_via1_7
* cell instance $11841 r0 *1 15.105,28.77
X$11841 719 VIA_via1_4
* cell instance $11842 r0 *1 18.335,28.77
X$11842 720 VIA_via1_4
* cell instance $11843 r0 *1 18.335,28.91
X$11843 720 VIA_via2_5
* cell instance $11844 r0 *1 21.945,28.91
X$11844 720 VIA_via1_4
* cell instance $11845 r0 *1 21.945,28.91
X$11845 720 VIA_via2_5
* cell instance $11846 r0 *1 86.545,30.03
X$11846 721 VIA_via1_4
* cell instance $11847 r0 *1 87.495,30.03
X$11847 721 VIA_via1_4
* cell instance $11848 r0 *1 85.215,29.61
X$11848 722 VIA_via1_7
* cell instance $11849 r0 *1 85.215,29.61
X$11849 722 VIA_via2_5
* cell instance $11850 r0 *1 84.835,29.61
X$11850 722 VIA_via2_5
* cell instance $11851 r0 *1 84.835,28.77
X$11851 722 VIA_via1_4
* cell instance $11852 r0 *1 29.925,29.19
X$11852 723 VIA_via1_7
* cell instance $11853 r0 *1 29.925,30.03
X$11853 723 VIA_via1_4
* cell instance $11854 r0 *1 84.455,67.83
X$11854 724 VIA_via1_7
* cell instance $11855 r0 *1 66.785,31.43
X$11855 724 VIA_via1_7
* cell instance $11856 r0 *1 66.975,62.23
X$11856 724 VIA_via1_7
* cell instance $11857 r0 *1 66.975,62.23
X$11857 724 VIA_via2_5
* cell instance $11858 r0 *1 43.035,62.23
X$11858 724 VIA_via1_7
* cell instance $11859 r0 *1 43.035,62.23
X$11859 724 VIA_via2_5
* cell instance $11860 r0 *1 53.675,88.69
X$11860 724 VIA_via2_5
* cell instance $11861 r0 *1 84.455,62.51
X$11861 724 VIA_via2_5
* cell instance $11862 r0 *1 84.375,62.51
X$11862 724 VIA_via3_2
* cell instance $11863 r0 *1 66.785,30.59
X$11863 724 VIA_via2_5
* cell instance $11864 r0 *1 85.405,29.47
X$11864 724 VIA_via2_5
* cell instance $11865 r0 *1 82.175,39.97
X$11865 724 VIA_via1_4
* cell instance $11866 r0 *1 82.175,39.97
X$11866 724 VIA_via2_5
* cell instance $11867 r0 *1 82.135,39.97
X$11867 724 VIA_via3_2
* cell instance $11868 r0 *1 85.405,25.97
X$11868 724 VIA_via1_4
* cell instance $11869 r0 *1 53.675,86.03
X$11869 724 VIA_via1_4
* cell instance $11870 r0 *1 53.675,90.37
X$11870 724 VIA_via1_4
* cell instance $11871 r0 *1 42.465,88.83
X$11871 724 VIA_via1_4
* cell instance $11872 r0 *1 42.465,88.69
X$11872 724 VIA_via2_5
* cell instance $11873 r0 *1 84.835,62.37
X$11873 724 VIA_via1_4
* cell instance $11874 r0 *1 84.835,62.51
X$11874 724 VIA_via2_5
* cell instance $11875 r0 *1 43.605,30.45
X$11875 724 VIA_via1_4
* cell instance $11876 r0 *1 43.605,30.45
X$11876 724 VIA_via2_5
* cell instance $11877 r0 *1 67.295,61.95
X$11877 724 VIA_via4_0
* cell instance $11878 r0 *1 43.775,61.95
X$11878 724 VIA_via4_0
* cell instance $11879 r0 *1 84.375,61.95
X$11879 724 VIA_via4_0
* cell instance $11880 r0 *1 43.775,30.45
X$11880 724 VIA_via3_2
* cell instance $11881 r0 *1 43.775,62.23
X$11881 724 VIA_via3_2
* cell instance $11882 r0 *1 67.295,62.23
X$11882 724 VIA_via3_2
* cell instance $11883 r0 *1 82.135,30.59
X$11883 724 VIA_via3_2
* cell instance $11884 r0 *1 43.775,88.69
X$11884 724 VIA_via3_2
* cell instance $11885 r0 *1 82.135,29.47
X$11885 724 VIA_via3_2
* cell instance $11886 r0 *1 34.105,28.77
X$11886 725 VIA_via2_5
* cell instance $11887 r0 *1 34.675,28.77
X$11887 725 VIA_via1_4
* cell instance $11888 r0 *1 34.675,28.77
X$11888 725 VIA_via2_5
* cell instance $11889 r0 *1 31.825,28.77
X$11889 725 VIA_via1_4
* cell instance $11890 r0 *1 31.825,28.77
X$11890 725 VIA_via2_5
* cell instance $11891 r0 *1 34.105,27.65
X$11891 725 VIA_via1_4
* cell instance $11892 r0 *1 38.855,28.77
X$11892 726 VIA_via1_4
* cell instance $11893 r0 *1 38.855,28.77
X$11893 726 VIA_via2_5
* cell instance $11894 r0 *1 37.715,28.77
X$11894 726 VIA_via1_4
* cell instance $11895 r0 *1 37.715,28.77
X$11895 726 VIA_via2_5
* cell instance $11896 r0 *1 41.515,30.03
X$11896 727 VIA_via1_4
* cell instance $11897 r0 *1 41.515,30.03
X$11897 727 VIA_via2_5
* cell instance $11898 r0 *1 37.905,30.03
X$11898 727 VIA_via1_4
* cell instance $11899 r0 *1 37.905,30.03
X$11899 727 VIA_via2_5
* cell instance $11900 r0 *1 74.765,29.89
X$11900 728 VIA_via1_4
* cell instance $11901 r0 *1 74.765,29.89
X$11901 728 VIA_via2_5
* cell instance $11902 r0 *1 71.155,30.03
X$11902 728 VIA_via1_4
* cell instance $11903 r0 *1 71.155,29.89
X$11903 728 VIA_via2_5
* cell instance $11904 r0 *1 53.675,29.19
X$11904 729 VIA_via1_7
* cell instance $11905 r0 *1 53.675,29.33
X$11905 729 VIA_via2_5
* cell instance $11906 r0 *1 52.535,29.33
X$11906 729 VIA_via2_5
* cell instance $11907 r0 *1 52.535,30.03
X$11907 729 VIA_via1_4
* cell instance $11908 r0 *1 69.635,28.77
X$11908 730 VIA_via1_4
* cell instance $11909 r0 *1 70.585,28.77
X$11909 730 VIA_via1_4
* cell instance $11910 r0 *1 68.115,29.61
X$11910 731 VIA_via1_7
* cell instance $11911 r0 *1 68.115,29.61
X$11911 731 VIA_via2_5
* cell instance $11912 r0 *1 66.025,29.61
X$11912 731 VIA_via2_5
* cell instance $11913 r0 *1 66.025,28.77
X$11913 731 VIA_via1_4
* cell instance $11914 r0 *1 4.655,30.45
X$11914 732 VIA_via2_5
* cell instance $11915 r0 *1 7.695,30.45
X$11915 732 VIA_via2_5
* cell instance $11916 r0 *1 7.695,35.63
X$11916 732 VIA_via1_4
* cell instance $11917 r0 *1 8.265,30.45
X$11917 732 VIA_via1_4
* cell instance $11918 r0 *1 8.265,30.45
X$11918 732 VIA_via2_5
* cell instance $11919 r0 *1 4.655,30.03
X$11919 732 VIA_via1_4
* cell instance $11920 r0 *1 18.525,31.85
X$11920 733 VIA_via2_5
* cell instance $11921 r0 *1 16.625,31.85
X$11921 733 VIA_via2_5
* cell instance $11922 r0 *1 18.715,31.85
X$11922 733 VIA_via1_4
* cell instance $11923 r0 *1 18.715,31.85
X$11923 733 VIA_via2_5
* cell instance $11924 r0 *1 18.525,34.37
X$11924 733 VIA_via1_4
* cell instance $11925 r0 *1 16.435,30.03
X$11925 733 VIA_via1_4
* cell instance $11926 r0 *1 23.085,30.59
X$11926 734 VIA_via1_7
* cell instance $11927 r0 *1 22.705,31.57
X$11927 734 VIA_via1_4
* cell instance $11928 r0 *1 29.545,30.45
X$11928 735 VIA_via2_5
* cell instance $11929 r0 *1 31.635,30.45
X$11929 735 VIA_via2_5
* cell instance $11930 r0 *1 31.635,34.37
X$11930 735 VIA_via1_4
* cell instance $11931 r0 *1 29.545,28.77
X$11931 735 VIA_via1_4
* cell instance $11932 r0 *1 32.205,30.45
X$11932 735 VIA_via1_4
* cell instance $11933 r0 *1 32.205,30.45
X$11933 735 VIA_via2_5
* cell instance $11934 r0 *1 40.375,31.85
X$11934 736 VIA_via2_5
* cell instance $11935 r0 *1 38.475,31.85
X$11935 736 VIA_via2_5
* cell instance $11936 r0 *1 38.475,31.57
X$11936 736 VIA_via1_4
* cell instance $11937 r0 *1 41.135,30.03
X$11937 736 VIA_via1_4
* cell instance $11938 r0 *1 40.185,30.45
X$11938 736 VIA_via1_4
* cell instance $11939 r0 *1 47.785,31.57
X$11939 737 VIA_via2_5
* cell instance $11940 r0 *1 45.315,31.57
X$11940 737 VIA_via2_5
* cell instance $11941 r0 *1 47.025,31.57
X$11941 737 VIA_via1_4
* cell instance $11942 r0 *1 47.025,31.57
X$11942 737 VIA_via2_5
* cell instance $11943 r0 *1 47.785,32.83
X$11943 737 VIA_via1_4
* cell instance $11944 r0 *1 45.505,30.03
X$11944 737 VIA_via1_4
* cell instance $11945 r0 *1 50.635,31.85
X$11945 738 VIA_via2_5
* cell instance $11946 r0 *1 52.155,31.85
X$11946 738 VIA_via2_5
* cell instance $11947 r0 *1 50.635,30.03
X$11947 738 VIA_via1_4
* cell instance $11948 r0 *1 52.155,34.37
X$11948 738 VIA_via1_4
* cell instance $11949 r0 *1 52.345,31.85
X$11949 738 VIA_via1_4
* cell instance $11950 r0 *1 67.355,33.95
X$11950 739 VIA_via1_4
* cell instance $11951 r0 *1 66.975,31.57
X$11951 739 VIA_via1_4
* cell instance $11952 r0 *1 67.735,34.37
X$11952 739 VIA_via1_4
* cell instance $11953 r0 *1 66.975,32.69
X$11953 740 VIA_via1_4
* cell instance $11954 r0 *1 66.975,32.69
X$11954 740 VIA_via2_5
* cell instance $11955 r0 *1 67.545,31.57
X$11955 740 VIA_via1_4
* cell instance $11956 r0 *1 67.735,32.83
X$11956 740 VIA_via1_4
* cell instance $11957 r0 *1 67.735,32.69
X$11957 740 VIA_via2_5
* cell instance $11958 r0 *1 69.445,30.59
X$11958 741 VIA_via1_7
* cell instance $11959 r0 *1 72.865,31.85
X$11959 741 VIA_via2_5
* cell instance $11960 r0 *1 69.635,31.85
X$11960 741 VIA_via2_5
* cell instance $11961 r0 *1 72.865,32.83
X$11961 741 VIA_via1_4
* cell instance $11962 r0 *1 72.485,31.57
X$11962 742 VIA_via1_4
* cell instance $11963 r0 *1 72.485,31.57
X$11963 742 VIA_via2_5
* cell instance $11964 r0 *1 72.675,32.55
X$11964 742 VIA_via1_4
* cell instance $11965 r0 *1 71.155,31.57
X$11965 742 VIA_via1_4
* cell instance $11966 r0 *1 71.155,31.57
X$11966 742 VIA_via2_5
* cell instance $11967 r0 *1 73.815,30.03
X$11967 743 VIA_via1_4
* cell instance $11968 r0 *1 73.435,30.45
X$11968 743 VIA_via1_4
* cell instance $11969 r0 *1 73.055,31.57
X$11969 743 VIA_via1_4
* cell instance $11970 r0 *1 69.825,33.53
X$11970 744 VIA_via2_5
* cell instance $11971 r0 *1 68.495,33.53
X$11971 744 VIA_via2_5
* cell instance $11972 r0 *1 56.335,37.17
X$11972 744 VIA_via2_5
* cell instance $11973 r0 *1 74.005,33.53
X$11973 744 VIA_via2_5
* cell instance $11974 r0 *1 74.385,31.57
X$11974 744 VIA_via2_5
* cell instance $11975 r0 *1 92.245,33.11
X$11975 744 VIA_via2_5
* cell instance $11976 r0 *1 68.115,46.83
X$11976 744 VIA_via2_5
* cell instance $11977 r0 *1 83.695,38.57
X$11977 744 VIA_via2_5
* cell instance $11978 r0 *1 83.885,42.63
X$11978 744 VIA_via2_5
* cell instance $11979 r0 *1 83.125,33.11
X$11979 744 VIA_via2_5
* cell instance $11980 r0 *1 83.125,31.57
X$11980 744 VIA_via2_5
* cell instance $11981 r0 *1 83.695,33.11
X$11981 744 VIA_via2_5
* cell instance $11982 r0 *1 56.335,33.53
X$11982 744 VIA_via2_5
* cell instance $11983 r0 *1 55.575,33.53
X$11983 744 VIA_via2_5
* cell instance $11984 r0 *1 52.725,37.17
X$11984 744 VIA_via1_4
* cell instance $11985 r0 *1 52.725,37.17
X$11985 744 VIA_via2_5
* cell instance $11986 r0 *1 77.425,38.43
X$11986 744 VIA_via1_4
* cell instance $11987 r0 *1 77.425,38.43
X$11987 744 VIA_via2_5
* cell instance $11988 r0 *1 83.695,45.57
X$11988 744 VIA_via1_4
* cell instance $11989 r0 *1 68.305,42.77
X$11989 744 VIA_via1_4
* cell instance $11990 r0 *1 92.435,42.77
X$11990 744 VIA_via1_4
* cell instance $11991 r0 *1 92.435,42.63
X$11991 744 VIA_via2_5
* cell instance $11992 r0 *1 83.125,28.77
X$11992 744 VIA_via1_4
* cell instance $11993 r0 *1 74.005,32.83
X$11993 744 VIA_via1_4
* cell instance $11994 r0 *1 74.385,31.85
X$11994 744 VIA_via1_4
* cell instance $11995 r0 *1 92.245,31.57
X$11995 744 VIA_via1_4
* cell instance $11996 r0 *1 58.425,46.83
X$11996 744 VIA_via1_4
* cell instance $11997 r0 *1 58.425,46.83
X$11997 744 VIA_via2_5
* cell instance $11998 r0 *1 55.575,30.03
X$11998 744 VIA_via1_4
* cell instance $11999 r0 *1 70.015,31.57
X$11999 744 VIA_via1_4
* cell instance $12000 r0 *1 86.735,32.55
X$12000 745 VIA_via2_5
* cell instance $12001 r0 *1 84.265,32.55
X$12001 745 VIA_via2_5
* cell instance $12002 r0 *1 82.745,32.41
X$12002 745 VIA_via2_5
* cell instance $12003 r0 *1 82.935,31.57
X$12003 745 VIA_via1_4
* cell instance $12004 r0 *1 84.265,32.83
X$12004 745 VIA_via1_4
* cell instance $12005 r0 *1 86.735,31.85
X$12005 745 VIA_via1_4
* cell instance $12006 r0 *1 84.645,32.41
X$12006 746 VIA_via1_7
* cell instance $12007 r0 *1 84.455,31.57
X$12007 746 VIA_via1_4
* cell instance $12008 r0 *1 69.825,31.01
X$12008 747 VIA_via1_7
* cell instance $12009 r0 *1 69.825,31.01
X$12009 747 VIA_via2_5
* cell instance $12010 r0 *1 90.915,31.57
X$12010 747 VIA_via1_4
* cell instance $12011 r0 *1 90.915,31.57
X$12011 747 VIA_via2_5
* cell instance $12012 r0 *1 91.105,31.71
X$12012 748 VIA_via1_4
* cell instance $12013 r0 *1 91.105,31.71
X$12013 748 VIA_via2_5
* cell instance $12014 r0 *1 89.775,56.77
X$12014 748 VIA_via1_4
* cell instance $12015 r0 *1 89.775,56.63
X$12015 748 VIA_via2_5
* cell instance $12016 r0 *1 90.725,56.77
X$12016 748 VIA_via1_4
* cell instance $12017 r0 *1 90.725,56.63
X$12017 748 VIA_via2_5
* cell instance $12018 r0 *1 91.375,31.71
X$12018 748 VIA_via3_2
* cell instance $12019 r0 *1 91.375,56.49
X$12019 748 VIA_via3_2
* cell instance $12020 r0 *1 16.815,30.59
X$12020 749 VIA_via1_7
* cell instance $12021 r0 *1 16.815,31.71
X$12021 749 VIA_via2_5
* cell instance $12022 r0 *1 16.435,31.57
X$12022 749 VIA_via1_4
* cell instance $12023 r0 *1 16.435,31.71
X$12023 749 VIA_via2_5
* cell instance $12024 r0 *1 29.545,31.57
X$12024 750 VIA_via1_4
* cell instance $12025 r0 *1 29.545,31.57
X$12025 750 VIA_via2_5
* cell instance $12026 r0 *1 29.925,32.55
X$12026 750 VIA_via1_4
* cell instance $12027 r0 *1 28.595,31.57
X$12027 750 VIA_via1_4
* cell instance $12028 r0 *1 28.595,31.57
X$12028 750 VIA_via2_5
* cell instance $12029 r0 *1 83.695,30.59
X$12029 751 VIA_via1_7
* cell instance $12030 r0 *1 82.935,34.37
X$12030 751 VIA_via2_5
* cell instance $12031 r0 *1 82.935,31.85
X$12031 751 VIA_via2_5
* cell instance $12032 r0 *1 83.695,31.85
X$12032 751 VIA_via2_5
* cell instance $12033 r0 *1 77.995,34.37
X$12033 751 VIA_via1_4
* cell instance $12034 r0 *1 77.995,34.37
X$12034 751 VIA_via2_5
* cell instance $12035 r0 *1 34.865,30.59
X$12035 752 VIA_via1_7
* cell instance $12036 r0 *1 34.865,30.59
X$12036 752 VIA_via2_5
* cell instance $12037 r0 *1 33.725,30.59
X$12037 752 VIA_via2_5
* cell instance $12038 r0 *1 33.725,31.57
X$12038 752 VIA_via1_4
* cell instance $12039 r0 *1 82.365,32.55
X$12039 753 VIA_via2_5
* cell instance $12040 r0 *1 82.365,31.57
X$12040 753 VIA_via1_4
* cell instance $12041 r0 *1 82.365,31.71
X$12041 753 VIA_via2_5
* cell instance $12042 r0 *1 83.315,32.55
X$12042 753 VIA_via1_4
* cell instance $12043 r0 *1 83.315,32.55
X$12043 753 VIA_via2_5
* cell instance $12044 r0 *1 81.225,31.57
X$12044 753 VIA_via1_4
* cell instance $12045 r0 *1 81.225,31.71
X$12045 753 VIA_via2_5
* cell instance $12046 r0 *1 77.235,31.85
X$12046 754 VIA_via2_5
* cell instance $12047 r0 *1 77.235,32.83
X$12047 754 VIA_via1_4
* cell instance $12048 r0 *1 78.375,31.85
X$12048 754 VIA_via1_4
* cell instance $12049 r0 *1 78.375,31.85
X$12049 754 VIA_via2_5
* cell instance $12050 r0 *1 77.235,30.03
X$12050 754 VIA_via1_4
* cell instance $12051 r0 *1 78.185,30.59
X$12051 755 VIA_via1_7
* cell instance $12052 r0 *1 78.185,31.71
X$12052 755 VIA_via2_5
* cell instance $12053 r0 *1 76.095,31.57
X$12053 755 VIA_via1_4
* cell instance $12054 r0 *1 76.095,31.71
X$12054 755 VIA_via2_5
* cell instance $12055 r0 *1 45.885,30.59
X$12055 756 VIA_via1_7
* cell instance $12056 r0 *1 45.885,30.59
X$12056 756 VIA_via2_5
* cell instance $12057 r0 *1 44.745,30.59
X$12057 756 VIA_via2_5
* cell instance $12058 r0 *1 44.745,31.57
X$12058 756 VIA_via1_4
* cell instance $12059 r0 *1 51.015,30.59
X$12059 757 VIA_via1_7
* cell instance $12060 r0 *1 51.015,31.57
X$12060 757 VIA_via2_5
* cell instance $12061 r0 *1 50.065,31.57
X$12061 757 VIA_via1_4
* cell instance $12062 r0 *1 50.065,31.57
X$12062 757 VIA_via2_5
* cell instance $12063 r0 *1 70.395,31.71
X$12063 758 VIA_via2_5
* cell instance $12064 r0 *1 72.105,31.71
X$12064 758 VIA_via2_5
* cell instance $12065 r0 *1 72.105,31.43
X$12065 758 VIA_via1_4
* cell instance $12066 r0 *1 70.395,32.83
X$12066 758 VIA_via1_4
* cell instance $12067 r0 *1 57.855,32.41
X$12067 759 VIA_via1_7
* cell instance $12068 r0 *1 57.855,31.57
X$12068 759 VIA_via2_5
* cell instance $12069 r0 *1 55.195,31.57
X$12069 759 VIA_via1_4
* cell instance $12070 r0 *1 55.195,31.57
X$12070 759 VIA_via2_5
* cell instance $12071 r0 *1 69.445,31.57
X$12071 760 VIA_via1_4
* cell instance $12072 r0 *1 69.445,31.57
X$12072 760 VIA_via2_5
* cell instance $12073 r0 *1 67.925,31.57
X$12073 760 VIA_via1_4
* cell instance $12074 r0 *1 67.925,31.57
X$12074 760 VIA_via2_5
* cell instance $12075 r0 *1 62.415,32.41
X$12075 761 VIA_via1_7
* cell instance $12076 r0 *1 62.415,31.57
X$12076 761 VIA_via2_5
* cell instance $12077 r0 *1 60.325,31.57
X$12077 761 VIA_via1_4
* cell instance $12078 r0 *1 60.325,31.57
X$12078 761 VIA_via2_5
* cell instance $12079 r0 *1 23.465,34.23
X$12079 762 VIA_via1_7
* cell instance $12080 r0 *1 23.465,34.09
X$12080 762 VIA_via2_5
* cell instance $12081 r0 *1 32.395,34.23
X$12081 762 VIA_via1_7
* cell instance $12082 r0 *1 32.395,34.09
X$12082 762 VIA_via2_5
* cell instance $12083 r0 *1 26.315,34.23
X$12083 762 VIA_via1_7
* cell instance $12084 r0 *1 26.315,34.09
X$12084 762 VIA_via2_5
* cell instance $12085 r0 *1 42.465,32.97
X$12085 762 VIA_via1_7
* cell instance $12086 r0 *1 4.275,32.83
X$12086 762 VIA_via2_5
* cell instance $12087 r0 *1 48.355,35.63
X$12087 762 VIA_via2_5
* cell instance $12088 r0 *1 42.465,34.09
X$12088 762 VIA_via2_5
* cell instance $12089 r0 *1 42.465,34.51
X$12089 762 VIA_via2_5
* cell instance $12090 r0 *1 36.195,34.09
X$12090 762 VIA_via2_5
* cell instance $12091 r0 *1 49.305,35.63
X$12091 762 VIA_via2_5
* cell instance $12092 r0 *1 23.275,33.11
X$12092 762 VIA_via2_5
* cell instance $12093 r0 *1 49.305,36.75
X$12093 762 VIA_via1_4
* cell instance $12094 r0 *1 4.085,35.63
X$12094 762 VIA_via1_4
* cell instance $12095 r0 *1 8.835,32.83
X$12095 762 VIA_via1_4
* cell instance $12096 r0 *1 8.835,32.83
X$12096 762 VIA_via2_5
* cell instance $12097 r0 *1 3.705,32.83
X$12097 762 VIA_via1_4
* cell instance $12098 r0 *1 3.705,32.83
X$12098 762 VIA_via2_5
* cell instance $12099 r0 *1 5.985,32.83
X$12099 762 VIA_via1_4
* cell instance $12100 r0 *1 5.985,32.83
X$12100 762 VIA_via2_5
* cell instance $12101 r0 *1 48.165,34.37
X$12101 762 VIA_via1_4
* cell instance $12102 r0 *1 48.165,34.51
X$12102 762 VIA_via2_5
* cell instance $12103 r0 *1 36.385,35.63
X$12103 762 VIA_via1_4
* cell instance $12104 r0 *1 27.265,35.21
X$12104 763 VIA_via1_7
* cell instance $12105 r0 *1 29.165,33.53
X$12105 763 VIA_via2_5
* cell instance $12106 r0 *1 30.305,32.83
X$12106 763 VIA_via2_5
* cell instance $12107 r0 *1 30.305,33.53
X$12107 763 VIA_via2_5
* cell instance $12108 r0 *1 28.405,33.53
X$12108 763 VIA_via2_5
* cell instance $12109 r0 *1 27.265,33.53
X$12109 763 VIA_via2_5
* cell instance $12110 r0 *1 22.515,33.53
X$12110 763 VIA_via2_5
* cell instance $12111 r0 *1 23.085,33.53
X$12111 763 VIA_via2_5
* cell instance $12112 r0 *1 22.895,37.17
X$12112 763 VIA_via1_4
* cell instance $12113 r0 *1 22.515,35.63
X$12113 763 VIA_via1_4
* cell instance $12114 r0 *1 23.465,31.57
X$12114 763 VIA_via1_4
* cell instance $12115 r0 *1 23.085,32.83
X$12115 763 VIA_via1_4
* cell instance $12116 r0 *1 28.405,32.83
X$12116 763 VIA_via1_4
* cell instance $12117 r0 *1 31.825,32.83
X$12117 763 VIA_via1_4
* cell instance $12118 r0 *1 31.825,32.83
X$12118 763 VIA_via2_5
* cell instance $12119 r0 *1 29.165,34.37
X$12119 763 VIA_via1_4
* cell instance $12120 r0 *1 27.455,35.63
X$12120 763 VIA_via1_4
* cell instance $12121 r0 *1 30.305,37.17
X$12121 763 VIA_via1_4
* cell instance $12122 r0 *1 24.225,34.37
X$12122 764 VIA_via1_4
* cell instance $12123 r0 *1 24.605,33.25
X$12123 764 VIA_via1_4
* cell instance $12124 r0 *1 24.985,34.37
X$12124 764 VIA_via1_4
* cell instance $12125 r0 *1 28.975,31.99
X$12125 765 VIA_via1_7
* cell instance $12126 r0 *1 27.645,32.83
X$12126 765 VIA_via1_4
* cell instance $12127 r0 *1 33.535,33.81
X$12127 766 VIA_via1_7
* cell instance $12128 r0 *1 33.535,33.67
X$12128 766 VIA_via2_5
* cell instance $12129 r0 *1 31.065,33.39
X$12129 766 VIA_via2_5
* cell instance $12130 r0 *1 31.065,32.83
X$12130 766 VIA_via1_4
* cell instance $12131 r0 *1 33.345,33.25
X$12131 767 VIA_via1_4
* cell instance $12132 r0 *1 34.105,34.37
X$12132 767 VIA_via1_4
* cell instance $12133 r0 *1 34.105,34.37
X$12133 767 VIA_via2_5
* cell instance $12134 r0 *1 33.155,34.37
X$12134 767 VIA_via1_4
* cell instance $12135 r0 *1 33.155,34.37
X$12135 767 VIA_via2_5
* cell instance $12136 r0 *1 38.475,32.55
X$12136 768 VIA_via2_5
* cell instance $12137 r0 *1 39.805,32.55
X$12137 768 VIA_via2_5
* cell instance $12138 r0 *1 38.475,35.63
X$12138 768 VIA_via1_4
* cell instance $12139 r0 *1 39.805,31.57
X$12139 768 VIA_via1_4
* cell instance $12140 r0 *1 41.515,32.55
X$12140 768 VIA_via1_4
* cell instance $12141 r0 *1 41.515,32.55
X$12141 768 VIA_via2_5
* cell instance $12142 r0 *1 46.835,32.97
X$12142 769 VIA_via1_4
* cell instance $12143 r0 *1 46.835,32.97
X$12143 769 VIA_via2_5
* cell instance $12144 r0 *1 43.225,32.83
X$12144 769 VIA_via1_4
* cell instance $12145 r0 *1 43.225,32.97
X$12145 769 VIA_via2_5
* cell instance $12146 r0 *1 47.215,32.83
X$12146 769 VIA_via1_4
* cell instance $12147 r0 *1 47.215,32.97
X$12147 769 VIA_via2_5
* cell instance $12148 r0 *1 48.165,33.39
X$12148 770 VIA_via1_7
* cell instance $12149 r0 *1 47.975,37.17
X$12149 770 VIA_via1_4
* cell instance $12150 r0 *1 63.745,81.55
X$12150 771 VIA_via1_7
* cell instance $12151 r0 *1 74.765,80.85
X$12151 771 VIA_via2_5
* cell instance $12152 r0 *1 63.745,80.99
X$12152 771 VIA_via2_5
* cell instance $12153 r0 *1 63.745,80.29
X$12153 771 VIA_via2_5
* cell instance $12154 r0 *1 68.875,33.11
X$12154 771 VIA_via2_5
* cell instance $12155 r0 *1 52.535,32.69
X$12155 771 VIA_via2_5
* cell instance $12156 r0 *1 56.715,32.83
X$12156 771 VIA_via1_4
* cell instance $12157 r0 *1 56.715,32.69
X$12157 771 VIA_via2_5
* cell instance $12158 r0 *1 74.765,83.23
X$12158 771 VIA_via1_4
* cell instance $12159 r0 *1 57.095,80.43
X$12159 771 VIA_via1_4
* cell instance $12160 r0 *1 57.095,80.29
X$12160 771 VIA_via2_5
* cell instance $12161 r0 *1 58.805,32.83
X$12161 771 VIA_via1_4
* cell instance $12162 r0 *1 58.805,32.69
X$12162 771 VIA_via2_5
* cell instance $12163 r0 *1 58.805,32.97
X$12163 771 VIA_via2_5
* cell instance $12164 r0 *1 52.535,31.57
X$12164 771 VIA_via1_4
* cell instance $12165 r0 *1 68.875,34.37
X$12165 771 VIA_via1_4
* cell instance $12166 r0 *1 57.775,80.29
X$12166 771 VIA_via3_2
* cell instance $12167 r0 *1 58.055,32.69
X$12167 771 VIA_via3_2
* cell instance $12168 r0 *1 57.855,34.37
X$12168 772 VIA_via2_5
* cell instance $12169 r0 *1 57.475,32.83
X$12169 772 VIA_via1_4
* cell instance $12170 r0 *1 57.475,31.85
X$12170 772 VIA_via1_4
* cell instance $12171 r0 *1 56.145,34.37
X$12171 772 VIA_via1_4
* cell instance $12172 r0 *1 56.145,34.37
X$12172 772 VIA_via2_5
* cell instance $12173 r0 *1 62.035,33.39
X$12173 773 VIA_via2_5
* cell instance $12174 r0 *1 60.895,32.83
X$12174 773 VIA_via2_5
* cell instance $12175 r0 *1 61.085,33.39
X$12175 773 VIA_via2_5
* cell instance $12176 r0 *1 59.565,32.83
X$12176 773 VIA_via1_4
* cell instance $12177 r0 *1 59.565,32.83
X$12177 773 VIA_via2_5
* cell instance $12178 r0 *1 61.085,33.95
X$12178 773 VIA_via1_4
* cell instance $12179 r0 *1 62.035,34.37
X$12179 773 VIA_via1_4
* cell instance $12180 r0 *1 61.655,32.83
X$12180 774 VIA_via2_5
* cell instance $12181 r0 *1 62.605,31.85
X$12181 774 VIA_via1_4
* cell instance $12182 r0 *1 61.465,34.37
X$12182 774 VIA_via1_4
* cell instance $12183 r0 *1 62.035,32.83
X$12183 774 VIA_via1_4
* cell instance $12184 r0 *1 62.035,32.83
X$12184 774 VIA_via2_5
* cell instance $12185 r0 *1 81.605,31.99
X$12185 775 VIA_via1_7
* cell instance $12186 r0 *1 81.035,32.83
X$12186 775 VIA_via1_4
* cell instance $12187 r0 *1 90.535,32.83
X$12187 776 VIA_via2_5
* cell instance $12188 r0 *1 85.785,32.83
X$12188 776 VIA_via1_4
* cell instance $12189 r0 *1 85.785,32.83
X$12189 776 VIA_via2_5
* cell instance $12190 r0 *1 89.965,32.83
X$12190 776 VIA_via1_4
* cell instance $12191 r0 *1 89.965,32.83
X$12191 776 VIA_via2_5
* cell instance $12192 r0 *1 90.535,34.37
X$12192 776 VIA_via1_4
* cell instance $12193 r0 *1 90.915,32.41
X$12193 777 VIA_via1_7
* cell instance $12194 r0 *1 90.725,31.57
X$12194 777 VIA_via1_4
* cell instance $12195 r0 *1 94.715,32.83
X$12195 778 VIA_via2_5
* cell instance $12196 r0 *1 92.435,32.83
X$12196 778 VIA_via1_4
* cell instance $12197 r0 *1 92.435,32.83
X$12197 778 VIA_via2_5
* cell instance $12198 r0 *1 94.715,31.43
X$12198 778 VIA_via1_4
* cell instance $12199 r0 *1 92.625,32.41
X$12199 779 VIA_via1_7
* cell instance $12200 r0 *1 92.625,32.41
X$12200 779 VIA_via2_5
* cell instance $12201 r0 *1 91.675,32.41
X$12201 779 VIA_via2_5
* cell instance $12202 r0 *1 91.675,31.57
X$12202 779 VIA_via1_4
* cell instance $12203 r0 *1 87.685,32.83
X$12203 780 VIA_via1_4
* cell instance $12204 r0 *1 86.735,32.83
X$12204 780 VIA_via1_4
* cell instance $12205 r0 *1 17.575,33.81
X$12205 781 VIA_via1_7
* cell instance $12206 r0 *1 17.575,32.83
X$12206 781 VIA_via2_5
* cell instance $12207 r0 *1 15.485,32.83
X$12207 781 VIA_via1_4
* cell instance $12208 r0 *1 15.485,32.83
X$12208 781 VIA_via2_5
* cell instance $12209 r0 *1 24.605,33.81
X$12209 782 VIA_via1_7
* cell instance $12210 r0 *1 24.795,33.25
X$12210 782 VIA_via2_5
* cell instance $12211 r0 *1 22.325,33.25
X$12211 782 VIA_via2_5
* cell instance $12212 r0 *1 22.325,32.83
X$12212 782 VIA_via1_4
* cell instance $12213 r0 *1 80.845,30.59
X$12213 783 VIA_via1_7
* cell instance $12214 r0 *1 80.845,32.83
X$12214 783 VIA_via2_5
* cell instance $12215 r0 *1 79.705,32.83
X$12215 783 VIA_via1_4
* cell instance $12216 r0 *1 79.705,32.83
X$12216 783 VIA_via2_5
* cell instance $12217 r0 *1 77.805,33.95
X$12217 784 VIA_via1_4
* cell instance $12218 r0 *1 77.805,32.83
X$12218 784 VIA_via1_4
* cell instance $12219 r0 *1 77.805,32.83
X$12219 784 VIA_via2_5
* cell instance $12220 r0 *1 75.335,32.83
X$12220 784 VIA_via1_4
* cell instance $12221 r0 *1 75.335,32.83
X$12221 784 VIA_via2_5
* cell instance $12222 r0 *1 40.185,32.83
X$12222 785 VIA_via2_5
* cell instance $12223 r0 *1 39.235,32.83
X$12223 785 VIA_via1_4
* cell instance $12224 r0 *1 39.235,32.83
X$12224 785 VIA_via2_5
* cell instance $12225 r0 *1 40.185,31.43
X$12225 785 VIA_via1_4
* cell instance $12226 r0 *1 44.555,32.83
X$12226 786 VIA_via1_4
* cell instance $12227 r0 *1 44.555,32.69
X$12227 786 VIA_via2_5
* cell instance $12228 r0 *1 43.605,32.69
X$12228 786 VIA_via1_4
* cell instance $12229 r0 *1 43.605,32.69
X$12229 786 VIA_via2_5
* cell instance $12230 r0 *1 73.435,31.99
X$12230 787 VIA_via1_7
* cell instance $12231 r0 *1 73.435,32.83
X$12231 787 VIA_via1_4
* cell instance $12232 r0 *1 64.695,32.83
X$12232 788 VIA_via1_4
* cell instance $12233 r0 *1 64.695,32.97
X$12233 788 VIA_via2_5
* cell instance $12234 r0 *1 68.685,32.97
X$12234 788 VIA_via1_4
* cell instance $12235 r0 *1 68.685,32.97
X$12235 788 VIA_via2_5
* cell instance $12236 r0 *1 8.645,37.59
X$12236 789 VIA_via1_7
* cell instance $12237 r0 *1 8.645,38.43
X$12237 789 VIA_via2_5
* cell instance $12238 r0 *1 9.975,38.43
X$12238 789 VIA_via2_5
* cell instance $12239 r0 *1 8.455,38.43
X$12239 789 VIA_via2_5
* cell instance $12240 r0 *1 6.555,35.77
X$12240 789 VIA_via2_5
* cell instance $12241 r0 *1 3.515,35.77
X$12241 789 VIA_via2_5
* cell instance $12242 r0 *1 9.975,35.77
X$12242 789 VIA_via2_5
* cell instance $12243 r0 *1 4.845,35.91
X$12243 789 VIA_via2_5
* cell instance $12244 r0 *1 9.975,34.37
X$12244 789 VIA_via1_4
* cell instance $12245 r0 *1 6.555,34.37
X$12245 789 VIA_via1_4
* cell instance $12246 r0 *1 3.135,34.37
X$12246 789 VIA_via1_4
* cell instance $12247 r0 *1 8.455,39.97
X$12247 789 VIA_via1_4
* cell instance $12248 r0 *1 7.885,38.43
X$12248 789 VIA_via1_4
* cell instance $12249 r0 *1 7.885,38.43
X$12249 789 VIA_via2_5
* cell instance $12250 r0 *1 3.325,38.43
X$12250 789 VIA_via1_4
* cell instance $12251 r0 *1 4.085,39.97
X$12251 789 VIA_via1_4
* cell instance $12252 r0 *1 4.845,37.17
X$12252 789 VIA_via1_4
* cell instance $12253 r0 *1 12.635,38.43
X$12253 789 VIA_via1_4
* cell instance $12254 r0 *1 12.635,38.43
X$12254 789 VIA_via2_5
* cell instance $12255 r0 *1 7.125,34.79
X$12255 790 VIA_via2_5
* cell instance $12256 r0 *1 7.125,35.63
X$12256 790 VIA_via1_4
* cell instance $12257 r0 *1 4.465,32.83
X$12257 790 VIA_via1_4
* cell instance $12258 r0 *1 4.655,34.65
X$12258 790 VIA_via1_4
* cell instance $12259 r0 *1 4.655,34.79
X$12259 790 VIA_via2_5
* cell instance $12260 r0 *1 17.765,33.25
X$12260 791 VIA_via1_4
* cell instance $12261 r0 *1 17.955,34.37
X$12261 791 VIA_via1_4
* cell instance $12262 r0 *1 17.195,34.37
X$12262 791 VIA_via1_4
* cell instance $12263 r0 *1 17.765,34.23
X$12263 792 VIA_via1_7
* cell instance $12264 r0 *1 17.765,34.09
X$12264 792 VIA_via2_5
* cell instance $12265 r0 *1 15.105,34.23
X$12265 792 VIA_via1_7
* cell instance $12266 r0 *1 15.105,34.09
X$12266 792 VIA_via2_5
* cell instance $12267 r0 *1 29.545,80.57
X$12267 792 VIA_via1_7
* cell instance $12268 r0 *1 29.545,80.57
X$12268 792 VIA_via2_5
* cell instance $12269 r0 *1 18.145,59.43
X$12269 792 VIA_via1_7
* cell instance $12270 r0 *1 18.145,59.29
X$12270 792 VIA_via2_5
* cell instance $12271 r0 *1 25.555,79.87
X$12271 792 VIA_via2_5
* cell instance $12272 r0 *1 29.545,80.29
X$12272 792 VIA_via2_5
* cell instance $12273 r0 *1 16.625,79.17
X$12273 792 VIA_via2_5
* cell instance $12274 r0 *1 16.815,79.87
X$12274 792 VIA_via2_5
* cell instance $12275 r0 *1 38.285,80.29
X$12275 792 VIA_via2_5
* cell instance $12276 r0 *1 39.235,57.47
X$12276 792 VIA_via2_5
* cell instance $12277 r0 *1 38.285,81.97
X$12277 792 VIA_via1_4
* cell instance $12278 r0 *1 39.235,55.65
X$12278 792 VIA_via1_4
* cell instance $12279 r0 *1 25.555,80.43
X$12279 792 VIA_via1_4
* cell instance $12280 r0 *1 25.555,80.57
X$12280 792 VIA_via2_5
* cell instance $12281 r0 *1 16.055,79.17
X$12281 792 VIA_via1_4
* cell instance $12282 r0 *1 16.055,79.17
X$12282 792 VIA_via2_5
* cell instance $12283 r0 *1 16.625,80.43
X$12283 792 VIA_via1_4
* cell instance $12284 r0 *1 15.865,35.63
X$12284 792 VIA_via1_4
* cell instance $12285 r0 *1 15.865,35.63
X$12285 792 VIA_via2_5
* cell instance $12286 r0 *1 37.895,57.47
X$12286 792 VIA_via4_0
* cell instance $12287 r0 *1 37.895,57.47
X$12287 792 VIA_via3_2
* cell instance $12288 r0 *1 26.135,57.47
X$12288 792 VIA_via4_0
* cell instance $12289 r0 *1 17.735,58.03
X$12289 792 VIA_via4_0
* cell instance $12290 r0 *1 17.455,34.09
X$12290 792 VIA_via3_2
* cell instance $12291 r0 *1 17.455,35.63
X$12291 792 VIA_via3_2
* cell instance $12292 r0 *1 26.135,58.03
X$12292 792 VIA_via3_2
* cell instance $12293 r0 *1 26.125,58.03
X$12293 792 VIA_via2_5
* cell instance $12294 r0 *1 26.135,58.03
X$12294 792 VIA_via4_0
* cell instance $12295 r0 *1 26.125,58.03
X$12295 792 VIA_via1_4
* cell instance $12296 r0 *1 17.735,59.29
X$12296 792 VIA_via3_2
* cell instance $12297 r0 *1 30.685,34.37
X$12297 793 VIA_via1_4
* cell instance $12298 r0 *1 30.685,34.37
X$12298 793 VIA_via2_5
* cell instance $12299 r0 *1 27.075,34.37
X$12299 793 VIA_via1_4
* cell instance $12300 r0 *1 27.075,34.37
X$12300 793 VIA_via2_5
* cell instance $12301 r0 *1 31.065,34.37
X$12301 793 VIA_via1_4
* cell instance $12302 r0 *1 31.065,34.37
X$12302 793 VIA_via2_5
* cell instance $12303 r0 *1 39.045,41.23
X$12303 794 VIA_via1_4
* cell instance $12304 r0 *1 38.855,31.43
X$12304 794 VIA_via1_4
* cell instance $12305 r0 *1 52.155,37.17
X$12305 795 VIA_via1_4
* cell instance $12306 r0 *1 52.535,34.37
X$12306 795 VIA_via1_4
* cell instance $12307 r0 *1 54.055,34.23
X$12307 796 VIA_via1_7
* cell instance $12308 r0 *1 61.275,32.97
X$12308 796 VIA_via1_7
* cell instance $12309 r0 *1 62.605,56.21
X$12309 796 VIA_via1_7
* cell instance $12310 r0 *1 62.605,56.21
X$12310 796 VIA_via2_5
* cell instance $12311 r0 *1 52.155,56.21
X$12311 796 VIA_via2_5
* cell instance $12312 r0 *1 54.055,33.95
X$12312 796 VIA_via2_5
* cell instance $12313 r0 *1 61.275,33.95
X$12313 796 VIA_via2_5
* cell instance $12314 r0 *1 50.445,33.95
X$12314 796 VIA_via2_5
* cell instance $12315 r0 *1 62.795,48.37
X$12315 796 VIA_via1_4
* cell instance $12316 r0 *1 62.795,48.37
X$12316 796 VIA_via2_5
* cell instance $12317 r0 *1 50.445,34.37
X$12317 796 VIA_via1_4
* cell instance $12318 r0 *1 52.155,56.77
X$12318 796 VIA_via1_4
* cell instance $12319 r0 *1 62.535,33.95
X$12319 796 VIA_via3_2
* cell instance $12320 r0 *1 62.535,48.37
X$12320 796 VIA_via3_2
* cell instance $12321 r0 *1 56.525,33.25
X$12321 797 VIA_via1_4
* cell instance $12322 r0 *1 54.815,34.37
X$12322 797 VIA_via1_4
* cell instance $12323 r0 *1 54.815,34.37
X$12323 797 VIA_via2_5
* cell instance $12324 r0 *1 55.575,34.37
X$12324 797 VIA_via1_4
* cell instance $12325 r0 *1 55.575,34.37
X$12325 797 VIA_via2_5
* cell instance $12326 r0 *1 57.475,46.83
X$12326 798 VIA_via1_4
* cell instance $12327 r0 *1 57.095,33.95
X$12327 798 VIA_via1_4
* cell instance $12328 r0 *1 84.835,40.81
X$12328 799 VIA_via1_7
* cell instance $12329 r0 *1 84.835,40.67
X$12329 799 VIA_via2_5
* cell instance $12330 r0 *1 68.875,40.53
X$12330 799 VIA_via2_5
* cell instance $12331 r0 *1 85.975,40.67
X$12331 799 VIA_via2_5
* cell instance $12332 r0 *1 64.695,41.79
X$12332 799 VIA_via2_5
* cell instance $12333 r0 *1 64.315,41.79
X$12333 799 VIA_via2_5
* cell instance $12334 r0 *1 68.115,38.43
X$12334 799 VIA_via2_5
* cell instance $12335 r0 *1 68.305,45.57
X$12335 799 VIA_via2_5
* cell instance $12336 r0 *1 68.875,38.43
X$12336 799 VIA_via2_5
* cell instance $12337 r0 *1 67.165,38.43
X$12337 799 VIA_via1_4
* cell instance $12338 r0 *1 67.165,38.43
X$12338 799 VIA_via2_5
* cell instance $12339 r0 *1 64.315,39.97
X$12339 799 VIA_via1_4
* cell instance $12340 r0 *1 64.315,40.11
X$12340 799 VIA_via2_5
* cell instance $12341 r0 *1 64.505,42.77
X$12341 799 VIA_via1_4
* cell instance $12342 r0 *1 86.355,32.83
X$12342 799 VIA_via1_4
* cell instance $12343 r0 *1 85.975,34.37
X$12343 799 VIA_via1_4
* cell instance $12344 r0 *1 67.925,45.57
X$12344 799 VIA_via1_4
* cell instance $12345 r0 *1 67.925,45.57
X$12345 799 VIA_via2_5
* cell instance $12346 r0 *1 68.305,44.03
X$12346 799 VIA_via1_4
* cell instance $12347 r0 *1 68.875,39.97
X$12347 799 VIA_via1_4
* cell instance $12348 r0 *1 68.875,40.11
X$12348 799 VIA_via2_5
* cell instance $12349 r0 *1 68.305,32.83
X$12349 799 VIA_via1_4
* cell instance $12350 r0 *1 68.305,34.37
X$12350 799 VIA_via1_4
* cell instance $12351 r0 *1 71.345,37.17
X$12351 800 VIA_via1_4
* cell instance $12352 r0 *1 71.535,35.63
X$12352 800 VIA_via1_4
* cell instance $12353 r0 *1 71.155,34.37
X$12353 800 VIA_via1_4
* cell instance $12354 r0 *1 77.615,39.83
X$12354 801 VIA_via2_5
* cell instance $12355 r0 *1 73.625,39.83
X$12355 801 VIA_via2_5
* cell instance $12356 r0 *1 78.185,38.15
X$12356 801 VIA_via2_5
* cell instance $12357 r0 *1 74.005,39.83
X$12357 801 VIA_via2_5
* cell instance $12358 r0 *1 74.575,39.83
X$12358 801 VIA_via2_5
* cell instance $12359 r0 *1 76.665,38.15
X$12359 801 VIA_via2_5
* cell instance $12360 r0 *1 77.615,38.15
X$12360 801 VIA_via2_5
* cell instance $12361 r0 *1 81.415,38.43
X$12361 801 VIA_via1_4
* cell instance $12362 r0 *1 81.415,38.43
X$12362 801 VIA_via2_5
* cell instance $12363 r0 *1 78.185,38.43
X$12363 801 VIA_via1_4
* cell instance $12364 r0 *1 78.185,38.43
X$12364 801 VIA_via2_5
* cell instance $12365 r0 *1 73.625,40.04
X$12365 801 VIA_via1_4
* cell instance $12366 r0 *1 77.615,40.04
X$12366 801 VIA_via1_4
* cell instance $12367 r0 *1 77.615,41.23
X$12367 801 VIA_via1_4
* cell instance $12368 r0 *1 74.575,42.77
X$12368 801 VIA_via1_4
* cell instance $12369 r0 *1 74.005,37.17
X$12369 801 VIA_via1_4
* cell instance $12370 r0 *1 76.285,34.37
X$12370 801 VIA_via1_4
* cell instance $12371 r0 *1 76.855,31.57
X$12371 801 VIA_via1_4
* cell instance $12372 r0 *1 78.185,33.39
X$12372 802 VIA_via1_7
* cell instance $12373 r0 *1 78.755,34.37
X$12373 802 VIA_via1_4
* cell instance $12374 r0 *1 80.085,33.39
X$12374 803 VIA_via1_7
* cell instance $12375 r0 *1 80.085,33.39
X$12375 803 VIA_via2_5
* cell instance $12376 r0 *1 79.325,33.39
X$12376 803 VIA_via2_5
* cell instance $12377 r0 *1 78.945,35.63
X$12377 803 VIA_via1_4
* cell instance $12378 r0 *1 85.405,34.37
X$12378 804 VIA_via1_4
* cell instance $12379 r0 *1 85.405,34.37
X$12379 804 VIA_via2_5
* cell instance $12380 r0 *1 89.965,34.37
X$12380 804 VIA_via1_4
* cell instance $12381 r0 *1 89.965,34.37
X$12381 804 VIA_via2_5
* cell instance $12382 r0 *1 89.585,34.37
X$12382 804 VIA_via1_4
* cell instance $12383 r0 *1 89.585,34.37
X$12383 804 VIA_via2_5
* cell instance $12384 r0 *1 90.915,33.81
X$12384 805 VIA_via1_7
* cell instance $12385 r0 *1 90.725,32.83
X$12385 805 VIA_via1_4
* cell instance $12386 r0 *1 94.715,40.95
X$12386 806 VIA_via2_5
* cell instance $12387 r0 *1 96.615,40.95
X$12387 806 VIA_via2_5
* cell instance $12388 r0 *1 94.715,40.11
X$12388 806 VIA_via2_5
* cell instance $12389 r0 *1 92.055,40.95
X$12389 806 VIA_via2_5
* cell instance $12390 r0 *1 81.985,44.03
X$12390 806 VIA_via2_5
* cell instance $12391 r0 *1 86.355,44.03
X$12391 806 VIA_via2_5
* cell instance $12392 r0 *1 90.535,35.35
X$12392 806 VIA_via2_5
* cell instance $12393 r0 *1 94.715,35.35
X$12393 806 VIA_via2_5
* cell instance $12394 r0 *1 83.695,44.03
X$12394 806 VIA_via1_4
* cell instance $12395 r0 *1 83.695,44.03
X$12395 806 VIA_via2_5
* cell instance $12396 r0 *1 81.795,45.57
X$12396 806 VIA_via1_4
* cell instance $12397 r0 *1 93.385,39.97
X$12397 806 VIA_via1_4
* cell instance $12398 r0 *1 93.385,40.11
X$12398 806 VIA_via2_5
* cell instance $12399 r0 *1 90.535,35.63
X$12399 806 VIA_via1_4
* cell instance $12400 r0 *1 94.525,34.37
X$12400 806 VIA_via1_4
* cell instance $12401 r0 *1 96.615,45.15
X$12401 806 VIA_via1_4
* cell instance $12402 r0 *1 86.355,41.23
X$12402 806 VIA_via1_4
* cell instance $12403 r0 *1 86.355,41.37
X$12403 806 VIA_via2_5
* cell instance $12404 r0 *1 92.055,41.23
X$12404 806 VIA_via1_4
* cell instance $12405 r0 *1 92.055,41.37
X$12405 806 VIA_via2_5
* cell instance $12406 r0 *1 4.845,33.39
X$12406 807 VIA_via1_7
* cell instance $12407 r0 *1 4.845,33.39
X$12407 807 VIA_via2_5
* cell instance $12408 r0 *1 2.375,33.39
X$12408 807 VIA_via2_5
* cell instance $12409 r0 *1 2.375,34.37
X$12409 807 VIA_via1_4
* cell instance $12410 r0 *1 7.125,33.39
X$12410 808 VIA_via1_7
* cell instance $12411 r0 *1 7.125,34.37
X$12411 808 VIA_via2_5
* cell instance $12412 r0 *1 5.795,34.37
X$12412 808 VIA_via1_4
* cell instance $12413 r0 *1 5.795,34.37
X$12413 808 VIA_via2_5
* cell instance $12414 r0 *1 9.975,33.39
X$12414 809 VIA_via1_7
* cell instance $12415 r0 *1 9.975,33.39
X$12415 809 VIA_via2_5
* cell instance $12416 r0 *1 9.215,33.39
X$12416 809 VIA_via2_5
* cell instance $12417 r0 *1 9.215,34.37
X$12417 809 VIA_via1_4
* cell instance $12418 r0 *1 10.925,33.95
X$12418 810 VIA_via2_5
* cell instance $12419 r0 *1 9.595,33.95
X$12419 810 VIA_via2_5
* cell instance $12420 r0 *1 11.495,33.95
X$12420 810 VIA_via1_4
* cell instance $12421 r0 *1 11.495,33.95
X$12421 810 VIA_via2_5
* cell instance $12422 r0 *1 9.595,32.83
X$12422 810 VIA_via1_4
* cell instance $12423 r0 *1 10.925,35.63
X$12423 810 VIA_via1_4
* cell instance $12424 r0 *1 91.485,35.21
X$12424 811 VIA_via1_7
* cell instance $12425 r0 *1 91.485,34.37
X$12425 811 VIA_via2_5
* cell instance $12426 r0 *1 91.865,34.37
X$12426 811 VIA_via1_4
* cell instance $12427 r0 *1 91.865,34.37
X$12427 811 VIA_via2_5
* cell instance $12428 r0 *1 14.535,34.37
X$12428 812 VIA_via2_5
* cell instance $12429 r0 *1 13.585,34.37
X$12429 812 VIA_via2_5
* cell instance $12430 r0 *1 14.535,33.25
X$12430 812 VIA_via1_4
* cell instance $12431 r0 *1 15.295,34.37
X$12431 812 VIA_via1_4
* cell instance $12432 r0 *1 15.295,34.37
X$12432 812 VIA_via2_5
* cell instance $12433 r0 *1 13.585,35.63
X$12433 812 VIA_via1_4
* cell instance $12434 r0 *1 9.785,81.83
X$12434 813 VIA_via1_7
* cell instance $12435 r0 *1 24.795,34.23
X$12435 813 VIA_via1_7
* cell instance $12436 r0 *1 24.795,34.23
X$12436 813 VIA_via2_5
* cell instance $12437 r0 *1 11.685,58.17
X$12437 813 VIA_via1_7
* cell instance $12438 r0 *1 11.685,58.17
X$12438 813 VIA_via2_5
* cell instance $12439 r0 *1 10.545,79.87
X$12439 813 VIA_via2_5
* cell instance $12440 r0 *1 14.535,77.49
X$12440 813 VIA_via2_5
* cell instance $12441 r0 *1 10.545,77.63
X$12441 813 VIA_via2_5
* cell instance $12442 r0 *1 20.995,80.01
X$12442 813 VIA_via2_5
* cell instance $12443 r0 *1 10.735,35.35
X$12443 813 VIA_via2_5
* cell instance $12444 r0 *1 8.455,35.35
X$12444 813 VIA_via2_5
* cell instance $12445 r0 *1 6.935,35.35
X$12445 813 VIA_via2_5
* cell instance $12446 r0 *1 16.055,45.15
X$12446 813 VIA_via2_5
* cell instance $12447 r0 *1 24.035,45.15
X$12447 813 VIA_via2_5
* cell instance $12448 r0 *1 15.295,46.13
X$12448 813 VIA_via2_5
* cell instance $12449 r0 *1 16.055,46.13
X$12449 813 VIA_via2_5
* cell instance $12450 r0 *1 14.725,58.17
X$12450 813 VIA_via2_5
* cell instance $12451 r0 *1 13.585,58.17
X$12451 813 VIA_via2_5
* cell instance $12452 r0 *1 23.845,34.23
X$12452 813 VIA_via2_5
* cell instance $12453 r0 *1 23.845,35.35
X$12453 813 VIA_via2_5
* cell instance $12454 r0 *1 13.585,62.37
X$12454 813 VIA_via1_4
* cell instance $12455 r0 *1 9.975,77.63
X$12455 813 VIA_via1_4
* cell instance $12456 r0 *1 9.975,77.63
X$12456 813 VIA_via2_5
* cell instance $12457 r0 *1 20.995,80.43
X$12457 813 VIA_via1_4
* cell instance $12458 r0 *1 6.935,35.63
X$12458 813 VIA_via1_4
* cell instance $12459 r0 *1 8.455,35.63
X$12459 813 VIA_via1_4
* cell instance $12460 r0 *1 10.735,35.63
X$12460 813 VIA_via1_4
* cell instance $12461 r0 *1 6.555,37.17
X$12461 813 VIA_via1_4
* cell instance $12462 r0 *1 25.365,45.15
X$12462 813 VIA_via1_4
* cell instance $12463 r0 *1 25.365,45.15
X$12463 813 VIA_via2_5
* cell instance $12464 r0 *1 78.565,33.95
X$12464 814 VIA_via2_5
* cell instance $12465 r0 *1 78.755,35.63
X$12465 814 VIA_via1_4
* cell instance $12466 r0 *1 79.135,33.95
X$12466 814 VIA_via1_4
* cell instance $12467 r0 *1 79.135,33.95
X$12467 814 VIA_via2_5
* cell instance $12468 r0 *1 27.455,34.37
X$12468 815 VIA_via1_4
* cell instance $12469 r0 *1 28.405,34.37
X$12469 815 VIA_via1_4
* cell instance $12470 r0 *1 76.285,33.39
X$12470 816 VIA_via1_7
* cell instance $12471 r0 *1 76.285,33.67
X$12471 816 VIA_via2_5
* cell instance $12472 r0 *1 75.525,33.67
X$12472 816 VIA_via2_5
* cell instance $12473 r0 *1 75.525,34.37
X$12473 816 VIA_via1_4
* cell instance $12474 r0 *1 37.525,35.21
X$12474 817 VIA_via1_7
* cell instance $12475 r0 *1 37.525,34.37
X$12475 817 VIA_via2_5
* cell instance $12476 r0 *1 36.385,34.37
X$12476 817 VIA_via1_4
* cell instance $12477 r0 *1 36.385,34.37
X$12477 817 VIA_via2_5
* cell instance $12478 r0 *1 73.245,33.39
X$12478 818 VIA_via1_7
* cell instance $12479 r0 *1 73.245,33.39
X$12479 818 VIA_via2_5
* cell instance $12480 r0 *1 73.815,33.39
X$12480 818 VIA_via2_5
* cell instance $12481 r0 *1 73.815,35.63
X$12481 818 VIA_via1_4
* cell instance $12482 r0 *1 65.265,34.37
X$12482 819 VIA_via2_5
* cell instance $12483 r0 *1 65.075,34.37
X$12483 819 VIA_via1_4
* cell instance $12484 r0 *1 68.685,34.37
X$12484 819 VIA_via1_4
* cell instance $12485 r0 *1 68.685,34.37
X$12485 819 VIA_via2_5
* cell instance $12486 r0 *1 51.395,35.35
X$12486 820 VIA_via1_4
* cell instance $12487 r0 *1 51.585,34.37
X$12487 820 VIA_via1_4
* cell instance $12488 r0 *1 51.585,34.37
X$12488 820 VIA_via2_5
* cell instance $12489 r0 *1 48.925,34.37
X$12489 820 VIA_via1_4
* cell instance $12490 r0 *1 48.925,34.37
X$12490 820 VIA_via2_5
* cell instance $12491 r0 *1 64.125,57.61
X$12491 821 VIA_via1_7
* cell instance $12492 r0 *1 64.125,57.61
X$12492 821 VIA_via2_5
* cell instance $12493 r0 *1 65.075,57.61
X$12493 821 VIA_via2_5
* cell instance $12494 r0 *1 64.505,35.49
X$12494 821 VIA_via2_5
* cell instance $12495 r0 *1 51.015,33.39
X$12495 821 VIA_via2_5
* cell instance $12496 r0 *1 57.665,35.49
X$12496 821 VIA_via2_5
* cell instance $12497 r0 *1 57.665,33.39
X$12497 821 VIA_via2_5
* cell instance $12498 r0 *1 51.015,32.83
X$12498 821 VIA_via1_4
* cell instance $12499 r0 *1 53.865,58.03
X$12499 821 VIA_via1_4
* cell instance $12500 r0 *1 53.865,57.89
X$12500 821 VIA_via2_5
* cell instance $12501 r0 *1 59.185,35.63
X$12501 821 VIA_via1_4
* cell instance $12502 r0 *1 59.185,35.49
X$12502 821 VIA_via2_5
* cell instance $12503 r0 *1 56.715,35.63
X$12503 821 VIA_via1_4
* cell instance $12504 r0 *1 56.715,35.49
X$12504 821 VIA_via2_5
* cell instance $12505 r0 *1 65.075,55.23
X$12505 821 VIA_via1_4
* cell instance $12506 r0 *1 55.195,33.81
X$12506 822 VIA_via1_7
* cell instance $12507 r0 *1 55.195,33.81
X$12507 822 VIA_via2_5
* cell instance $12508 r0 *1 54.245,33.81
X$12508 822 VIA_via2_5
* cell instance $12509 r0 *1 54.245,32.83
X$12509 822 VIA_via1_4
* cell instance $12510 r0 *1 56.715,34.37
X$12510 823 VIA_via1_4
* cell instance $12511 r0 *1 56.525,34.37
X$12511 823 VIA_via1_4
* cell instance $12512 r0 *1 59.945,33.39
X$12512 824 VIA_via1_7
* cell instance $12513 r0 *1 59.945,33.39
X$12513 824 VIA_via2_5
* cell instance $12514 r0 *1 58.805,33.39
X$12514 824 VIA_via2_5
* cell instance $12515 r0 *1 58.805,34.37
X$12515 824 VIA_via1_4
* cell instance $12516 r0 *1 6.745,34.65
X$12516 825 VIA_via2_5
* cell instance $12517 r0 *1 8.645,34.65
X$12517 825 VIA_via2_5
* cell instance $12518 r0 *1 6.745,32.83
X$12518 825 VIA_via1_4
* cell instance $12519 r0 *1 8.645,35.63
X$12519 825 VIA_via1_4
* cell instance $12520 r0 *1 8.075,34.65
X$12520 825 VIA_via1_4
* cell instance $12521 r0 *1 8.075,34.65
X$12521 825 VIA_via2_5
* cell instance $12522 r0 *1 16.055,35.63
X$12522 826 VIA_via1_4
* cell instance $12523 r0 *1 14.915,34.65
X$12523 826 VIA_via1_4
* cell instance $12524 r0 *1 14.915,35.63
X$12524 826 VIA_via1_4
* cell instance $12525 r0 *1 18.905,34.79
X$12525 827 VIA_via1_7
* cell instance $12526 r0 *1 18.715,37.17
X$12526 827 VIA_via1_4
* cell instance $12527 r0 *1 30.495,31.43
X$12527 828 VIA_via1_4
* cell instance $12528 r0 *1 31.255,35.63
X$12528 828 VIA_via1_4
* cell instance $12529 r0 *1 37.145,41.23
X$12529 829 VIA_via2_5
* cell instance $12530 r0 *1 37.525,57.05
X$12530 829 VIA_via2_5
* cell instance $12531 r0 *1 26.315,35.77
X$12531 829 VIA_via2_5
* cell instance $12532 r0 *1 28.025,59.43
X$12532 829 VIA_via2_5
* cell instance $12533 r0 *1 19.095,35.77
X$12533 829 VIA_via2_5
* cell instance $12534 r0 *1 28.025,57.19
X$12534 829 VIA_via2_5
* cell instance $12535 r0 *1 28.025,58.03
X$12535 829 VIA_via1_4
* cell instance $12536 r0 *1 39.425,41.23
X$12536 829 VIA_via1_4
* cell instance $12537 r0 *1 39.425,41.23
X$12537 829 VIA_via2_5
* cell instance $12538 r0 *1 23.085,59.57
X$12538 829 VIA_via1_4
* cell instance $12539 r0 *1 23.085,59.43
X$12539 829 VIA_via2_5
* cell instance $12540 r0 *1 36.575,57.05
X$12540 829 VIA_via1_4
* cell instance $12541 r0 *1 36.575,57.05
X$12541 829 VIA_via2_5
* cell instance $12542 r0 *1 19.095,37.17
X$12542 829 VIA_via1_4
* cell instance $12543 r0 *1 19.095,37.03
X$12543 829 VIA_via2_5
* cell instance $12544 r0 *1 18.145,37.17
X$12544 829 VIA_via1_4
* cell instance $12545 r0 *1 18.145,37.03
X$12545 829 VIA_via2_5
* cell instance $12546 r0 *1 19.665,37.17
X$12546 829 VIA_via1_4
* cell instance $12547 r0 *1 19.665,37.03
X$12547 829 VIA_via2_5
* cell instance $12548 r0 *1 17.955,35.63
X$12548 829 VIA_via1_4
* cell instance $12549 r0 *1 17.955,35.77
X$12549 829 VIA_via2_5
* cell instance $12550 r0 *1 35.815,35.63
X$12550 829 VIA_via1_4
* cell instance $12551 r0 *1 35.815,35.63
X$12551 829 VIA_via2_5
* cell instance $12552 r0 *1 35.935,35.63
X$12552 829 VIA_via3_2
* cell instance $12553 r0 *1 26.315,37.17
X$12553 829 VIA_via1_4
* cell instance $12554 r0 *1 26.315,37.03
X$12554 829 VIA_via2_5
* cell instance $12555 r0 *1 31.635,35.63
X$12555 829 VIA_via1_4
* cell instance $12556 r0 *1 31.635,35.63
X$12556 829 VIA_via2_5
* cell instance $12557 r0 *1 35.935,41.23
X$12557 829 VIA_via3_2
* cell instance $12558 r0 *1 32.015,34.79
X$12558 830 VIA_via1_7
* cell instance $12559 r0 *1 31.825,35.63
X$12559 830 VIA_via1_4
* cell instance $12560 r0 *1 24.415,62.09
X$12560 831 VIA_via2_5
* cell instance $12561 r0 *1 20.995,62.09
X$12561 831 VIA_via2_5
* cell instance $12562 r0 *1 38.285,58.59
X$12562 831 VIA_via2_5
* cell instance $12563 r0 *1 38.175,58.59
X$12563 831 VIA_via3_2
* cell instance $12564 r0 *1 27.265,36.89
X$12564 831 VIA_via2_5
* cell instance $12565 r0 *1 16.435,36.89
X$12565 831 VIA_via2_5
* cell instance $12566 r0 *1 17.575,36.89
X$12566 831 VIA_via2_5
* cell instance $12567 r0 *1 17.005,36.89
X$12567 831 VIA_via2_5
* cell instance $12568 r0 *1 32.015,36.89
X$12568 831 VIA_via2_5
* cell instance $12569 r0 *1 24.415,58.45
X$12569 831 VIA_via2_5
* cell instance $12570 r0 *1 38.285,59.15
X$12570 831 VIA_via1_4
* cell instance $12571 r0 *1 39.235,42.77
X$12571 831 VIA_via1_4
* cell instance $12572 r0 *1 39.235,42.77
X$12572 831 VIA_via2_5
* cell instance $12573 r0 *1 20.995,62.37
X$12573 831 VIA_via1_4
* cell instance $12574 r0 *1 24.415,58.03
X$12574 831 VIA_via1_4
* cell instance $12575 r0 *1 17.005,37.17
X$12575 831 VIA_via1_4
* cell instance $12576 r0 *1 17.005,38.5
X$12576 831 VIA_via1_4
* cell instance $12577 r0 *1 17.575,37.17
X$12577 831 VIA_via1_4
* cell instance $12578 r0 *1 16.435,37.17
X$12578 831 VIA_via1_4
* cell instance $12579 r0 *1 35.245,35.63
X$12579 831 VIA_via1_4
* cell instance $12580 r0 *1 35.245,35.49
X$12580 831 VIA_via2_5
* cell instance $12581 r0 *1 32.205,35.63
X$12581 831 VIA_via1_4
* cell instance $12582 r0 *1 32.205,35.49
X$12582 831 VIA_via2_5
* cell instance $12583 r0 *1 27.265,37.17
X$12583 831 VIA_via1_4
* cell instance $12584 r0 *1 38.175,35.49
X$12584 831 VIA_via3_2
* cell instance $12585 r0 *1 38.175,42.77
X$12585 831 VIA_via3_2
* cell instance $12586 r0 *1 35.055,34.79
X$12586 832 VIA_via1_7
* cell instance $12587 r0 *1 34.865,35.63
X$12587 832 VIA_via1_4
* cell instance $12588 r0 *1 38.665,35.63
X$12588 833 VIA_via2_5
* cell instance $12589 r0 *1 37.905,35.63
X$12589 833 VIA_via1_4
* cell instance $12590 r0 *1 37.905,35.63
X$12590 833 VIA_via2_5
* cell instance $12591 r0 *1 38.665,34.65
X$12591 833 VIA_via1_4
* cell instance $12592 r0 *1 37.145,35.63
X$12592 833 VIA_via1_4
* cell instance $12593 r0 *1 37.145,35.63
X$12593 833 VIA_via2_5
* cell instance $12594 r0 *1 43.985,35.63
X$12594 834 VIA_via2_5
* cell instance $12595 r0 *1 42.845,35.63
X$12595 834 VIA_via2_5
* cell instance $12596 r0 *1 44.175,37.17
X$12596 834 VIA_via1_4
* cell instance $12597 r0 *1 42.845,36.75
X$12597 834 VIA_via1_4
* cell instance $12598 r0 *1 40.375,35.63
X$12598 834 VIA_via1_4
* cell instance $12599 r0 *1 40.375,35.63
X$12599 834 VIA_via2_5
* cell instance $12600 r0 *1 44.745,38.01
X$12600 835 VIA_via1_7
* cell instance $12601 r0 *1 44.175,35.63
X$12601 835 VIA_via1_4
* cell instance $12602 r0 *1 43.795,37.03
X$12602 836 VIA_via2_5
* cell instance $12603 r0 *1 46.265,37.03
X$12603 836 VIA_via2_5
* cell instance $12604 r0 *1 44.745,37.17
X$12604 836 VIA_via1_4
* cell instance $12605 r0 *1 44.745,37.03
X$12605 836 VIA_via2_5
* cell instance $12606 r0 *1 43.795,38.43
X$12606 836 VIA_via1_4
* cell instance $12607 r0 *1 46.455,35.35
X$12607 836 VIA_via1_4
* cell instance $12608 r0 *1 46.645,30.59
X$12608 837 VIA_via1_7
* cell instance $12609 r0 *1 46.265,38.43
X$12609 837 VIA_via1_4
* cell instance $12610 r0 *1 49.305,34.79
X$12610 838 VIA_via1_7
* cell instance $12611 r0 *1 49.115,35.63
X$12611 838 VIA_via1_4
* cell instance $12612 r0 *1 55.005,37.03
X$12612 839 VIA_via2_5
* cell instance $12613 r0 *1 49.875,37.03
X$12613 839 VIA_via2_5
* cell instance $12614 r0 *1 55.385,37.03
X$12614 839 VIA_via2_5
* cell instance $12615 r0 *1 56.525,37.17
X$12615 839 VIA_via1_4
* cell instance $12616 r0 *1 56.525,37.03
X$12616 839 VIA_via2_5
* cell instance $12617 r0 *1 49.495,38.43
X$12617 839 VIA_via1_4
* cell instance $12618 r0 *1 50.065,39.97
X$12618 839 VIA_via1_4
* cell instance $12619 r0 *1 53.105,37.03
X$12619 839 VIA_via1_4
* cell instance $12620 r0 *1 53.105,37.03
X$12620 839 VIA_via2_5
* cell instance $12621 r0 *1 59.755,37.17
X$12621 839 VIA_via1_4
* cell instance $12622 r0 *1 59.755,37.03
X$12622 839 VIA_via2_5
* cell instance $12623 r0 *1 55.005,38.43
X$12623 839 VIA_via1_4
* cell instance $12624 r0 *1 49.875,35.63
X$12624 839 VIA_via1_4
* cell instance $12625 r0 *1 55.385,35.63
X$12625 839 VIA_via1_4
* cell instance $12626 r0 *1 55.005,32.83
X$12626 839 VIA_via1_4
* cell instance $12627 r0 *1 50.635,38.43
X$12627 840 VIA_via2_5
* cell instance $12628 r0 *1 50.635,39.13
X$12628 840 VIA_via2_5
* cell instance $12629 r0 *1 38.475,39.97
X$12629 840 VIA_via2_5
* cell instance $12630 r0 *1 55.955,46.83
X$12630 840 VIA_via2_5
* cell instance $12631 r0 *1 56.145,39.13
X$12631 840 VIA_via2_5
* cell instance $12632 r0 *1 38.475,60.13
X$12632 840 VIA_via2_5
* cell instance $12633 r0 *1 72.675,35.35
X$12633 840 VIA_via2_5
* cell instance $12634 r0 *1 56.145,45.71
X$12634 840 VIA_via2_5
* cell instance $12635 r0 *1 75.905,35.35
X$12635 840 VIA_via2_5
* cell instance $12636 r0 *1 78.375,35.35
X$12636 840 VIA_via2_5
* cell instance $12637 r0 *1 61.845,45.01
X$12637 840 VIA_via2_5
* cell instance $12638 r0 *1 72.485,45.01
X$12638 840 VIA_via2_5
* cell instance $12639 r0 *1 51.585,38.43
X$12639 840 VIA_via1_4
* cell instance $12640 r0 *1 51.585,38.43
X$12640 840 VIA_via2_5
* cell instance $12641 r0 *1 75.905,35.63
X$12641 840 VIA_via1_4
* cell instance $12642 r0 *1 78.375,34.37
X$12642 840 VIA_via1_4
* cell instance $12643 r0 *1 61.845,45.57
X$12643 840 VIA_via1_4
* cell instance $12644 r0 *1 61.845,45.71
X$12644 840 VIA_via2_5
* cell instance $12645 r0 *1 61.975,45.71
X$12645 840 VIA_via3_2
* cell instance $12646 r0 *1 56.145,46.9
X$12646 840 VIA_via1_4
* cell instance $12647 r0 *1 56.145,46.83
X$12647 840 VIA_via2_5
* cell instance $12648 r0 *1 38.475,59.57
X$12648 840 VIA_via1_4
* cell instance $12649 r0 *1 46.075,37.17
X$12649 840 VIA_via1_4
* cell instance $12650 r0 *1 46.075,37.31
X$12650 840 VIA_via2_5
* cell instance $12651 r0 *1 38.285,39.97
X$12651 840 VIA_via1_4
* cell instance $12652 r0 *1 38.475,42.77
X$12652 840 VIA_via1_4
* cell instance $12653 r0 *1 62.795,59.85
X$12653 840 VIA_via1_4
* cell instance $12654 r0 *1 62.795,59.99
X$12654 840 VIA_via2_5
* cell instance $12655 r0 *1 72.675,35.63
X$12655 840 VIA_via1_4
* cell instance $12656 r0 *1 61.975,59.99
X$12656 840 VIA_via3_2
* cell instance $12657 r0 *1 44.615,37.31
X$12657 840 VIA_via3_2
* cell instance $12658 r0 *1 44.615,39.97
X$12658 840 VIA_via3_2
* cell instance $12659 r0 *1 44.615,39.13
X$12659 840 VIA_via3_2
* cell instance $12660 r0 *1 83.505,52.71
X$12660 841 VIA_via2_5
* cell instance $12661 r0 *1 82.935,52.57
X$12661 841 VIA_via2_5
* cell instance $12662 r0 *1 83.505,53.83
X$12662 841 VIA_via2_5
* cell instance $12663 r0 *1 82.745,37.87
X$12663 841 VIA_via2_5
* cell instance $12664 r0 *1 74.385,37.87
X$12664 841 VIA_via2_5
* cell instance $12665 r0 *1 74.005,35.35
X$12665 841 VIA_via1_4
* cell instance $12666 r0 *1 84.455,53.97
X$12666 841 VIA_via1_4
* cell instance $12667 r0 *1 84.455,53.83
X$12667 841 VIA_via2_5
* cell instance $12668 r0 *1 84.455,54.11
X$12668 841 VIA_via2_5
* cell instance $12669 r0 *1 85.595,53.97
X$12669 841 VIA_via1_4
* cell instance $12670 r0 *1 85.595,54.11
X$12670 841 VIA_via2_5
* cell instance $12671 r0 *1 96.235,35.35
X$12671 842 VIA_via2_5
* cell instance $12672 r0 *1 96.235,35.63
X$12672 842 VIA_via1_4
* cell instance $12673 r0 *1 97.255,35.35
X$12673 842 VIA_via3_2
* cell instance $12674 r0 *1 97.255,35.35
X$12674 842 VIA_via4_0
* cell instance $12675 r0 *1 95.095,35.49
X$12675 843 VIA_via2_5
* cell instance $12676 r0 *1 91.865,35.63
X$12676 843 VIA_via1_4
* cell instance $12677 r0 *1 91.865,35.49
X$12677 843 VIA_via2_5
* cell instance $12678 r0 *1 95.095,34.37
X$12678 843 VIA_via1_4
* cell instance $12679 r0 *1 96.045,35.49
X$12679 843 VIA_via1_4
* cell instance $12680 r0 *1 96.045,35.49
X$12680 843 VIA_via2_5
* cell instance $12681 r0 *1 95.475,34.79
X$12681 844 VIA_via1_7
* cell instance $12682 r0 *1 95.475,34.79
X$12682 844 VIA_via2_5
* cell instance $12683 r0 *1 93.765,34.79
X$12683 844 VIA_via2_5
* cell instance $12684 r0 *1 93.765,35.63
X$12684 844 VIA_via1_4
* cell instance $12685 r0 *1 6.365,35.63
X$12685 845 VIA_via2_5
* cell instance $12686 r0 *1 6.745,37.17
X$12686 845 VIA_via1_4
* cell instance $12687 r0 *1 4.845,35.63
X$12687 845 VIA_via1_4
* cell instance $12688 r0 *1 4.845,35.63
X$12688 845 VIA_via2_5
* cell instance $12689 r0 *1 6.365,36.75
X$12689 845 VIA_via1_4
* cell instance $12690 r0 *1 92.435,34.65
X$12690 846 VIA_via2_5
* cell instance $12691 r0 *1 91.105,35.63
X$12691 846 VIA_via1_4
* cell instance $12692 r0 *1 91.105,35.63
X$12692 846 VIA_via2_5
* cell instance $12693 r0 *1 94.145,34.65
X$12693 846 VIA_via1_4
* cell instance $12694 r0 *1 94.145,34.65
X$12694 846 VIA_via2_5
* cell instance $12695 r0 *1 92.435,35.63
X$12695 846 VIA_via1_4
* cell instance $12696 r0 *1 92.435,35.63
X$12696 846 VIA_via2_5
* cell instance $12697 r0 *1 13.965,35.21
X$12697 847 VIA_via1_7
* cell instance $12698 r0 *1 13.965,35.21
X$12698 847 VIA_via2_5
* cell instance $12699 r0 *1 12.255,35.21
X$12699 847 VIA_via2_5
* cell instance $12700 r0 *1 12.255,32.83
X$12700 847 VIA_via1_4
* cell instance $12701 r0 *1 86.355,34.51
X$12701 848 VIA_via1_4
* cell instance $12702 r0 *1 86.355,34.51
X$12702 848 VIA_via2_5
* cell instance $12703 r0 *1 87.305,34.37
X$12703 848 VIA_via1_4
* cell instance $12704 r0 *1 87.305,34.51
X$12704 848 VIA_via2_5
* cell instance $12705 r0 *1 16.245,34.79
X$12705 849 VIA_via1_7
* cell instance $12706 r0 *1 16.245,34.79
X$12706 849 VIA_via2_5
* cell instance $12707 r0 *1 17.575,34.79
X$12707 849 VIA_via2_5
* cell instance $12708 r0 *1 17.575,35.63
X$12708 849 VIA_via1_4
* cell instance $12709 r0 *1 78.185,34.79
X$12709 850 VIA_via1_7
* cell instance $12710 r0 *1 78.185,35.63
X$12710 850 VIA_via1_4
* cell instance $12711 r0 *1 23.275,35.63
X$12711 851 VIA_via2_5
* cell instance $12712 r0 *1 23.275,38.43
X$12712 851 VIA_via1_4
* cell instance $12713 r0 *1 24.035,35.63
X$12713 851 VIA_via1_4
* cell instance $12714 r0 *1 24.035,35.63
X$12714 851 VIA_via2_5
* cell instance $12715 r0 *1 19.855,35.63
X$12715 851 VIA_via1_4
* cell instance $12716 r0 *1 19.855,35.63
X$12716 851 VIA_via2_5
* cell instance $12717 r0 *1 25.935,34.79
X$12717 852 VIA_via1_7
* cell instance $12718 r0 *1 25.935,34.79
X$12718 852 VIA_via2_5
* cell instance $12719 r0 *1 26.885,34.79
X$12719 852 VIA_via2_5
* cell instance $12720 r0 *1 26.885,37.17
X$12720 852 VIA_via1_4
* cell instance $12721 r0 *1 73.625,35.63
X$12721 853 VIA_via1_4
* cell instance $12722 r0 *1 73.625,33.11
X$12722 853 VIA_via1_4
* cell instance $12723 r0 *1 71.535,34.79
X$12723 854 VIA_via1_7
* cell instance $12724 r0 *1 71.535,34.79
X$12724 854 VIA_via2_5
* cell instance $12725 r0 *1 69.255,34.79
X$12725 854 VIA_via2_5
* cell instance $12726 r0 *1 69.255,35.63
X$12726 854 VIA_via1_4
* cell instance $12727 r0 *1 62.415,34.79
X$12727 855 VIA_via1_7
* cell instance $12728 r0 *1 62.415,35.63
X$12728 855 VIA_via1_4
* cell instance $12729 r0 *1 61.275,35.63
X$12729 856 VIA_via2_5
* cell instance $12730 r0 *1 61.275,36.75
X$12730 856 VIA_via1_4
* cell instance $12731 r0 *1 61.275,38.43
X$12731 856 VIA_via1_4
* cell instance $12732 r0 *1 59.945,35.63
X$12732 856 VIA_via1_4
* cell instance $12733 r0 *1 59.945,35.63
X$12733 856 VIA_via2_5
* cell instance $12734 r0 *1 17.005,36.19
X$12734 857 VIA_via1_7
* cell instance $12735 r0 *1 17.765,37.17
X$12735 857 VIA_via1_4
* cell instance $12736 r0 *1 37.715,45.43
X$12736 858 VIA_via1_7
* cell instance $12737 r0 *1 37.715,45.43
X$12737 858 VIA_via2_5
* cell instance $12738 r0 *1 37.615,45.43
X$12738 858 VIA_via3_2
* cell instance $12739 r0 *1 48.355,41.37
X$12739 858 VIA_via1_7
* cell instance $12740 r0 *1 48.355,41.37
X$12740 858 VIA_via2_5
* cell instance $12741 r0 *1 13.775,45.43
X$12741 858 VIA_via1_7
* cell instance $12742 r0 *1 16.815,41.37
X$12742 858 VIA_via1_7
* cell instance $12743 r0 *1 16.815,41.37
X$12743 858 VIA_via2_5
* cell instance $12744 r0 *1 40.185,35.77
X$12744 858 VIA_via1_7
* cell instance $12745 r0 *1 48.545,43.75
X$12745 858 VIA_via2_5
* cell instance $12746 r0 *1 48.925,43.75
X$12746 858 VIA_via2_5
* cell instance $12747 r0 *1 48.545,45.43
X$12747 858 VIA_via2_5
* cell instance $12748 r0 *1 27.455,36.75
X$12748 858 VIA_via2_5
* cell instance $12749 r0 *1 48.925,41.37
X$12749 858 VIA_via2_5
* cell instance $12750 r0 *1 40.185,36.05
X$12750 858 VIA_via2_5
* cell instance $12751 r0 *1 14.345,41.37
X$12751 858 VIA_via2_5
* cell instance $12752 r0 *1 19.665,36.75
X$12752 858 VIA_via2_5
* cell instance $12753 r0 *1 14.345,36.75
X$12753 858 VIA_via2_5
* cell instance $12754 r0 *1 27.455,37.73
X$12754 858 VIA_via2_5
* cell instance $12755 r0 *1 13.775,41.37
X$12755 858 VIA_via2_5
* cell instance $12756 r0 *1 35.625,37.73
X$12756 858 VIA_via2_5
* cell instance $12757 r0 *1 48.545,45.15
X$12757 858 VIA_via1_4
* cell instance $12758 r0 *1 19.665,35.63
X$12758 858 VIA_via1_4
* cell instance $12759 r0 *1 27.455,37.17
X$12759 858 VIA_via1_4
* cell instance $12760 r0 *1 35.625,38.43
X$12760 858 VIA_via1_4
* cell instance $12761 r0 *1 13.395,46.83
X$12761 858 VIA_via1_4
* cell instance $12762 r0 *1 14.345,38.43
X$12762 858 VIA_via1_4
* cell instance $12763 r0 *1 37.615,36.05
X$12763 858 VIA_via3_2
* cell instance $12764 r0 *1 37.615,37.73
X$12764 858 VIA_via3_2
* cell instance $12765 r0 *1 35.815,36.19
X$12765 859 VIA_via1_7
* cell instance $12766 r0 *1 36.005,39.97
X$12766 859 VIA_via1_4
* cell instance $12767 r0 *1 41.325,36.19
X$12767 860 VIA_via1_7
* cell instance $12768 r0 *1 40.565,37.17
X$12768 860 VIA_via1_4
* cell instance $12769 r0 *1 52.915,36.19
X$12769 861 VIA_via1_7
* cell instance $12770 r0 *1 52.915,38.43
X$12770 861 VIA_via1_4
* cell instance $12771 r0 *1 43.415,41.37
X$12771 862 VIA_via1_7
* cell instance $12772 r0 *1 49.685,42.63
X$12772 862 VIA_via1_7
* cell instance $12773 r0 *1 52.535,49.63
X$12773 862 VIA_via2_5
* cell instance $12774 r0 *1 52.345,49.91
X$12774 862 VIA_via2_5
* cell instance $12775 r0 *1 42.275,44.03
X$12775 862 VIA_via2_5
* cell instance $12776 r0 *1 72.295,38.85
X$12776 862 VIA_via2_5
* cell instance $12777 r0 *1 53.485,38.85
X$12777 862 VIA_via2_5
* cell instance $12778 r0 *1 50.255,38.85
X$12778 862 VIA_via2_5
* cell instance $12779 r0 *1 43.415,42.07
X$12779 862 VIA_via2_5
* cell instance $12780 r0 *1 42.275,42.07
X$12780 862 VIA_via2_5
* cell instance $12781 r0 *1 49.685,42.07
X$12781 862 VIA_via2_5
* cell instance $12782 r0 *1 41.705,49.91
X$12782 862 VIA_via2_5
* cell instance $12783 r0 *1 77.995,38.29
X$12783 862 VIA_via2_5
* cell instance $12784 r0 *1 52.535,48.37
X$12784 862 VIA_via1_4
* cell instance $12785 r0 *1 78.185,37.17
X$12785 862 VIA_via1_4
* cell instance $12786 r0 *1 72.295,38.43
X$12786 862 VIA_via1_4
* cell instance $12787 r0 *1 72.295,38.29
X$12787 862 VIA_via2_5
* cell instance $12788 r0 *1 41.705,53.97
X$12788 862 VIA_via1_4
* cell instance $12789 r0 *1 41.895,48.37
X$12789 862 VIA_via1_4
* cell instance $12790 r0 *1 40.375,44.03
X$12790 862 VIA_via1_4
* cell instance $12791 r0 *1 40.375,44.03
X$12791 862 VIA_via2_5
* cell instance $12792 r0 *1 54.055,35.63
X$12792 862 VIA_via1_4
* cell instance $12793 r0 *1 52.345,50.75
X$12793 862 VIA_via1_4
* cell instance $12794 r0 *1 60.135,49.63
X$12794 862 VIA_via1_4
* cell instance $12795 r0 *1 60.135,49.63
X$12795 862 VIA_via2_5
* cell instance $12796 r0 *1 60.135,57.61
X$12796 863 VIA_via1_7
* cell instance $12797 r0 *1 60.135,57.61
X$12797 863 VIA_via2_5
* cell instance $12798 r0 *1 59.945,58.59
X$12798 863 VIA_via1_7
* cell instance $12799 r0 *1 59.945,58.59
X$12799 863 VIA_via2_5
* cell instance $12800 r0 *1 59.185,38.57
X$12800 863 VIA_via1_7
* cell instance $12801 r0 *1 59.185,38.57
X$12801 863 VIA_via2_5
* cell instance $12802 r0 *1 60.895,57.61
X$12802 863 VIA_via2_5
* cell instance $12803 r0 *1 51.585,58.59
X$12803 863 VIA_via2_5
* cell instance $12804 r0 *1 60.705,49.63
X$12804 863 VIA_via2_5
* cell instance $12805 r0 *1 48.925,37.59
X$12805 863 VIA_via2_5
* cell instance $12806 r0 *1 53.675,37.59
X$12806 863 VIA_via2_5
* cell instance $12807 r0 *1 53.675,37.17
X$12807 863 VIA_via1_4
* cell instance $12808 r0 *1 53.675,37.31
X$12808 863 VIA_via2_5
* cell instance $12809 r0 *1 48.925,37.17
X$12809 863 VIA_via1_4
* cell instance $12810 r0 *1 61.655,49.63
X$12810 863 VIA_via1_4
* cell instance $12811 r0 *1 61.655,49.63
X$12811 863 VIA_via2_5
* cell instance $12812 r0 *1 51.585,58.03
X$12812 863 VIA_via1_4
* cell instance $12813 r0 *1 59.735,37.31
X$12813 863 VIA_via3_2
* cell instance $12814 r0 *1 59.735,38.57
X$12814 863 VIA_via3_2
* cell instance $12815 r0 *1 59.735,49.49
X$12815 863 VIA_via3_2
* cell instance $12816 r0 *1 71.535,49.21
X$12816 864 VIA_via1_7
* cell instance $12817 r0 *1 62.415,48.23
X$12817 864 VIA_via2_5
* cell instance $12818 r0 *1 73.055,48.23
X$12818 864 VIA_via2_5
* cell instance $12819 r0 *1 71.535,48.23
X$12819 864 VIA_via2_5
* cell instance $12820 r0 *1 57.095,42.77
X$12820 864 VIA_via1_4
* cell instance $12821 r0 *1 57.095,42.77
X$12821 864 VIA_via2_5
* cell instance $12822 r0 *1 55.575,42.77
X$12822 864 VIA_via1_4
* cell instance $12823 r0 *1 55.575,42.77
X$12823 864 VIA_via2_5
* cell instance $12824 r0 *1 62.415,46.83
X$12824 864 VIA_via1_4
* cell instance $12825 r0 *1 55.385,48.37
X$12825 864 VIA_via1_4
* cell instance $12826 r0 *1 55.385,48.37
X$12826 864 VIA_via2_5
* cell instance $12827 r0 *1 73.245,35.63
X$12827 864 VIA_via1_4
* cell instance $12828 r0 *1 56.935,48.23
X$12828 864 VIA_via3_2
* cell instance $12829 r0 *1 56.935,42.77
X$12829 864 VIA_via3_2
* cell instance $12830 r0 *1 72.675,36.05
X$12830 865 VIA_via1_4
* cell instance $12831 r0 *1 73.055,35.63
X$12831 865 VIA_via1_4
* cell instance $12832 r0 *1 76.475,37.17
X$12832 866 VIA_via1_4
* cell instance $12833 r0 *1 76.475,37.17
X$12833 866 VIA_via2_5
* cell instance $12834 r0 *1 75.525,37.17
X$12834 866 VIA_via1_4
* cell instance $12835 r0 *1 75.525,37.17
X$12835 866 VIA_via2_5
* cell instance $12836 r0 *1 71.915,37.17
X$12836 866 VIA_via1_4
* cell instance $12837 r0 *1 71.915,37.17
X$12837 866 VIA_via2_5
* cell instance $12838 r0 *1 82.935,37.17
X$12838 867 VIA_via2_5
* cell instance $12839 r0 *1 80.655,37.17
X$12839 867 VIA_via1_4
* cell instance $12840 r0 *1 80.655,37.17
X$12840 867 VIA_via2_5
* cell instance $12841 r0 *1 82.935,38.15
X$12841 867 VIA_via1_4
* cell instance $12842 r0 *1 78.945,37.17
X$12842 867 VIA_via1_4
* cell instance $12843 r0 *1 78.945,37.17
X$12843 867 VIA_via2_5
* cell instance $12844 r0 *1 86.165,37.03
X$12844 868 VIA_via2_5
* cell instance $12845 r0 *1 83.885,37.17
X$12845 868 VIA_via1_4
* cell instance $12846 r0 *1 83.885,37.03
X$12846 868 VIA_via2_5
* cell instance $12847 r0 *1 78.375,37.17
X$12847 868 VIA_via1_4
* cell instance $12848 r0 *1 78.375,37.03
X$12848 868 VIA_via2_5
* cell instance $12849 r0 *1 86.165,38.29
X$12849 868 VIA_via1_4
* cell instance $12850 r0 *1 87.495,38.01
X$12850 869 VIA_via1_7
* cell instance $12851 r0 *1 87.115,37.17
X$12851 869 VIA_via1_4
* cell instance $12852 r0 *1 5.225,36.19
X$12852 870 VIA_via1_7
* cell instance $12853 r0 *1 5.225,36.19
X$12853 870 VIA_via2_5
* cell instance $12854 r0 *1 4.085,36.19
X$12854 870 VIA_via2_5
* cell instance $12855 r0 *1 4.085,37.17
X$12855 870 VIA_via1_4
* cell instance $12856 r0 *1 8.075,36.19
X$12856 871 VIA_via1_7
* cell instance $12857 r0 *1 8.075,36.61
X$12857 871 VIA_via2_5
* cell instance $12858 r0 *1 17.195,36.61
X$12858 871 VIA_via2_5
* cell instance $12859 r0 *1 17.195,37.17
X$12859 871 VIA_via1_4
* cell instance $12860 r0 *1 92.815,36.19
X$12860 872 VIA_via1_7
* cell instance $12861 r0 *1 92.815,36.19
X$12861 872 VIA_via2_5
* cell instance $12862 r0 *1 92.245,36.19
X$12862 872 VIA_via2_5
* cell instance $12863 r0 *1 92.245,37.17
X$12863 872 VIA_via1_4
* cell instance $12864 r0 *1 9.595,36.19
X$12864 873 VIA_via1_7
* cell instance $12865 r0 *1 9.595,37.17
X$12865 873 VIA_via2_5
* cell instance $12866 r0 *1 16.055,37.17
X$12866 873 VIA_via1_4
* cell instance $12867 r0 *1 16.055,37.17
X$12867 873 VIA_via2_5
* cell instance $12868 r0 *1 12.635,35.77
X$12868 874 VIA_via2_5
* cell instance $12869 r0 *1 15.295,35.77
X$12869 874 VIA_via1_4
* cell instance $12870 r0 *1 15.295,35.77
X$12870 874 VIA_via2_5
* cell instance $12871 r0 *1 12.635,34.37
X$12871 874 VIA_via1_4
* cell instance $12872 r0 *1 11.875,36.19
X$12872 875 VIA_via1_7
* cell instance $12873 r0 *1 11.875,36.19
X$12873 875 VIA_via2_5
* cell instance $12874 r0 *1 16.625,36.19
X$12874 875 VIA_via2_5
* cell instance $12875 r0 *1 16.625,37.17
X$12875 875 VIA_via1_4
* cell instance $12876 r0 *1 94.905,45.57
X$12876 876 VIA_via2_5
* cell instance $12877 r0 *1 95.475,45.57
X$12877 876 VIA_via2_5
* cell instance $12878 r0 *1 94.715,42.77
X$12878 876 VIA_via2_5
* cell instance $12879 r0 *1 89.205,42.77
X$12879 876 VIA_via2_5
* cell instance $12880 r0 *1 89.205,37.17
X$12880 876 VIA_via2_5
* cell instance $12881 r0 *1 91.865,42.77
X$12881 876 VIA_via1_4
* cell instance $12882 r0 *1 91.865,42.77
X$12882 876 VIA_via2_5
* cell instance $12883 r0 *1 93.195,42.77
X$12883 876 VIA_via1_4
* cell instance $12884 r0 *1 93.195,42.77
X$12884 876 VIA_via2_5
* cell instance $12885 r0 *1 94.905,42.77
X$12885 876 VIA_via1_4
* cell instance $12886 r0 *1 94.905,42.77
X$12886 876 VIA_via2_5
* cell instance $12887 r0 *1 94.715,41.23
X$12887 876 VIA_via1_4
* cell instance $12888 r0 *1 93.765,45.57
X$12888 876 VIA_via1_4
* cell instance $12889 r0 *1 93.765,45.57
X$12889 876 VIA_via2_5
* cell instance $12890 r0 *1 95.475,48.37
X$12890 876 VIA_via1_4
* cell instance $12891 r0 *1 87.875,37.17
X$12891 876 VIA_via1_4
* cell instance $12892 r0 *1 87.875,37.17
X$12892 876 VIA_via2_5
* cell instance $12893 r0 *1 95.095,38.43
X$12893 876 VIA_via1_4
* cell instance $12894 r0 *1 89.205,39.97
X$12894 876 VIA_via1_4
* cell instance $12895 r0 *1 17.955,46.83
X$12895 877 VIA_via1_4
* cell instance $12896 r0 *1 17.955,46.83
X$12896 877 VIA_via2_5
* cell instance $12897 r0 *1 18.145,36.75
X$12897 877 VIA_via1_4
* cell instance $12898 r0 *1 18.145,36.75
X$12898 877 VIA_via2_5
* cell instance $12899 r0 *1 18.295,36.75
X$12899 877 VIA_via3_2
* cell instance $12900 r0 *1 18.295,46.83
X$12900 877 VIA_via3_2
* cell instance $12901 r0 *1 21.375,30.59
X$12901 878 VIA_via1_7
* cell instance $12902 r0 *1 21.375,37.17
X$12902 878 VIA_via2_5
* cell instance $12903 r0 *1 19.285,37.17
X$12903 878 VIA_via1_4
* cell instance $12904 r0 *1 19.285,37.17
X$12904 878 VIA_via2_5
* cell instance $12905 r0 *1 20.805,35.77
X$12905 879 VIA_via1_4
* cell instance $12906 r0 *1 20.805,35.77
X$12906 879 VIA_via2_5
* cell instance $12907 r0 *1 21.755,35.63
X$12907 879 VIA_via1_4
* cell instance $12908 r0 *1 21.755,35.77
X$12908 879 VIA_via2_5
* cell instance $12909 r0 *1 29.545,37.17
X$12909 880 VIA_via1_4
* cell instance $12910 r0 *1 29.545,37.17
X$12910 880 VIA_via2_5
* cell instance $12911 r0 *1 28.595,37.17
X$12911 880 VIA_via1_4
* cell instance $12912 r0 *1 28.595,37.17
X$12912 880 VIA_via2_5
* cell instance $12913 r0 *1 57.285,55.51
X$12913 881 VIA_via2_5
* cell instance $12914 r0 *1 57.285,52.85
X$12914 881 VIA_via2_5
* cell instance $12915 r0 *1 73.815,52.71
X$12915 881 VIA_via2_5
* cell instance $12916 r0 *1 39.995,42.91
X$12916 881 VIA_via2_5
* cell instance $12917 r0 *1 45.315,42.91
X$12917 881 VIA_via2_5
* cell instance $12918 r0 *1 45.315,42.49
X$12918 881 VIA_via2_5
* cell instance $12919 r0 *1 35.435,42.91
X$12919 881 VIA_via2_5
* cell instance $12920 r0 *1 55.195,48.65
X$12920 881 VIA_via2_5
* cell instance $12921 r0 *1 57.285,48.65
X$12921 881 VIA_via2_5
* cell instance $12922 r0 *1 61.655,48.65
X$12922 881 VIA_via2_5
* cell instance $12923 r0 *1 34.485,55.93
X$12923 881 VIA_via2_5
* cell instance $12924 r0 *1 51.395,42.77
X$12924 881 VIA_via1_4
* cell instance $12925 r0 *1 51.395,42.77
X$12925 881 VIA_via2_5
* cell instance $12926 r0 *1 77.995,37.17
X$12926 881 VIA_via1_4
* cell instance $12927 r0 *1 77.995,37.17
X$12927 881 VIA_via2_5
* cell instance $12928 r0 *1 61.655,48.37
X$12928 881 VIA_via1_4
* cell instance $12929 r0 *1 55.195,48.37
X$12929 881 VIA_via1_4
* cell instance $12930 r0 *1 45.315,39.97
X$12930 881 VIA_via1_4
* cell instance $12931 r0 *1 39.995,44.03
X$12931 881 VIA_via1_4
* cell instance $12932 r0 *1 34.485,56.77
X$12932 881 VIA_via1_4
* cell instance $12933 r0 *1 58.235,55.51
X$12933 881 VIA_via1_4
* cell instance $12934 r0 *1 58.235,55.51
X$12934 881 VIA_via2_5
* cell instance $12935 r0 *1 35.435,41.23
X$12935 881 VIA_via1_4
* cell instance $12936 r0 *1 32.395,42.77
X$12936 881 VIA_via1_4
* cell instance $12937 r0 *1 32.395,42.77
X$12937 881 VIA_via2_5
* cell instance $12938 r0 *1 73.815,53.97
X$12938 881 VIA_via1_4
* cell instance $12939 r0 *1 73.815,53.97
X$12939 881 VIA_via2_5
* cell instance $12940 r0 *1 54.975,42.77
X$12940 881 VIA_via3_2
* cell instance $12941 r0 *1 54.975,48.65
X$12941 881 VIA_via3_2
* cell instance $12942 r0 *1 78.215,53.97
X$12942 881 VIA_via3_2
* cell instance $12943 r0 *1 78.215,37.17
X$12943 881 VIA_via3_2
* cell instance $12944 r0 *1 77.995,36.61
X$12944 882 VIA_via1_7
* cell instance $12945 r0 *1 77.995,35.63
X$12945 882 VIA_via1_4
* cell instance $12946 r0 *1 72.295,36.61
X$12946 883 VIA_via1_7
* cell instance $12947 r0 *1 72.295,35.63
X$12947 883 VIA_via1_4
* cell instance $12948 r0 *1 60.325,36.19
X$12948 884 VIA_via1_7
* cell instance $12949 r0 *1 60.325,36.19
X$12949 884 VIA_via2_5
* cell instance $12950 r0 *1 58.995,36.19
X$12950 884 VIA_via2_5
* cell instance $12951 r0 *1 58.995,37.17
X$12951 884 VIA_via1_4
* cell instance $12952 r0 *1 45.695,37.17
X$12952 885 VIA_via1_4
* cell instance $12953 r0 *1 45.695,37.17
X$12953 885 VIA_via2_5
* cell instance $12954 r0 *1 45.125,37.17
X$12954 885 VIA_via1_4
* cell instance $12955 r0 *1 45.125,37.17
X$12955 885 VIA_via2_5
* cell instance $12956 r0 *1 57.855,36.19
X$12956 886 VIA_via1_7
* cell instance $12957 r0 *1 57.855,36.19
X$12957 886 VIA_via2_5
* cell instance $12958 r0 *1 55.765,36.19
X$12958 886 VIA_via2_5
* cell instance $12959 r0 *1 55.765,37.17
X$12959 886 VIA_via1_4
* cell instance $12960 r0 *1 7.315,40.11
X$12960 887 VIA_via2_5
* cell instance $12961 r0 *1 5.225,40.11
X$12961 887 VIA_via2_5
* cell instance $12962 r0 *1 7.315,41.23
X$12962 887 VIA_via1_4
* cell instance $12963 r0 *1 4.845,38.29
X$12963 887 VIA_via1_4
* cell instance $12964 r0 *1 5.225,38.43
X$12964 887 VIA_via1_4
* cell instance $12965 r0 *1 16.625,39.41
X$12965 888 VIA_via1_7
* cell instance $12966 r0 *1 16.625,39.41
X$12966 888 VIA_via2_5
* cell instance $12967 r0 *1 17.575,39.41
X$12967 888 VIA_via2_5
* cell instance $12968 r0 *1 17.575,38.43
X$12968 888 VIA_via1_4
* cell instance $12969 r0 *1 17.955,36.19
X$12969 889 VIA_via1_7
* cell instance $12970 r0 *1 18.335,38.43
X$12970 889 VIA_via1_4
* cell instance $12971 r0 *1 16.055,51.03
X$12971 890 VIA_via1_7
* cell instance $12972 r0 *1 16.055,50.75
X$12972 890 VIA_via2_5
* cell instance $12973 r0 *1 18.525,52.15
X$12973 890 VIA_via2_5
* cell instance $12974 r0 *1 19.855,52.15
X$12974 890 VIA_via2_5
* cell instance $12975 r0 *1 18.525,50.75
X$12975 890 VIA_via2_5
* cell instance $12976 r0 *1 19.855,53.97
X$12976 890 VIA_via1_4
* cell instance $12977 r0 *1 18.335,38.15
X$12977 890 VIA_via1_4
* cell instance $12978 r0 *1 52.535,38.15
X$12978 891 VIA_via2_5
* cell instance $12979 r0 *1 45.885,40.53
X$12979 891 VIA_via2_5
* cell instance $12980 r0 *1 45.885,38.01
X$12980 891 VIA_via2_5
* cell instance $12981 r0 *1 39.235,40.25
X$12981 891 VIA_via2_5
* cell instance $12982 r0 *1 56.335,46.55
X$12982 891 VIA_via2_5
* cell instance $12983 r0 *1 57.095,46.55
X$12983 891 VIA_via2_5
* cell instance $12984 r0 *1 17.765,42.35
X$12984 891 VIA_via2_5
* cell instance $12985 r0 *1 17.735,42.35
X$12985 891 VIA_via3_2
* cell instance $12986 r0 *1 26.695,38.99
X$12986 891 VIA_via2_5
* cell instance $12987 r0 *1 25.365,38.99
X$12987 891 VIA_via2_5
* cell instance $12988 r0 *1 25.365,37.87
X$12988 891 VIA_via2_5
* cell instance $12989 r0 *1 35.625,41.09
X$12989 891 VIA_via2_5
* cell instance $12990 r0 *1 26.695,41.09
X$12990 891 VIA_via2_5
* cell instance $12991 r0 *1 35.625,40.25
X$12991 891 VIA_via2_5
* cell instance $12992 r0 *1 17.955,38.01
X$12992 891 VIA_via2_5
* cell instance $12993 r0 *1 56.335,38.01
X$12993 891 VIA_via2_5
* cell instance $12994 r0 *1 56.335,42.35
X$12994 891 VIA_via1_4
* cell instance $12995 r0 *1 56.335,43.19
X$12995 891 VIA_via1_7
* cell instance $12996 r0 *1 52.535,38.43
X$12996 891 VIA_via1_4
* cell instance $12997 r0 *1 57.095,46.83
X$12997 891 VIA_via1_4
* cell instance $12998 r0 *1 39.045,44.03
X$12998 891 VIA_via1_4
* cell instance $12999 r0 *1 45.885,38.43
X$12999 891 VIA_via1_4
* cell instance $13000 r0 *1 17.955,38.43
X$13000 891 VIA_via1_4
* cell instance $13001 r0 *1 17.955,38.43
X$13001 891 VIA_via2_5
* cell instance $13002 r0 *1 35.625,39.97
X$13002 891 VIA_via1_4
* cell instance $13003 r0 *1 26.505,38.43
X$13003 891 VIA_via1_4
* cell instance $13004 r0 *1 31.255,41.23
X$13004 891 VIA_via1_4
* cell instance $13005 r0 *1 31.255,41.09
X$13005 891 VIA_via2_5
* cell instance $13006 r0 *1 17.765,39.97
X$13006 891 VIA_via1_4
* cell instance $13007 r0 *1 17.765,39.97
X$13007 891 VIA_via2_5
* cell instance $13008 r0 *1 17.735,39.97
X$13008 891 VIA_via3_2
* cell instance $13009 r0 *1 17.765,44.03
X$13009 891 VIA_via1_4
* cell instance $13010 r0 *1 17.735,38.43
X$13010 891 VIA_via3_2
* cell instance $13011 r0 *1 19.475,37.59
X$13011 892 VIA_via1_7
* cell instance $13012 r0 *1 18.905,39.83
X$13012 892 VIA_via2_5
* cell instance $13013 r0 *1 18.145,39.97
X$13013 892 VIA_via1_4
* cell instance $13014 r0 *1 18.145,39.97
X$13014 892 VIA_via2_5
* cell instance $13015 r0 *1 19.095,70.49
X$13015 893 VIA_via2_5
* cell instance $13016 r0 *1 20.235,70.49
X$13016 893 VIA_via2_5
* cell instance $13017 r0 *1 20.425,70.49
X$13017 893 VIA_via2_5
* cell instance $13018 r0 *1 17.005,45.85
X$13018 893 VIA_via2_5
* cell instance $13019 r0 *1 16.895,45.85
X$13019 893 VIA_via3_2
* cell instance $13020 r0 *1 24.795,39.83
X$13020 893 VIA_via2_5
* cell instance $13021 r0 *1 19.475,39.13
X$13021 893 VIA_via2_5
* cell instance $13022 r0 *1 20.425,60.69
X$13022 893 VIA_via2_5
* cell instance $13023 r0 *1 28.215,60.69
X$13023 893 VIA_via2_5
* cell instance $13024 r0 *1 27.835,57.47
X$13024 893 VIA_via2_5
* cell instance $13025 r0 *1 28.215,57.61
X$13025 893 VIA_via2_5
* cell instance $13026 r0 *1 31.635,59.15
X$13026 893 VIA_via1_4
* cell instance $13027 r0 *1 31.635,59.15
X$13027 893 VIA_via2_5
* cell instance $13028 r0 *1 27.835,56.77
X$13028 893 VIA_via1_4
* cell instance $13029 r0 *1 20.425,62.37
X$13029 893 VIA_via1_4
* cell instance $13030 r0 *1 19.095,72.03
X$13030 893 VIA_via1_4
* cell instance $13031 r0 *1 20.425,74.83
X$13031 893 VIA_via1_4
* cell instance $13032 r0 *1 19.475,38.43
X$13032 893 VIA_via1_4
* cell instance $13033 r0 *1 19.475,38.29
X$13033 893 VIA_via2_5
* cell instance $13034 r0 *1 24.795,38.43
X$13034 893 VIA_via1_4
* cell instance $13035 r0 *1 24.795,38.29
X$13035 893 VIA_via2_5
* cell instance $13036 r0 *1 30.115,39.97
X$13036 893 VIA_via1_4
* cell instance $13037 r0 *1 30.115,39.83
X$13037 893 VIA_via2_5
* cell instance $13038 r0 *1 16.625,48.37
X$13038 893 VIA_via1_4
* cell instance $13039 r0 *1 16.625,48.37
X$13039 893 VIA_via2_5
* cell instance $13040 r0 *1 16.625,39.97
X$13040 893 VIA_via1_4
* cell instance $13041 r0 *1 16.625,39.97
X$13041 893 VIA_via2_5
* cell instance $13042 r0 *1 17.005,45.57
X$13042 893 VIA_via1_4
* cell instance $13043 r0 *1 29.775,57.47
X$13043 893 VIA_via3_2
* cell instance $13044 r0 *1 29.775,58.59
X$13044 893 VIA_via3_2
* cell instance $13045 r0 *1 29.775,39.83
X$13045 893 VIA_via3_2
* cell instance $13046 r0 *1 16.895,48.37
X$13046 893 VIA_via3_2
* cell instance $13047 r0 *1 17.175,39.97
X$13047 893 VIA_via3_2
* cell instance $13048 r0 *1 21.945,38.15
X$13048 894 VIA_via2_5
* cell instance $13049 r0 *1 24.415,38.15
X$13049 894 VIA_via2_5
* cell instance $13050 r0 *1 23.845,38.15
X$13050 894 VIA_via2_5
* cell instance $13051 r0 *1 24.415,37.45
X$13051 894 VIA_via1_4
* cell instance $13052 r0 *1 23.845,38.43
X$13052 894 VIA_via1_4
* cell instance $13053 r0 *1 21.945,38.43
X$13053 894 VIA_via1_4
* cell instance $13054 r0 *1 26.125,37.59
X$13054 895 VIA_via1_7
* cell instance $13055 r0 *1 26.125,38.15
X$13055 895 VIA_via2_5
* cell instance $13056 r0 *1 26.885,38.43
X$13056 895 VIA_via1_4
* cell instance $13057 r0 *1 26.885,38.43
X$13057 895 VIA_via2_5
* cell instance $13058 r0 *1 27.075,37.59
X$13058 896 VIA_via1_7
* cell instance $13059 r0 *1 26.695,38.395
X$13059 896 VIA_via1_4
* cell instance $13060 r0 *1 26.695,42.77
X$13060 897 VIA_via2_5
* cell instance $13061 r0 *1 27.075,42.77
X$13061 897 VIA_via2_5
* cell instance $13062 r0 *1 25.555,49.63
X$13062 897 VIA_via1_4
* cell instance $13063 r0 *1 26.885,38.15
X$13063 897 VIA_via1_4
* cell instance $13064 r0 *1 25.935,46.97
X$13064 897 VIA_via1_4
* cell instance $13065 r0 *1 26.505,46.97
X$13065 897 VIA_via1_7
* cell instance $13066 r0 *1 27.645,37.45
X$13066 898 VIA_via2_5
* cell instance $13067 r0 *1 29.165,37.45
X$13067 898 VIA_via2_5
* cell instance $13068 r0 *1 27.645,37.17
X$13068 898 VIA_via1_4
* cell instance $13069 r0 *1 29.165,38.43
X$13069 898 VIA_via1_4
* cell instance $13070 r0 *1 31.825,37.45
X$13070 898 VIA_via1_4
* cell instance $13071 r0 *1 31.825,37.45
X$13071 898 VIA_via2_5
* cell instance $13072 r0 *1 37.145,38.43
X$13072 899 VIA_via1_4
* cell instance $13073 r0 *1 37.145,38.29
X$13073 899 VIA_via2_5
* cell instance $13074 r0 *1 41.895,38.29
X$13074 899 VIA_via1_4
* cell instance $13075 r0 *1 41.895,38.29
X$13075 899 VIA_via2_5
* cell instance $13076 r0 *1 35.815,38.43
X$13076 899 VIA_via1_4
* cell instance $13077 r0 *1 35.815,38.29
X$13077 899 VIA_via2_5
* cell instance $13078 r0 *1 36.955,38.57
X$13078 900 VIA_via1_7
* cell instance $13079 r0 *1 28.975,38.57
X$13079 900 VIA_via1_7
* cell instance $13080 r0 *1 36.575,42.63
X$13080 900 VIA_via1_7
* cell instance $13081 r0 *1 14.725,39.83
X$13081 900 VIA_via1_7
* cell instance $13082 r0 *1 59.565,45.43
X$13082 900 VIA_via1_7
* cell instance $13083 r0 *1 23.085,38.57
X$13083 900 VIA_via1_7
* cell instance $13084 r0 *1 36.955,38.85
X$13084 900 VIA_via2_5
* cell instance $13085 r0 *1 44.175,37.87
X$13085 900 VIA_via2_5
* cell instance $13086 r0 *1 44.175,39.83
X$13086 900 VIA_via2_5
* cell instance $13087 r0 *1 48.925,41.09
X$13087 900 VIA_via2_5
* cell instance $13088 r0 *1 48.925,37.87
X$13088 900 VIA_via2_5
* cell instance $13089 r0 *1 59.565,46.69
X$13089 900 VIA_via2_5
* cell instance $13090 r0 *1 14.725,40.39
X$13090 900 VIA_via2_5
* cell instance $13091 r0 *1 18.335,40.39
X$13091 900 VIA_via2_5
* cell instance $13092 r0 *1 50.065,46.69
X$13092 900 VIA_via2_5
* cell instance $13093 r0 *1 23.275,38.85
X$13093 900 VIA_via2_5
* cell instance $13094 r0 *1 28.975,38.85
X$13094 900 VIA_via2_5
* cell instance $13095 r0 *1 36.765,39.83
X$13095 900 VIA_via2_5
* cell instance $13096 r0 *1 23.275,40.39
X$13096 900 VIA_via2_5
* cell instance $13097 r0 *1 36.765,38.85
X$13097 900 VIA_via2_5
* cell instance $13098 r0 *1 50.065,41.23
X$13098 900 VIA_via1_4
* cell instance $13099 r0 *1 50.065,41.09
X$13099 900 VIA_via2_5
* cell instance $13100 r0 *1 53.675,46.83
X$13100 900 VIA_via1_4
* cell instance $13101 r0 *1 53.675,46.69
X$13101 900 VIA_via2_5
* cell instance $13102 r0 *1 59.565,43.05
X$13102 900 VIA_via1_4
* cell instance $13103 r0 *1 43.985,37.17
X$13103 900 VIA_via1_4
* cell instance $13104 r0 *1 18.335,39.97
X$13104 900 VIA_via1_4
* cell instance $13105 r0 *1 45.315,48.51
X$13105 901 VIA_via2_5
* cell instance $13106 r0 *1 45.505,38.71
X$13106 901 VIA_via2_5
* cell instance $13107 r0 *1 46.075,38.15
X$13107 901 VIA_via2_5
* cell instance $13108 r0 *1 46.265,38.15
X$13108 901 VIA_via1_4
* cell instance $13109 r0 *1 44.555,49.49
X$13109 901 VIA_via1_4
* cell instance $13110 r0 *1 44.555,48.37
X$13110 901 VIA_via1_4
* cell instance $13111 r0 *1 44.555,48.51
X$13111 901 VIA_via2_5
* cell instance $13112 r0 *1 51.395,42.21
X$13112 902 VIA_via1_7
* cell instance $13113 r0 *1 51.965,38.43
X$13113 902 VIA_via1_4
* cell instance $13114 r0 *1 52.345,37.59
X$13114 903 VIA_via1_7
* cell instance $13115 r0 *1 52.725,38.43
X$13115 903 VIA_via1_4
* cell instance $13116 r0 *1 54.435,37.73
X$13116 904 VIA_via2_5
* cell instance $13117 r0 *1 56.525,37.73
X$13117 904 VIA_via2_5
* cell instance $13118 r0 *1 56.905,38.43
X$13118 904 VIA_via1_4
* cell instance $13119 r0 *1 54.435,37.17
X$13119 904 VIA_via1_4
* cell instance $13120 r0 *1 56.525,38.15
X$13120 904 VIA_via1_4
* cell instance $13121 r0 *1 57.475,38.43
X$13121 905 VIA_via1_4
* cell instance $13122 r0 *1 58.045,37.45
X$13122 905 VIA_via1_4
* cell instance $13123 r0 *1 57.475,35.63
X$13123 905 VIA_via1_4
* cell instance $13124 r0 *1 66.215,38.43
X$13124 906 VIA_via1_4
* cell instance $13125 r0 *1 66.215,38.43
X$13125 906 VIA_via2_5
* cell instance $13126 r0 *1 66.785,39.97
X$13126 906 VIA_via1_4
* cell instance $13127 r0 *1 66.595,38.43
X$13127 906 VIA_via1_4
* cell instance $13128 r0 *1 66.595,38.43
X$13128 906 VIA_via2_5
* cell instance $13129 r0 *1 86.735,40.81
X$13129 907 VIA_via1_7
* cell instance $13130 r0 *1 86.735,41.79
X$13130 907 VIA_via1_7
* cell instance $13131 r0 *1 86.735,42.49
X$13131 907 VIA_via2_5
* cell instance $13132 r0 *1 86.735,38.43
X$13132 907 VIA_via2_5
* cell instance $13133 r0 *1 77.045,43.89
X$13133 907 VIA_via2_5
* cell instance $13134 r0 *1 76.285,43.89
X$13134 907 VIA_via2_5
* cell instance $13135 r0 *1 77.045,42.49
X$13135 907 VIA_via2_5
* cell instance $13136 r0 *1 73.245,46.55
X$13136 907 VIA_via2_5
* cell instance $13137 r0 *1 75.905,46.55
X$13137 907 VIA_via2_5
* cell instance $13138 r0 *1 76.285,46.55
X$13138 907 VIA_via2_5
* cell instance $13139 r0 *1 81.225,42.49
X$13139 907 VIA_via2_5
* cell instance $13140 r0 *1 80.655,42.49
X$13140 907 VIA_via2_5
* cell instance $13141 r0 *1 77.045,42.77
X$13141 907 VIA_via1_4
* cell instance $13142 r0 *1 76.855,38.43
X$13142 907 VIA_via1_4
* cell instance $13143 r0 *1 81.225,42.77
X$13143 907 VIA_via1_4
* cell instance $13144 r0 *1 80.655,39.97
X$13144 907 VIA_via1_4
* cell instance $13145 r0 *1 74.765,44.03
X$13145 907 VIA_via1_4
* cell instance $13146 r0 *1 74.765,43.89
X$13146 907 VIA_via2_5
* cell instance $13147 r0 *1 76.285,45.57
X$13147 907 VIA_via1_4
* cell instance $13148 r0 *1 75.905,48.37
X$13148 907 VIA_via1_4
* cell instance $13149 r0 *1 73.245,46.83
X$13149 907 VIA_via1_4
* cell instance $13150 r0 *1 87.115,38.43
X$13150 907 VIA_via1_4
* cell instance $13151 r0 *1 87.115,38.43
X$13151 907 VIA_via2_5
* cell instance $13152 r0 *1 88.445,38.43
X$13152 907 VIA_via1_4
* cell instance $13153 r0 *1 88.445,38.29
X$13153 907 VIA_via2_5
* cell instance $13154 r0 *1 81.035,37.59
X$13154 908 VIA_via1_7
* cell instance $13155 r0 *1 80.655,38.43
X$13155 908 VIA_via1_4
* cell instance $13156 r0 *1 84.265,37.59
X$13156 909 VIA_via1_7
* cell instance $13157 r0 *1 83.885,38.43
X$13157 909 VIA_via1_4
* cell instance $13158 r0 *1 89.395,37.87
X$13158 910 VIA_via2_5
* cell instance $13159 r0 *1 90.345,37.87
X$13159 910 VIA_via2_5
* cell instance $13160 r0 *1 86.545,37.87
X$13160 910 VIA_via2_5
* cell instance $13161 r0 *1 86.545,38.395
X$13161 910 VIA_via1_4
* cell instance $13162 r0 *1 90.345,38.43
X$13162 910 VIA_via1_4
* cell instance $13163 r0 *1 89.395,37.45
X$13163 910 VIA_via1_4
* cell instance $13164 r0 *1 90.725,38.43
X$13164 911 VIA_via2_5
* cell instance $13165 r0 *1 87.875,38.43
X$13165 911 VIA_via1_4
* cell instance $13166 r0 *1 87.875,38.43
X$13166 911 VIA_via2_5
* cell instance $13167 r0 *1 89.775,38.43
X$13167 911 VIA_via1_4
* cell instance $13168 r0 *1 89.775,38.43
X$13168 911 VIA_via2_5
* cell instance $13169 r0 *1 90.725,39.55
X$13169 911 VIA_via1_4
* cell instance $13170 r0 *1 90.725,38.01
X$13170 912 VIA_via1_7
* cell instance $13171 r0 *1 90.535,37.17
X$13171 912 VIA_via1_4
* cell instance $13172 r0 *1 90.725,37.59
X$13172 913 VIA_via1_7
* cell instance $13173 r0 *1 91.105,38.43
X$13173 913 VIA_via1_4
* cell instance $13174 r0 *1 92.435,55.23
X$13174 914 VIA_via2_5
* cell instance $13175 r0 *1 93.385,54.95
X$13175 914 VIA_via2_5
* cell instance $13176 r0 *1 92.435,54.95
X$13176 914 VIA_via2_5
* cell instance $13177 r0 *1 92.055,38.15
X$13177 914 VIA_via1_4
* cell instance $13178 r0 *1 92.055,38.15
X$13178 914 VIA_via2_5
* cell instance $13179 r0 *1 92.055,56.77
X$13179 914 VIA_via1_4
* cell instance $13180 r0 *1 92.055,56.77
X$13180 914 VIA_via2_5
* cell instance $13181 r0 *1 93.385,55.16
X$13181 914 VIA_via1_4
* cell instance $13182 r0 *1 92.215,56.77
X$13182 914 VIA_via3_2
* cell instance $13183 r0 *1 92.215,55.23
X$13183 914 VIA_via3_2
* cell instance $13184 r0 *1 92.215,38.15
X$13184 914 VIA_via3_2
* cell instance $13185 r0 *1 7.695,37.59
X$13185 915 VIA_via1_7
* cell instance $13186 r0 *1 7.695,38.01
X$13186 915 VIA_via2_5
* cell instance $13187 r0 *1 16.625,38.01
X$13187 915 VIA_via2_5
* cell instance $13188 r0 *1 16.625,38.43
X$13188 915 VIA_via1_4
* cell instance $13189 r0 *1 11.875,38.43
X$13189 916 VIA_via1_4
* cell instance $13190 r0 *1 11.875,38.29
X$13190 916 VIA_via2_5
* cell instance $13191 r0 *1 15.485,38.29
X$13191 916 VIA_via1_4
* cell instance $13192 r0 *1 15.485,38.29
X$13192 916 VIA_via2_5
* cell instance $13193 r0 *1 16.245,37.59
X$13193 917 VIA_via1_7
* cell instance $13194 r0 *1 18.145,37.87
X$13194 917 VIA_via2_5
* cell instance $13195 r0 *1 16.245,37.87
X$13195 917 VIA_via2_5
* cell instance $13196 r0 *1 18.145,38.43
X$13196 917 VIA_via1_4
* cell instance $13197 r0 *1 17.385,37.59
X$13197 918 VIA_via1_7
* cell instance $13198 r0 *1 17.385,37.59
X$13198 918 VIA_via2_5
* cell instance $13199 r0 *1 17.955,42.07
X$13199 918 VIA_via2_5
* cell instance $13200 r0 *1 17.955,44.03
X$13200 918 VIA_via1_4
* cell instance $13201 r0 *1 16.895,42.07
X$13201 918 VIA_via3_2
* cell instance $13202 r0 *1 16.895,37.59
X$13202 918 VIA_via3_2
* cell instance $13203 r0 *1 77.615,37.17
X$13203 919 VIA_via1_4
* cell instance $13204 r0 *1 77.615,37.31
X$13204 919 VIA_via2_5
* cell instance $13205 r0 *1 79.325,37.31
X$13205 919 VIA_via1_4
* cell instance $13206 r0 *1 79.325,37.31
X$13206 919 VIA_via2_5
* cell instance $13207 r0 *1 17.385,38.36
X$13207 920 VIA_via1_4
* cell instance $13208 r0 *1 17.385,38.29
X$13208 920 VIA_via2_5
* cell instance $13209 r0 *1 16.245,38.29
X$13209 920 VIA_via1_4
* cell instance $13210 r0 *1 16.245,38.29
X$13210 920 VIA_via2_5
* cell instance $13211 r0 *1 73.245,37.17
X$13211 921 VIA_via1_4
* cell instance $13212 r0 *1 73.245,37.31
X$13212 921 VIA_via2_5
* cell instance $13213 r0 *1 76.855,37.31
X$13213 921 VIA_via1_4
* cell instance $13214 r0 *1 76.855,37.31
X$13214 921 VIA_via2_5
* cell instance $13215 r0 *1 18.905,37.59
X$13215 922 VIA_via1_7
* cell instance $13216 r0 *1 18.905,37.59
X$13216 922 VIA_via2_5
* cell instance $13217 r0 *1 18.335,43.05
X$13217 922 VIA_via2_5
* cell instance $13218 r0 *1 20.235,43.05
X$13218 922 VIA_via2_5
* cell instance $13219 r0 *1 20.235,37.59
X$13219 922 VIA_via2_5
* cell instance $13220 r0 *1 18.145,44.03
X$13220 922 VIA_via1_4
* cell instance $13221 r0 *1 63.935,38.43
X$13221 923 VIA_via1_4
* cell instance $13222 r0 *1 63.935,38.29
X$13222 923 VIA_via2_5
* cell instance $13223 r0 *1 67.545,38.29
X$13223 923 VIA_via1_4
* cell instance $13224 r0 *1 67.545,38.29
X$13224 923 VIA_via2_5
* cell instance $13225 r0 *1 22.895,38.01
X$13225 924 VIA_via1_7
* cell instance $13226 r0 *1 22.895,38.01
X$13226 924 VIA_via2_5
* cell instance $13227 r0 *1 22.135,38.01
X$13227 924 VIA_via2_5
* cell instance $13228 r0 *1 22.135,37.17
X$13228 924 VIA_via1_4
* cell instance $13229 r0 *1 55.955,51.31
X$13229 925 VIA_via2_5
* cell instance $13230 r0 *1 53.485,51.31
X$13230 925 VIA_via2_5
* cell instance $13231 r0 *1 53.295,38.15
X$13231 925 VIA_via2_5
* cell instance $13232 r0 *1 52.915,38.15
X$13232 925 VIA_via1_4
* cell instance $13233 r0 *1 52.915,38.15
X$13233 925 VIA_via2_5
* cell instance $13234 r0 *1 53.865,51.17
X$13234 925 VIA_via1_4
* cell instance $13235 r0 *1 53.865,51.31
X$13235 925 VIA_via2_5
* cell instance $13236 r0 *1 55.955,52.43
X$13236 925 VIA_via1_4
* cell instance $13237 r0 *1 35.435,38.01
X$13237 926 VIA_via1_7
* cell instance $13238 r0 *1 35.435,38.01
X$13238 926 VIA_via2_5
* cell instance $13239 r0 *1 35.815,38.01
X$13239 926 VIA_via2_5
* cell instance $13240 r0 *1 35.815,37.17
X$13240 926 VIA_via1_4
* cell instance $13241 r0 *1 45.885,37.59
X$13241 927 VIA_via1_7
* cell instance $13242 r0 *1 45.885,37.73
X$13242 927 VIA_via2_5
* cell instance $13243 r0 *1 45.505,37.73
X$13243 927 VIA_via2_5
* cell instance $13244 r0 *1 45.505,38.43
X$13244 927 VIA_via1_4
* cell instance $13245 r0 *1 10.355,39.97
X$13245 928 VIA_via1_4
* cell instance $13246 r0 *1 9.405,41.23
X$13246 928 VIA_via1_4
* cell instance $13247 r0 *1 9.405,38.85
X$13247 928 VIA_via1_4
* cell instance $13248 r0 *1 34.295,38.57
X$13248 929 VIA_via1_7
* cell instance $13249 r0 *1 34.295,38.71
X$13249 929 VIA_via2_5
* cell instance $13250 r0 *1 46.645,38.57
X$13250 929 VIA_via1_7
* cell instance $13251 r0 *1 43.605,38.57
X$13251 929 VIA_via1_7
* cell instance $13252 r0 *1 43.605,38.71
X$13252 929 VIA_via2_5
* cell instance $13253 r0 *1 27.265,38.57
X$13253 929 VIA_via1_7
* cell instance $13254 r0 *1 21.755,38.57
X$13254 929 VIA_via1_7
* cell instance $13255 r0 *1 21.755,38.71
X$13255 929 VIA_via2_5
* cell instance $13256 r0 *1 12.445,39.83
X$13256 929 VIA_via1_7
* cell instance $13257 r0 *1 46.455,38.99
X$13257 929 VIA_via2_5
* cell instance $13258 r0 *1 46.645,38.99
X$13258 929 VIA_via2_5
* cell instance $13259 r0 *1 14.725,48.51
X$13259 929 VIA_via2_5
* cell instance $13260 r0 *1 27.455,38.71
X$13260 929 VIA_via2_5
* cell instance $13261 r0 *1 12.635,39.13
X$13261 929 VIA_via2_5
* cell instance $13262 r0 *1 15.105,39.13
X$13262 929 VIA_via2_5
* cell instance $13263 r0 *1 19.855,38.99
X$13263 929 VIA_via2_5
* cell instance $13264 r0 *1 35.815,46.83
X$13264 929 VIA_via1_4
* cell instance $13265 r0 *1 35.815,46.83
X$13265 929 VIA_via2_5
* cell instance $13266 r0 *1 46.455,45.15
X$13266 929 VIA_via1_4
* cell instance $13267 r0 *1 19.665,39.97
X$13267 929 VIA_via1_4
* cell instance $13268 r0 *1 14.915,44.03
X$13268 929 VIA_via1_4
* cell instance $13269 r0 *1 12.635,48.37
X$13269 929 VIA_via1_4
* cell instance $13270 r0 *1 12.635,48.51
X$13270 929 VIA_via2_5
* cell instance $13271 r0 *1 36.775,46.83
X$13271 929 VIA_via3_2
* cell instance $13272 r0 *1 36.775,38.71
X$13272 929 VIA_via3_2
* cell instance $13273 r0 *1 14.535,38.85
X$13273 930 VIA_via2_5
* cell instance $13274 r0 *1 14.155,38.85
X$13274 930 VIA_via1_4
* cell instance $13275 r0 *1 14.155,38.85
X$13275 930 VIA_via2_5
* cell instance $13276 r0 *1 14.535,38.43
X$13276 930 VIA_via1_4
* cell instance $13277 r0 *1 14.915,39.97
X$13277 930 VIA_via1_4
* cell instance $13278 r0 *1 17.005,38.99
X$13278 931 VIA_via1_7
* cell instance $13279 r0 *1 16.815,44.73
X$13279 931 VIA_via2_5
* cell instance $13280 r0 *1 17.765,44.73
X$13280 931 VIA_via2_5
* cell instance $13281 r0 *1 17.765,46.83
X$13281 931 VIA_via1_4
* cell instance $13282 r0 *1 45.125,39.97
X$13282 932 VIA_via2_5
* cell instance $13283 r0 *1 37.715,40.11
X$13283 932 VIA_via2_5
* cell instance $13284 r0 *1 16.815,45.01
X$13284 932 VIA_via2_5
* cell instance $13285 r0 *1 17.005,44.87
X$13285 932 VIA_via2_5
* cell instance $13286 r0 *1 30.495,40.81
X$13286 932 VIA_via2_5
* cell instance $13287 r0 *1 34.865,40.81
X$13287 932 VIA_via2_5
* cell instance $13288 r0 *1 25.745,41.23
X$13288 932 VIA_via2_5
* cell instance $13289 r0 *1 51.775,39.97
X$13289 932 VIA_via2_5
* cell instance $13290 r0 *1 51.775,38.43
X$13290 932 VIA_via1_4
* cell instance $13291 r0 *1 51.775,46.55
X$13291 932 VIA_via1_4
* cell instance $13292 r0 *1 38.285,44.03
X$13292 932 VIA_via1_4
* cell instance $13293 r0 *1 45.125,38.43
X$13293 932 VIA_via1_4
* cell instance $13294 r0 *1 17.195,38.43
X$13294 932 VIA_via1_4
* cell instance $13295 r0 *1 17.195,38.57
X$13295 932 VIA_via2_5
* cell instance $13296 r0 *1 25.745,38.43
X$13296 932 VIA_via1_4
* cell instance $13297 r0 *1 25.745,38.57
X$13297 932 VIA_via2_5
* cell instance $13298 r0 *1 30.495,41.23
X$13298 932 VIA_via1_4
* cell instance $13299 r0 *1 30.495,41.23
X$13299 932 VIA_via2_5
* cell instance $13300 r0 *1 34.865,39.97
X$13300 932 VIA_via1_4
* cell instance $13301 r0 *1 34.865,40.11
X$13301 932 VIA_via2_5
* cell instance $13302 r0 *1 16.815,46.83
X$13302 932 VIA_via1_4
* cell instance $13303 r0 *1 17.005,39.97
X$13303 932 VIA_via1_4
* cell instance $13304 r0 *1 17.005,44.03
X$13304 932 VIA_via1_4
* cell instance $13305 r0 *1 19.475,39.55
X$13305 933 VIA_via1_4
* cell instance $13306 r0 *1 19.095,38.43
X$13306 933 VIA_via1_4
* cell instance $13307 r0 *1 21.565,39.97
X$13307 934 VIA_via2_5
* cell instance $13308 r0 *1 21.565,40.95
X$13308 934 VIA_via1_4
* cell instance $13309 r0 *1 19.095,39.97
X$13309 934 VIA_via1_4
* cell instance $13310 r0 *1 19.095,39.97
X$13310 934 VIA_via2_5
* cell instance $13311 r0 *1 19.855,39.97
X$13311 934 VIA_via1_4
* cell instance $13312 r0 *1 19.855,39.97
X$13312 934 VIA_via2_5
* cell instance $13313 r0 *1 26.125,39.69
X$13313 935 VIA_via1_4
* cell instance $13314 r0 *1 25.935,38.43
X$13314 935 VIA_via1_4
* cell instance $13315 r0 *1 26.125,42.21
X$13315 936 VIA_via1_7
* cell instance $13316 r0 *1 25.935,39.97
X$13316 936 VIA_via1_4
* cell instance $13317 r0 *1 26.885,39.97
X$13317 937 VIA_via2_5
* cell instance $13318 r0 *1 22.325,60.55
X$13318 937 VIA_via2_5
* cell instance $13319 r0 *1 21.755,60.55
X$13319 937 VIA_via2_5
* cell instance $13320 r0 *1 26.695,57.19
X$13320 937 VIA_via2_5
* cell instance $13321 r0 *1 28.405,60.55
X$13321 937 VIA_via2_5
* cell instance $13322 r0 *1 28.405,59.29
X$13322 937 VIA_via2_5
* cell instance $13323 r0 *1 28.405,57.05
X$13323 937 VIA_via2_5
* cell instance $13324 r0 *1 33.915,59.29
X$13324 937 VIA_via1_4
* cell instance $13325 r0 *1 33.915,59.29
X$13325 937 VIA_via2_5
* cell instance $13326 r0 *1 28.405,56.77
X$13326 937 VIA_via1_4
* cell instance $13327 r0 *1 21.565,67.97
X$13327 937 VIA_via1_4
* cell instance $13328 r0 *1 22.325,60.83
X$13328 937 VIA_via1_4
* cell instance $13329 r0 *1 16.435,38.43
X$13329 937 VIA_via1_4
* cell instance $13330 r0 *1 26.315,39.97
X$13330 937 VIA_via1_4
* cell instance $13331 r0 *1 26.315,39.97
X$13331 937 VIA_via2_5
* cell instance $13332 r0 *1 21.945,73.57
X$13332 937 VIA_via1_4
* cell instance $13333 r0 *1 21.945,73.57
X$13333 937 VIA_via2_5
* cell instance $13334 r0 *1 26.695,73.57
X$13334 937 VIA_via1_4
* cell instance $13335 r0 *1 26.695,73.57
X$13335 937 VIA_via2_5
* cell instance $13336 r0 *1 16.625,46.83
X$13336 937 VIA_via1_4
* cell instance $13337 r0 *1 16.245,41.23
X$13337 937 VIA_via1_4
* cell instance $13338 r0 *1 16.245,41.23
X$13338 937 VIA_via2_5
* cell instance $13339 r0 *1 16.335,41.23
X$13339 937 VIA_via3_2
* cell instance $13340 r0 *1 16.625,44.03
X$13340 937 VIA_via1_4
* cell instance $13341 r0 *1 26.135,40.39
X$13341 937 VIA_via4_0
* cell instance $13342 r0 *1 16.335,40.39
X$13342 937 VIA_via4_0
* cell instance $13343 r0 *1 26.135,39.97
X$13343 937 VIA_via3_2
* cell instance $13344 r0 *1 28.405,38.99
X$13344 938 VIA_via1_7
* cell instance $13345 r0 *1 27.265,39.97
X$13345 938 VIA_via1_4
* cell instance $13346 r0 *1 27.455,38.43
X$13346 939 VIA_via1_4
* cell instance $13347 r0 *1 27.455,38.43
X$13347 939 VIA_via2_5
* cell instance $13348 r0 *1 29.735,38.43
X$13348 939 VIA_via1_4
* cell instance $13349 r0 *1 29.735,38.43
X$13349 939 VIA_via2_5
* cell instance $13350 r0 *1 29.545,39.55
X$13350 939 VIA_via1_4
* cell instance $13351 r0 *1 30.115,38.99
X$13351 940 VIA_via1_7
* cell instance $13352 r0 *1 29.735,39.97
X$13352 940 VIA_via1_4
* cell instance $13353 r0 *1 3.515,45.43
X$13353 941 VIA_via1_7
* cell instance $13354 r0 *1 5.225,41.37
X$13354 941 VIA_via1_7
* cell instance $13355 r0 *1 7.505,42.63
X$13355 941 VIA_via1_7
* cell instance $13356 r0 *1 7.505,42.49
X$13356 941 VIA_via2_5
* cell instance $13357 r0 *1 10.165,39.83
X$13357 941 VIA_via1_7
* cell instance $13358 r0 *1 39.425,45.43
X$13358 941 VIA_via1_7
* cell instance $13359 r0 *1 31.255,38.57
X$13359 941 VIA_via1_7
* cell instance $13360 r0 *1 39.615,41.37
X$13360 941 VIA_via1_7
* cell instance $13361 r0 *1 21.185,42.63
X$13361 941 VIA_via1_7
* cell instance $13362 r0 *1 48.355,45.15
X$13362 941 VIA_via2_5
* cell instance $13363 r0 *1 39.615,43.61
X$13363 941 VIA_via2_5
* cell instance $13364 r0 *1 39.425,45.15
X$13364 941 VIA_via2_5
* cell instance $13365 r0 *1 47.025,45.15
X$13365 941 VIA_via2_5
* cell instance $13366 r0 *1 8.455,43.33
X$13366 941 VIA_via2_5
* cell instance $13367 r0 *1 5.225,42.49
X$13367 941 VIA_via2_5
* cell instance $13368 r0 *1 8.455,42.49
X$13368 941 VIA_via2_5
* cell instance $13369 r0 *1 39.425,44.31
X$13369 941 VIA_via2_5
* cell instance $13370 r0 *1 3.515,42.49
X$13370 941 VIA_via2_5
* cell instance $13371 r0 *1 39.615,42.21
X$13371 941 VIA_via2_5
* cell instance $13372 r0 *1 20.995,43.33
X$13372 941 VIA_via2_5
* cell instance $13373 r0 *1 29.355,42.49
X$13373 941 VIA_via2_5
* cell instance $13374 r0 *1 30.115,42.49
X$13374 941 VIA_via2_5
* cell instance $13375 r0 *1 10.165,43.33
X$13375 941 VIA_via2_5
* cell instance $13376 r0 *1 29.355,43.33
X$13376 941 VIA_via2_5
* cell instance $13377 r0 *1 48.355,42.77
X$13377 941 VIA_via1_4
* cell instance $13378 r0 *1 47.025,46.55
X$13378 941 VIA_via1_4
* cell instance $13379 r0 *1 29.355,42.77
X$13379 941 VIA_via1_4
* cell instance $13380 r0 *1 33.345,42.91
X$13380 942 VIA_via1_7
* cell instance $13381 r0 *1 36.005,44.03
X$13381 942 VIA_via2_5
* cell instance $13382 r0 *1 36.385,44.03
X$13382 942 VIA_via2_5
* cell instance $13383 r0 *1 33.345,44.03
X$13383 942 VIA_via2_5
* cell instance $13384 r0 *1 33.345,39.97
X$13384 942 VIA_via2_5
* cell instance $13385 r0 *1 36.005,45.57
X$13385 942 VIA_via1_4
* cell instance $13386 r0 *1 31.255,44.03
X$13386 942 VIA_via1_4
* cell instance $13387 r0 *1 31.255,44.03
X$13387 942 VIA_via2_5
* cell instance $13388 r0 *1 36.575,44.03
X$13388 942 VIA_via1_4
* cell instance $13389 r0 *1 36.575,44.03
X$13389 942 VIA_via2_5
* cell instance $13390 r0 *1 28.025,39.97
X$13390 942 VIA_via1_4
* cell instance $13391 r0 *1 28.025,39.97
X$13391 942 VIA_via2_5
* cell instance $13392 r0 *1 27.835,44.03
X$13392 942 VIA_via1_4
* cell instance $13393 r0 *1 27.835,44.03
X$13393 942 VIA_via2_5
* cell instance $13394 r0 *1 36.575,37.17
X$13394 942 VIA_via1_4
* cell instance $13395 r0 *1 33.345,41.23
X$13395 942 VIA_via1_4
* cell instance $13396 r0 *1 33.725,42.77
X$13396 942 VIA_via1_4
* cell instance $13397 r0 *1 31.825,39.97
X$13397 942 VIA_via1_4
* cell instance $13398 r0 *1 31.825,39.97
X$13398 942 VIA_via2_5
* cell instance $13399 r0 *1 33.535,38.43
X$13399 943 VIA_via2_5
* cell instance $13400 r0 *1 31.445,38.43
X$13400 943 VIA_via1_4
* cell instance $13401 r0 *1 31.445,38.43
X$13401 943 VIA_via2_5
* cell instance $13402 r0 *1 33.345,39.55
X$13402 943 VIA_via1_4
* cell instance $13403 r0 *1 33.725,39.97
X$13403 943 VIA_via1_4
* cell instance $13404 r0 *1 33.725,38.99
X$13404 944 VIA_via1_7
* cell instance $13405 r0 *1 33.915,41.23
X$13405 944 VIA_via2_5
* cell instance $13406 r0 *1 32.585,41.23
X$13406 944 VIA_via1_4
* cell instance $13407 r0 *1 32.585,41.23
X$13407 944 VIA_via2_5
* cell instance $13408 r0 *1 34.295,39.13
X$13408 945 VIA_via2_5
* cell instance $13409 r0 *1 32.775,39.13
X$13409 945 VIA_via2_5
* cell instance $13410 r0 *1 34.295,39.97
X$13410 945 VIA_via1_4
* cell instance $13411 r0 *1 34.865,41.51
X$13411 945 VIA_via1_4
* cell instance $13412 r0 *1 32.775,38.43
X$13412 945 VIA_via1_4
* cell instance $13413 r0 *1 35.245,36.19
X$13413 946 VIA_via1_7
* cell instance $13414 r0 *1 35.815,39.97
X$13414 946 VIA_via1_4
* cell instance $13415 r0 *1 38.095,38.57
X$13415 947 VIA_via2_5
* cell instance $13416 r0 *1 38.095,37.45
X$13416 947 VIA_via1_4
* cell instance $13417 r0 *1 37.715,38.43
X$13417 947 VIA_via1_4
* cell instance $13418 r0 *1 37.715,38.57
X$13418 947 VIA_via2_5
* cell instance $13419 r0 *1 34.485,38.43
X$13419 947 VIA_via1_4
* cell instance $13420 r0 *1 34.485,38.57
X$13420 947 VIA_via2_5
* cell instance $13421 r0 *1 38.095,38.99
X$13421 948 VIA_via1_7
* cell instance $13422 r0 *1 37.905,39.97
X$13422 948 VIA_via1_4
* cell instance $13423 r0 *1 40.755,40.81
X$13423 949 VIA_via1_7
* cell instance $13424 r0 *1 41.135,39.97
X$13424 949 VIA_via1_4
* cell instance $13425 r0 *1 57.855,38.99
X$13425 950 VIA_via1_7
* cell instance $13426 r0 *1 57.475,39.97
X$13426 950 VIA_via1_4
* cell instance $13427 r0 *1 60.705,39.97
X$13427 951 VIA_via2_5
* cell instance $13428 r0 *1 59.945,38.43
X$13428 951 VIA_via1_4
* cell instance $13429 r0 *1 60.705,38.43
X$13429 951 VIA_via1_4
* cell instance $13430 r0 *1 61.845,39.97
X$13430 951 VIA_via1_4
* cell instance $13431 r0 *1 61.845,39.97
X$13431 951 VIA_via2_5
* cell instance $13432 r0 *1 60.325,38.99
X$13432 952 VIA_via1_7
* cell instance $13433 r0 *1 59.565,39.97
X$13433 952 VIA_via1_4
* cell instance $13434 r0 *1 61.655,38.99
X$13434 953 VIA_via1_7
* cell instance $13435 r0 *1 62.225,39.97
X$13435 953 VIA_via1_4
* cell instance $13436 r0 *1 66.595,41.23
X$13436 954 VIA_via2_5
* cell instance $13437 r0 *1 66.595,43.89
X$13437 954 VIA_via2_5
* cell instance $13438 r0 *1 68.495,48.37
X$13438 954 VIA_via2_5
* cell instance $13439 r0 *1 68.685,43.89
X$13439 954 VIA_via2_5
* cell instance $13440 r0 *1 64.885,41.23
X$13440 954 VIA_via2_5
* cell instance $13441 r0 *1 69.065,43.89
X$13441 954 VIA_via2_5
* cell instance $13442 r0 *1 65.455,41.23
X$13442 954 VIA_via1_4
* cell instance $13443 r0 *1 65.455,41.23
X$13443 954 VIA_via2_5
* cell instance $13444 r0 *1 66.595,42.77
X$13444 954 VIA_via1_4
* cell instance $13445 r0 *1 69.065,42.35
X$13445 954 VIA_via1_4
* cell instance $13446 r0 *1 69.065,43.19
X$13446 954 VIA_via1_7
* cell instance $13447 r0 *1 72.105,48.37
X$13447 954 VIA_via1_4
* cell instance $13448 r0 *1 72.105,48.37
X$13448 954 VIA_via2_5
* cell instance $13449 r0 *1 70.395,44.03
X$13449 954 VIA_via1_4
* cell instance $13450 r0 *1 70.395,43.89
X$13450 954 VIA_via2_5
* cell instance $13451 r0 *1 68.495,46.83
X$13451 954 VIA_via1_4
* cell instance $13452 r0 *1 66.595,45.57
X$13452 954 VIA_via1_4
* cell instance $13453 r0 *1 64.695,38.43
X$13453 954 VIA_via1_4
* cell instance $13454 r0 *1 69.255,41.23
X$13454 954 VIA_via1_4
* cell instance $13455 r0 *1 66.975,39.97
X$13455 955 VIA_via2_5
* cell instance $13456 r0 *1 66.215,39.97
X$13456 955 VIA_via1_4
* cell instance $13457 r0 *1 66.215,39.97
X$13457 955 VIA_via2_5
* cell instance $13458 r0 *1 66.975,40.95
X$13458 955 VIA_via1_4
* cell instance $13459 r0 *1 63.745,39.97
X$13459 955 VIA_via1_4
* cell instance $13460 r0 *1 63.745,39.97
X$13460 955 VIA_via2_5
* cell instance $13461 r0 *1 88.825,38.99
X$13461 956 VIA_via1_7
* cell instance $13462 r0 *1 88.445,39.97
X$13462 956 VIA_via1_4
* cell instance $13463 r0 *1 92.435,39.41
X$13463 957 VIA_via1_7
* cell instance $13464 r0 *1 92.625,38.43
X$13464 957 VIA_via1_4
* cell instance $13465 r0 *1 96.615,39.97
X$13465 958 VIA_via2_5
* cell instance $13466 r0 *1 92.055,39.97
X$13466 958 VIA_via1_4
* cell instance $13467 r0 *1 92.055,39.97
X$13467 958 VIA_via2_5
* cell instance $13468 r0 *1 93.955,39.97
X$13468 958 VIA_via1_4
* cell instance $13469 r0 *1 93.955,39.97
X$13469 958 VIA_via2_5
* cell instance $13470 r0 *1 96.615,38.85
X$13470 958 VIA_via1_4
* cell instance $13471 r0 *1 94.335,39.41
X$13471 959 VIA_via1_7
* cell instance $13472 r0 *1 94.335,38.43
X$13472 959 VIA_via1_4
* cell instance $13473 r0 *1 2.565,38.43
X$13473 960 VIA_via1_4
* cell instance $13474 r0 *1 2.565,38.43
X$13474 960 VIA_via2_5
* cell instance $13475 r0 *1 6.175,38.43
X$13475 960 VIA_via1_4
* cell instance $13476 r0 *1 6.175,38.43
X$13476 960 VIA_via2_5
* cell instance $13477 r0 *1 6.365,40.81
X$13477 961 VIA_via1_7
* cell instance $13478 r0 *1 6.365,39.97
X$13478 961 VIA_via2_5
* cell instance $13479 r0 *1 3.325,39.97
X$13479 961 VIA_via1_4
* cell instance $13480 r0 *1 3.325,39.97
X$13480 961 VIA_via2_5
* cell instance $13481 r0 *1 11.305,39.41
X$13481 962 VIA_via1_7
* cell instance $13482 r0 *1 11.305,39.41
X$13482 962 VIA_via2_5
* cell instance $13483 r0 *1 7.125,39.41
X$13483 962 VIA_via2_5
* cell instance $13484 r0 *1 7.125,38.43
X$13484 962 VIA_via1_4
* cell instance $13485 r0 *1 92.815,38.43
X$13485 963 VIA_via1_4
* cell instance $13486 r0 *1 92.815,38.43
X$13486 963 VIA_via2_5
* cell instance $13487 r0 *1 91.865,38.43
X$13487 963 VIA_via1_4
* cell instance $13488 r0 *1 91.865,38.43
X$13488 963 VIA_via2_5
* cell instance $13489 r0 *1 92.435,37.59
X$13489 964 VIA_via1_7
* cell instance $13490 r0 *1 92.435,38.57
X$13490 964 VIA_via2_5
* cell instance $13491 r0 *1 92.055,38.43
X$13491 964 VIA_via1_4
* cell instance $13492 r0 *1 92.055,38.57
X$13492 964 VIA_via2_5
* cell instance $13493 r0 *1 9.025,40.81
X$13493 965 VIA_via1_7
* cell instance $13494 r0 *1 9.025,39.97
X$13494 965 VIA_via2_5
* cell instance $13495 r0 *1 7.695,39.97
X$13495 965 VIA_via1_4
* cell instance $13496 r0 *1 7.695,39.97
X$13496 965 VIA_via2_5
* cell instance $13497 r0 *1 86.545,39.41
X$13497 966 VIA_via1_7
* cell instance $13498 r0 *1 86.545,39.41
X$13498 966 VIA_via2_5
* cell instance $13499 r0 *1 91.295,39.41
X$13499 966 VIA_via2_5
* cell instance $13500 r0 *1 91.295,38.43
X$13500 966 VIA_via1_4
* cell instance $13501 r0 *1 7.695,40.81
X$13501 967 VIA_via1_7
* cell instance $13502 r0 *1 7.885,38.71
X$13502 967 VIA_via2_5
* cell instance $13503 r0 *1 16.055,38.71
X$13503 967 VIA_via2_5
* cell instance $13504 r0 *1 16.055,38.43
X$13504 967 VIA_via1_4
* cell instance $13505 r0 *1 12.635,39.97
X$13505 968 VIA_via1_4
* cell instance $13506 r0 *1 12.635,39.97
X$13506 968 VIA_via2_5
* cell instance $13507 r0 *1 15.485,39.97
X$13507 968 VIA_via1_4
* cell instance $13508 r0 *1 15.485,39.97
X$13508 968 VIA_via2_5
* cell instance $13509 r0 *1 15.485,40.95
X$13509 968 VIA_via1_4
* cell instance $13510 r0 *1 16.245,39.97
X$13510 969 VIA_via1_4
* cell instance $13511 r0 *1 15.865,39.97
X$13511 969 VIA_via1_4
* cell instance $13512 r0 *1 16.815,37.59
X$13512 970 VIA_via1_7
* cell instance $13513 r0 *1 17.955,38.99
X$13513 970 VIA_via2_5
* cell instance $13514 r0 *1 16.815,38.99
X$13514 970 VIA_via2_5
* cell instance $13515 r0 *1 17.955,39.97
X$13515 970 VIA_via1_4
* cell instance $13516 r0 *1 83.315,39.83
X$13516 971 VIA_via1_4
* cell instance $13517 r0 *1 83.315,39.83
X$13517 971 VIA_via2_5
* cell instance $13518 r0 *1 86.165,39.97
X$13518 971 VIA_via1_4
* cell instance $13519 r0 *1 86.165,39.83
X$13519 971 VIA_via2_5
* cell instance $13520 r0 *1 20.045,40.11
X$13520 972 VIA_via2_5
* cell instance $13521 r0 *1 20.045,38.71
X$13521 972 VIA_via2_5
* cell instance $13522 r0 *1 19.285,38.71
X$13522 972 VIA_via1_4
* cell instance $13523 r0 *1 19.285,38.71
X$13523 972 VIA_via2_5
* cell instance $13524 r0 *1 17.385,40.04
X$13524 972 VIA_via1_4
* cell instance $13525 r0 *1 17.385,40.11
X$13525 972 VIA_via2_5
* cell instance $13526 r0 *1 24.225,38.43
X$13526 973 VIA_via1_4
* cell instance $13527 r0 *1 24.415,38.43
X$13527 973 VIA_via1_4
* cell instance $13528 r0 *1 76.285,39.55
X$13528 974 VIA_via2_5
* cell instance $13529 r0 *1 82.365,40.25
X$13529 974 VIA_via2_5
* cell instance $13530 r0 *1 79.135,39.55
X$13530 974 VIA_via2_5
* cell instance $13531 r0 *1 82.365,39.97
X$13531 974 VIA_via1_4
* cell instance $13532 r0 *1 79.135,40.25
X$13532 974 VIA_via1_4
* cell instance $13533 r0 *1 79.135,40.25
X$13533 974 VIA_via2_5
* cell instance $13534 r0 *1 76.285,38.43
X$13534 974 VIA_via1_4
* cell instance $13535 r0 *1 24.605,38.43
X$13535 975 VIA_via1_4
* cell instance $13536 r0 *1 24.605,38.43
X$13536 975 VIA_via2_5
* cell instance $13537 r0 *1 26.125,38.43
X$13537 975 VIA_via1_4
* cell instance $13538 r0 *1 26.125,38.43
X$13538 975 VIA_via2_5
* cell instance $13539 r0 *1 77.235,38.99
X$13539 976 VIA_via1_7
* cell instance $13540 r0 *1 77.235,38.99
X$13540 976 VIA_via2_5
* cell instance $13541 r0 *1 76.855,38.99
X$13541 976 VIA_via2_5
* cell instance $13542 r0 *1 76.855,39.97
X$13542 976 VIA_via1_4
* cell instance $13543 r0 *1 71.725,39.97
X$13543 977 VIA_via2_5
* cell instance $13544 r0 *1 71.535,39.97
X$13544 977 VIA_via1_4
* cell instance $13545 r0 *1 71.535,39.97
X$13545 977 VIA_via2_5
* cell instance $13546 r0 *1 71.725,41.23
X$13546 977 VIA_via1_4
* cell instance $13547 r0 *1 75.145,39.97
X$13547 977 VIA_via1_4
* cell instance $13548 r0 *1 75.145,39.97
X$13548 977 VIA_via2_5
* cell instance $13549 r0 *1 70.585,39.55
X$13549 978 VIA_via2_5
* cell instance $13550 r0 *1 70.585,46.83
X$13550 978 VIA_via1_4
* cell instance $13551 r0 *1 68.495,39.55
X$13551 978 VIA_via1_4
* cell instance $13552 r0 *1 68.495,39.55
X$13552 978 VIA_via2_5
* cell instance $13553 r0 *1 67.165,39.83
X$13553 979 VIA_via1_4
* cell instance $13554 r0 *1 67.165,39.83
X$13554 979 VIA_via2_5
* cell instance $13555 r0 *1 68.115,39.97
X$13555 979 VIA_via1_4
* cell instance $13556 r0 *1 68.115,39.83
X$13556 979 VIA_via2_5
* cell instance $13557 r0 *1 39.615,38.43
X$13557 980 VIA_via1_4
* cell instance $13558 r0 *1 39.615,38.43
X$13558 980 VIA_via2_5
* cell instance $13559 r0 *1 36.765,38.43
X$13559 980 VIA_via1_4
* cell instance $13560 r0 *1 36.765,38.43
X$13560 980 VIA_via2_5
* cell instance $13561 r0 *1 38.095,39.97
X$13561 981 VIA_via1_4
* cell instance $13562 r0 *1 38.095,39.97
X$13562 981 VIA_via2_5
* cell instance $13563 r0 *1 35.245,39.97
X$13563 981 VIA_via1_4
* cell instance $13564 r0 *1 35.245,39.97
X$13564 981 VIA_via2_5
* cell instance $13565 r0 *1 45.315,39.41
X$13565 982 VIA_via1_7
* cell instance $13566 r0 *1 45.315,38.43
X$13566 982 VIA_via1_4
* cell instance $13567 r0 *1 48.165,37.59
X$13567 983 VIA_via1_7
* cell instance $13568 r0 *1 48.165,38.85
X$13568 983 VIA_via2_5
* cell instance $13569 r0 *1 46.075,38.85
X$13569 983 VIA_via2_5
* cell instance $13570 r0 *1 46.075,38.43
X$13570 983 VIA_via1_4
* cell instance $13571 r0 *1 50.825,38.57
X$13571 984 VIA_via2_5
* cell instance $13572 r0 *1 51.015,38.57
X$13572 984 VIA_via1_4
* cell instance $13573 r0 *1 51.015,38.57
X$13573 984 VIA_via2_5
* cell instance $13574 r0 *1 50.825,41.23
X$13574 984 VIA_via1_4
* cell instance $13575 r0 *1 46.835,38.43
X$13575 984 VIA_via1_4
* cell instance $13576 r0 *1 46.835,38.57
X$13576 984 VIA_via2_5
* cell instance $13577 r0 *1 54.815,37.59
X$13577 985 VIA_via1_7
* cell instance $13578 r0 *1 54.815,38.43
X$13578 985 VIA_via2_5
* cell instance $13579 r0 *1 54.245,38.43
X$13579 985 VIA_via1_4
* cell instance $13580 r0 *1 54.245,38.43
X$13580 985 VIA_via2_5
* cell instance $13581 r0 *1 47.785,38.43
X$13581 986 VIA_via1_4
* cell instance $13582 r0 *1 47.785,38.43
X$13582 986 VIA_via2_5
* cell instance $13583 r0 *1 48.735,38.43
X$13583 986 VIA_via1_4
* cell instance $13584 r0 *1 48.735,38.43
X$13584 986 VIA_via2_5
* cell instance $13585 r0 *1 52.155,38.71
X$13585 987 VIA_via2_5
* cell instance $13586 r0 *1 52.155,38.43
X$13586 987 VIA_via1_4
* cell instance $13587 r0 *1 51.585,38.85
X$13587 987 VIA_via1_4
* cell instance $13588 r0 *1 51.585,38.71
X$13588 987 VIA_via2_5
* cell instance $13589 r0 *1 55.765,59.57
X$13589 988 VIA_via2_5
* cell instance $13590 r0 *1 55.005,41.23
X$13590 988 VIA_via2_5
* cell instance $13591 r0 *1 43.035,52.29
X$13591 988 VIA_via2_5
* cell instance $13592 r0 *1 36.005,60.69
X$13592 988 VIA_via2_5
* cell instance $13593 r0 *1 31.255,60.69
X$13593 988 VIA_via2_5
* cell instance $13594 r0 *1 36.005,52.29
X$13594 988 VIA_via2_5
* cell instance $13595 r0 *1 36.385,59.57
X$13595 988 VIA_via2_5
* cell instance $13596 r0 *1 36.385,60.69
X$13596 988 VIA_via2_5
* cell instance $13597 r0 *1 55.385,41.23
X$13597 988 VIA_via2_5
* cell instance $13598 r0 *1 53.485,39.97
X$13598 988 VIA_via1_4
* cell instance $13599 r0 *1 53.485,39.97
X$13599 988 VIA_via2_5
* cell instance $13600 r0 *1 55.955,41.23
X$13600 988 VIA_via1_4
* cell instance $13601 r0 *1 55.955,41.23
X$13601 988 VIA_via2_5
* cell instance $13602 r0 *1 55.005,39.97
X$13602 988 VIA_via1_4
* cell instance $13603 r0 *1 55.005,39.97
X$13603 988 VIA_via2_5
* cell instance $13604 r0 *1 37.525,59.57
X$13604 988 VIA_via1_4
* cell instance $13605 r0 *1 37.525,59.57
X$13605 988 VIA_via2_5
* cell instance $13606 r0 *1 31.255,59.57
X$13606 988 VIA_via1_4
* cell instance $13607 r0 *1 33.915,52.43
X$13607 988 VIA_via1_4
* cell instance $13608 r0 *1 33.915,52.29
X$13608 988 VIA_via2_5
* cell instance $13609 r0 *1 43.225,48.37
X$13609 988 VIA_via1_4
* cell instance $13610 r0 *1 31.445,62.37
X$13610 988 VIA_via1_4
* cell instance $13611 r0 *1 36.005,62.37
X$13611 988 VIA_via1_4
* cell instance $13612 r0 *1 36.005,62.37
X$13612 988 VIA_via2_5
* cell instance $13613 r0 *1 38.665,62.37
X$13613 988 VIA_via1_4
* cell instance $13614 r0 *1 38.665,62.37
X$13614 988 VIA_via2_5
* cell instance $13615 r0 *1 57.665,59.57
X$13615 988 VIA_via1_4
* cell instance $13616 r0 *1 57.665,59.57
X$13616 988 VIA_via2_5
* cell instance $13617 r0 *1 13.585,40.39
X$13617 989 VIA_via1_7
* cell instance $13618 r0 *1 13.205,41.23
X$13618 989 VIA_via1_4
* cell instance $13619 r0 *1 17.955,41.79
X$13619 990 VIA_via1_7
* cell instance $13620 r0 *1 18.145,42.77
X$13620 990 VIA_via1_4
* cell instance $13621 r0 *1 22.325,44.03
X$13621 991 VIA_via2_5
* cell instance $13622 r0 *1 23.465,44.03
X$13622 991 VIA_via2_5
* cell instance $13623 r0 *1 23.845,47.25
X$13623 991 VIA_via2_5
* cell instance $13624 r0 *1 22.325,47.25
X$13624 991 VIA_via2_5
* cell instance $13625 r0 *1 18.905,42.07
X$13625 991 VIA_via2_5
* cell instance $13626 r0 *1 23.465,42.07
X$13626 991 VIA_via2_5
* cell instance $13627 r0 *1 20.045,42.07
X$13627 991 VIA_via2_5
* cell instance $13628 r0 *1 13.965,41.65
X$13628 991 VIA_via2_5
* cell instance $13629 r0 *1 18.905,41.65
X$13629 991 VIA_via2_5
* cell instance $13630 r0 *1 18.905,42.77
X$13630 991 VIA_via1_4
* cell instance $13631 r0 *1 20.045,41.23
X$13631 991 VIA_via1_4
* cell instance $13632 r0 *1 23.655,41.23
X$13632 991 VIA_via1_4
* cell instance $13633 r0 *1 24.605,44.03
X$13633 991 VIA_via1_4
* cell instance $13634 r0 *1 24.605,44.03
X$13634 991 VIA_via2_5
* cell instance $13635 r0 *1 21.945,44.03
X$13635 991 VIA_via1_4
* cell instance $13636 r0 *1 22.135,44.03
X$13636 991 VIA_via1_4
* cell instance $13637 r0 *1 13.965,41.23
X$13637 991 VIA_via1_4
* cell instance $13638 r0 *1 22.325,46.83
X$13638 991 VIA_via1_4
* cell instance $13639 r0 *1 23.845,48.37
X$13639 991 VIA_via1_4
* cell instance $13640 r0 *1 5.035,38.57
X$13640 992 VIA_via1_7
* cell instance $13641 r0 *1 7.885,41.37
X$13641 992 VIA_via1_7
* cell instance $13642 r0 *1 40.945,45.43
X$13642 992 VIA_via1_7
* cell instance $13643 r0 *1 32.585,38.57
X$13643 992 VIA_via1_7
* cell instance $13644 r0 *1 42.085,41.37
X$13644 992 VIA_via1_7
* cell instance $13645 r0 *1 27.835,42.63
X$13645 992 VIA_via1_7
* cell instance $13646 r0 *1 47.215,47.95
X$13646 992 VIA_via2_5
* cell instance $13647 r0 *1 7.885,42.35
X$13647 992 VIA_via2_5
* cell instance $13648 r0 *1 47.025,41.93
X$13648 992 VIA_via2_5
* cell instance $13649 r0 *1 5.035,44.03
X$13649 992 VIA_via2_5
* cell instance $13650 r0 *1 42.085,41.93
X$13650 992 VIA_via2_5
* cell instance $13651 r0 *1 40.945,41.93
X$13651 992 VIA_via2_5
* cell instance $13652 r0 *1 5.035,42.35
X$13652 992 VIA_via2_5
* cell instance $13653 r0 *1 27.835,42.35
X$13653 992 VIA_via2_5
* cell instance $13654 r0 *1 6.365,44.03
X$13654 992 VIA_via2_5
* cell instance $13655 r0 *1 6.365,42.35
X$13655 992 VIA_via2_5
* cell instance $13656 r0 *1 23.085,42.35
X$13656 992 VIA_via2_5
* cell instance $13657 r0 *1 32.775,41.79
X$13657 992 VIA_via2_5
* cell instance $13658 r0 *1 22.325,42.77
X$13658 992 VIA_via2_5
* cell instance $13659 r0 *1 48.545,47.95
X$13659 992 VIA_via1_4
* cell instance $13660 r0 *1 48.545,47.95
X$13660 992 VIA_via2_5
* cell instance $13661 r0 *1 47.025,44.03
X$13661 992 VIA_via1_4
* cell instance $13662 r0 *1 22.515,42.77
X$13662 992 VIA_via1_4
* cell instance $13663 r0 *1 5.035,46.83
X$13663 992 VIA_via1_4
* cell instance $13664 r0 *1 6.555,44.03
X$13664 992 VIA_via1_4
* cell instance $13665 r0 *1 31.635,36.19
X$13665 993 VIA_via1_7
* cell instance $13666 r0 *1 31.635,41.23
X$13666 993 VIA_via1_4
* cell instance $13667 r0 *1 6.555,41.37
X$13667 994 VIA_via1_7
* cell instance $13668 r0 *1 9.215,41.37
X$13668 994 VIA_via1_7
* cell instance $13669 r0 *1 32.395,49.49
X$13669 994 VIA_via2_5
* cell instance $13670 r0 *1 33.345,49.35
X$13670 994 VIA_via2_5
* cell instance $13671 r0 *1 7.125,43.61
X$13671 994 VIA_via2_5
* cell instance $13672 r0 *1 7.885,43.61
X$13672 994 VIA_via2_5
* cell instance $13673 r0 *1 24.985,43.05
X$13673 994 VIA_via2_5
* cell instance $13674 r0 *1 30.685,43.05
X$13674 994 VIA_via2_5
* cell instance $13675 r0 *1 6.555,43.61
X$13675 994 VIA_via2_5
* cell instance $13676 r0 *1 9.215,43.61
X$13676 994 VIA_via2_5
* cell instance $13677 r0 *1 24.985,43.89
X$13677 994 VIA_via2_5
* cell instance $13678 r0 *1 33.725,42.35
X$13678 994 VIA_via2_5
* cell instance $13679 r0 *1 33.155,42.63
X$13679 994 VIA_via2_5
* cell instance $13680 r0 *1 23.465,60.41
X$13680 994 VIA_via2_5
* cell instance $13681 r0 *1 20.045,60.41
X$13681 994 VIA_via2_5
* cell instance $13682 r0 *1 32.395,60.41
X$13682 994 VIA_via2_5
* cell instance $13683 r0 *1 32.395,56.77
X$13683 994 VIA_via2_5
* cell instance $13684 r0 *1 42.465,56.91
X$13684 994 VIA_via1_4
* cell instance $13685 r0 *1 42.465,56.91
X$13685 994 VIA_via2_5
* cell instance $13686 r0 *1 31.825,56.77
X$13686 994 VIA_via1_4
* cell instance $13687 r0 *1 31.825,56.77
X$13687 994 VIA_via2_5
* cell instance $13688 r0 *1 20.045,66.43
X$13688 994 VIA_via1_4
* cell instance $13689 r0 *1 23.465,60.83
X$13689 994 VIA_via1_4
* cell instance $13690 r0 *1 7.885,44.03
X$13690 994 VIA_via1_4
* cell instance $13691 r0 *1 7.315,46.83
X$13691 994 VIA_via1_4
* cell instance $13692 r0 *1 24.985,42.77
X$13692 994 VIA_via1_4
* cell instance $13693 r0 *1 30.685,42.77
X$13693 994 VIA_via1_4
* cell instance $13694 r0 *1 30.685,42.63
X$13694 994 VIA_via2_5
* cell instance $13695 r0 *1 33.535,39.97
X$13695 994 VIA_via1_4
* cell instance $13696 r0 *1 34.675,40.39
X$13696 995 VIA_via1_7
* cell instance $13697 r0 *1 35.055,41.23
X$13697 995 VIA_via1_4
* cell instance $13698 r0 *1 35.245,40.81
X$13698 996 VIA_via1_7
* cell instance $13699 r0 *1 35.055,39.97
X$13699 996 VIA_via1_4
* cell instance $13700 r0 *1 35.625,49.77
X$13700 997 VIA_via2_5
* cell instance $13701 r0 *1 36.955,49.77
X$13701 997 VIA_via2_5
* cell instance $13702 r0 *1 35.625,49.56
X$13702 997 VIA_via1_4
* cell instance $13703 r0 *1 36.195,48.51
X$13703 997 VIA_via1_4
* cell instance $13704 r0 *1 36.955,48.51
X$13704 997 VIA_via1_4
* cell instance $13705 r0 *1 36.005,40.25
X$13705 997 VIA_via1_4
* cell instance $13706 r0 *1 43.605,41.23
X$13706 998 VIA_via1_4
* cell instance $13707 r0 *1 43.605,41.09
X$13707 998 VIA_via2_5
* cell instance $13708 r0 *1 43.415,40.25
X$13708 998 VIA_via1_4
* cell instance $13709 r0 *1 39.805,41.23
X$13709 998 VIA_via1_4
* cell instance $13710 r0 *1 39.805,41.09
X$13710 998 VIA_via2_5
* cell instance $13711 r0 *1 44.935,41.23
X$13711 999 VIA_via2_5
* cell instance $13712 r0 *1 42.275,41.23
X$13712 999 VIA_via1_4
* cell instance $13713 r0 *1 42.275,41.23
X$13713 999 VIA_via2_5
* cell instance $13714 r0 *1 44.935,42.35
X$13714 999 VIA_via1_4
* cell instance $13715 r0 *1 44.175,41.23
X$13715 999 VIA_via1_4
* cell instance $13716 r0 *1 44.175,41.23
X$13716 999 VIA_via2_5
* cell instance $13717 r0 *1 44.555,40.81
X$13717 1000 VIA_via1_7
* cell instance $13718 r0 *1 44.935,39.97
X$13718 1000 VIA_via1_4
* cell instance $13719 r0 *1 49.495,40.81
X$13719 1001 VIA_via1_7
* cell instance $13720 r0 *1 49.305,39.97
X$13720 1001 VIA_via1_4
* cell instance $13721 r0 *1 51.585,41.23
X$13721 1002 VIA_via2_5
* cell instance $13722 r0 *1 50.255,41.23
X$13722 1002 VIA_via1_4
* cell instance $13723 r0 *1 50.255,41.23
X$13723 1002 VIA_via2_5
* cell instance $13724 r0 *1 51.585,40.25
X$13724 1002 VIA_via1_4
* cell instance $13725 r0 *1 48.545,41.23
X$13725 1002 VIA_via1_4
* cell instance $13726 r0 *1 48.545,41.23
X$13726 1002 VIA_via2_5
* cell instance $13727 r0 *1 57.665,39.83
X$13727 1003 VIA_via1_4
* cell instance $13728 r0 *1 57.285,46.83
X$13728 1003 VIA_via1_4
* cell instance $13729 r0 *1 62.415,39.83
X$13729 1004 VIA_via1_4
* cell instance $13730 r0 *1 62.605,46.83
X$13730 1004 VIA_via1_4
* cell instance $13731 r0 *1 69.445,40.95
X$13731 1005 VIA_via2_5
* cell instance $13732 r0 *1 70.775,40.95
X$13732 1005 VIA_via1_4
* cell instance $13733 r0 *1 70.775,40.95
X$13733 1005 VIA_via2_5
* cell instance $13734 r0 *1 69.445,39.97
X$13734 1005 VIA_via1_4
* cell instance $13735 r0 *1 71.155,41.23
X$13735 1005 VIA_via1_4
* cell instance $13736 r0 *1 72.105,41.79
X$13736 1006 VIA_via1_7
* cell instance $13737 r0 *1 71.535,42.77
X$13737 1006 VIA_via1_4
* cell instance $13738 r0 *1 81.035,40.39
X$13738 1007 VIA_via1_7
* cell instance $13739 r0 *1 80.845,41.23
X$13739 1007 VIA_via1_4
* cell instance $13740 r0 *1 83.125,40.95
X$13740 1008 VIA_via1_4
* cell instance $13741 r0 *1 82.935,39.97
X$13741 1008 VIA_via1_4
* cell instance $13742 r0 *1 82.935,40.11
X$13742 1008 VIA_via2_5
* cell instance $13743 r0 *1 80.085,39.97
X$13743 1008 VIA_via1_4
* cell instance $13744 r0 *1 80.085,40.11
X$13744 1008 VIA_via2_5
* cell instance $13745 r0 *1 91.485,41.23
X$13745 1009 VIA_via2_5
* cell instance $13746 r0 *1 96.235,41.23
X$13746 1009 VIA_via1_4
* cell instance $13747 r0 *1 96.235,41.23
X$13747 1009 VIA_via2_5
* cell instance $13748 r0 *1 92.625,41.23
X$13748 1009 VIA_via1_4
* cell instance $13749 r0 *1 92.625,41.23
X$13749 1009 VIA_via2_5
* cell instance $13750 r0 *1 91.485,39.97
X$13750 1009 VIA_via1_4
* cell instance $13751 r0 *1 87.685,41.51
X$13751 1010 VIA_via2_5
* cell instance $13752 r0 *1 87.685,41.23
X$13752 1010 VIA_via1_4
* cell instance $13753 r0 *1 96.975,41.51
X$13753 1010 VIA_via3_2
* cell instance $13754 r0 *1 96.975,41.51
X$13754 1010 VIA_via4_0
* cell instance $13755 r0 *1 5.605,41.23
X$13755 1011 VIA_via2_5
* cell instance $13756 r0 *1 5.415,41.23
X$13756 1011 VIA_via1_4
* cell instance $13757 r0 *1 5.415,41.23
X$13757 1011 VIA_via2_5
* cell instance $13758 r0 *1 6.745,41.23
X$13758 1011 VIA_via1_4
* cell instance $13759 r0 *1 6.745,41.23
X$13759 1011 VIA_via2_5
* cell instance $13760 r0 *1 5.605,40.25
X$13760 1011 VIA_via1_4
* cell instance $13761 r0 *1 9.975,41.23
X$13761 1012 VIA_via1_4
* cell instance $13762 r0 *1 9.975,41.23
X$13762 1012 VIA_via2_5
* cell instance $13763 r0 *1 8.075,41.23
X$13763 1012 VIA_via1_4
* cell instance $13764 r0 *1 8.075,41.23
X$13764 1012 VIA_via2_5
* cell instance $13765 r0 *1 9.975,40.25
X$13765 1012 VIA_via1_4
* cell instance $13766 r0 *1 16.055,40.81
X$13766 1013 VIA_via1_7
* cell instance $13767 r0 *1 16.055,40.25
X$13767 1013 VIA_via2_5
* cell instance $13768 r0 *1 17.195,40.25
X$13768 1013 VIA_via2_5
* cell instance $13769 r0 *1 17.195,40.04
X$13769 1013 VIA_via1_4
* cell instance $13770 r0 *1 93.005,41.23
X$13770 1014 VIA_via1_4
* cell instance $13771 r0 *1 93.955,41.23
X$13771 1014 VIA_via1_4
* cell instance $13772 r0 *1 10.355,41.23
X$13772 1015 VIA_via1_4
* cell instance $13773 r0 *1 10.355,41.23
X$13773 1015 VIA_via2_5
* cell instance $13774 r0 *1 15.865,41.23
X$13774 1015 VIA_via1_4
* cell instance $13775 r0 *1 15.865,41.23
X$13775 1015 VIA_via2_5
* cell instance $13776 r0 *1 18.525,41.23
X$13776 1016 VIA_via2_5
* cell instance $13777 r0 *1 18.525,40.81
X$13777 1016 VIA_via2_5
* cell instance $13778 r0 *1 20.425,40.81
X$13778 1016 VIA_via2_5
* cell instance $13779 r0 *1 20.425,42.35
X$13779 1016 VIA_via1_4
* cell instance $13780 r0 *1 17.005,41.23
X$13780 1016 VIA_via1_4
* cell instance $13781 r0 *1 17.005,41.23
X$13781 1016 VIA_via2_5
* cell instance $13782 r0 *1 18.525,39.97
X$13782 1016 VIA_via1_4
* cell instance $13783 r0 *1 18.145,41.51
X$13783 1017 VIA_via2_5
* cell instance $13784 r0 *1 19.285,41.51
X$13784 1017 VIA_via2_5
* cell instance $13785 r0 *1 21.375,51.17
X$13785 1017 VIA_via1_4
* cell instance $13786 r0 *1 21.375,51.17
X$13786 1017 VIA_via2_5
* cell instance $13787 r0 *1 19.665,51.03
X$13787 1017 VIA_via1_4
* cell instance $13788 r0 *1 19.665,51.17
X$13788 1017 VIA_via2_5
* cell instance $13789 r0 *1 18.145,40.25
X$13789 1017 VIA_via1_4
* cell instance $13790 r0 *1 20.805,40.39
X$13790 1018 VIA_via1_7
* cell instance $13791 r0 *1 20.805,41.23
X$13791 1018 VIA_via2_5
* cell instance $13792 r0 *1 19.285,41.23
X$13792 1018 VIA_via1_4
* cell instance $13793 r0 *1 19.285,41.23
X$13793 1018 VIA_via2_5
* cell instance $13794 r0 *1 32.395,38.99
X$13794 1019 VIA_via1_7
* cell instance $13795 r0 *1 32.395,40.11
X$13795 1019 VIA_via2_5
* cell instance $13796 r0 *1 31.065,39.97
X$13796 1019 VIA_via1_4
* cell instance $13797 r0 *1 31.065,40.11
X$13797 1019 VIA_via2_5
* cell instance $13798 r0 *1 29.925,40.39
X$13798 1020 VIA_via1_7
* cell instance $13799 r0 *1 29.925,40.39
X$13799 1020 VIA_via2_5
* cell instance $13800 r0 *1 30.875,40.39
X$13800 1020 VIA_via2_5
* cell instance $13801 r0 *1 30.875,41.23
X$13801 1020 VIA_via1_4
* cell instance $13802 r0 *1 32.015,49.63
X$13802 1021 VIA_via2_5
* cell instance $13803 r0 *1 30.305,41.51
X$13803 1021 VIA_via2_5
* cell instance $13804 r0 *1 30.495,48.51
X$13804 1021 VIA_via2_5
* cell instance $13805 r0 *1 32.775,49.63
X$13805 1021 VIA_via1_4
* cell instance $13806 r0 *1 32.775,49.63
X$13806 1021 VIA_via2_5
* cell instance $13807 r0 *1 32.015,48.37
X$13807 1021 VIA_via1_4
* cell instance $13808 r0 *1 32.015,48.51
X$13808 1021 VIA_via2_5
* cell instance $13809 r0 *1 31.065,41.51
X$13809 1021 VIA_via1_4
* cell instance $13810 r0 *1 31.065,41.51
X$13810 1021 VIA_via2_5
* cell instance $13811 r0 *1 32.395,42.21
X$13811 1022 VIA_via1_7
* cell instance $13812 r0 *1 30.685,41.65
X$13812 1022 VIA_via2_5
* cell instance $13813 r0 *1 32.395,41.65
X$13813 1022 VIA_via2_5
* cell instance $13814 r0 *1 30.685,41.23
X$13814 1022 VIA_via1_4
* cell instance $13815 r0 *1 32.205,36.19
X$13815 1023 VIA_via1_7
* cell instance $13816 r0 *1 32.205,41.23
X$13816 1023 VIA_via2_5
* cell instance $13817 r0 *1 31.445,41.23
X$13817 1023 VIA_via1_4
* cell instance $13818 r0 *1 31.445,41.23
X$13818 1023 VIA_via2_5
* cell instance $13819 r0 *1 72.865,39.97
X$13819 1024 VIA_via1_4
* cell instance $13820 r0 *1 72.865,40.11
X$13820 1024 VIA_via2_5
* cell instance $13821 r0 *1 71.915,40.11
X$13821 1024 VIA_via1_4
* cell instance $13822 r0 *1 71.915,40.11
X$13822 1024 VIA_via2_5
* cell instance $13823 r0 *1 69.825,40.39
X$13823 1025 VIA_via1_7
* cell instance $13824 r0 *1 69.825,41.23
X$13824 1025 VIA_via2_5
* cell instance $13825 r0 *1 68.495,41.23
X$13825 1025 VIA_via1_4
* cell instance $13826 r0 *1 68.495,41.23
X$13826 1025 VIA_via2_5
* cell instance $13827 r0 *1 64.695,40.39
X$13827 1026 VIA_via1_7
* cell instance $13828 r0 *1 64.695,41.23
X$13828 1026 VIA_via1_4
* cell instance $13829 r0 *1 51.205,40.81
X$13829 1027 VIA_via1_7
* cell instance $13830 r0 *1 51.205,38.43
X$13830 1027 VIA_via1_4
* cell instance $13831 r0 *1 7.695,42.77
X$13831 1028 VIA_via1_4
* cell instance $13832 r0 *1 7.315,42.91
X$13832 1028 VIA_via1_4
* cell instance $13833 r0 *1 8.075,44.03
X$13833 1028 VIA_via1_4
* cell instance $13834 r0 *1 22.325,42.21
X$13834 1029 VIA_via1_7
* cell instance $13835 r0 *1 22.895,41.23
X$13835 1029 VIA_via1_4
* cell instance $13836 r0 *1 23.655,43.19
X$13836 1030 VIA_via1_7
* cell instance $13837 r0 *1 23.845,44.03
X$13837 1030 VIA_via1_4
* cell instance $13838 r0 *1 21.375,42.77
X$13838 1031 VIA_via1_4
* cell instance $13839 r0 *1 21.375,42.63
X$13839 1031 VIA_via2_5
* cell instance $13840 r0 *1 25.175,42.77
X$13840 1031 VIA_via1_4
* cell instance $13841 r0 *1 25.175,42.63
X$13841 1031 VIA_via2_5
* cell instance $13842 r0 *1 25.175,41.65
X$13842 1031 VIA_via1_4
* cell instance $13843 r0 *1 32.775,43.19
X$13843 1032 VIA_via2_5
* cell instance $13844 r0 *1 30.875,43.19
X$13844 1032 VIA_via2_5
* cell instance $13845 r0 *1 29.545,43.19
X$13845 1032 VIA_via2_5
* cell instance $13846 r0 *1 32.775,43.75
X$13846 1032 VIA_via1_4
* cell instance $13847 r0 *1 29.545,42.77
X$13847 1032 VIA_via1_4
* cell instance $13848 r0 *1 30.875,42.77
X$13848 1032 VIA_via1_4
* cell instance $13849 r0 *1 39.045,43.19
X$13849 1033 VIA_via1_7
* cell instance $13850 r0 *1 39.235,44.03
X$13850 1033 VIA_via1_4
* cell instance $13851 r0 *1 43.225,41.79
X$13851 1034 VIA_via1_7
* cell instance $13852 r0 *1 42.655,42.77
X$13852 1034 VIA_via1_4
* cell instance $13853 r0 *1 46.645,43.89
X$13853 1035 VIA_via1_7
* cell instance $13854 r0 *1 46.645,44.03
X$13854 1035 VIA_via2_5
* cell instance $13855 r0 *1 48.925,44.03
X$13855 1035 VIA_via2_5
* cell instance $13856 r0 *1 41.895,42.77
X$13856 1035 VIA_via2_5
* cell instance $13857 r0 *1 53.485,44.03
X$13857 1035 VIA_via1_4
* cell instance $13858 r0 *1 53.485,44.03
X$13858 1035 VIA_via2_5
* cell instance $13859 r0 *1 49.875,44.03
X$13859 1035 VIA_via1_4
* cell instance $13860 r0 *1 49.875,44.03
X$13860 1035 VIA_via2_5
* cell instance $13861 r0 *1 49.305,46.83
X$13861 1035 VIA_via1_4
* cell instance $13862 r0 *1 46.645,42.77
X$13862 1035 VIA_via1_4
* cell instance $13863 r0 *1 46.645,42.77
X$13863 1035 VIA_via2_5
* cell instance $13864 r0 *1 43.415,42.77
X$13864 1035 VIA_via1_4
* cell instance $13865 r0 *1 43.415,42.77
X$13865 1035 VIA_via2_5
* cell instance $13866 r0 *1 41.895,39.97
X$13866 1035 VIA_via1_4
* cell instance $13867 r0 *1 48.925,45.57
X$13867 1035 VIA_via1_4
* cell instance $13868 r0 *1 47.215,43.05
X$13868 1036 VIA_via2_5
* cell instance $13869 r0 *1 50.445,43.05
X$13869 1036 VIA_via2_5
* cell instance $13870 r0 *1 50.445,42.77
X$13870 1036 VIA_via1_4
* cell instance $13871 r0 *1 48.165,43.05
X$13871 1036 VIA_via1_4
* cell instance $13872 r0 *1 48.165,43.05
X$13872 1036 VIA_via2_5
* cell instance $13873 r0 *1 47.215,44.03
X$13873 1036 VIA_via1_4
* cell instance $13874 r0 *1 49.495,43.19
X$13874 1037 VIA_via1_7
* cell instance $13875 r0 *1 49.115,44.03
X$13875 1037 VIA_via1_4
* cell instance $13876 r0 *1 58.615,47.11
X$13876 1038 VIA_via2_5
* cell instance $13877 r0 *1 58.425,47.11
X$13877 1038 VIA_via2_5
* cell instance $13878 r0 *1 52.915,47.11
X$13878 1038 VIA_via2_5
* cell instance $13879 r0 *1 52.345,47.11
X$13879 1038 VIA_via2_5
* cell instance $13880 r0 *1 64.315,42.77
X$13880 1038 VIA_via2_5
* cell instance $13881 r0 *1 60.325,42.77
X$13881 1038 VIA_via2_5
* cell instance $13882 r0 *1 58.615,42.77
X$13882 1038 VIA_via2_5
* cell instance $13883 r0 *1 52.915,45.57
X$13883 1038 VIA_via1_4
* cell instance $13884 r0 *1 60.325,39.97
X$13884 1038 VIA_via1_4
* cell instance $13885 r0 *1 64.315,44.03
X$13885 1038 VIA_via1_4
* cell instance $13886 r0 *1 61.845,42.77
X$13886 1038 VIA_via1_4
* cell instance $13887 r0 *1 61.845,42.77
X$13887 1038 VIA_via2_5
* cell instance $13888 r0 *1 58.995,45.57
X$13888 1038 VIA_via1_4
* cell instance $13889 r0 *1 58.805,47.11
X$13889 1038 VIA_via1_4
* cell instance $13890 r0 *1 58.805,47.11
X$13890 1038 VIA_via2_5
* cell instance $13891 r0 *1 58.235,44.03
X$13891 1038 VIA_via1_4
* cell instance $13892 r0 *1 52.345,49.63
X$13892 1038 VIA_via1_4
* cell instance $13893 r0 *1 58.425,49.63
X$13893 1038 VIA_via1_4
* cell instance $13894 r0 *1 68.685,43.61
X$13894 1039 VIA_via1_7
* cell instance $13895 r0 *1 66.025,44.17
X$13895 1039 VIA_via2_5
* cell instance $13896 r0 *1 68.495,44.17
X$13896 1039 VIA_via2_5
* cell instance $13897 r0 *1 65.835,42.77
X$13897 1039 VIA_via1_4
* cell instance $13898 r0 *1 70.015,44.03
X$13898 1040 VIA_via2_5
* cell instance $13899 r0 *1 70.205,44.03
X$13899 1040 VIA_via2_5
* cell instance $13900 r0 *1 70.395,42.77
X$13900 1040 VIA_via1_4
* cell instance $13901 r0 *1 70.015,45.57
X$13901 1040 VIA_via1_4
* cell instance $13902 r0 *1 71.915,44.03
X$13902 1040 VIA_via1_4
* cell instance $13903 r0 *1 71.915,44.03
X$13903 1040 VIA_via2_5
* cell instance $13904 r0 *1 83.315,42.77
X$13904 1041 VIA_via2_5
* cell instance $13905 r0 *1 81.795,42.77
X$13905 1041 VIA_via1_4
* cell instance $13906 r0 *1 81.795,42.77
X$13906 1041 VIA_via2_5
* cell instance $13907 r0 *1 82.555,42.77
X$13907 1041 VIA_via1_4
* cell instance $13908 r0 *1 82.555,42.77
X$13908 1041 VIA_via2_5
* cell instance $13909 r0 *1 83.315,43.75
X$13909 1041 VIA_via1_4
* cell instance $13910 r0 *1 84.645,43.05
X$13910 1042 VIA_via2_5
* cell instance $13911 r0 *1 84.455,43.05
X$13911 1042 VIA_via2_5
* cell instance $13912 r0 *1 85.215,43.05
X$13912 1042 VIA_via2_5
* cell instance $13913 r0 *1 81.415,46.83
X$13913 1042 VIA_via2_5
* cell instance $13914 r0 *1 84.075,46.83
X$13914 1042 VIA_via2_5
* cell instance $13915 r0 *1 88.635,43.05
X$13915 1042 VIA_via2_5
* cell instance $13916 r0 *1 86.925,43.05
X$13916 1042 VIA_via2_5
* cell instance $13917 r0 *1 84.645,38.43
X$13917 1042 VIA_via1_4
* cell instance $13918 r0 *1 85.215,42.77
X$13918 1042 VIA_via1_4
* cell instance $13919 r0 *1 81.605,41.23
X$13919 1042 VIA_via1_4
* cell instance $13920 r0 *1 84.455,45.15
X$13920 1042 VIA_via1_4
* cell instance $13921 r0 *1 84.075,45.85
X$13921 1042 VIA_via1_4
* cell instance $13922 r0 *1 81.795,44.03
X$13922 1042 VIA_via1_4
* cell instance $13923 r0 *1 82.745,46.83
X$13923 1042 VIA_via1_4
* cell instance $13924 r0 *1 82.745,46.83
X$13924 1042 VIA_via2_5
* cell instance $13925 r0 *1 76.855,46.83
X$13925 1042 VIA_via1_4
* cell instance $13926 r0 *1 76.855,46.83
X$13926 1042 VIA_via2_5
* cell instance $13927 r0 *1 88.635,42.77
X$13927 1042 VIA_via1_4
* cell instance $13928 r0 *1 86.925,44.03
X$13928 1042 VIA_via1_4
* cell instance $13929 r0 *1 8.645,42.77
X$13929 1043 VIA_via1_4
* cell instance $13930 r0 *1 8.645,42.77
X$13930 1043 VIA_via2_5
* cell instance $13931 r0 *1 5.035,42.77
X$13931 1043 VIA_via1_4
* cell instance $13932 r0 *1 5.035,42.77
X$13932 1043 VIA_via2_5
* cell instance $13933 r0 *1 84.645,43.61
X$13933 1044 VIA_via1_7
* cell instance $13934 r0 *1 84.835,42.77
X$13934 1044 VIA_via2_5
* cell instance $13935 r0 *1 84.455,42.77
X$13935 1044 VIA_via1_4
* cell instance $13936 r0 *1 84.455,42.77
X$13936 1044 VIA_via2_5
* cell instance $13937 r0 *1 22.705,42.77
X$13937 1045 VIA_via1_4
* cell instance $13938 r0 *1 22.705,42.77
X$13938 1045 VIA_via2_5
* cell instance $13939 r0 *1 25.745,42.77
X$13939 1045 VIA_via1_4
* cell instance $13940 r0 *1 25.745,42.77
X$13940 1045 VIA_via2_5
* cell instance $13941 r0 *1 26.125,43.75
X$13941 1045 VIA_via1_4
* cell instance $13942 r0 *1 77.425,42.21
X$13942 1046 VIA_via1_7
* cell instance $13943 r0 *1 77.425,42.21
X$13943 1046 VIA_via2_5
* cell instance $13944 r0 *1 76.855,42.21
X$13944 1046 VIA_via2_5
* cell instance $13945 r0 *1 76.855,41.23
X$13945 1046 VIA_via1_4
* cell instance $13946 r0 *1 79.135,42.77
X$13946 1047 VIA_via2_5
* cell instance $13947 r0 *1 76.475,42.77
X$13947 1047 VIA_via1_4
* cell instance $13948 r0 *1 76.475,42.77
X$13948 1047 VIA_via2_5
* cell instance $13949 r0 *1 76.095,44.03
X$13949 1047 VIA_via1_4
* cell instance $13950 r0 *1 79.135,41.65
X$13950 1047 VIA_via1_4
* cell instance $13951 r0 *1 75.525,43.05
X$13951 1048 VIA_via2_5
* cell instance $13952 r0 *1 76.095,43.05
X$13952 1048 VIA_via1_4
* cell instance $13953 r0 *1 76.095,43.05
X$13953 1048 VIA_via2_5
* cell instance $13954 r0 *1 74.195,44.03
X$13954 1048 VIA_via1_4
* cell instance $13955 r0 *1 74.195,44.03
X$13955 1048 VIA_via2_5
* cell instance $13956 r0 *1 75.525,44.03
X$13956 1048 VIA_via1_4
* cell instance $13957 r0 *1 75.525,44.03
X$13957 1048 VIA_via2_5
* cell instance $13958 r0 *1 75.145,43.61
X$13958 1049 VIA_via1_7
* cell instance $13959 r0 *1 75.145,43.05
X$13959 1049 VIA_via2_5
* cell instance $13960 r0 *1 73.815,43.05
X$13960 1049 VIA_via2_5
* cell instance $13961 r0 *1 73.815,42.77
X$13961 1049 VIA_via1_4
* cell instance $13962 r0 *1 32.015,42.77
X$13962 1050 VIA_via1_4
* cell instance $13963 r0 *1 31.825,42.77
X$13963 1050 VIA_via1_4
* cell instance $13964 r0 *1 67.735,42.49
X$13964 1051 VIA_via2_5
* cell instance $13965 r0 *1 68.115,42.49
X$13965 1051 VIA_via1_4
* cell instance $13966 r0 *1 68.115,42.49
X$13966 1051 VIA_via2_5
* cell instance $13967 r0 *1 67.735,44.03
X$13967 1051 VIA_via1_4
* cell instance $13968 r0 *1 67.735,44.03
X$13968 1051 VIA_via2_5
* cell instance $13969 r0 *1 66.975,44.03
X$13969 1051 VIA_via1_4
* cell instance $13970 r0 *1 66.975,44.03
X$13970 1051 VIA_via2_5
* cell instance $13971 r0 *1 37.715,42.63
X$13971 1052 VIA_via1_4
* cell instance $13972 r0 *1 37.715,42.63
X$13972 1052 VIA_via2_5
* cell instance $13973 r0 *1 38.095,42.77
X$13973 1052 VIA_via1_4
* cell instance $13974 r0 *1 38.095,42.63
X$13974 1052 VIA_via2_5
* cell instance $13975 r0 *1 38.855,36.19
X$13975 1053 VIA_via1_7
* cell instance $13976 r0 *1 38.855,42.7
X$13976 1053 VIA_via1_4
* cell instance $13977 r0 *1 50.825,42.77
X$13977 1054 VIA_via1_4
* cell instance $13978 r0 *1 51.015,42.77
X$13978 1054 VIA_via1_4
* cell instance $13979 r0 *1 49.875,43.75
X$13979 1055 VIA_via2_5
* cell instance $13980 r0 *1 51.395,43.75
X$13980 1055 VIA_via1_4
* cell instance $13981 r0 *1 51.395,43.75
X$13981 1055 VIA_via2_5
* cell instance $13982 r0 *1 49.875,42.77
X$13982 1055 VIA_via1_4
* cell instance $13983 r0 *1 49.875,42.77
X$13983 1055 VIA_via2_5
* cell instance $13984 r0 *1 48.545,42.785
X$13984 1055 VIA_via1_4
* cell instance $13985 r0 *1 48.545,42.77
X$13985 1055 VIA_via2_5
* cell instance $13986 r0 *1 8.265,44.03
X$13986 1056 VIA_via2_5
* cell instance $13987 r0 *1 8.265,45.15
X$13987 1056 VIA_via1_4
* cell instance $13988 r0 *1 8.645,44.03
X$13988 1056 VIA_via1_4
* cell instance $13989 r0 *1 6.745,44.03
X$13989 1056 VIA_via1_4
* cell instance $13990 r0 *1 6.745,44.03
X$13990 1056 VIA_via2_5
* cell instance $13991 r0 *1 15.105,44.45
X$13991 1057 VIA_via2_5
* cell instance $13992 r0 *1 15.105,44.03
X$13992 1057 VIA_via1_4
* cell instance $13993 r0 *1 14.725,44.45
X$13993 1057 VIA_via1_4
* cell instance $13994 r0 *1 14.725,44.45
X$13994 1057 VIA_via2_5
* cell instance $13995 r0 *1 15.865,45.57
X$13995 1057 VIA_via1_4
* cell instance $13996 r0 *1 17.575,44.31
X$13996 1058 VIA_via2_5
* cell instance $13997 r0 *1 18.525,44.31
X$13997 1058 VIA_via2_5
* cell instance $13998 r0 *1 19.475,44.31
X$13998 1058 VIA_via2_5
* cell instance $13999 r0 *1 18.525,46.83
X$13999 1058 VIA_via1_4
* cell instance $14000 r0 *1 19.475,45.57
X$14000 1058 VIA_via1_4
* cell instance $14001 r0 *1 17.575,44.03
X$14001 1058 VIA_via1_4
* cell instance $14002 r0 *1 31.445,43.75
X$14002 1059 VIA_via2_5
* cell instance $14003 r0 *1 28.025,43.75
X$14003 1059 VIA_via2_5
* cell instance $14004 r0 *1 28.025,42.77
X$14004 1059 VIA_via1_4
* cell instance $14005 r0 *1 29.355,43.75
X$14005 1059 VIA_via1_4
* cell instance $14006 r0 *1 29.355,43.75
X$14006 1059 VIA_via2_5
* cell instance $14007 r0 *1 31.445,42.77
X$14007 1059 VIA_via1_4
* cell instance $14008 r0 *1 38.855,45.01
X$14008 1060 VIA_via1_7
* cell instance $14009 r0 *1 38.095,44.03
X$14009 1060 VIA_via2_5
* cell instance $14010 r0 *1 35.815,44.03
X$14010 1060 VIA_via1_4
* cell instance $14011 r0 *1 35.815,43.89
X$14011 1060 VIA_via2_5
* cell instance $14012 r0 *1 38.285,43.19
X$14012 1061 VIA_via1_7
* cell instance $14013 r0 *1 38.665,44.03
X$14013 1061 VIA_via1_4
* cell instance $14014 r0 *1 39.805,43.61
X$14014 1062 VIA_via1_7
* cell instance $14015 r0 *1 39.805,43.47
X$14015 1062 VIA_via2_5
* cell instance $14016 r0 *1 38.475,43.75
X$14016 1062 VIA_via2_5
* cell instance $14017 r0 *1 38.475,44.03
X$14017 1062 VIA_via1_4
* cell instance $14018 r0 *1 40.565,53.97
X$14018 1063 VIA_via1_4
* cell instance $14019 r0 *1 39.425,51.31
X$14019 1063 VIA_via1_4
* cell instance $14020 r0 *1 40.185,51.31
X$14020 1063 VIA_via1_4
* cell instance $14021 r0 *1 38.855,44.31
X$14021 1063 VIA_via1_4
* cell instance $14022 r0 *1 46.265,44.17
X$14022 1064 VIA_via2_5
* cell instance $14023 r0 *1 45.885,42.77
X$14023 1064 VIA_via1_4
* cell instance $14024 r0 *1 48.165,44.17
X$14024 1064 VIA_via1_4
* cell instance $14025 r0 *1 48.165,44.17
X$14025 1064 VIA_via2_5
* cell instance $14026 r0 *1 54.625,45.43
X$14026 1065 VIA_via1_7
* cell instance $14027 r0 *1 54.625,45.29
X$14027 1065 VIA_via2_5
* cell instance $14028 r0 *1 61.085,52.43
X$14028 1065 VIA_via2_5
* cell instance $14029 r0 *1 45.885,45.29
X$14029 1065 VIA_via2_5
* cell instance $14030 r0 *1 61.085,48.09
X$14030 1065 VIA_via2_5
* cell instance $14031 r0 *1 54.625,44.17
X$14031 1065 VIA_via2_5
* cell instance $14032 r0 *1 61.085,44.17
X$14032 1065 VIA_via2_5
* cell instance $14033 r0 *1 61.845,48.09
X$14033 1065 VIA_via2_5
* cell instance $14034 r0 *1 59.945,44.03
X$14034 1065 VIA_via1_4
* cell instance $14035 r0 *1 59.945,44.17
X$14035 1065 VIA_via2_5
* cell instance $14036 r0 *1 45.315,53.97
X$14036 1065 VIA_via1_4
* cell instance $14037 r0 *1 45.885,45.57
X$14037 1065 VIA_via1_4
* cell instance $14038 r0 *1 61.085,55.23
X$14038 1065 VIA_via1_4
* cell instance $14039 r0 *1 61.845,52.43
X$14039 1065 VIA_via1_4
* cell instance $14040 r0 *1 61.845,52.43
X$14040 1065 VIA_via2_5
* cell instance $14041 r0 *1 63.935,43.75
X$14041 1066 VIA_via2_5
* cell instance $14042 r0 *1 66.405,43.75
X$14042 1066 VIA_via2_5
* cell instance $14043 r0 *1 63.935,42.77
X$14043 1066 VIA_via1_4
* cell instance $14044 r0 *1 65.835,43.75
X$14044 1066 VIA_via1_4
* cell instance $14045 r0 *1 65.835,43.75
X$14045 1066 VIA_via2_5
* cell instance $14046 r0 *1 66.405,44.03
X$14046 1066 VIA_via1_4
* cell instance $14047 r0 *1 67.355,44.59
X$14047 1067 VIA_via1_7
* cell instance $14048 r0 *1 67.165,45.57
X$14048 1067 VIA_via1_4
* cell instance $14049 r0 *1 84.265,43.75
X$14049 1068 VIA_via2_5
* cell instance $14050 r0 *1 86.735,43.75
X$14050 1068 VIA_via2_5
* cell instance $14051 r0 *1 83.125,43.75
X$14051 1068 VIA_via2_5
* cell instance $14052 r0 *1 83.125,42.77
X$14052 1068 VIA_via1_4
* cell instance $14053 r0 *1 84.265,44.03
X$14053 1068 VIA_via1_4
* cell instance $14054 r0 *1 86.735,43.05
X$14054 1068 VIA_via1_4
* cell instance $14055 r0 *1 86.735,44.03
X$14055 1069 VIA_via2_5
* cell instance $14056 r0 *1 88.445,44.03
X$14056 1069 VIA_via1_4
* cell instance $14057 r0 *1 88.445,44.03
X$14057 1069 VIA_via2_5
* cell instance $14058 r0 *1 86.925,45.57
X$14058 1069 VIA_via1_4
* cell instance $14059 r0 *1 88.825,44.03
X$14059 1069 VIA_via1_4
* cell instance $14060 r0 *1 88.825,44.03
X$14060 1069 VIA_via2_5
* cell instance $14061 r0 *1 89.395,45.57
X$14061 1070 VIA_via2_5
* cell instance $14062 r0 *1 88.255,45.57
X$14062 1070 VIA_via1_4
* cell instance $14063 r0 *1 88.255,45.57
X$14063 1070 VIA_via2_5
* cell instance $14064 r0 *1 89.395,44.03
X$14064 1070 VIA_via1_4
* cell instance $14065 r0 *1 90.155,43.05
X$14065 1070 VIA_via1_4
* cell instance $14066 r0 *1 91.675,44.59
X$14066 1071 VIA_via1_7
* cell instance $14067 r0 *1 91.485,45.57
X$14067 1071 VIA_via1_4
* cell instance $14068 r0 *1 95.285,44.03
X$14068 1072 VIA_via2_5
* cell instance $14069 r0 *1 95.285,45.15
X$14069 1072 VIA_via1_4
* cell instance $14070 r0 *1 92.625,44.03
X$14070 1072 VIA_via1_4
* cell instance $14071 r0 *1 92.625,44.03
X$14071 1072 VIA_via2_5
* cell instance $14072 r0 *1 90.725,44.03
X$14072 1072 VIA_via1_4
* cell instance $14073 r0 *1 90.725,44.03
X$14073 1072 VIA_via2_5
* cell instance $14074 r0 *1 88.445,54.39
X$14074 1073 VIA_via2_5
* cell instance $14075 r0 *1 88.445,58.31
X$14075 1073 VIA_via2_5
* cell instance $14076 r0 *1 94.715,54.25
X$14076 1073 VIA_via2_5
* cell instance $14077 r0 *1 79.515,58.31
X$14077 1073 VIA_via2_5
* cell instance $14078 r0 *1 82.935,58.31
X$14078 1073 VIA_via2_5
* cell instance $14079 r0 *1 76.855,57.75
X$14079 1073 VIA_via2_5
* cell instance $14080 r0 *1 79.515,57.75
X$14080 1073 VIA_via2_5
* cell instance $14081 r0 *1 92.055,43.75
X$14081 1073 VIA_via2_5
* cell instance $14082 r0 *1 94.525,43.75
X$14082 1073 VIA_via2_5
* cell instance $14083 r0 *1 92.055,44.03
X$14083 1073 VIA_via1_4
* cell instance $14084 r0 *1 94.525,44.03
X$14084 1073 VIA_via1_4
* cell instance $14085 r0 *1 94.905,54.25
X$14085 1073 VIA_via1_4
* cell instance $14086 r0 *1 94.905,54.25
X$14086 1073 VIA_via2_5
* cell instance $14087 r0 *1 79.515,59.57
X$14087 1073 VIA_via1_4
* cell instance $14088 r0 *1 82.935,58.03
X$14088 1073 VIA_via1_4
* cell instance $14089 r0 *1 77.045,52.43
X$14089 1073 VIA_via1_4
* cell instance $14090 r0 *1 76.855,58.03
X$14090 1073 VIA_via1_4
* cell instance $14091 r0 *1 76.855,55.23
X$14091 1073 VIA_via1_4
* cell instance $14092 r0 *1 96.425,43.89
X$14092 1074 VIA_via2_5
* cell instance $14093 r0 *1 95.095,44.03
X$14093 1074 VIA_via1_4
* cell instance $14094 r0 *1 95.095,43.89
X$14094 1074 VIA_via2_5
* cell instance $14095 r0 *1 96.425,43.05
X$14095 1074 VIA_via1_4
* cell instance $14096 r0 *1 91.295,44.03
X$14096 1074 VIA_via1_4
* cell instance $14097 r0 *1 91.295,43.89
X$14097 1074 VIA_via2_5
* cell instance $14098 r0 *1 7.695,44.59
X$14098 1075 VIA_via1_7
* cell instance $14099 r0 *1 7.695,44.59
X$14099 1075 VIA_via2_5
* cell instance $14100 r0 *1 5.985,44.59
X$14100 1075 VIA_via2_5
* cell instance $14101 r0 *1 5.985,45.57
X$14101 1075 VIA_via1_4
* cell instance $14102 r0 *1 94.145,44.17
X$14102 1076 VIA_via2_5
* cell instance $14103 r0 *1 94.145,42.77
X$14103 1076 VIA_via1_4
* cell instance $14104 r0 *1 95.475,44.17
X$14104 1076 VIA_via1_4
* cell instance $14105 r0 *1 95.475,44.17
X$14105 1076 VIA_via2_5
* cell instance $14106 r0 *1 12.445,44.03
X$14106 1077 VIA_via1_4
* cell instance $14107 r0 *1 12.445,43.89
X$14107 1077 VIA_via2_5
* cell instance $14108 r0 *1 16.055,43.89
X$14108 1077 VIA_via1_4
* cell instance $14109 r0 *1 16.055,43.89
X$14109 1077 VIA_via2_5
* cell instance $14110 r0 *1 16.245,43.75
X$14110 1078 VIA_via2_5
* cell instance $14111 r0 *1 9.025,43.75
X$14111 1078 VIA_via1_4
* cell instance $14112 r0 *1 9.025,43.75
X$14112 1078 VIA_via2_5
* cell instance $14113 r0 *1 16.245,44.03
X$14113 1078 VIA_via1_4
* cell instance $14114 r0 *1 17.195,44.03
X$14114 1079 VIA_via1_4
* cell instance $14115 r0 *1 17.195,44.17
X$14115 1079 VIA_via2_5
* cell instance $14116 r0 *1 16.435,44.17
X$14116 1079 VIA_via1_4
* cell instance $14117 r0 *1 16.435,44.17
X$14117 1079 VIA_via2_5
* cell instance $14118 r0 *1 28.975,43.19
X$14118 1080 VIA_via1_7
* cell instance $14119 r0 *1 28.975,43.19
X$14119 1080 VIA_via2_5
* cell instance $14120 r0 *1 27.075,43.19
X$14120 1080 VIA_via2_5
* cell instance $14121 r0 *1 27.075,44.03
X$14121 1080 VIA_via1_4
* cell instance $14122 r0 *1 30.495,43.19
X$14122 1081 VIA_via1_7
* cell instance $14123 r0 *1 30.495,44.03
X$14123 1081 VIA_via1_4
* cell instance $14124 r0 *1 83.505,43.19
X$14124 1082 VIA_via1_7
* cell instance $14125 r0 *1 83.505,43.33
X$14125 1082 VIA_via2_5
* cell instance $14126 r0 *1 79.515,43.33
X$14126 1082 VIA_via2_5
* cell instance $14127 r0 *1 79.515,44.03
X$14127 1082 VIA_via1_4
* cell instance $14128 r0 *1 37.905,43.75
X$14128 1083 VIA_via2_5
* cell instance $14129 r0 *1 36.765,43.75
X$14129 1083 VIA_via2_5
* cell instance $14130 r0 *1 38.095,43.75
X$14130 1083 VIA_via1_4
* cell instance $14131 r0 *1 38.095,43.75
X$14131 1083 VIA_via2_5
* cell instance $14132 r0 *1 37.905,45.57
X$14132 1083 VIA_via1_4
* cell instance $14133 r0 *1 36.765,42.77
X$14133 1083 VIA_via1_4
* cell instance $14134 r0 *1 82.175,43.19
X$14134 1084 VIA_via1_7
* cell instance $14135 r0 *1 82.175,43.19
X$14135 1084 VIA_via2_5
* cell instance $14136 r0 *1 81.035,43.19
X$14136 1084 VIA_via2_5
* cell instance $14137 r0 *1 81.035,44.03
X$14137 1084 VIA_via1_4
* cell instance $14138 r0 *1 41.515,43.89
X$14138 1085 VIA_via1_4
* cell instance $14139 r0 *1 41.515,43.89
X$14139 1085 VIA_via2_5
* cell instance $14140 r0 *1 39.615,44.03
X$14140 1085 VIA_via1_4
* cell instance $14141 r0 *1 39.615,43.89
X$14141 1085 VIA_via2_5
* cell instance $14142 r0 *1 39.425,41.79
X$14142 1086 VIA_via1_7
* cell instance $14143 r0 *1 39.425,44.03
X$14143 1086 VIA_via1_4
* cell instance $14144 r0 *1 39.805,46.13
X$14144 1087 VIA_via2_5
* cell instance $14145 r0 *1 39.805,44.73
X$14145 1087 VIA_via2_5
* cell instance $14146 r0 *1 40.565,44.73
X$14146 1087 VIA_via2_5
* cell instance $14147 r0 *1 40.185,46.13
X$14147 1087 VIA_via2_5
* cell instance $14148 r0 *1 39.615,45.57
X$14148 1087 VIA_via1_4
* cell instance $14149 r0 *1 40.565,44.03
X$14149 1087 VIA_via1_4
* cell instance $14150 r0 *1 40.185,46.55
X$14150 1087 VIA_via1_4
* cell instance $14151 r0 *1 80.465,53.27
X$14151 1088 VIA_via2_5
* cell instance $14152 r0 *1 84.645,53.27
X$14152 1088 VIA_via2_5
* cell instance $14153 r0 *1 85.405,53.27
X$14153 1088 VIA_via2_5
* cell instance $14154 r0 *1 80.275,44.17
X$14154 1088 VIA_via2_5
* cell instance $14155 r0 *1 78.565,44.17
X$14155 1088 VIA_via2_5
* cell instance $14156 r0 *1 78.565,35.91
X$14156 1088 VIA_via1_4
* cell instance $14157 r0 *1 84.645,53.97
X$14157 1088 VIA_via1_4
* cell instance $14158 r0 *1 85.405,53.97
X$14158 1088 VIA_via1_4
* cell instance $14159 r0 *1 76.475,44.59
X$14159 1089 VIA_via1_7
* cell instance $14160 r0 *1 76.475,44.59
X$14160 1089 VIA_via2_5
* cell instance $14161 r0 *1 75.525,44.59
X$14161 1089 VIA_via2_5
* cell instance $14162 r0 *1 75.525,45.57
X$14162 1089 VIA_via1_4
* cell instance $14163 r0 *1 70.775,43.19
X$14163 1090 VIA_via1_7
* cell instance $14164 r0 *1 70.775,43.19
X$14164 1090 VIA_via2_5
* cell instance $14165 r0 *1 69.635,43.19
X$14165 1090 VIA_via2_5
* cell instance $14166 r0 *1 69.635,44.03
X$14166 1090 VIA_via1_4
* cell instance $14167 r0 *1 61.085,43.61
X$14167 1091 VIA_via1_7
* cell instance $14168 r0 *1 61.085,42.77
X$14168 1091 VIA_via1_4
* cell instance $14169 r0 *1 60.325,44.03
X$14169 1092 VIA_via2_5
* cell instance $14170 r0 *1 63.365,44.03
X$14170 1092 VIA_via2_5
* cell instance $14171 r0 *1 63.365,43.05
X$14171 1092 VIA_via1_4
* cell instance $14172 r0 *1 60.135,44.03
X$14172 1092 VIA_via1_4
* cell instance $14173 r0 *1 60.135,44.03
X$14173 1092 VIA_via2_5
* cell instance $14174 r0 *1 60.325,45.57
X$14174 1092 VIA_via1_4
* cell instance $14175 r0 *1 64.885,43.19
X$14175 1093 VIA_via1_7
* cell instance $14176 r0 *1 64.885,43.19
X$14176 1093 VIA_via2_5
* cell instance $14177 r0 *1 63.555,43.19
X$14177 1093 VIA_via2_5
* cell instance $14178 r0 *1 63.555,44.03
X$14178 1093 VIA_via1_4
* cell instance $14179 r0 *1 5.795,46.27
X$14179 1094 VIA_via2_5
* cell instance $14180 r0 *1 3.325,46.55
X$14180 1094 VIA_via2_5
* cell instance $14181 r0 *1 6.365,46.83
X$14181 1094 VIA_via2_5
* cell instance $14182 r0 *1 6.745,46.83
X$14182 1094 VIA_via2_5
* cell instance $14183 r0 *1 6.745,46.27
X$14183 1094 VIA_via2_5
* cell instance $14184 r0 *1 3.325,46.83
X$14184 1094 VIA_via1_4
* cell instance $14185 r0 *1 6.365,48.37
X$14185 1094 VIA_via1_4
* cell instance $14186 r0 *1 5.795,42.77
X$14186 1094 VIA_via1_4
* cell instance $14187 r0 *1 12.065,45.57
X$14187 1094 VIA_via1_4
* cell instance $14188 r0 *1 11.685,46.83
X$14188 1094 VIA_via1_4
* cell instance $14189 r0 *1 11.685,46.83
X$14189 1094 VIA_via2_5
* cell instance $14190 r0 *1 9.595,46.83
X$14190 1094 VIA_via1_4
* cell instance $14191 r0 *1 9.595,46.83
X$14191 1094 VIA_via2_5
* cell instance $14192 r0 *1 9.405,46.83
X$14192 1094 VIA_via1_4
* cell instance $14193 r0 *1 6.745,45.57
X$14193 1094 VIA_via1_4
* cell instance $14194 r0 *1 13.205,44.03
X$14194 1094 VIA_via1_4
* cell instance $14195 r0 *1 13.585,45.57
X$14195 1095 VIA_via1_4
* cell instance $14196 r0 *1 13.585,45.57
X$14196 1095 VIA_via2_5
* cell instance $14197 r0 *1 13.965,45.57
X$14197 1095 VIA_via1_4
* cell instance $14198 r0 *1 13.965,45.57
X$14198 1095 VIA_via2_5
* cell instance $14199 r0 *1 15.295,45.57
X$14199 1095 VIA_via1_4
* cell instance $14200 r0 *1 15.295,45.57
X$14200 1095 VIA_via2_5
* cell instance $14201 r0 *1 17.385,44.03
X$14201 1096 VIA_via1_4
* cell instance $14202 r0 *1 17.005,45.15
X$14202 1096 VIA_via1_4
* cell instance $14203 r0 *1 16.435,46.69
X$14203 1097 VIA_via2_5
* cell instance $14204 r0 *1 21.185,46.41
X$14204 1097 VIA_via2_5
* cell instance $14205 r0 *1 16.625,49.63
X$14205 1097 VIA_via1_4
* cell instance $14206 r0 *1 20.235,46.83
X$14206 1097 VIA_via1_4
* cell instance $14207 r0 *1 20.235,46.83
X$14207 1097 VIA_via2_5
* cell instance $14208 r0 *1 20.995,45.57
X$14208 1097 VIA_via1_4
* cell instance $14209 r0 *1 23.845,46.83
X$14209 1097 VIA_via1_4
* cell instance $14210 r0 *1 23.845,46.83
X$14210 1097 VIA_via2_5
* cell instance $14211 r0 *1 41.135,45.57
X$14211 1098 VIA_via1_4
* cell instance $14212 r0 *1 41.135,45.71
X$14212 1098 VIA_via2_5
* cell instance $14213 r0 *1 41.135,44.03
X$14213 1098 VIA_via1_4
* cell instance $14214 r0 *1 45.315,45.71
X$14214 1098 VIA_via1_4
* cell instance $14215 r0 *1 45.315,45.71
X$14215 1098 VIA_via2_5
* cell instance $14216 r0 *1 47.975,62.23
X$14216 1099 VIA_via1_7
* cell instance $14217 r0 *1 47.975,62.23
X$14217 1099 VIA_via2_5
* cell instance $14218 r0 *1 77.805,45.43
X$14218 1099 VIA_via1_7
* cell instance $14219 r0 *1 77.805,45.43
X$14219 1099 VIA_via2_5
* cell instance $14220 r0 *1 34.485,80.57
X$14220 1099 VIA_via1_7
* cell instance $14221 r0 *1 34.485,80.57
X$14221 1099 VIA_via2_5
* cell instance $14222 r0 *1 41.895,80.57
X$14222 1099 VIA_via1_7
* cell instance $14223 r0 *1 41.895,80.57
X$14223 1099 VIA_via2_5
* cell instance $14224 r0 *1 47.215,79.03
X$14224 1099 VIA_via1_7
* cell instance $14225 r0 *1 47.215,79.03
X$14225 1099 VIA_via2_5
* cell instance $14226 r0 *1 69.255,45.43
X$14226 1099 VIA_via1_7
* cell instance $14227 r0 *1 69.255,45.43
X$14227 1099 VIA_via2_5
* cell instance $14228 r0 *1 66.975,73.43
X$14228 1099 VIA_via1_7
* cell instance $14229 r0 *1 47.215,80.57
X$14229 1099 VIA_via2_5
* cell instance $14230 r0 *1 47.215,79.87
X$14230 1099 VIA_via2_5
* cell instance $14231 r0 *1 55.385,80.01
X$14231 1099 VIA_via2_5
* cell instance $14232 r0 *1 67.355,71.47
X$14232 1099 VIA_via2_5
* cell instance $14233 r0 *1 74.575,57.89
X$14233 1099 VIA_via2_5
* cell instance $14234 r0 *1 79.325,71.75
X$14234 1099 VIA_via2_5
* cell instance $14235 r0 *1 41.895,46.27
X$14235 1099 VIA_via2_5
* cell instance $14236 r0 *1 47.405,46.27
X$14236 1099 VIA_via2_5
* cell instance $14237 r0 *1 74.385,45.43
X$14237 1099 VIA_via2_5
* cell instance $14238 r0 *1 55.385,80.43
X$14238 1099 VIA_via1_4
* cell instance $14239 r0 *1 41.895,46.55
X$14239 1099 VIA_via1_4
* cell instance $14240 r0 *1 79.325,72.03
X$14240 1099 VIA_via1_4
* cell instance $14241 r0 *1 75.335,58.03
X$14241 1099 VIA_via1_4
* cell instance $14242 r0 *1 75.335,57.89
X$14242 1099 VIA_via2_5
* cell instance $14243 r0 *1 47.415,79.03
X$14243 1099 VIA_via3_2
* cell instance $14244 r0 *1 75.135,71.47
X$14244 1099 VIA_via3_2
* cell instance $14245 r0 *1 75.135,71.75
X$14245 1099 VIA_via3_2
* cell instance $14246 r0 *1 47.135,62.23
X$14246 1099 VIA_via3_2
* cell instance $14247 r0 *1 75.135,57.89
X$14247 1099 VIA_via3_2
* cell instance $14248 r0 *1 54.435,45.85
X$14248 1100 VIA_via1_4
* cell instance $14249 r0 *1 52.535,46.83
X$14249 1100 VIA_via1_4
* cell instance $14250 r0 *1 52.535,46.83
X$14250 1100 VIA_via2_5
* cell instance $14251 r0 *1 53.865,46.83
X$14251 1100 VIA_via1_4
* cell instance $14252 r0 *1 53.865,46.83
X$14252 1100 VIA_via2_5
* cell instance $14253 r0 *1 55.005,44.45
X$14253 1101 VIA_via1_4
* cell instance $14254 r0 *1 54.815,45.57
X$14254 1101 VIA_via1_4
* cell instance $14255 r0 *1 54.435,46.83
X$14255 1101 VIA_via1_4
* cell instance $14256 r0 *1 61.655,45.99
X$14256 1102 VIA_via1_7
* cell instance $14257 r0 *1 62.035,46.83
X$14257 1102 VIA_via1_4
* cell instance $14258 r0 *1 70.015,45.85
X$14258 1103 VIA_via2_5
* cell instance $14259 r0 *1 68.495,45.85
X$14259 1103 VIA_via2_5
* cell instance $14260 r0 *1 69.445,45.85
X$14260 1103 VIA_via2_5
* cell instance $14261 r0 *1 69.445,45.57
X$14261 1103 VIA_via1_4
* cell instance $14262 r0 *1 68.495,45.57
X$14262 1103 VIA_via1_4
* cell instance $14263 r0 *1 70.015,46.55
X$14263 1103 VIA_via1_4
* cell instance $14264 r0 *1 70.965,45.99
X$14264 1104 VIA_via1_7
* cell instance $14265 r0 *1 71.155,46.83
X$14265 1104 VIA_via1_4
* cell instance $14266 r0 *1 54.435,72.31
X$14266 1105 VIA_via2_5
* cell instance $14267 r0 *1 66.975,70.35
X$14267 1105 VIA_via2_5
* cell instance $14268 r0 *1 66.975,71.75
X$14268 1105 VIA_via2_5
* cell instance $14269 r0 *1 66.025,72.31
X$14269 1105 VIA_via2_5
* cell instance $14270 r0 *1 77.235,53.41
X$14270 1105 VIA_via2_5
* cell instance $14271 r0 *1 76.285,53.41
X$14271 1105 VIA_via2_5
* cell instance $14272 r0 *1 76.475,70.35
X$14272 1105 VIA_via2_5
* cell instance $14273 r0 *1 47.975,72.31
X$14273 1105 VIA_via2_5
* cell instance $14274 r0 *1 77.425,45.71
X$14274 1105 VIA_via2_5
* cell instance $14275 r0 *1 66.025,72.03
X$14275 1105 VIA_via1_4
* cell instance $14276 r0 *1 66.025,71.89
X$14276 1105 VIA_via2_5
* cell instance $14277 r0 *1 54.435,72.03
X$14277 1105 VIA_via1_4
* cell instance $14278 r0 *1 75.905,45.57
X$14278 1105 VIA_via1_4
* cell instance $14279 r0 *1 75.905,45.71
X$14279 1105 VIA_via2_5
* cell instance $14280 r0 *1 67.545,45.57
X$14280 1105 VIA_via1_4
* cell instance $14281 r0 *1 67.545,45.71
X$14281 1105 VIA_via2_5
* cell instance $14282 r0 *1 44.365,58.45
X$14282 1105 VIA_via1_4
* cell instance $14283 r0 *1 44.365,58.45
X$14283 1105 VIA_via2_5
* cell instance $14284 r0 *1 44.335,58.45
X$14284 1105 VIA_via3_2
* cell instance $14285 r0 *1 43.985,59.57
X$14285 1105 VIA_via1_4
* cell instance $14286 r0 *1 43.985,59.57
X$14286 1105 VIA_via2_5
* cell instance $14287 r0 *1 37.335,72.03
X$14287 1105 VIA_via1_4
* cell instance $14288 r0 *1 37.335,72.03
X$14288 1105 VIA_via2_5
* cell instance $14289 r0 *1 47.785,70.77
X$14289 1105 VIA_via1_4
* cell instance $14290 r0 *1 41.515,72.03
X$14290 1105 VIA_via1_4
* cell instance $14291 r0 *1 41.515,72.03
X$14291 1105 VIA_via2_5
* cell instance $14292 r0 *1 76.475,62.37
X$14292 1105 VIA_via1_4
* cell instance $14293 r0 *1 76.665,69.23
X$14293 1105 VIA_via1_4
* cell instance $14294 r0 *1 44.335,72.31
X$14294 1105 VIA_via3_2
* cell instance $14295 r0 *1 44.335,59.57
X$14295 1105 VIA_via3_2
* cell instance $14296 r0 *1 77.235,45.99
X$14296 1106 VIA_via1_7
* cell instance $14297 r0 *1 76.095,46.83
X$14297 1106 VIA_via1_4
* cell instance $14298 r0 *1 78.375,45.71
X$14298 1107 VIA_via2_5
* cell instance $14299 r0 *1 76.855,45.57
X$14299 1107 VIA_via1_4
* cell instance $14300 r0 *1 76.855,45.57
X$14300 1107 VIA_via2_5
* cell instance $14301 r0 *1 77.995,45.57
X$14301 1107 VIA_via1_4
* cell instance $14302 r0 *1 77.995,45.71
X$14302 1107 VIA_via2_5
* cell instance $14303 r0 *1 78.375,46.55
X$14303 1107 VIA_via1_4
* cell instance $14304 r0 *1 79.325,45.99
X$14304 1108 VIA_via1_7
* cell instance $14305 r0 *1 79.515,46.83
X$14305 1108 VIA_via1_4
* cell instance $14306 r0 *1 84.265,45.57
X$14306 1109 VIA_via2_5
* cell instance $14307 r0 *1 78.565,45.57
X$14307 1109 VIA_via1_4
* cell instance $14308 r0 *1 78.565,45.57
X$14308 1109 VIA_via2_5
* cell instance $14309 r0 *1 84.265,46.55
X$14309 1109 VIA_via1_4
* cell instance $14310 r0 *1 82.365,45.57
X$14310 1109 VIA_via1_4
* cell instance $14311 r0 *1 82.365,45.57
X$14311 1109 VIA_via2_5
* cell instance $14312 r0 *1 82.745,45.99
X$14312 1110 VIA_via1_7
* cell instance $14313 r0 *1 81.985,46.83
X$14313 1110 VIA_via1_4
* cell instance $14314 r0 *1 95.285,71.61
X$14314 1111 VIA_via1_7
* cell instance $14315 r0 *1 80.845,50.75
X$14315 1111 VIA_via2_5
* cell instance $14316 r0 *1 80.735,50.75
X$14316 1111 VIA_via3_2
* cell instance $14317 r0 *1 84.835,70.49
X$14317 1111 VIA_via2_5
* cell instance $14318 r0 *1 81.225,70.49
X$14318 1111 VIA_via2_5
* cell instance $14319 r0 *1 86.355,70.49
X$14319 1111 VIA_via2_5
* cell instance $14320 r0 *1 95.285,70.77
X$14320 1111 VIA_via2_5
* cell instance $14321 r0 *1 86.355,45.85
X$14321 1111 VIA_via2_5
* cell instance $14322 r0 *1 81.035,45.85
X$14322 1111 VIA_via2_5
* cell instance $14323 r0 *1 87.685,45.85
X$14323 1111 VIA_via2_5
* cell instance $14324 r0 *1 81.035,48.37
X$14324 1111 VIA_via1_4
* cell instance $14325 r0 *1 86.355,45.57
X$14325 1111 VIA_via1_4
* cell instance $14326 r0 *1 87.685,45.57
X$14326 1111 VIA_via1_4
* cell instance $14327 r0 *1 86.355,70.77
X$14327 1111 VIA_via1_4
* cell instance $14328 r0 *1 86.355,70.77
X$14328 1111 VIA_via2_5
* cell instance $14329 r0 *1 80.845,72.03
X$14329 1111 VIA_via1_4
* cell instance $14330 r0 *1 84.835,70.77
X$14330 1111 VIA_via1_4
* cell instance $14331 r0 *1 80.845,51.17
X$14331 1111 VIA_via1_4
* cell instance $14332 r0 *1 80.735,57.47
X$14332 1111 VIA_via3_2
* cell instance $14333 r0 *1 80.655,57.47
X$14333 1111 VIA_via2_5
* cell instance $14334 r0 *1 89.775,44.59
X$14334 1112 VIA_via1_7
* cell instance $14335 r0 *1 90.155,45.57
X$14335 1112 VIA_via1_4
* cell instance $14336 r0 *1 96.235,45.57
X$14336 1113 VIA_via1_4
* cell instance $14337 r0 *1 96.235,45.57
X$14337 1113 VIA_via2_5
* cell instance $14338 r0 *1 97.255,47.11
X$14338 1113 VIA_via4_0
* cell instance $14339 r0 *1 97.255,45.57
X$14339 1113 VIA_via3_2
* cell instance $14340 r0 *1 93.005,44.59
X$14340 1114 VIA_via1_7
* cell instance $14341 r0 *1 93.005,45.57
X$14341 1114 VIA_via1_4
* cell instance $14342 r0 *1 11.305,45.57
X$14342 1115 VIA_via1_4
* cell instance $14343 r0 *1 11.305,45.71
X$14343 1115 VIA_via2_5
* cell instance $14344 r0 *1 14.915,45.71
X$14344 1115 VIA_via1_4
* cell instance $14345 r0 *1 14.915,45.71
X$14345 1115 VIA_via2_5
* cell instance $14346 r0 *1 88.635,45.01
X$14346 1116 VIA_via1_7
* cell instance $14347 r0 *1 88.635,45.01
X$14347 1116 VIA_via2_5
* cell instance $14348 r0 *1 87.875,45.01
X$14348 1116 VIA_via2_5
* cell instance $14349 r0 *1 87.875,42.77
X$14349 1116 VIA_via1_4
* cell instance $14350 r0 *1 16.245,45.57
X$14350 1117 VIA_via1_4
* cell instance $14351 r0 *1 16.245,45.57
X$14351 1117 VIA_via2_5
* cell instance $14352 r0 *1 16.625,45.57
X$14352 1117 VIA_via1_4
* cell instance $14353 r0 *1 16.625,45.57
X$14353 1117 VIA_via2_5
* cell instance $14354 r0 *1 87.305,45.01
X$14354 1118 VIA_via1_7
* cell instance $14355 r0 *1 87.305,45.01
X$14355 1118 VIA_via2_5
* cell instance $14356 r0 *1 86.165,45.01
X$14356 1118 VIA_via2_5
* cell instance $14357 r0 *1 86.165,44.03
X$14357 1118 VIA_via1_4
* cell instance $14358 r0 *1 21.375,45.71
X$14358 1119 VIA_via2_5
* cell instance $14359 r0 *1 21.375,48.37
X$14359 1119 VIA_via1_4
* cell instance $14360 r0 *1 20.235,45.71
X$14360 1119 VIA_via1_4
* cell instance $14361 r0 *1 20.235,45.71
X$14361 1119 VIA_via2_5
* cell instance $14362 r0 *1 78.945,45.57
X$14362 1120 VIA_via1_4
* cell instance $14363 r0 *1 79.135,45.57
X$14363 1120 VIA_via1_4
* cell instance $14364 r0 *1 18.335,45.85
X$14364 1121 VIA_via2_5
* cell instance $14365 r0 *1 17.955,47.25
X$14365 1121 VIA_via2_5
* cell instance $14366 r0 *1 18.335,47.25
X$14366 1121 VIA_via2_5
* cell instance $14367 r0 *1 17.955,49.63
X$14367 1121 VIA_via1_4
* cell instance $14368 r0 *1 21.945,45.71
X$14368 1121 VIA_via1_4
* cell instance $14369 r0 *1 21.945,45.85
X$14369 1121 VIA_via2_5
* cell instance $14370 r0 *1 35.435,49.35
X$14370 1122 VIA_via2_5
* cell instance $14371 r0 *1 35.375,49.35
X$14371 1122 VIA_via3_2
* cell instance $14372 r0 *1 44.745,52.71
X$14372 1122 VIA_via2_5
* cell instance $14373 r0 *1 38.665,52.71
X$14373 1122 VIA_via2_5
* cell instance $14374 r0 *1 28.595,48.51
X$14374 1122 VIA_via2_5
* cell instance $14375 r0 *1 17.195,50.19
X$14375 1122 VIA_via2_5
* cell instance $14376 r0 *1 22.895,50.33
X$14376 1122 VIA_via2_5
* cell instance $14377 r0 *1 28.595,50.33
X$14377 1122 VIA_via2_5
* cell instance $14378 r0 *1 32.015,51.31
X$14378 1122 VIA_via2_5
* cell instance $14379 r0 *1 28.595,51.31
X$14379 1122 VIA_via2_5
* cell instance $14380 r0 *1 38.095,51.17
X$14380 1122 VIA_via1_4
* cell instance $14381 r0 *1 38.095,51.17
X$14381 1122 VIA_via2_5
* cell instance $14382 r0 *1 38.665,51.17
X$14382 1122 VIA_via1_4
* cell instance $14383 r0 *1 38.665,51.17
X$14383 1122 VIA_via2_5
* cell instance $14384 r0 *1 35.435,46.83
X$14384 1122 VIA_via1_4
* cell instance $14385 r0 *1 44.745,53.55
X$14385 1122 VIA_via1_4
* cell instance $14386 r0 *1 17.005,49.63
X$14386 1122 VIA_via1_4
* cell instance $14387 r0 *1 17.955,53.97
X$14387 1122 VIA_via1_4
* cell instance $14388 r0 *1 22.895,51.17
X$14388 1122 VIA_via1_4
* cell instance $14389 r0 *1 31.825,55.23
X$14389 1122 VIA_via1_4
* cell instance $14390 r0 *1 28.405,48.37
X$14390 1122 VIA_via1_4
* cell instance $14391 r0 *1 29.355,48.37
X$14391 1122 VIA_via1_4
* cell instance $14392 r0 *1 29.355,48.51
X$14392 1122 VIA_via2_5
* cell instance $14393 r0 *1 22.135,45.57
X$14393 1122 VIA_via1_4
* cell instance $14394 r0 *1 22.135,45.57
X$14394 1122 VIA_via2_5
* cell instance $14395 r0 *1 35.375,51.31
X$14395 1122 VIA_via3_2
* cell instance $14396 r0 *1 21.935,45.57
X$14396 1122 VIA_via3_2
* cell instance $14397 r0 *1 21.935,50.33
X$14397 1122 VIA_via3_2
* cell instance $14398 r0 *1 70.775,45.57
X$14398 1123 VIA_via1_4
* cell instance $14399 r0 *1 70.775,45.57
X$14399 1123 VIA_via2_5
* cell instance $14400 r0 *1 70.395,45.57
X$14400 1123 VIA_via1_4
* cell instance $14401 r0 *1 70.395,45.57
X$14401 1123 VIA_via2_5
* cell instance $14402 r0 *1 37.335,45.85
X$14402 1124 VIA_via2_5
* cell instance $14403 r0 *1 36.005,45.85
X$14403 1124 VIA_via2_5
* cell instance $14404 r0 *1 37.335,42.77
X$14404 1124 VIA_via1_4
* cell instance $14405 r0 *1 36.005,46.83
X$14405 1124 VIA_via1_4
* cell instance $14406 r0 *1 37.525,45.85
X$14406 1124 VIA_via1_4
* cell instance $14407 r0 *1 37.525,45.85
X$14407 1124 VIA_via2_5
* cell instance $14408 r0 *1 36.955,46.41
X$14408 1125 VIA_via1_7
* cell instance $14409 r0 *1 36.955,45.57
X$14409 1125 VIA_via2_5
* cell instance $14410 r0 *1 35.245,45.57
X$14410 1125 VIA_via1_4
* cell instance $14411 r0 *1 35.245,45.57
X$14411 1125 VIA_via2_5
* cell instance $14412 r0 *1 43.035,45.57
X$14412 1126 VIA_via1_4
* cell instance $14413 r0 *1 43.035,45.57
X$14413 1126 VIA_via2_5
* cell instance $14414 r0 *1 42.085,45.57
X$14414 1126 VIA_via1_4
* cell instance $14415 r0 *1 42.085,45.57
X$14415 1126 VIA_via2_5
* cell instance $14416 r0 *1 61.465,45.57
X$14416 1127 VIA_via1_4
* cell instance $14417 r0 *1 61.465,45.57
X$14417 1127 VIA_via2_5
* cell instance $14418 r0 *1 60.705,45.57
X$14418 1127 VIA_via1_4
* cell instance $14419 r0 *1 60.705,45.57
X$14419 1127 VIA_via2_5
* cell instance $14420 r0 *1 59.755,44.45
X$14420 1128 VIA_via1_4
* cell instance $14421 r0 *1 59.755,45.57
X$14421 1128 VIA_via1_4
* cell instance $14422 r0 *1 59.755,45.57
X$14422 1128 VIA_via2_5
* cell instance $14423 r0 *1 57.855,45.57
X$14423 1128 VIA_via1_4
* cell instance $14424 r0 *1 57.855,45.57
X$14424 1128 VIA_via2_5
* cell instance $14425 r0 *1 58.805,45.01
X$14425 1129 VIA_via1_7
* cell instance $14426 r0 *1 58.805,45.01
X$14426 1129 VIA_via2_5
* cell instance $14427 r0 *1 57.475,45.01
X$14427 1129 VIA_via2_5
* cell instance $14428 r0 *1 57.475,44.03
X$14428 1129 VIA_via1_4
* cell instance $14429 r0 *1 59.375,54.81
X$14429 1130 VIA_via1_7
* cell instance $14430 r0 *1 59.375,54.95
X$14430 1130 VIA_via2_5
* cell instance $14431 r0 *1 60.515,54.95
X$14431 1130 VIA_via2_5
* cell instance $14432 r0 *1 57.665,46.27
X$14432 1130 VIA_via2_5
* cell instance $14433 r0 *1 59.755,46.41
X$14433 1130 VIA_via2_5
* cell instance $14434 r0 *1 47.595,54.81
X$14434 1130 VIA_via2_5
* cell instance $14435 r0 *1 52.725,46.27
X$14435 1130 VIA_via2_5
* cell instance $14436 r0 *1 52.535,45.57
X$14436 1130 VIA_via2_5
* cell instance $14437 r0 *1 52.345,46.83
X$14437 1130 VIA_via1_4
* cell instance $14438 r0 *1 57.665,45.57
X$14438 1130 VIA_via1_4
* cell instance $14439 r0 *1 47.595,58.03
X$14439 1130 VIA_via1_4
* cell instance $14440 r0 *1 47.595,45.57
X$14440 1130 VIA_via1_4
* cell instance $14441 r0 *1 47.595,45.57
X$14441 1130 VIA_via2_5
* cell instance $14442 r0 *1 60.515,52.43
X$14442 1130 VIA_via1_4
* cell instance $14443 r0 *1 55.765,45.01
X$14443 1131 VIA_via1_7
* cell instance $14444 r0 *1 55.765,45.01
X$14444 1131 VIA_via2_5
* cell instance $14445 r0 *1 52.725,45.01
X$14445 1131 VIA_via2_5
* cell instance $14446 r0 *1 52.725,44.03
X$14446 1131 VIA_via1_4
* cell instance $14447 r0 *1 4.845,46.13
X$14447 1132 VIA_via2_5
* cell instance $14448 r0 *1 3.705,46.13
X$14448 1132 VIA_via2_5
* cell instance $14449 r0 *1 7.505,46.13
X$14449 1132 VIA_via2_5
* cell instance $14450 r0 *1 3.705,45.57
X$14450 1132 VIA_via1_4
* cell instance $14451 r0 *1 4.845,46.55
X$14451 1132 VIA_via1_4
* cell instance $14452 r0 *1 7.505,46.83
X$14452 1132 VIA_via1_4
* cell instance $14453 r0 *1 13.585,47.11
X$14453 1133 VIA_via2_5
* cell instance $14454 r0 *1 14.535,47.11
X$14454 1133 VIA_via2_5
* cell instance $14455 r0 *1 13.205,47.11
X$14455 1133 VIA_via1_4
* cell instance $14456 r0 *1 14.535,48.37
X$14456 1133 VIA_via1_4
* cell instance $14457 r0 *1 13.585,46.83
X$14457 1133 VIA_via1_4
* cell instance $14458 r0 *1 17.005,46.83
X$14458 1134 VIA_via1_4
* cell instance $14459 r0 *1 16.625,47.25
X$14459 1134 VIA_via1_4
* cell instance $14460 r0 *1 18.145,48.23
X$14460 1135 VIA_via1_4
* cell instance $14461 r0 *1 18.145,48.37
X$14461 1135 VIA_via2_5
* cell instance $14462 r0 *1 17.955,46.55
X$14462 1135 VIA_via1_4
* cell instance $14463 r0 *1 19.855,48.37
X$14463 1135 VIA_via1_4
* cell instance $14464 r0 *1 19.855,48.37
X$14464 1135 VIA_via2_5
* cell instance $14465 r0 *1 27.265,46.97
X$14465 1136 VIA_via1_7
* cell instance $14466 r0 *1 27.265,46.83
X$14466 1136 VIA_via2_5
* cell instance $14467 r0 *1 38.475,48.51
X$14467 1136 VIA_via1_7
* cell instance $14468 r0 *1 34.105,49.77
X$14468 1136 VIA_via1_7
* cell instance $14469 r0 *1 45.505,49.49
X$14469 1136 VIA_via1_7
* cell instance $14470 r0 *1 41.135,51.31
X$14470 1136 VIA_via1_7
* cell instance $14471 r0 *1 55.955,50.47
X$14471 1136 VIA_via2_5
* cell instance $14472 r0 *1 45.505,50.47
X$14472 1136 VIA_via2_5
* cell instance $14473 r0 *1 34.105,50.05
X$14473 1136 VIA_via2_5
* cell instance $14474 r0 *1 38.665,50.05
X$14474 1136 VIA_via2_5
* cell instance $14475 r0 *1 41.135,50.61
X$14475 1136 VIA_via2_5
* cell instance $14476 r0 *1 41.135,50.05
X$14476 1136 VIA_via2_5
* cell instance $14477 r0 *1 19.665,48.51
X$14477 1136 VIA_via2_5
* cell instance $14478 r0 *1 19.285,47.25
X$14478 1136 VIA_via2_5
* cell instance $14479 r0 *1 19.665,47.25
X$14479 1136 VIA_via2_5
* cell instance $14480 r0 *1 34.105,46.83
X$14480 1136 VIA_via2_5
* cell instance $14481 r0 *1 20.425,49.35
X$14481 1136 VIA_via2_5
* cell instance $14482 r0 *1 19.665,49.35
X$14482 1136 VIA_via2_5
* cell instance $14483 r0 *1 16.245,49.21
X$14483 1136 VIA_via2_5
* cell instance $14484 r0 *1 20.425,51.17
X$14484 1136 VIA_via1_4
* cell instance $14485 r0 *1 16.245,51.17
X$14485 1136 VIA_via1_4
* cell instance $14486 r0 *1 55.955,50.75
X$14486 1136 VIA_via1_4
* cell instance $14487 r0 *1 56.715,51.45
X$14487 1136 VIA_via1_4
* cell instance $14488 r0 *1 56.715,52.43
X$14488 1136 VIA_via1_4
* cell instance $14489 r0 *1 19.285,46.83
X$14489 1136 VIA_via1_4
* cell instance $14490 r0 *1 19.285,46.97
X$14490 1136 VIA_via2_5
* cell instance $14491 r0 *1 18.715,48.37
X$14491 1136 VIA_via1_4
* cell instance $14492 r0 *1 18.715,48.51
X$14492 1136 VIA_via2_5
* cell instance $14493 r0 *1 38.285,47.95
X$14493 1137 VIA_via2_5
* cell instance $14494 r0 *1 35.625,51.03
X$14494 1137 VIA_via2_5
* cell instance $14495 r0 *1 41.515,50.89
X$14495 1137 VIA_via2_5
* cell instance $14496 r0 *1 45.125,50.89
X$14496 1137 VIA_via2_5
* cell instance $14497 r0 *1 19.095,46.27
X$14497 1137 VIA_via2_5
* cell instance $14498 r0 *1 19.665,46.27
X$14498 1137 VIA_via2_5
* cell instance $14499 r0 *1 27.645,46.69
X$14499 1137 VIA_via2_5
* cell instance $14500 r0 *1 27.645,46.97
X$14500 1137 VIA_via2_5
* cell instance $14501 r0 *1 27.075,46.27
X$14501 1137 VIA_via2_5
* cell instance $14502 r0 *1 33.915,46.97
X$14502 1137 VIA_via2_5
* cell instance $14503 r0 *1 33.915,47.95
X$14503 1137 VIA_via2_5
* cell instance $14504 r0 *1 20.805,50.61
X$14504 1137 VIA_via2_5
* cell instance $14505 r0 *1 16.625,50.61
X$14505 1137 VIA_via2_5
* cell instance $14506 r0 *1 19.285,50.33
X$14506 1137 VIA_via2_5
* cell instance $14507 r0 *1 33.915,51.03
X$14507 1137 VIA_via2_5
* cell instance $14508 r0 *1 35.625,54.95
X$14508 1137 VIA_via2_5
* cell instance $14509 r0 *1 30.305,55.37
X$14509 1137 VIA_via2_5
* cell instance $14510 r0 *1 35.625,55.37
X$14510 1137 VIA_via2_5
* cell instance $14511 r0 *1 37.145,54.95
X$14511 1137 VIA_via1_4
* cell instance $14512 r0 *1 37.145,54.95
X$14512 1137 VIA_via2_5
* cell instance $14513 r0 *1 33.915,49.63
X$14513 1137 VIA_via1_4
* cell instance $14514 r0 *1 30.305,56.77
X$14514 1137 VIA_via1_4
* cell instance $14515 r0 *1 38.285,48.37
X$14515 1137 VIA_via1_4
* cell instance $14516 r0 *1 45.125,49.63
X$14516 1137 VIA_via1_4
* cell instance $14517 r0 *1 41.515,51.17
X$14517 1137 VIA_via1_4
* cell instance $14518 r0 *1 16.625,51.17
X$14518 1137 VIA_via1_4
* cell instance $14519 r0 *1 20.805,51.17
X$14519 1137 VIA_via1_4
* cell instance $14520 r0 *1 27.075,46.83
X$14520 1137 VIA_via1_4
* cell instance $14521 r0 *1 27.075,46.69
X$14521 1137 VIA_via2_5
* cell instance $14522 r0 *1 19.095,48.37
X$14522 1137 VIA_via1_4
* cell instance $14523 r0 *1 19.665,46.83
X$14523 1137 VIA_via1_4
* cell instance $14524 r0 *1 54.245,50.33
X$14524 1138 VIA_via2_5
* cell instance $14525 r0 *1 53.295,50.33
X$14525 1138 VIA_via2_5
* cell instance $14526 r0 *1 36.005,50.33
X$14526 1138 VIA_via2_5
* cell instance $14527 r0 *1 36.005,49.21
X$14527 1138 VIA_via2_5
* cell instance $14528 r0 *1 40.945,50.33
X$14528 1138 VIA_via2_5
* cell instance $14529 r0 *1 44.935,50.33
X$14529 1138 VIA_via2_5
* cell instance $14530 r0 *1 20.995,50.75
X$14530 1138 VIA_via2_5
* cell instance $14531 r0 *1 21.755,50.61
X$14531 1138 VIA_via2_5
* cell instance $14532 r0 *1 20.235,50.75
X$14532 1138 VIA_via2_5
* cell instance $14533 r0 *1 25.935,49.21
X$14533 1138 VIA_via2_5
* cell instance $14534 r0 *1 32.395,49.21
X$14534 1138 VIA_via2_5
* cell instance $14535 r0 *1 26.315,51.03
X$14535 1138 VIA_via2_5
* cell instance $14536 r0 *1 26.315,49.21
X$14536 1138 VIA_via2_5
* cell instance $14537 r0 *1 40.945,53.97
X$14537 1138 VIA_via1_4
* cell instance $14538 r0 *1 36.005,49.63
X$14538 1138 VIA_via1_4
* cell instance $14539 r0 *1 25.935,49.63
X$14539 1138 VIA_via1_4
* cell instance $14540 r0 *1 32.395,48.37
X$14540 1138 VIA_via1_4
* cell instance $14541 r0 *1 44.935,48.37
X$14541 1138 VIA_via1_4
* cell instance $14542 r0 *1 20.235,53.97
X$14542 1138 VIA_via1_4
* cell instance $14543 r0 *1 21.755,51.17
X$14543 1138 VIA_via1_4
* cell instance $14544 r0 *1 21.755,51.03
X$14544 1138 VIA_via2_5
* cell instance $14545 r0 *1 53.295,50.75
X$14545 1138 VIA_via1_4
* cell instance $14546 r0 *1 54.245,51.17
X$14546 1138 VIA_via1_4
* cell instance $14547 r0 *1 20.235,48.37
X$14547 1138 VIA_via1_4
* cell instance $14548 r0 *1 19.855,45.57
X$14548 1138 VIA_via1_4
* cell instance $14549 r0 *1 65.835,61.67
X$14549 1139 VIA_via2_5
* cell instance $14550 r0 *1 45.505,48.93
X$14550 1139 VIA_via2_5
* cell instance $14551 r0 *1 40.755,48.93
X$14551 1139 VIA_via2_5
* cell instance $14552 r0 *1 40.755,51.59
X$14552 1139 VIA_via2_5
* cell instance $14553 r0 *1 41.515,51.59
X$14553 1139 VIA_via2_5
* cell instance $14554 r0 *1 41.325,59.99
X$14554 1139 VIA_via2_5
* cell instance $14555 r0 *1 36.575,48.93
X$14555 1139 VIA_via2_5
* cell instance $14556 r0 *1 32.965,48.79
X$14556 1139 VIA_via2_5
* cell instance $14557 r0 *1 26.505,48.79
X$14557 1139 VIA_via2_5
* cell instance $14558 r0 *1 41.325,61.67
X$14558 1139 VIA_via2_5
* cell instance $14559 r0 *1 20.805,50.05
X$14559 1139 VIA_via2_5
* cell instance $14560 r0 *1 22.135,50.05
X$14560 1139 VIA_via2_5
* cell instance $14561 r0 *1 21.375,50.05
X$14561 1139 VIA_via2_5
* cell instance $14562 r0 *1 30.305,59.99
X$14562 1139 VIA_via2_5
* cell instance $14563 r0 *1 26.505,51.17
X$14563 1139 VIA_via2_5
* cell instance $14564 r0 *1 65.835,61.95
X$14564 1139 VIA_via1_4
* cell instance $14565 r0 *1 41.515,53.97
X$14565 1139 VIA_via1_4
* cell instance $14566 r0 *1 30.305,59.57
X$14566 1139 VIA_via1_4
* cell instance $14567 r0 *1 36.575,49.63
X$14567 1139 VIA_via1_4
* cell instance $14568 r0 *1 26.505,49.63
X$14568 1139 VIA_via1_4
* cell instance $14569 r0 *1 32.965,48.37
X$14569 1139 VIA_via1_4
* cell instance $14570 r0 *1 45.505,48.37
X$14570 1139 VIA_via1_4
* cell instance $14571 r0 *1 20.805,53.97
X$14571 1139 VIA_via1_4
* cell instance $14572 r0 *1 22.325,51.17
X$14572 1139 VIA_via1_4
* cell instance $14573 r0 *1 22.325,51.17
X$14573 1139 VIA_via2_5
* cell instance $14574 r0 *1 20.805,48.37
X$14574 1139 VIA_via1_4
* cell instance $14575 r0 *1 20.425,45.57
X$14575 1139 VIA_via1_4
* cell instance $14576 r0 *1 57.475,54.81
X$14576 1140 VIA_via1_7
* cell instance $14577 r0 *1 57.475,54.81
X$14577 1140 VIA_via2_5
* cell instance $14578 r0 *1 57.095,55.37
X$14578 1140 VIA_via1_4
* cell instance $14579 r0 *1 57.095,55.37
X$14579 1140 VIA_via2_5
* cell instance $14580 r0 *1 58.045,54.81
X$14580 1140 VIA_via2_5
* cell instance $14581 r0 *1 20.805,45.99
X$14581 1140 VIA_via2_5
* cell instance $14582 r0 *1 23.465,45.99
X$14582 1140 VIA_via2_5
* cell instance $14583 r0 *1 23.465,51.31
X$14583 1140 VIA_via2_5
* cell instance $14584 r0 *1 44.555,59.57
X$14584 1140 VIA_via1_4
* cell instance $14585 r0 *1 44.555,59.57
X$14585 1140 VIA_via2_5
* cell instance $14586 r0 *1 44.615,59.57
X$14586 1140 VIA_via3_2
* cell instance $14587 r0 *1 37.335,51.17
X$14587 1140 VIA_via1_4
* cell instance $14588 r0 *1 37.335,51.17
X$14588 1140 VIA_via2_5
* cell instance $14589 r0 *1 31.825,51.17
X$14589 1140 VIA_via1_4
* cell instance $14590 r0 *1 31.825,51.17
X$14590 1140 VIA_via2_5
* cell instance $14591 r0 *1 28.215,51.17
X$14591 1140 VIA_via1_4
* cell instance $14592 r0 *1 28.215,51.17
X$14592 1140 VIA_via2_5
* cell instance $14593 r0 *1 23.465,52.43
X$14593 1140 VIA_via1_4
* cell instance $14594 r0 *1 23.465,49.63
X$14594 1140 VIA_via1_4
* cell instance $14595 r0 *1 23.275,55.23
X$14595 1140 VIA_via1_4
* cell instance $14596 r0 *1 36.575,55.23
X$14596 1140 VIA_via1_4
* cell instance $14597 r0 *1 36.575,55.09
X$14597 1140 VIA_via2_5
* cell instance $14598 r0 *1 36.495,55.09
X$14598 1140 VIA_via3_2
* cell instance $14599 r0 *1 36.575,55.37
X$14599 1140 VIA_via2_5
* cell instance $14600 r0 *1 58.045,52.43
X$14600 1140 VIA_via1_4
* cell instance $14601 r0 *1 20.615,46.83
X$14601 1140 VIA_via1_4
* cell instance $14602 r0 *1 36.495,51.17
X$14602 1140 VIA_via3_2
* cell instance $14603 r0 *1 44.615,55.37
X$14603 1140 VIA_via3_2
* cell instance $14604 r0 *1 20.995,45.99
X$14604 1141 VIA_via1_7
* cell instance $14605 r0 *1 21.185,48.37
X$14605 1141 VIA_via1_4
* cell instance $14606 r0 *1 34.865,75.95
X$14606 1142 VIA_via2_5
* cell instance $14607 r0 *1 53.865,49.07
X$14607 1142 VIA_via2_5
* cell instance $14608 r0 *1 55.955,49.07
X$14608 1142 VIA_via2_5
* cell instance $14609 r0 *1 21.185,73.99
X$14609 1142 VIA_via2_5
* cell instance $14610 r0 *1 22.135,73.99
X$14610 1142 VIA_via2_5
* cell instance $14611 r0 *1 20.615,73.99
X$14611 1142 VIA_via2_5
* cell instance $14612 r0 *1 49.115,74.55
X$14612 1142 VIA_via2_5
* cell instance $14613 r0 *1 40.565,75.95
X$14613 1142 VIA_via2_5
* cell instance $14614 r0 *1 54.625,74.55
X$14614 1142 VIA_via2_5
* cell instance $14615 r0 *1 53.865,47.25
X$14615 1142 VIA_via2_5
* cell instance $14616 r0 *1 17.575,47.11
X$14616 1142 VIA_via2_5
* cell instance $14617 r0 *1 29.355,58.73
X$14617 1142 VIA_via2_5
* cell instance $14618 r0 *1 54.625,74.83
X$14618 1142 VIA_via1_4
* cell instance $14619 r0 *1 55.955,48.65
X$14619 1142 VIA_via1_4
* cell instance $14620 r0 *1 40.535,76.3
X$14620 1142 VIA_via1_4
* cell instance $14621 r0 *1 34.865,76.37
X$14621 1142 VIA_via1_4
* cell instance $14622 r0 *1 48.735,76.37
X$14622 1142 VIA_via1_4
* cell instance $14623 r0 *1 48.735,76.23
X$14623 1142 VIA_via2_5
* cell instance $14624 r0 *1 29.355,58.03
X$14624 1142 VIA_via1_4
* cell instance $14625 r0 *1 26.885,76.37
X$14625 1142 VIA_via1_4
* cell instance $14626 r0 *1 26.885,76.37
X$14626 1142 VIA_via2_5
* cell instance $14627 r0 *1 26.975,76.37
X$14627 1142 VIA_via3_2
* cell instance $14628 r0 *1 26.975,76.51
X$14628 1142 VIA_via4_0
* cell instance $14629 r0 *1 21.945,62.37
X$14629 1142 VIA_via1_4
* cell instance $14630 r0 *1 21.945,62.23
X$14630 1142 VIA_via2_5
* cell instance $14631 r0 *1 21.375,76.37
X$14631 1142 VIA_via1_4
* cell instance $14632 r0 *1 21.375,76.37
X$14632 1142 VIA_via2_5
* cell instance $14633 r0 *1 21.375,76.37
X$14633 1142 VIA_via3_2
* cell instance $14634 r0 *1 21.375,76.51
X$14634 1142 VIA_via4_0
* cell instance $14635 r0 *1 20.615,73.57
X$14635 1142 VIA_via1_4
* cell instance $14636 r0 *1 17.575,46.83
X$14636 1142 VIA_via1_4
* cell instance $14637 r0 *1 54.415,74.55
X$14637 1142 VIA_via3_2
* cell instance $14638 r0 *1 34.815,76.65
X$14638 1142 VIA_via3_2
* cell instance $14639 r0 *1 34.815,76.51
X$14639 1142 VIA_via4_0
* cell instance $14640 r0 *1 34.865,76.65
X$14640 1142 VIA_via2_5
* cell instance $14641 r0 *1 27.535,58.73
X$14641 1142 VIA_via3_2
* cell instance $14642 r0 *1 27.535,62.23
X$14642 1142 VIA_via3_2
* cell instance $14643 r0 *1 54.415,49.07
X$14643 1142 VIA_via3_2
* cell instance $14644 r0 *1 35.055,50.75
X$14644 1143 VIA_via2_5
* cell instance $14645 r0 *1 33.535,50.75
X$14645 1143 VIA_via2_5
* cell instance $14646 r0 *1 36.765,50.75
X$14646 1143 VIA_via1_4
* cell instance $14647 r0 *1 36.765,50.75
X$14647 1143 VIA_via2_5
* cell instance $14648 r0 *1 36.955,51.17
X$14648 1143 VIA_via1_4
* cell instance $14649 r0 *1 33.535,51.17
X$14649 1143 VIA_via1_4
* cell instance $14650 r0 *1 35.055,46.83
X$14650 1143 VIA_via1_4
* cell instance $14651 r0 *1 52.725,48.37
X$14651 1144 VIA_via1_4
* cell instance $14652 r0 *1 52.725,48.37
X$14652 1144 VIA_via2_5
* cell instance $14653 r0 *1 50.825,47.25
X$14653 1144 VIA_via1_4
* cell instance $14654 r0 *1 51.205,48.37
X$14654 1144 VIA_via1_4
* cell instance $14655 r0 *1 51.205,48.37
X$14655 1144 VIA_via2_5
* cell instance $14656 r0 *1 67.545,50.75
X$14656 1145 VIA_via2_5
* cell instance $14657 r0 *1 68.685,47.11
X$14657 1145 VIA_via2_5
* cell instance $14658 r0 *1 61.655,46.83
X$14658 1145 VIA_via1_4
* cell instance $14659 r0 *1 61.655,46.97
X$14659 1145 VIA_via2_5
* cell instance $14660 r0 *1 51.395,46.83
X$14660 1145 VIA_via1_4
* cell instance $14661 r0 *1 51.395,46.97
X$14661 1145 VIA_via2_5
* cell instance $14662 r0 *1 56.335,46.83
X$14662 1145 VIA_via1_4
* cell instance $14663 r0 *1 56.335,46.97
X$14663 1145 VIA_via2_5
* cell instance $14664 r0 *1 68.685,50.75
X$14664 1145 VIA_via1_4
* cell instance $14665 r0 *1 68.685,50.75
X$14665 1145 VIA_via2_5
* cell instance $14666 r0 *1 67.545,52.43
X$14666 1145 VIA_via1_4
* cell instance $14667 r0 *1 51.775,52.43
X$14667 1145 VIA_via1_4
* cell instance $14668 r0 *1 90.535,56.35
X$14668 1146 VIA_via2_5
* cell instance $14669 r0 *1 70.965,55.79
X$14669 1146 VIA_via2_5
* cell instance $14670 r0 *1 89.775,56.35
X$14670 1146 VIA_via2_5
* cell instance $14671 r0 *1 89.585,55.79
X$14671 1146 VIA_via2_5
* cell instance $14672 r0 *1 70.775,47.11
X$14672 1146 VIA_via1_4
* cell instance $14673 r0 *1 89.585,56.77
X$14673 1146 VIA_via1_4
* cell instance $14674 r0 *1 90.535,56.77
X$14674 1146 VIA_via1_4
* cell instance $14675 r0 *1 71.725,43.19
X$14675 1147 VIA_via1_7
* cell instance $14676 r0 *1 71.345,46.83
X$14676 1147 VIA_via1_4
* cell instance $14677 r0 *1 79.895,44.59
X$14677 1148 VIA_via1_7
* cell instance $14678 r0 *1 79.705,46.83
X$14678 1148 VIA_via1_4
* cell instance $14679 r0 *1 4.655,45.99
X$14679 1149 VIA_via1_7
* cell instance $14680 r0 *1 4.655,45.99
X$14680 1149 VIA_via2_5
* cell instance $14681 r0 *1 2.565,45.99
X$14681 1149 VIA_via2_5
* cell instance $14682 r0 *1 2.565,46.83
X$14682 1149 VIA_via1_4
* cell instance $14683 r0 *1 7.885,46.97
X$14683 1150 VIA_via2_5
* cell instance $14684 r0 *1 5.225,46.83
X$14684 1150 VIA_via1_4
* cell instance $14685 r0 *1 5.225,46.97
X$14685 1150 VIA_via2_5
* cell instance $14686 r0 *1 7.885,47.95
X$14686 1150 VIA_via1_4
* cell instance $14687 r0 *1 8.075,46.83
X$14687 1150 VIA_via1_4
* cell instance $14688 r0 *1 8.075,46.97
X$14688 1150 VIA_via2_5
* cell instance $14689 r0 *1 10.925,46.83
X$14689 1151 VIA_via1_4
* cell instance $14690 r0 *1 10.925,46.69
X$14690 1151 VIA_via2_5
* cell instance $14691 r0 *1 14.535,46.69
X$14691 1151 VIA_via1_4
* cell instance $14692 r0 *1 14.535,46.69
X$14692 1151 VIA_via2_5
* cell instance $14693 r0 *1 91.675,45.99
X$14693 1152 VIA_via1_7
* cell instance $14694 r0 *1 91.675,45.99
X$14694 1152 VIA_via2_5
* cell instance $14695 r0 *1 89.395,60.9
X$14695 1152 VIA_via1_4
* cell instance $14696 r0 *1 89.395,60.97
X$14696 1152 VIA_via2_5
* cell instance $14697 r0 *1 89.415,60.69
X$14697 1152 VIA_via3_2
* cell instance $14698 r0 *1 89.415,45.99
X$14698 1152 VIA_via3_2
* cell instance $14699 r0 *1 90.345,45.99
X$14699 1153 VIA_via1_7
* cell instance $14700 r0 *1 90.345,46.41
X$14700 1153 VIA_via2_5
* cell instance $14701 r0 *1 89.775,62.37
X$14701 1153 VIA_via1_4
* cell instance $14702 r0 *1 89.775,62.51
X$14702 1153 VIA_via2_5
* cell instance $14703 r0 *1 89.975,62.51
X$14703 1153 VIA_via3_2
* cell instance $14704 r0 *1 89.975,46.41
X$14704 1153 VIA_via3_2
* cell instance $14705 r0 *1 88.255,55.09
X$14705 1154 VIA_via2_5
* cell instance $14706 r0 *1 91.865,57.75
X$14706 1154 VIA_via2_5
* cell instance $14707 r0 *1 88.255,48.93
X$14707 1154 VIA_via2_5
* cell instance $14708 r0 *1 88.635,46.55
X$14708 1154 VIA_via2_5
* cell instance $14709 r0 *1 88.635,48.93
X$14709 1154 VIA_via2_5
* cell instance $14710 r0 *1 79.705,46.55
X$14710 1154 VIA_via1_4
* cell instance $14711 r0 *1 79.705,46.55
X$14711 1154 VIA_via2_5
* cell instance $14712 r0 *1 91.865,56.77
X$14712 1154 VIA_via1_4
* cell instance $14713 r0 *1 93.195,55.23
X$14713 1154 VIA_via1_4
* cell instance $14714 r0 *1 93.195,55.09
X$14714 1154 VIA_via2_5
* cell instance $14715 r0 *1 91.655,55.09
X$14715 1154 VIA_via3_2
* cell instance $14716 r0 *1 91.655,57.75
X$14716 1154 VIA_via3_2
* cell instance $14717 r0 *1 8.455,46.97
X$14717 1155 VIA_via1_4
* cell instance $14718 r0 *1 8.455,46.97
X$14718 1155 VIA_via2_5
* cell instance $14719 r0 *1 16.245,46.83
X$14719 1155 VIA_via1_4
* cell instance $14720 r0 *1 16.245,46.97
X$14720 1155 VIA_via2_5
* cell instance $14721 r0 *1 75.715,45.99
X$14721 1156 VIA_via1_7
* cell instance $14722 r0 *1 78.755,46.27
X$14722 1156 VIA_via2_5
* cell instance $14723 r0 *1 75.715,46.27
X$14723 1156 VIA_via2_5
* cell instance $14724 r0 *1 78.755,46.83
X$14724 1156 VIA_via1_4
* cell instance $14725 r0 *1 31.255,74.27
X$14725 1157 VIA_via2_5
* cell instance $14726 r0 *1 28.405,74.55
X$14726 1157 VIA_via2_5
* cell instance $14727 r0 *1 28.785,74.55
X$14727 1157 VIA_via2_5
* cell instance $14728 r0 *1 29.355,74.55
X$14728 1157 VIA_via2_5
* cell instance $14729 r0 *1 62.225,73.99
X$14729 1157 VIA_via2_5
* cell instance $14730 r0 *1 20.045,46.13
X$14730 1157 VIA_via2_5
* cell instance $14731 r0 *1 21.565,54.11
X$14731 1157 VIA_via2_5
* cell instance $14732 r0 *1 21.945,51.87
X$14732 1157 VIA_via2_5
* cell instance $14733 r0 *1 21.565,51.87
X$14733 1157 VIA_via2_5
* cell instance $14734 r0 *1 29.355,61.25
X$14734 1157 VIA_via2_5
* cell instance $14735 r0 *1 29.925,61.25
X$14735 1157 VIA_via2_5
* cell instance $14736 r0 *1 26.125,51.87
X$14736 1157 VIA_via2_5
* cell instance $14737 r0 *1 29.925,51.87
X$14737 1157 VIA_via2_5
* cell instance $14738 r0 *1 28.785,67.13
X$14738 1157 VIA_via2_5
* cell instance $14739 r0 *1 29.925,67.13
X$14739 1157 VIA_via2_5
* cell instance $14740 r0 *1 29.545,62.93
X$14740 1157 VIA_via2_5
* cell instance $14741 r0 *1 30.495,62.93
X$14741 1157 VIA_via2_5
* cell instance $14742 r0 *1 62.225,74.55
X$14742 1157 VIA_via1_4
* cell instance $14743 r0 *1 29.925,59.57
X$14743 1157 VIA_via1_4
* cell instance $14744 r0 *1 26.125,49.63
X$14744 1157 VIA_via1_4
* cell instance $14745 r0 *1 29.355,74.83
X$14745 1157 VIA_via1_4
* cell instance $14746 r0 *1 28.405,76.37
X$14746 1157 VIA_via1_4
* cell instance $14747 r0 *1 20.425,53.97
X$14747 1157 VIA_via1_4
* cell instance $14748 r0 *1 20.425,54.11
X$14748 1157 VIA_via2_5
* cell instance $14749 r0 *1 21.945,51.17
X$14749 1157 VIA_via1_4
* cell instance $14750 r0 *1 29.925,66.43
X$14750 1157 VIA_via1_4
* cell instance $14751 r0 *1 31.255,73.57
X$14751 1157 VIA_via1_4
* cell instance $14752 r0 *1 20.425,48.37
X$14752 1157 VIA_via1_4
* cell instance $14753 r0 *1 20.045,45.57
X$14753 1157 VIA_via1_4
* cell instance $14754 r0 *1 20.255,46.13
X$14754 1157 VIA_via3_2
* cell instance $14755 r0 *1 20.535,48.65
X$14755 1157 VIA_via3_2
* cell instance $14756 r0 *1 20.425,48.65
X$14756 1157 VIA_via2_5
* cell instance $14757 r0 *1 20.535,51.87
X$14757 1157 VIA_via3_2
* cell instance $14758 r0 *1 54.245,51.87
X$14758 1158 VIA_via2_5
* cell instance $14759 r0 *1 55.955,54.53
X$14759 1158 VIA_via2_5
* cell instance $14760 r0 *1 54.245,54.53
X$14760 1158 VIA_via2_5
* cell instance $14761 r0 *1 33.155,51.45
X$14761 1158 VIA_via2_5
* cell instance $14762 r0 *1 42.085,51.87
X$14762 1158 VIA_via2_5
* cell instance $14763 r0 *1 37.905,51.45
X$14763 1158 VIA_via2_5
* cell instance $14764 r0 *1 42.085,51.45
X$14764 1158 VIA_via2_5
* cell instance $14765 r0 *1 20.615,46.13
X$14765 1158 VIA_via2_5
* cell instance $14766 r0 *1 21.375,52.71
X$14766 1158 VIA_via2_5
* cell instance $14767 r0 *1 21.185,49.91
X$14767 1158 VIA_via2_5
* cell instance $14768 r0 *1 21.375,51.45
X$14768 1158 VIA_via2_5
* cell instance $14769 r0 *1 23.085,51.45
X$14769 1158 VIA_via2_5
* cell instance $14770 r0 *1 23.085,49.91
X$14770 1158 VIA_via2_5
* cell instance $14771 r0 *1 18.145,52.71
X$14771 1158 VIA_via2_5
* cell instance $14772 r0 *1 29.925,51.45
X$14772 1158 VIA_via2_5
* cell instance $14773 r0 *1 27.265,51.45
X$14773 1158 VIA_via2_5
* cell instance $14774 r0 *1 42.085,51.17
X$14774 1158 VIA_via1_4
* cell instance $14775 r0 *1 38.095,56.77
X$14775 1158 VIA_via1_4
* cell instance $14776 r0 *1 33.155,51.17
X$14776 1158 VIA_via1_4
* cell instance $14777 r0 *1 27.265,51.17
X$14777 1158 VIA_via1_4
* cell instance $14778 r0 *1 21.375,52.43
X$14778 1158 VIA_via1_4
* cell instance $14779 r0 *1 18.145,53.97
X$14779 1158 VIA_via1_4
* cell instance $14780 r0 *1 21.185,49.63
X$14780 1158 VIA_via1_4
* cell instance $14781 r0 *1 54.245,52.43
X$14781 1158 VIA_via1_4
* cell instance $14782 r0 *1 55.955,54.95
X$14782 1158 VIA_via1_4
* cell instance $14783 r0 *1 30.305,48.37
X$14783 1158 VIA_via1_4
* cell instance $14784 r0 *1 20.615,45.57
X$14784 1158 VIA_via1_4
* cell instance $14785 r0 *1 20.815,46.13
X$14785 1158 VIA_via3_2
* cell instance $14786 r0 *1 20.815,49.91
X$14786 1158 VIA_via3_2
* cell instance $14787 r0 *1 67.355,45.99
X$14787 1159 VIA_via1_7
* cell instance $14788 r0 *1 70.395,46.27
X$14788 1159 VIA_via2_5
* cell instance $14789 r0 *1 67.355,46.27
X$14789 1159 VIA_via2_5
* cell instance $14790 r0 *1 70.395,46.83
X$14790 1159 VIA_via1_4
* cell instance $14791 r0 *1 40.565,45.99
X$14791 1160 VIA_via1_7
* cell instance $14792 r0 *1 40.565,45.99
X$14792 1160 VIA_via2_5
* cell instance $14793 r0 *1 37.905,45.99
X$14793 1160 VIA_via2_5
* cell instance $14794 r0 *1 37.905,46.83
X$14794 1160 VIA_via1_4
* cell instance $14795 r0 *1 68.875,45.99
X$14795 1161 VIA_via1_7
* cell instance $14796 r0 *1 67.735,46.41
X$14796 1161 VIA_via2_5
* cell instance $14797 r0 *1 68.875,46.41
X$14797 1161 VIA_via2_5
* cell instance $14798 r0 *1 67.735,46.83
X$14798 1161 VIA_via1_4
* cell instance $14799 r0 *1 67.355,49.49
X$14799 1162 VIA_via2_5
* cell instance $14800 r0 *1 83.125,52.01
X$14800 1162 VIA_via2_5
* cell instance $14801 r0 *1 79.705,52.01
X$14801 1162 VIA_via2_5
* cell instance $14802 r0 *1 79.705,49.49
X$14802 1162 VIA_via2_5
* cell instance $14803 r0 *1 67.355,46.55
X$14803 1162 VIA_via2_5
* cell instance $14804 r0 *1 57.475,46.55
X$14804 1162 VIA_via1_4
* cell instance $14805 r0 *1 57.475,46.55
X$14805 1162 VIA_via2_5
* cell instance $14806 r0 *1 79.705,52.43
X$14806 1162 VIA_via1_4
* cell instance $14807 r0 *1 83.125,52.43
X$14807 1162 VIA_via1_4
* cell instance $14808 r0 *1 62.795,36.19
X$14808 1163 VIA_via1_7
* cell instance $14809 r0 *1 62.795,46.83
X$14809 1163 VIA_via1_4
* cell instance $14810 r0 *1 52.155,47.81
X$14810 1164 VIA_via1_7
* cell instance $14811 r0 *1 52.155,46.83
X$14811 1164 VIA_via2_5
* cell instance $14812 r0 *1 48.545,46.83
X$14812 1164 VIA_via1_4
* cell instance $14813 r0 *1 48.545,46.83
X$14813 1164 VIA_via2_5
* cell instance $14814 r0 *1 53.485,46.41
X$14814 1165 VIA_via1_7
* cell instance $14815 r0 *1 53.485,46.41
X$14815 1165 VIA_via2_5
* cell instance $14816 r0 *1 52.155,46.41
X$14816 1165 VIA_via2_5
* cell instance $14817 r0 *1 52.155,45.57
X$14817 1165 VIA_via1_4
* cell instance $14818 r0 *1 55.765,46.55
X$14818 1166 VIA_via2_5
* cell instance $14819 r0 *1 54.815,46.55
X$14819 1166 VIA_via1_4
* cell instance $14820 r0 *1 54.815,46.55
X$14820 1166 VIA_via2_5
* cell instance $14821 r0 *1 55.765,46.83
X$14821 1166 VIA_via1_4
* cell instance $14822 r0 *1 5.035,49.21
X$14822 1167 VIA_via1_7
* cell instance $14823 r0 *1 5.035,48.23
X$14823 1167 VIA_via2_5
* cell instance $14824 r0 *1 4.575,48.23
X$14824 1167 VIA_via4_0
* cell instance $14825 r0 *1 4.575,48.23
X$14825 1167 VIA_via3_2
* cell instance $14826 r0 *1 6.175,47.39
X$14826 1168 VIA_via1_7
* cell instance $14827 r0 *1 5.605,48.37
X$14827 1168 VIA_via1_4
* cell instance $14828 r0 *1 22.705,49.91
X$14828 1169 VIA_via1_4
* cell instance $14829 r0 *1 23.085,48.37
X$14829 1169 VIA_via1_4
* cell instance $14830 r0 *1 27.645,51.17
X$14830 1170 VIA_via1_4
* cell instance $14831 r0 *1 27.645,51.17
X$14831 1170 VIA_via2_5
* cell instance $14832 r0 *1 26.885,51.17
X$14832 1170 VIA_via1_4
* cell instance $14833 r0 *1 26.885,51.17
X$14833 1170 VIA_via2_5
* cell instance $14834 r0 *1 27.835,51.17
X$14834 1170 VIA_via1_4
* cell instance $14835 r0 *1 28.025,48.37
X$14835 1170 VIA_via1_4
* cell instance $14836 r0 *1 31.445,50.61
X$14836 1171 VIA_via2_5
* cell instance $14837 r0 *1 32.585,50.61
X$14837 1171 VIA_via2_5
* cell instance $14838 r0 *1 32.585,48.65
X$14838 1171 VIA_via2_5
* cell instance $14839 r0 *1 32.585,49.35
X$14839 1171 VIA_via1_4
* cell instance $14840 r0 *1 31.445,51.17
X$14840 1171 VIA_via1_4
* cell instance $14841 r0 *1 30.685,48.37
X$14841 1171 VIA_via1_4
* cell instance $14842 r0 *1 30.685,48.37
X$14842 1171 VIA_via2_5
* cell instance $14843 r0 *1 28.975,48.37
X$14843 1171 VIA_via1_4
* cell instance $14844 r0 *1 28.975,48.37
X$14844 1171 VIA_via2_5
* cell instance $14845 r0 *1 32.395,48.09
X$14845 1172 VIA_via1_7
* cell instance $14846 r0 *1 32.395,48.09
X$14846 1172 VIA_via2_5
* cell instance $14847 r0 *1 31.255,48.37
X$14847 1172 VIA_via1_4
* cell instance $14848 r0 *1 31.255,48.37
X$14848 1172 VIA_via2_5
* cell instance $14849 r0 *1 35.245,47.39
X$14849 1173 VIA_via1_7
* cell instance $14850 r0 *1 35.055,48.37
X$14850 1173 VIA_via1_4
* cell instance $14851 r0 *1 38.475,54.81
X$14851 1174 VIA_via1_7
* cell instance $14852 r0 *1 38.475,55.65
X$14852 1174 VIA_via1_4
* cell instance $14853 r0 *1 38.475,55.65
X$14853 1174 VIA_via2_5
* cell instance $14854 r0 *1 43.415,48.37
X$14854 1174 VIA_via2_5
* cell instance $14855 r0 *1 46.075,48.37
X$14855 1174 VIA_via2_5
* cell instance $14856 r0 *1 39.045,48.37
X$14856 1174 VIA_via2_5
* cell instance $14857 r0 *1 38.665,48.37
X$14857 1174 VIA_via2_5
* cell instance $14858 r0 *1 40.185,48.37
X$14858 1174 VIA_via2_5
* cell instance $14859 r0 *1 40.185,55.65
X$14859 1174 VIA_via2_5
* cell instance $14860 r0 *1 34.485,55.65
X$14860 1174 VIA_via2_5
* cell instance $14861 r0 *1 38.855,53.97
X$14861 1174 VIA_via1_4
* cell instance $14862 r0 *1 40.185,49.63
X$14862 1174 VIA_via1_4
* cell instance $14863 r0 *1 40.185,56.77
X$14863 1174 VIA_via1_4
* cell instance $14864 r0 *1 40.375,58.03
X$14864 1174 VIA_via1_4
* cell instance $14865 r0 *1 46.075,52.43
X$14865 1174 VIA_via1_4
* cell instance $14866 r0 *1 43.795,45.57
X$14866 1174 VIA_via1_4
* cell instance $14867 r0 *1 38.665,46.83
X$14867 1174 VIA_via1_4
* cell instance $14868 r0 *1 34.485,55.23
X$14868 1174 VIA_via1_4
* cell instance $14869 r0 *1 62.605,57.61
X$14869 1175 VIA_via1_7
* cell instance $14870 r0 *1 60.515,57.19
X$14870 1175 VIA_via2_5
* cell instance $14871 r0 *1 62.605,57.19
X$14871 1175 VIA_via2_5
* cell instance $14872 r0 *1 60.325,49.91
X$14872 1175 VIA_via2_5
* cell instance $14873 r0 *1 58.045,49.21
X$14873 1175 VIA_via2_5
* cell instance $14874 r0 *1 58.045,49.91
X$14874 1175 VIA_via2_5
* cell instance $14875 r0 *1 51.015,49.21
X$14875 1175 VIA_via2_5
* cell instance $14876 r0 *1 46.455,48.37
X$14876 1175 VIA_via2_5
* cell instance $14877 r0 *1 47.025,48.37
X$14877 1175 VIA_via2_5
* cell instance $14878 r0 *1 47.025,59.57
X$14878 1175 VIA_via2_5
* cell instance $14879 r0 *1 50.825,48.37
X$14879 1175 VIA_via2_5
* cell instance $14880 r0 *1 51.015,48.37
X$14880 1175 VIA_via1_4
* cell instance $14881 r0 *1 58.045,48.37
X$14881 1175 VIA_via1_4
* cell instance $14882 r0 *1 48.165,59.57
X$14882 1175 VIA_via1_4
* cell instance $14883 r0 *1 48.165,59.57
X$14883 1175 VIA_via2_5
* cell instance $14884 r0 *1 46.455,46.83
X$14884 1175 VIA_via1_4
* cell instance $14885 r0 *1 60.705,53.97
X$14885 1175 VIA_via1_4
* cell instance $14886 r0 *1 61.655,47.81
X$14886 1176 VIA_via1_7
* cell instance $14887 r0 *1 61.845,46.83
X$14887 1176 VIA_via1_4
* cell instance $14888 r0 *1 53.865,59.85
X$14888 1177 VIA_via2_5
* cell instance $14889 r0 *1 53.855,59.85
X$14889 1177 VIA_via3_2
* cell instance $14890 r0 *1 65.075,67.69
X$14890 1177 VIA_via2_5
* cell instance $14891 r0 *1 65.055,67.69
X$14891 1177 VIA_via3_2
* cell instance $14892 r0 *1 77.615,60.41
X$14892 1177 VIA_via2_5
* cell instance $14893 r0 *1 26.885,71.47
X$14893 1177 VIA_via2_5
* cell instance $14894 r0 *1 34.865,70.91
X$14894 1177 VIA_via2_5
* cell instance $14895 r0 *1 32.775,71.47
X$14895 1177 VIA_via2_5
* cell instance $14896 r0 *1 32.775,70.91
X$14896 1177 VIA_via2_5
* cell instance $14897 r0 *1 46.265,70.91
X$14897 1177 VIA_via2_5
* cell instance $14898 r0 *1 65.075,67.97
X$14898 1177 VIA_via1_4
* cell instance $14899 r0 *1 53.295,70.77
X$14899 1177 VIA_via1_4
* cell instance $14900 r0 *1 53.295,70.77
X$14900 1177 VIA_via2_5
* cell instance $14901 r0 *1 76.855,48.37
X$14901 1177 VIA_via1_4
* cell instance $14902 r0 *1 46.265,74.83
X$14902 1177 VIA_via1_4
* cell instance $14903 r0 *1 34.865,52.85
X$14903 1177 VIA_via1_4
* cell instance $14904 r0 *1 26.695,74.83
X$14904 1177 VIA_via1_4
* cell instance $14905 r0 *1 39.995,67.97
X$14905 1177 VIA_via1_4
* cell instance $14906 r0 *1 39.995,67.97
X$14906 1177 VIA_via2_5
* cell instance $14907 r0 *1 40.135,67.97
X$14907 1177 VIA_via3_2
* cell instance $14908 r0 *1 34.485,70.77
X$14908 1177 VIA_via1_4
* cell instance $14909 r0 *1 34.485,70.91
X$14909 1177 VIA_via2_5
* cell instance $14910 r0 *1 76.095,69.23
X$14910 1177 VIA_via1_4
* cell instance $14911 r0 *1 76.095,69.09
X$14911 1177 VIA_via2_5
* cell instance $14912 r0 *1 75.975,69.09
X$14912 1177 VIA_via3_2
* cell instance $14913 r0 *1 53.675,59.57
X$14913 1177 VIA_via1_4
* cell instance $14914 r0 *1 77.615,60.83
X$14914 1177 VIA_via1_4
* cell instance $14915 r0 *1 65.055,68.11
X$14915 1177 VIA_via4_0
* cell instance $14916 r0 *1 75.975,68.11
X$14916 1177 VIA_via4_0
* cell instance $14917 r0 *1 52.735,67.83
X$14917 1177 VIA_via3_2
* cell instance $14918 r0 *1 53.855,67.69
X$14918 1177 VIA_via3_2
* cell instance $14919 r0 *1 52.735,70.91
X$14919 1177 VIA_via3_2
* cell instance $14920 r0 *1 75.975,60.41
X$14920 1177 VIA_via3_2
* cell instance $14921 r0 *1 75.905,60.41
X$14921 1177 VIA_via2_5
* cell instance $14922 r0 *1 40.135,70.91
X$14922 1177 VIA_via3_2
* cell instance $14923 r0 *1 88.065,49.35
X$14923 1178 VIA_via2_5
* cell instance $14924 r0 *1 88.065,48.37
X$14924 1178 VIA_via1_4
* cell instance $14925 r0 *1 87.875,48.37
X$14925 1178 VIA_via1_4
* cell instance $14926 r0 *1 88.635,49.35
X$14926 1178 VIA_via1_4
* cell instance $14927 r0 *1 88.635,49.35
X$14927 1178 VIA_via2_5
* cell instance $14928 r0 *1 88.825,49.63
X$14928 1178 VIA_via1_4
* cell instance $14929 r0 *1 94.715,48.09
X$14929 1179 VIA_via2_5
* cell instance $14930 r0 *1 93.765,48.09
X$14930 1179 VIA_via1_4
* cell instance $14931 r0 *1 93.765,48.09
X$14931 1179 VIA_via2_5
* cell instance $14932 r0 *1 94.715,48.37
X$14932 1179 VIA_via1_4
* cell instance $14933 r0 *1 92.245,48.23
X$14933 1180 VIA_via1_4
* cell instance $14934 r0 *1 92.245,48.23
X$14934 1180 VIA_via2_5
* cell instance $14935 r0 *1 93.195,48.37
X$14935 1180 VIA_via1_4
* cell instance $14936 r0 *1 93.195,48.23
X$14936 1180 VIA_via2_5
* cell instance $14937 r0 *1 86.545,47.95
X$14937 1181 VIA_via2_5
* cell instance $14938 r0 *1 87.685,47.95
X$14938 1181 VIA_via1_4
* cell instance $14939 r0 *1 87.685,47.95
X$14939 1181 VIA_via2_5
* cell instance $14940 r0 *1 86.545,48.37
X$14940 1181 VIA_via1_4
* cell instance $14941 r0 *1 85.975,48.23
X$14941 1182 VIA_via1_4
* cell instance $14942 r0 *1 85.975,48.23
X$14942 1182 VIA_via2_5
* cell instance $14943 r0 *1 86.735,48.37
X$14943 1182 VIA_via1_4
* cell instance $14944 r0 *1 86.735,48.23
X$14944 1182 VIA_via2_5
* cell instance $14945 r0 *1 76.855,47.81
X$14945 1183 VIA_via1_7
* cell instance $14946 r0 *1 76.855,47.81
X$14946 1183 VIA_via2_5
* cell instance $14947 r0 *1 78.945,47.81
X$14947 1183 VIA_via2_5
* cell instance $14948 r0 *1 78.945,46.83
X$14948 1183 VIA_via1_4
* cell instance $14949 r0 *1 27.265,55.37
X$14949 1184 VIA_via1_7
* cell instance $14950 r0 *1 39.045,66.57
X$14950 1184 VIA_via1_7
* cell instance $14951 r0 *1 39.045,66.71
X$14951 1184 VIA_via2_5
* cell instance $14952 r0 *1 24.225,76.23
X$14952 1184 VIA_via1_7
* cell instance $14953 r0 *1 17.575,74.97
X$14953 1184 VIA_via1_7
* cell instance $14954 r0 *1 14.345,48.23
X$14954 1184 VIA_via1_7
* cell instance $14955 r0 *1 16.435,72.17
X$14955 1184 VIA_via1_7
* cell instance $14956 r0 *1 16.435,72.17
X$14956 1184 VIA_via2_5
* cell instance $14957 r0 *1 18.335,63.77
X$14957 1184 VIA_via1_7
* cell instance $14958 r0 *1 18.335,63.77
X$14958 1184 VIA_via2_5
* cell instance $14959 r0 *1 17.575,72.31
X$14959 1184 VIA_via2_5
* cell instance $14960 r0 *1 17.575,75.53
X$14960 1184 VIA_via2_5
* cell instance $14961 r0 *1 24.415,75.53
X$14961 1184 VIA_via2_5
* cell instance $14962 r0 *1 39.615,55.79
X$14962 1184 VIA_via2_5
* cell instance $14963 r0 *1 14.345,47.67
X$14963 1184 VIA_via2_5
* cell instance $14964 r0 *1 15.105,47.67
X$14964 1184 VIA_via2_5
* cell instance $14965 r0 *1 28.785,47.67
X$14965 1184 VIA_via2_5
* cell instance $14966 r0 *1 39.615,66.71
X$14966 1184 VIA_via2_5
* cell instance $14967 r0 *1 28.785,55.79
X$14967 1184 VIA_via2_5
* cell instance $14968 r0 *1 27.455,55.79
X$14968 1184 VIA_via2_5
* cell instance $14969 r0 *1 29.165,66.99
X$14969 1184 VIA_via2_5
* cell instance $14970 r0 *1 40.375,48.65
X$14970 1184 VIA_via1_4
* cell instance $14971 r0 *1 40.375,48.65
X$14971 1184 VIA_via2_5
* cell instance $14972 r0 *1 40.415,48.65
X$14972 1184 VIA_via3_2
* cell instance $14973 r0 *1 29.165,67.97
X$14973 1184 VIA_via1_4
* cell instance $14974 r0 *1 29.165,68.11
X$14974 1184 VIA_via2_5
* cell instance $14975 r0 *1 42.465,73.57
X$14975 1184 VIA_via1_4
* cell instance $14976 r0 *1 42.465,73.71
X$14976 1184 VIA_via2_5
* cell instance $14977 r0 *1 15.105,45.57
X$14977 1184 VIA_via1_4
* cell instance $14978 r0 *1 23.335,63.77
X$14978 1184 VIA_via3_2
* cell instance $14979 r0 *1 23.335,75.53
X$14979 1184 VIA_via3_2
* cell instance $14980 r0 *1 42.095,66.71
X$14980 1184 VIA_via3_2
* cell instance $14981 r0 *1 23.335,68.11
X$14981 1184 VIA_via3_2
* cell instance $14982 r0 *1 40.415,55.79
X$14982 1184 VIA_via3_2
* cell instance $14983 r0 *1 42.095,73.71
X$14983 1184 VIA_via3_2
* cell instance $14984 r0 *1 75.525,48.23
X$14984 1185 VIA_via2_5
* cell instance $14985 r0 *1 76.285,48.23
X$14985 1185 VIA_via1_4
* cell instance $14986 r0 *1 76.285,48.23
X$14986 1185 VIA_via2_5
* cell instance $14987 r0 *1 75.145,49.63
X$14987 1185 VIA_via1_4
* cell instance $14988 r0 *1 73.625,47.39
X$14988 1186 VIA_via1_7
* cell instance $14989 r0 *1 73.625,47.39
X$14989 1186 VIA_via2_5
* cell instance $14990 r0 *1 71.345,47.39
X$14990 1186 VIA_via2_5
* cell instance $14991 r0 *1 71.345,48.37
X$14991 1186 VIA_via1_4
* cell instance $14992 r0 *1 16.625,47.81
X$14992 1187 VIA_via1_7
* cell instance $14993 r0 *1 16.625,47.81
X$14993 1187 VIA_via2_5
* cell instance $14994 r0 *1 17.195,47.81
X$14994 1187 VIA_via2_5
* cell instance $14995 r0 *1 17.195,46.83
X$14995 1187 VIA_via1_4
* cell instance $14996 r0 *1 18.335,47.81
X$14996 1188 VIA_via1_7
* cell instance $14997 r0 *1 17.195,48.09
X$14997 1188 VIA_via2_5
* cell instance $14998 r0 *1 18.335,48.09
X$14998 1188 VIA_via2_5
* cell instance $14999 r0 *1 17.195,49.63
X$14999 1188 VIA_via1_4
* cell instance $15000 r0 *1 56.715,47.25
X$15000 1189 VIA_via2_5
* cell instance $15001 r0 *1 56.715,46.83
X$15001 1189 VIA_via1_4
* cell instance $15002 r0 *1 55.955,47.11
X$15002 1189 VIA_via1_4
* cell instance $15003 r0 *1 55.955,47.25
X$15003 1189 VIA_via2_5
* cell instance $15004 r0 *1 55.195,47.81
X$15004 1190 VIA_via1_7
* cell instance $15005 r0 *1 55.195,47.81
X$15005 1190 VIA_via2_5
* cell instance $15006 r0 *1 56.525,47.81
X$15006 1190 VIA_via2_5
* cell instance $15007 r0 *1 56.525,46.83
X$15007 1190 VIA_via1_4
* cell instance $15008 r0 *1 47.785,48.09
X$15008 1191 VIA_via2_5
* cell instance $15009 r0 *1 48.165,52.43
X$15009 1191 VIA_via1_4
* cell instance $15010 r0 *1 45.505,48.09
X$15010 1191 VIA_via1_4
* cell instance $15011 r0 *1 45.505,48.09
X$15011 1191 VIA_via2_5
* cell instance $15012 r0 *1 21.565,48.09
X$15012 1192 VIA_via1_7
* cell instance $15013 r0 *1 21.565,46.83
X$15013 1192 VIA_via1_4
* cell instance $15014 r0 *1 22.135,48.09
X$15014 1193 VIA_via2_5
* cell instance $15015 r0 *1 22.135,49.63
X$15015 1193 VIA_via1_4
* cell instance $15016 r0 *1 20.805,48.09
X$15016 1193 VIA_via1_4
* cell instance $15017 r0 *1 20.805,48.09
X$15017 1193 VIA_via2_5
* cell instance $15018 r0 *1 36.005,48.09
X$15018 1194 VIA_via1_7
* cell instance $15019 r0 *1 36.005,48.09
X$15019 1194 VIA_via2_5
* cell instance $15020 r0 *1 33.535,48.09
X$15020 1194 VIA_via2_5
* cell instance $15021 r0 *1 33.535,48.37
X$15021 1194 VIA_via1_4
* cell instance $15022 r0 *1 20.425,47.39
X$15022 1195 VIA_via1_7
* cell instance $15023 r0 *1 20.425,47.39
X$15023 1195 VIA_via2_5
* cell instance $15024 r0 *1 21.945,47.39
X$15024 1195 VIA_via2_5
* cell instance $15025 r0 *1 21.945,48.37
X$15025 1195 VIA_via1_4
* cell instance $15026 r0 *1 33.725,47.95
X$15026 1196 VIA_via1_4
* cell instance $15027 r0 *1 4.275,48.37
X$15027 1196 VIA_via1_4
* cell instance $15028 r0 *1 4.275,48.37
X$15028 1196 VIA_via2_5
* cell instance $15029 r0 *1 6.255,47.39
X$15029 1196 VIA_via4_0
* cell instance $15030 r0 *1 33.695,47.39
X$15030 1196 VIA_via4_0
* cell instance $15031 r0 *1 33.695,47.39
X$15031 1196 VIA_via3_2
* cell instance $15032 r0 *1 33.725,47.39
X$15032 1196 VIA_via2_5
* cell instance $15033 r0 *1 6.255,48.37
X$15033 1196 VIA_via3_2
* cell instance $15034 r0 *1 8.075,47.95
X$15034 1197 VIA_via2_5
* cell instance $15035 r0 *1 25.745,47.95
X$15035 1197 VIA_via1_4
* cell instance $15036 r0 *1 25.745,47.95
X$15036 1197 VIA_via2_5
* cell instance $15037 r0 *1 8.075,48.37
X$15037 1197 VIA_via1_4
* cell instance $15038 r0 *1 82.175,74.97
X$15038 1198 VIA_via2_5
* cell instance $15039 r0 *1 82.555,52.43
X$15039 1198 VIA_via2_5
* cell instance $15040 r0 *1 82.555,52.85
X$15040 1198 VIA_via2_5
* cell instance $15041 r0 *1 81.985,59.57
X$15041 1198 VIA_via2_5
* cell instance $15042 r0 *1 83.695,52.85
X$15042 1198 VIA_via2_5
* cell instance $15043 r0 *1 44.175,48.79
X$15043 1198 VIA_via2_5
* cell instance $15044 r0 *1 36.195,50.19
X$15044 1198 VIA_via2_5
* cell instance $15045 r0 *1 41.135,55.23
X$15045 1198 VIA_via2_5
* cell instance $15046 r0 *1 41.325,50.19
X$15046 1198 VIA_via2_5
* cell instance $15047 r0 *1 44.175,50.19
X$15047 1198 VIA_via2_5
* cell instance $15048 r0 *1 59.375,74.83
X$15048 1198 VIA_via1_4
* cell instance $15049 r0 *1 59.375,74.97
X$15049 1198 VIA_via2_5
* cell instance $15050 r0 *1 82.365,75.95
X$15050 1198 VIA_via1_4
* cell instance $15051 r0 *1 41.135,53.97
X$15051 1198 VIA_via1_4
* cell instance $15052 r0 *1 36.195,49.63
X$15052 1198 VIA_via1_4
* cell instance $15053 r0 *1 32.585,48.37
X$15053 1198 VIA_via1_4
* cell instance $15054 r0 *1 32.585,48.23
X$15054 1198 VIA_via2_5
* cell instance $15055 r0 *1 32.575,48.23
X$15055 1198 VIA_via3_2
* cell instance $15056 r0 *1 45.125,48.37
X$15056 1198 VIA_via1_4
* cell instance $15057 r0 *1 36.765,55.23
X$15057 1198 VIA_via1_4
* cell instance $15058 r0 *1 36.765,55.23
X$15058 1198 VIA_via2_5
* cell instance $15059 r0 *1 54.435,51.17
X$15059 1198 VIA_via1_4
* cell instance $15060 r0 *1 83.885,59.57
X$15060 1198 VIA_via1_4
* cell instance $15061 r0 *1 83.885,59.57
X$15061 1198 VIA_via2_5
* cell instance $15062 r0 *1 80.275,52.43
X$15062 1198 VIA_via1_4
* cell instance $15063 r0 *1 80.275,52.43
X$15063 1198 VIA_via2_5
* cell instance $15064 r0 *1 82.555,51.17
X$15064 1198 VIA_via1_4
* cell instance $15065 r0 *1 74.295,48.51
X$15065 1198 VIA_via4_0
* cell instance $15066 r0 *1 45.175,48.51
X$15066 1198 VIA_via4_0
* cell instance $15067 r0 *1 35.935,48.51
X$15067 1198 VIA_via4_0
* cell instance $15068 r0 *1 32.575,48.51
X$15068 1198 VIA_via4_0
* cell instance $15069 r0 *1 45.175,48.79
X$15069 1198 VIA_via3_2
* cell instance $15070 r0 *1 45.125,48.79
X$15070 1198 VIA_via2_5
* cell instance $15071 r0 *1 35.935,50.19
X$15071 1198 VIA_via3_2
* cell instance $15072 r0 *1 74.295,52.29
X$15072 1198 VIA_via3_2
* cell instance $15073 r0 *1 54.415,48.51
X$15073 1198 VIA_via3_2
* cell instance $15074 r0 *1 54.415,48.51
X$15074 1198 VIA_via4_0
* cell instance $15075 r0 *1 54.435,48.51
X$15075 1198 VIA_via2_5
* cell instance $15076 r0 *1 26.315,47.39
X$15076 1199 VIA_via1_7
* cell instance $15077 r0 *1 26.315,47.39
X$15077 1199 VIA_via2_5
* cell instance $15078 r0 *1 25.935,47.39
X$15078 1199 VIA_via2_5
* cell instance $15079 r0 *1 25.935,48.37
X$15079 1199 VIA_via1_4
* cell instance $15080 r0 *1 8.455,48.79
X$15080 1200 VIA_via1_7
* cell instance $15081 r0 *1 8.455,48.79
X$15081 1200 VIA_via2_5
* cell instance $15082 r0 *1 8.495,48.79
X$15082 1200 VIA_via3_2
* cell instance $15083 r0 *1 8.495,48.79
X$15083 1200 VIA_via4_0
* cell instance $15084 r0 *1 4.655,48.23
X$15084 1201 VIA_via1_4
* cell instance $15085 r0 *1 4.575,49.07
X$15085 1201 VIA_via3_2
* cell instance $15086 r0 *1 4.575,49.07
X$15086 1201 VIA_via4_0
* cell instance $15087 r0 *1 4.655,49.07
X$15087 1201 VIA_via2_5
* cell instance $15088 r0 *1 17.385,49.91
X$15088 1202 VIA_via1_7
* cell instance $15089 r0 *1 17.385,49.91
X$15089 1202 VIA_via2_5
* cell instance $15090 r0 *1 4.655,49.63
X$15090 1202 VIA_via1_4
* cell instance $15091 r0 *1 4.655,49.77
X$15091 1202 VIA_via2_5
* cell instance $15092 r0 *1 13.775,48.79
X$15092 1203 VIA_via1_7
* cell instance $15093 r0 *1 13.205,49.63
X$15093 1203 VIA_via1_4
* cell instance $15094 r0 *1 15.485,49.35
X$15094 1204 VIA_via1_4
* cell instance $15095 r0 *1 12.825,48.37
X$15095 1204 VIA_via1_4
* cell instance $15096 r0 *1 12.825,48.37
X$15096 1204 VIA_via2_5
* cell instance $15097 r0 *1 15.105,48.37
X$15097 1204 VIA_via1_4
* cell instance $15098 r0 *1 15.105,48.37
X$15098 1204 VIA_via2_5
* cell instance $15099 r0 *1 23.085,48.65
X$15099 1205 VIA_via2_5
* cell instance $15100 r0 *1 21.375,48.65
X$15100 1205 VIA_via2_5
* cell instance $15101 r0 *1 21.755,48.65
X$15101 1205 VIA_via2_5
* cell instance $15102 r0 *1 21.565,49.63
X$15102 1205 VIA_via1_4
* cell instance $15103 r0 *1 23.085,49.63
X$15103 1205 VIA_via1_4
* cell instance $15104 r0 *1 25.365,48.65
X$15104 1205 VIA_via1_4
* cell instance $15105 r0 *1 25.365,48.65
X$15105 1205 VIA_via2_5
* cell instance $15106 r0 *1 21.755,45.57
X$15106 1205 VIA_via1_4
* cell instance $15107 r0 *1 70.965,74.41
X$15107 1206 VIA_via1_7
* cell instance $15108 r0 *1 70.965,71.05
X$15108 1206 VIA_via2_5
* cell instance $15109 r0 *1 34.485,48.93
X$15109 1206 VIA_via2_5
* cell instance $15110 r0 *1 30.875,48.93
X$15110 1206 VIA_via2_5
* cell instance $15111 r0 *1 20.995,49.77
X$15111 1206 VIA_via2_5
* cell instance $15112 r0 *1 30.305,71.19
X$15112 1206 VIA_via2_5
* cell instance $15113 r0 *1 29.735,62.51
X$15113 1206 VIA_via2_5
* cell instance $15114 r0 *1 21.945,53.83
X$15114 1206 VIA_via2_5
* cell instance $15115 r0 *1 24.225,52.57
X$15115 1206 VIA_via2_5
* cell instance $15116 r0 *1 31.065,62.65
X$15116 1206 VIA_via2_5
* cell instance $15117 r0 *1 34.485,49.63
X$15117 1206 VIA_via1_4
* cell instance $15118 r0 *1 30.875,48.37
X$15118 1206 VIA_via1_4
* cell instance $15119 r0 *1 21.945,52.43
X$15119 1206 VIA_via1_4
* cell instance $15120 r0 *1 21.945,52.57
X$15120 1206 VIA_via2_5
* cell instance $15121 r0 *1 18.715,53.97
X$15121 1206 VIA_via1_4
* cell instance $15122 r0 *1 18.715,53.83
X$15122 1206 VIA_via2_5
* cell instance $15123 r0 *1 21.755,49.63
X$15123 1206 VIA_via1_4
* cell instance $15124 r0 *1 21.755,49.77
X$15124 1206 VIA_via2_5
* cell instance $15125 r0 *1 24.035,49.63
X$15125 1206 VIA_via1_4
* cell instance $15126 r0 *1 24.035,49.77
X$15126 1206 VIA_via2_5
* cell instance $15127 r0 *1 29.735,62.3
X$15127 1206 VIA_via1_4
* cell instance $15128 r0 *1 30.305,70.77
X$15128 1206 VIA_via1_4
* cell instance $15129 r0 *1 31.065,63.63
X$15129 1206 VIA_via1_4
* cell instance $15130 r0 *1 20.995,48.37
X$15130 1206 VIA_via1_4
* cell instance $15131 r0 *1 30.335,52.57
X$15131 1206 VIA_via3_2
* cell instance $15132 r0 *1 30.335,48.93
X$15132 1206 VIA_via3_2
* cell instance $15133 r0 *1 30.335,62.65
X$15133 1206 VIA_via3_2
* cell instance $15134 r0 *1 21.565,49.35
X$15134 1207 VIA_via1_4
* cell instance $15135 r0 *1 21.945,49.63
X$15135 1207 VIA_via1_4
* cell instance $15136 r0 *1 47.215,71.61
X$15136 1208 VIA_via1_7
* cell instance $15137 r0 *1 31.255,49.91
X$15137 1208 VIA_via2_5
* cell instance $15138 r0 *1 33.725,49.91
X$15138 1208 VIA_via2_5
* cell instance $15139 r0 *1 35.055,49.91
X$15139 1208 VIA_via2_5
* cell instance $15140 r0 *1 22.325,48.37
X$15140 1208 VIA_via2_5
* cell instance $15141 r0 *1 47.595,63.91
X$15141 1208 VIA_via2_5
* cell instance $15142 r0 *1 19.285,52.01
X$15142 1208 VIA_via2_5
* cell instance $15143 r0 *1 22.325,50.61
X$15143 1208 VIA_via2_5
* cell instance $15144 r0 *1 22.325,49.35
X$15144 1208 VIA_via2_5
* cell instance $15145 r0 *1 24.605,49.35
X$15145 1208 VIA_via2_5
* cell instance $15146 r0 *1 22.705,52.01
X$15146 1208 VIA_via2_5
* cell instance $15147 r0 *1 22.705,50.61
X$15147 1208 VIA_via2_5
* cell instance $15148 r0 *1 36.765,54.25
X$15148 1208 VIA_via2_5
* cell instance $15149 r0 *1 33.725,54.25
X$15149 1208 VIA_via2_5
* cell instance $15150 r0 *1 32.205,54.53
X$15150 1208 VIA_via2_5
* cell instance $15151 r0 *1 33.535,54.53
X$15151 1208 VIA_via2_5
* cell instance $15152 r0 *1 31.255,49.35
X$15152 1208 VIA_via2_5
* cell instance $15153 r0 *1 30.305,62.09
X$15153 1208 VIA_via2_5
* cell instance $15154 r0 *1 31.635,62.09
X$15154 1208 VIA_via2_5
* cell instance $15155 r0 *1 32.205,62.09
X$15155 1208 VIA_via2_5
* cell instance $15156 r0 *1 36.765,53.97
X$15156 1208 VIA_via1_4
* cell instance $15157 r0 *1 35.055,49.63
X$15157 1208 VIA_via1_4
* cell instance $15158 r0 *1 31.445,48.37
X$15158 1208 VIA_via1_4
* cell instance $15159 r0 *1 22.515,52.43
X$15159 1208 VIA_via1_4
* cell instance $15160 r0 *1 19.285,53.97
X$15160 1208 VIA_via1_4
* cell instance $15161 r0 *1 22.325,49.63
X$15161 1208 VIA_via1_4
* cell instance $15162 r0 *1 24.605,49.63
X$15162 1208 VIA_via1_4
* cell instance $15163 r0 *1 30.305,62.37
X$15163 1208 VIA_via1_4
* cell instance $15164 r0 *1 31.635,63.63
X$15164 1208 VIA_via1_4
* cell instance $15165 r0 *1 31.635,63.63
X$15165 1208 VIA_via2_5
* cell instance $15166 r0 *1 21.565,48.37
X$15166 1208 VIA_via1_4
* cell instance $15167 r0 *1 21.565,48.37
X$15167 1208 VIA_via2_5
* cell instance $15168 r0 *1 27.645,49.91
X$15168 1209 VIA_via2_5
* cell instance $15169 r0 *1 27.535,49.91
X$15169 1209 VIA_via3_2
* cell instance $15170 r0 *1 27.645,49.91
X$15170 1209 VIA_via1_7
* cell instance $15171 r0 *1 5.225,49.63
X$15171 1209 VIA_via1_4
* cell instance $15172 r0 *1 5.225,49.63
X$15172 1209 VIA_via2_5
* cell instance $15173 r0 *1 27.535,49.35
X$15173 1209 VIA_via4_0
* cell instance $15174 r0 *1 6.255,49.63
X$15174 1209 VIA_via3_2
* cell instance $15175 r0 *1 6.255,49.63
X$15175 1209 VIA_via4_0
* cell instance $15176 r0 *1 43.795,54.95
X$15176 1210 VIA_via1_7
* cell instance $15177 r0 *1 43.795,54.81
X$15177 1210 VIA_via2_5
* cell instance $15178 r0 *1 20.615,51.31
X$15178 1210 VIA_via2_5
* cell instance $15179 r0 *1 27.645,49.49
X$15179 1210 VIA_via2_5
* cell instance $15180 r0 *1 29.355,54.81
X$15180 1210 VIA_via2_5
* cell instance $15181 r0 *1 28.405,49.49
X$15181 1210 VIA_via1_4
* cell instance $15182 r0 *1 28.405,49.49
X$15182 1210 VIA_via2_5
* cell instance $15183 r0 *1 29.165,49.63
X$15183 1210 VIA_via1_7
* cell instance $15184 r0 *1 20.615,52.29
X$15184 1210 VIA_via1_4
* cell instance $15185 r0 *1 20.615,49.49
X$15185 1210 VIA_via1_4
* cell instance $15186 r0 *1 20.615,49.49
X$15186 1210 VIA_via2_5
* cell instance $15187 r0 *1 19.285,51.31
X$15187 1210 VIA_via1_4
* cell instance $15188 r0 *1 19.285,51.31
X$15188 1210 VIA_via2_5
* cell instance $15189 r0 *1 27.645,48.51
X$15189 1210 VIA_via1_4
* cell instance $15190 r0 *1 28.975,49.63
X$15190 1211 VIA_via1_4
* cell instance $15191 r0 *1 29.165,48.51
X$15191 1211 VIA_via1_4
* cell instance $15192 r0 *1 30.685,48.79
X$15192 1212 VIA_via1_7
* cell instance $15193 r0 *1 31.065,48.37
X$15193 1212 VIA_via1_4
* cell instance $15194 r0 *1 39.995,52.15
X$15194 1213 VIA_via1_7
* cell instance $15195 r0 *1 30.115,49.07
X$15195 1213 VIA_via2_5
* cell instance $15196 r0 *1 18.145,49.07
X$15196 1213 VIA_via2_5
* cell instance $15197 r0 *1 38.285,48.65
X$15197 1213 VIA_via2_5
* cell instance $15198 r0 *1 39.995,49.63
X$15198 1213 VIA_via2_5
* cell instance $15199 r0 *1 35.245,48.93
X$15199 1213 VIA_via2_5
* cell instance $15200 r0 *1 38.285,49.63
X$15200 1213 VIA_via1_4
* cell instance $15201 r0 *1 38.285,49.63
X$15201 1213 VIA_via2_5
* cell instance $15202 r0 *1 30.305,55.09
X$15202 1213 VIA_via1_4
* cell instance $15203 r0 *1 35.245,48.51
X$15203 1213 VIA_via1_4
* cell instance $15204 r0 *1 35.245,48.65
X$15204 1213 VIA_via2_5
* cell instance $15205 r0 *1 41.895,49.63
X$15205 1213 VIA_via1_4
* cell instance $15206 r0 *1 41.895,49.77
X$15206 1213 VIA_via2_5
* cell instance $15207 r0 *1 18.145,49.77
X$15207 1213 VIA_via1_4
* cell instance $15208 r0 *1 61.085,56.21
X$15208 1214 VIA_via1_7
* cell instance $15209 r0 *1 47.975,48.79
X$15209 1214 VIA_via2_5
* cell instance $15210 r0 *1 61.085,48.51
X$15210 1214 VIA_via2_5
* cell instance $15211 r0 *1 49.685,48.79
X$15211 1214 VIA_via2_5
* cell instance $15212 r0 *1 49.685,48.37
X$15212 1214 VIA_via1_4
* cell instance $15213 r0 *1 59.375,48.37
X$15213 1214 VIA_via1_4
* cell instance $15214 r0 *1 59.375,48.51
X$15214 1214 VIA_via2_5
* cell instance $15215 r0 *1 47.975,48.37
X$15215 1214 VIA_via1_4
* cell instance $15216 r0 *1 49.685,56.77
X$15216 1214 VIA_via1_4
* cell instance $15217 r0 *1 61.085,51.17
X$15217 1214 VIA_via1_4
* cell instance $15218 r0 *1 50.825,48.79
X$15218 1215 VIA_via1_7
* cell instance $15219 r0 *1 51.585,49.63
X$15219 1215 VIA_via1_4
* cell instance $15220 r0 *1 60.325,49.35
X$15220 1216 VIA_via2_5
* cell instance $15221 r0 *1 58.235,49.35
X$15221 1216 VIA_via2_5
* cell instance $15222 r0 *1 58.235,48.37
X$15222 1216 VIA_via1_4
* cell instance $15223 r0 *1 59.945,49.35
X$15223 1216 VIA_via1_4
* cell instance $15224 r0 *1 59.945,49.35
X$15224 1216 VIA_via2_5
* cell instance $15225 r0 *1 60.325,49.63
X$15225 1216 VIA_via1_4
* cell instance $15226 r0 *1 60.895,48.37
X$15226 1217 VIA_via2_5
* cell instance $15227 r0 *1 59.565,48.37
X$15227 1217 VIA_via1_4
* cell instance $15228 r0 *1 59.565,48.37
X$15228 1217 VIA_via2_5
* cell instance $15229 r0 *1 60.895,50.75
X$15229 1217 VIA_via1_4
* cell instance $15230 r0 *1 60.895,49.63
X$15230 1217 VIA_via1_4
* cell instance $15231 r0 *1 62.225,49.77
X$15231 1218 VIA_via2_5
* cell instance $15232 r0 *1 83.315,50.33
X$15232 1218 VIA_via2_5
* cell instance $15233 r0 *1 81.985,49.91
X$15233 1218 VIA_via2_5
* cell instance $15234 r0 *1 81.985,50.33
X$15234 1218 VIA_via2_5
* cell instance $15235 r0 *1 62.225,47.11
X$15235 1218 VIA_via1_4
* cell instance $15236 r0 *1 83.315,51.17
X$15236 1218 VIA_via1_4
* cell instance $15237 r0 *1 81.985,51.17
X$15237 1218 VIA_via1_4
* cell instance $15238 r0 *1 72.295,75.81
X$15238 1219 VIA_via1_7
* cell instance $15239 r0 *1 72.295,71.19
X$15239 1219 VIA_via2_5
* cell instance $15240 r0 *1 70.205,71.19
X$15240 1219 VIA_via2_5
* cell instance $15241 r0 *1 70.015,49.77
X$15241 1219 VIA_via2_5
* cell instance $15242 r0 *1 69.825,49.63
X$15242 1219 VIA_via1_4
* cell instance $15243 r0 *1 71.345,49.77
X$15243 1219 VIA_via1_4
* cell instance $15244 r0 *1 71.345,49.77
X$15244 1219 VIA_via2_5
* cell instance $15245 r0 *1 70.015,52.43
X$15245 1219 VIA_via1_4
* cell instance $15246 r0 *1 70.015,51.17
X$15246 1219 VIA_via1_4
* cell instance $15247 r0 *1 70.205,51.03
X$15247 1220 VIA_via2_5
* cell instance $15248 r0 *1 70.775,51.03
X$15248 1220 VIA_via1_4
* cell instance $15249 r0 *1 70.775,51.03
X$15249 1220 VIA_via2_5
* cell instance $15250 r0 *1 70.395,49.63
X$15250 1220 VIA_via1_4
* cell instance $15251 r0 *1 69.825,51.17
X$15251 1220 VIA_via1_4
* cell instance $15252 r0 *1 69.825,51.03
X$15252 1220 VIA_via2_5
* cell instance $15253 r0 *1 72.675,48.51
X$15253 1221 VIA_via2_5
* cell instance $15254 r0 *1 73.625,48.51
X$15254 1221 VIA_via1_4
* cell instance $15255 r0 *1 73.625,48.51
X$15255 1221 VIA_via2_5
* cell instance $15256 r0 *1 74.005,48.37
X$15256 1221 VIA_via1_4
* cell instance $15257 r0 *1 74.005,48.51
X$15257 1221 VIA_via2_5
* cell instance $15258 r0 *1 72.675,46.83
X$15258 1221 VIA_via1_4
* cell instance $15259 r0 *1 77.425,48.51
X$15259 1222 VIA_via2_5
* cell instance $15260 r0 *1 74.575,48.37
X$15260 1222 VIA_via1_4
* cell instance $15261 r0 *1 74.575,48.51
X$15261 1222 VIA_via2_5
* cell instance $15262 r0 *1 75.335,48.37
X$15262 1222 VIA_via1_4
* cell instance $15263 r0 *1 75.335,48.51
X$15263 1222 VIA_via2_5
* cell instance $15264 r0 *1 77.425,49.35
X$15264 1222 VIA_via1_4
* cell instance $15265 r0 *1 86.735,53.97
X$15265 1223 VIA_via2_5
* cell instance $15266 r0 *1 87.305,53.97
X$15266 1223 VIA_via2_5
* cell instance $15267 r0 *1 80.465,53.97
X$15267 1223 VIA_via2_5
* cell instance $15268 r0 *1 78.945,53.97
X$15268 1223 VIA_via2_5
* cell instance $15269 r0 *1 78.945,49.63
X$15269 1223 VIA_via2_5
* cell instance $15270 r0 *1 87.115,49.63
X$15270 1223 VIA_via1_4
* cell instance $15271 r0 *1 75.905,49.63
X$15271 1223 VIA_via1_4
* cell instance $15272 r0 *1 75.905,49.63
X$15272 1223 VIA_via2_5
* cell instance $15273 r0 *1 78.945,51.17
X$15273 1223 VIA_via1_4
* cell instance $15274 r0 *1 80.465,55.23
X$15274 1223 VIA_via1_4
* cell instance $15275 r0 *1 87.305,55.23
X$15275 1223 VIA_via1_4
* cell instance $15276 r0 *1 81.795,49.63
X$15276 1223 VIA_via1_4
* cell instance $15277 r0 *1 81.795,49.63
X$15277 1223 VIA_via2_5
* cell instance $15278 r0 *1 82.935,52.85
X$15278 1223 VIA_via1_4
* cell instance $15279 r0 *1 80.085,53.97
X$15279 1223 VIA_via1_4
* cell instance $15280 r0 *1 80.085,53.97
X$15280 1223 VIA_via2_5
* cell instance $15281 r0 *1 83.125,53.97
X$15281 1223 VIA_via1_4
* cell instance $15282 r0 *1 83.125,53.97
X$15282 1223 VIA_via2_5
* cell instance $15283 r0 *1 90.725,63.21
X$15283 1224 VIA_via1_7
* cell instance $15284 r0 *1 90.725,64.19
X$15284 1224 VIA_via1_7
* cell instance $15285 r0 *1 91.485,57.33
X$15285 1224 VIA_via2_5
* cell instance $15286 r0 *1 90.535,57.33
X$15286 1224 VIA_via2_5
* cell instance $15287 r0 *1 86.165,49.49
X$15287 1224 VIA_via2_5
* cell instance $15288 r0 *1 84.075,49.49
X$15288 1224 VIA_via2_5
* cell instance $15289 r0 *1 92.435,49.35
X$15289 1224 VIA_via2_5
* cell instance $15290 r0 *1 90.725,63.91
X$15290 1224 VIA_via2_5
* cell instance $15291 r0 *1 86.165,48.37
X$15291 1224 VIA_via1_4
* cell instance $15292 r0 *1 92.435,48.37
X$15292 1224 VIA_via1_4
* cell instance $15293 r0 *1 90.345,65.17
X$15293 1224 VIA_via1_4
* cell instance $15294 r0 *1 92.815,63.63
X$15294 1224 VIA_via1_4
* cell instance $15295 r0 *1 92.815,63.63
X$15295 1224 VIA_via2_5
* cell instance $15296 r0 *1 91.675,52.43
X$15296 1224 VIA_via1_4
* cell instance $15297 r0 *1 91.675,52.29
X$15297 1224 VIA_via2_5
* cell instance $15298 r0 *1 90.725,49.63
X$15298 1224 VIA_via1_4
* cell instance $15299 r0 *1 90.725,49.49
X$15299 1224 VIA_via2_5
* cell instance $15300 r0 *1 92.815,56.77
X$15300 1224 VIA_via1_4
* cell instance $15301 r0 *1 92.815,56.91
X$15301 1224 VIA_via2_5
* cell instance $15302 r0 *1 91.485,56.77
X$15302 1224 VIA_via1_4
* cell instance $15303 r0 *1 91.485,56.91
X$15303 1224 VIA_via2_5
* cell instance $15304 r0 *1 84.075,51.17
X$15304 1224 VIA_via1_4
* cell instance $15305 r0 *1 83.885,52.43
X$15305 1224 VIA_via1_4
* cell instance $15306 r0 *1 92.495,52.29
X$15306 1224 VIA_via3_2
* cell instance $15307 r0 *1 92.495,56.91
X$15307 1224 VIA_via3_2
* cell instance $15308 r0 *1 91.935,52.29
X$15308 1224 VIA_via3_2
* cell instance $15309 r0 *1 91.935,49.49
X$15309 1224 VIA_via3_2
* cell instance $15310 r0 *1 90.915,57.75
X$15310 1225 VIA_via2_5
* cell instance $15311 r0 *1 90.815,57.75
X$15311 1225 VIA_via3_2
* cell instance $15312 r0 *1 85.975,56.21
X$15312 1225 VIA_via2_5
* cell instance $15313 r0 *1 91.105,60.83
X$15313 1225 VIA_via2_5
* cell instance $15314 r0 *1 91.105,59.43
X$15314 1225 VIA_via2_5
* cell instance $15315 r0 *1 90.915,50.75
X$15315 1225 VIA_via2_5
* cell instance $15316 r0 *1 86.545,51.73
X$15316 1225 VIA_via2_5
* cell instance $15317 r0 *1 84.835,51.73
X$15317 1225 VIA_via2_5
* cell instance $15318 r0 *1 84.265,51.73
X$15318 1225 VIA_via2_5
* cell instance $15319 r0 *1 92.815,50.75
X$15319 1225 VIA_via2_5
* cell instance $15320 r0 *1 86.355,48.37
X$15320 1225 VIA_via1_4
* cell instance $15321 r0 *1 92.815,48.37
X$15321 1225 VIA_via1_4
* cell instance $15322 r0 *1 91.485,61.95
X$15322 1225 VIA_via1_4
* cell instance $15323 r0 *1 90.915,51.17
X$15323 1225 VIA_via1_4
* cell instance $15324 r0 *1 90.725,54.04
X$15324 1225 VIA_via1_4
* cell instance $15325 r0 *1 90.725,54.11
X$15325 1225 VIA_via2_5
* cell instance $15326 r0 *1 91.485,60.83
X$15326 1225 VIA_via1_4
* cell instance $15327 r0 *1 91.485,60.83
X$15327 1225 VIA_via2_5
* cell instance $15328 r0 *1 85.975,56.77
X$15328 1225 VIA_via1_4
* cell instance $15329 r0 *1 84.265,51.17
X$15329 1225 VIA_via1_4
* cell instance $15330 r0 *1 92.435,59.57
X$15330 1225 VIA_via1_4
* cell instance $15331 r0 *1 92.435,59.43
X$15331 1225 VIA_via2_5
* cell instance $15332 r0 *1 84.835,52.43
X$15332 1225 VIA_via1_4
* cell instance $15333 r0 *1 84.075,52.43
X$15333 1225 VIA_via1_4
* cell instance $15334 r0 *1 90.535,51.73
X$15334 1225 VIA_via3_2
* cell instance $15335 r0 *1 90.535,50.75
X$15335 1225 VIA_via3_2
* cell instance $15336 r0 *1 90.535,54.11
X$15336 1225 VIA_via3_2
* cell instance $15337 r0 *1 90.815,56.21
X$15337 1225 VIA_via3_2
* cell instance $15338 r0 *1 90.725,56.21
X$15338 1225 VIA_via2_5
* cell instance $15339 r0 *1 94.715,75.53
X$15339 1226 VIA_via2_5
* cell instance $15340 r0 *1 93.575,75.53
X$15340 1226 VIA_via2_5
* cell instance $15341 r0 *1 88.445,75.53
X$15341 1226 VIA_via2_5
* cell instance $15342 r0 *1 86.545,59.15
X$15342 1226 VIA_via2_5
* cell instance $15343 r0 *1 91.485,51.73
X$15343 1226 VIA_via2_5
* cell instance $15344 r0 *1 93.195,59.85
X$15344 1226 VIA_via2_5
* cell instance $15345 r0 *1 92.055,60.55
X$15345 1226 VIA_via2_5
* cell instance $15346 r0 *1 93.195,60.55
X$15346 1226 VIA_via2_5
* cell instance $15347 r0 *1 86.925,48.79
X$15347 1226 VIA_via2_5
* cell instance $15348 r0 *1 86.925,48.37
X$15348 1226 VIA_via1_4
* cell instance $15349 r0 *1 93.385,48.37
X$15349 1226 VIA_via1_4
* cell instance $15350 r0 *1 93.385,48.51
X$15350 1226 VIA_via2_5
* cell instance $15351 r0 *1 87.495,74.83
X$15351 1226 VIA_via1_4
* cell instance $15352 r0 *1 87.495,74.83
X$15352 1226 VIA_via2_5
* cell instance $15353 r0 *1 88.065,74.83
X$15353 1226 VIA_via1_4
* cell instance $15354 r0 *1 88.065,74.83
X$15354 1226 VIA_via2_5
* cell instance $15355 r0 *1 88.445,75.25
X$15355 1226 VIA_via1_4
* cell instance $15356 r0 *1 94.715,76.37
X$15356 1226 VIA_via1_4
* cell instance $15357 r0 *1 93.575,66.43
X$15357 1226 VIA_via1_4
* cell instance $15358 r0 *1 91.485,51.17
X$15358 1226 VIA_via1_4
* cell instance $15359 r0 *1 91.295,53.97
X$15359 1226 VIA_via1_4
* cell instance $15360 r0 *1 91.295,53.97
X$15360 1226 VIA_via2_5
* cell instance $15361 r0 *1 86.545,56.77
X$15361 1226 VIA_via1_4
* cell instance $15362 r0 *1 92.055,60.83
X$15362 1226 VIA_via1_4
* cell instance $15363 r0 *1 93.005,59.57
X$15363 1226 VIA_via1_4
* cell instance $15364 r0 *1 91.095,51.73
X$15364 1226 VIA_via3_2
* cell instance $15365 r0 *1 91.095,59.15
X$15365 1226 VIA_via3_2
* cell instance $15366 r0 *1 92.775,59.15
X$15366 1226 VIA_via3_2
* cell instance $15367 r0 *1 92.775,59.85
X$15367 1226 VIA_via3_2
* cell instance $15368 r0 *1 91.095,53.97
X$15368 1226 VIA_via3_2
* cell instance $15369 r0 *1 91.095,48.65
X$15369 1226 VIA_via3_2
* cell instance $15370 r0 *1 87.685,58.17
X$15370 1227 VIA_via2_5
* cell instance $15371 r0 *1 91.295,58.17
X$15371 1227 VIA_via2_5
* cell instance $15372 r0 *1 94.715,58.03
X$15372 1227 VIA_via2_5
* cell instance $15373 r0 *1 92.625,58.03
X$15373 1227 VIA_via2_5
* cell instance $15374 r0 *1 93.575,58.03
X$15374 1227 VIA_via1_4
* cell instance $15375 r0 *1 93.575,58.03
X$15375 1227 VIA_via2_5
* cell instance $15376 r0 *1 91.485,58.17
X$15376 1227 VIA_via1_4
* cell instance $15377 r0 *1 91.485,58.17
X$15377 1227 VIA_via2_5
* cell instance $15378 r0 *1 90.725,58.03
X$15378 1227 VIA_via1_4
* cell instance $15379 r0 *1 90.725,58.17
X$15379 1227 VIA_via2_5
* cell instance $15380 r0 *1 87.685,59.57
X$15380 1227 VIA_via1_4
* cell instance $15381 r0 *1 86.735,60.83
X$15381 1227 VIA_via1_4
* cell instance $15382 r0 *1 92.435,49.63
X$15382 1227 VIA_via1_4
* cell instance $15383 r0 *1 91.295,55.23
X$15383 1227 VIA_via1_4
* cell instance $15384 r0 *1 94.905,60.83
X$15384 1227 VIA_via1_4
* cell instance $15385 r0 *1 87.115,57.61
X$15385 1228 VIA_via2_5
* cell instance $15386 r0 *1 90.915,59.71
X$15386 1228 VIA_via2_5
* cell instance $15387 r0 *1 87.495,49.21
X$15387 1228 VIA_via2_5
* cell instance $15388 r0 *1 94.145,49.21
X$15388 1228 VIA_via2_5
* cell instance $15389 r0 *1 93.005,49.21
X$15389 1228 VIA_via2_5
* cell instance $15390 r0 *1 93.005,53.55
X$15390 1228 VIA_via2_5
* cell instance $15391 r0 *1 92.055,66.71
X$15391 1228 VIA_via2_5
* cell instance $15392 r0 *1 94.145,66.15
X$15392 1228 VIA_via2_5
* cell instance $15393 r0 *1 91.105,66.71
X$15393 1228 VIA_via2_5
* cell instance $15394 r0 *1 92.055,66.15
X$15394 1228 VIA_via2_5
* cell instance $15395 r0 *1 80.275,67.41
X$15395 1228 VIA_via2_5
* cell instance $15396 r0 *1 79.135,67.41
X$15396 1228 VIA_via2_5
* cell instance $15397 r0 *1 87.495,48.37
X$15397 1228 VIA_via1_4
* cell instance $15398 r0 *1 79.325,67.97
X$15398 1228 VIA_via1_4
* cell instance $15399 r0 *1 94.145,66.43
X$15399 1228 VIA_via1_4
* cell instance $15400 r0 *1 92.055,66.43
X$15400 1228 VIA_via1_4
* cell instance $15401 r0 *1 87.115,56.77
X$15401 1228 VIA_via1_4
* cell instance $15402 r0 *1 94.145,49.63
X$15402 1228 VIA_via1_4
* cell instance $15403 r0 *1 91.865,53.97
X$15403 1228 VIA_via1_4
* cell instance $15404 r0 *1 93.005,51.17
X$15404 1228 VIA_via1_4
* cell instance $15405 r0 *1 80.275,66.85
X$15405 1228 VIA_via1_4
* cell instance $15406 r0 *1 80.275,66.71
X$15406 1228 VIA_via2_5
* cell instance $15407 r0 *1 93.575,59.57
X$15407 1228 VIA_via1_4
* cell instance $15408 r0 *1 93.575,59.71
X$15408 1228 VIA_via2_5
* cell instance $15409 r0 *1 91.865,59.57
X$15409 1228 VIA_via1_4
* cell instance $15410 r0 *1 91.865,59.57
X$15410 1228 VIA_via2_5
* cell instance $15411 r0 *1 91.935,53.55
X$15411 1228 VIA_via3_2
* cell instance $15412 r0 *1 91.865,53.55
X$15412 1228 VIA_via2_5
* cell instance $15413 r0 *1 91.935,57.61
X$15413 1228 VIA_via3_2
* cell instance $15414 r0 *1 91.935,58.73
X$15414 1228 VIA_via3_2
* cell instance $15415 r0 *1 91.865,58.73
X$15415 1228 VIA_via2_5
* cell instance $15416 r0 *1 93.005,48.37
X$15416 1229 VIA_via1_4
* cell instance $15417 r0 *1 94.335,49.49
X$15417 1229 VIA_via1_4
* cell instance $15418 r0 *1 88.825,71.61
X$15418 1230 VIA_via1_7
* cell instance $15419 r0 *1 88.825,71.61
X$15419 1230 VIA_via2_5
* cell instance $15420 r0 *1 88.825,54.67
X$15420 1230 VIA_via2_5
* cell instance $15421 r0 *1 89.585,54.67
X$15421 1230 VIA_via2_5
* cell instance $15422 r0 *1 95.855,56.63
X$15422 1230 VIA_via2_5
* cell instance $15423 r0 *1 95.855,59.57
X$15423 1230 VIA_via2_5
* cell instance $15424 r0 *1 96.045,51.03
X$15424 1230 VIA_via2_5
* cell instance $15425 r0 *1 94.525,54.53
X$15425 1230 VIA_via2_5
* cell instance $15426 r0 *1 93.385,54.53
X$15426 1230 VIA_via2_5
* cell instance $15427 r0 *1 86.545,71.61
X$15427 1230 VIA_via2_5
* cell instance $15428 r0 *1 95.095,71.61
X$15428 1230 VIA_via2_5
* cell instance $15429 r0 *1 86.545,73.57
X$15429 1230 VIA_via1_4
* cell instance $15430 r0 *1 95.095,65.17
X$15430 1230 VIA_via1_4
* cell instance $15431 r0 *1 96.045,65.17
X$15431 1230 VIA_via1_4
* cell instance $15432 r0 *1 89.205,49.63
X$15432 1230 VIA_via1_4
* cell instance $15433 r0 *1 94.525,56.77
X$15433 1230 VIA_via1_4
* cell instance $15434 r0 *1 94.525,56.63
X$15434 1230 VIA_via2_5
* cell instance $15435 r0 *1 94.905,51.17
X$15435 1230 VIA_via1_4
* cell instance $15436 r0 *1 94.905,51.03
X$15436 1230 VIA_via2_5
* cell instance $15437 r0 *1 95.015,51.03
X$15437 1230 VIA_via3_2
* cell instance $15438 r0 *1 96.235,49.63
X$15438 1230 VIA_via1_4
* cell instance $15439 r0 *1 93.385,53.97
X$15439 1230 VIA_via1_4
* cell instance $15440 r0 *1 89.395,55.23
X$15440 1230 VIA_via1_4
* cell instance $15441 r0 *1 95.095,59.57
X$15441 1230 VIA_via1_4
* cell instance $15442 r0 *1 95.095,59.57
X$15442 1230 VIA_via2_5
* cell instance $15443 r0 *1 95.015,54.53
X$15443 1230 VIA_via3_2
* cell instance $15444 r0 *1 96.235,49.35
X$15444 1231 VIA_via1_4
* cell instance $15445 r0 *1 96.805,51.17
X$15445 1231 VIA_via1_4
* cell instance $15446 r0 *1 19.095,49.91
X$15446 1232 VIA_via1_7
* cell instance $15447 r0 *1 3.325,49.35
X$15447 1232 VIA_via2_5
* cell instance $15448 r0 *1 3.325,49.63
X$15448 1232 VIA_via1_4
* cell instance $15449 r0 *1 4.015,49.35
X$15449 1232 VIA_via4_0
* cell instance $15450 r0 *1 4.015,49.35
X$15450 1232 VIA_via3_2
* cell instance $15451 r0 *1 19.135,49.35
X$15451 1232 VIA_via3_2
* cell instance $15452 r0 *1 19.095,49.35
X$15452 1232 VIA_via2_5
* cell instance $15453 r0 *1 19.135,49.35
X$15453 1232 VIA_via4_0
* cell instance $15454 r0 *1 40.945,49.91
X$15454 1233 VIA_via1_7
* cell instance $15455 r0 *1 40.945,49.91
X$15455 1233 VIA_via2_5
* cell instance $15456 r0 *1 3.895,49.63
X$15456 1233 VIA_via1_4
* cell instance $15457 r0 *1 3.895,49.63
X$15457 1233 VIA_via2_5
* cell instance $15458 r0 *1 4.015,49.63
X$15458 1233 VIA_via3_2
* cell instance $15459 r0 *1 4.015,49.91
X$15459 1233 VIA_via4_0
* cell instance $15460 r0 *1 40.695,49.91
X$15460 1233 VIA_via3_2
* cell instance $15461 r0 *1 40.695,49.91
X$15461 1233 VIA_via4_0
* cell instance $15462 r0 *1 95.855,48.65
X$15462 1234 VIA_via2_5
* cell instance $15463 r0 *1 96.995,48.65
X$15463 1234 VIA_via1_4
* cell instance $15464 r0 *1 96.995,48.65
X$15464 1234 VIA_via2_5
* cell instance $15465 r0 *1 94.525,49.63
X$15465 1234 VIA_via1_4
* cell instance $15466 r0 *1 94.715,49.63
X$15466 1234 VIA_via1_4
* cell instance $15467 r0 *1 94.715,49.63
X$15467 1234 VIA_via2_5
* cell instance $15468 r0 *1 95.855,49.63
X$15468 1234 VIA_via1_4
* cell instance $15469 r0 *1 95.855,49.63
X$15469 1234 VIA_via2_5
* cell instance $15470 r0 *1 95.095,49.21
X$15470 1235 VIA_via1_7
* cell instance $15471 r0 *1 95.095,48.37
X$15471 1235 VIA_via2_5
* cell instance $15472 r0 *1 93.765,48.37
X$15472 1235 VIA_via1_4
* cell instance $15473 r0 *1 93.765,48.37
X$15473 1235 VIA_via2_5
* cell instance $15474 r0 *1 16.245,48.37
X$15474 1236 VIA_via1_4
* cell instance $15475 r0 *1 15.485,48.37
X$15475 1236 VIA_via1_4
* cell instance $15476 r0 *1 18.905,47.39
X$15476 1237 VIA_via1_7
* cell instance $15477 r0 *1 18.905,49.63
X$15477 1237 VIA_via1_4
* cell instance $15478 r0 *1 19.665,49.63
X$15478 1238 VIA_via1_4
* cell instance $15479 r0 *1 19.665,49.63
X$15479 1238 VIA_via2_5
* cell instance $15480 r0 *1 16.815,49.63
X$15480 1238 VIA_via1_4
* cell instance $15481 r0 *1 16.815,49.63
X$15481 1238 VIA_via2_5
* cell instance $15482 r0 *1 82.175,65.59
X$15482 1239 VIA_via1_7
* cell instance $15483 r0 *1 88.445,49.07
X$15483 1239 VIA_via2_5
* cell instance $15484 r0 *1 93.385,49.07
X$15484 1239 VIA_via2_5
* cell instance $15485 r0 *1 88.065,57.47
X$15485 1239 VIA_via2_5
* cell instance $15486 r0 *1 94.335,60.97
X$15486 1239 VIA_via2_5
* cell instance $15487 r0 *1 92.815,60.97
X$15487 1239 VIA_via2_5
* cell instance $15488 r0 *1 94.335,59.57
X$15488 1239 VIA_via2_5
* cell instance $15489 r0 *1 94.145,49.91
X$15489 1239 VIA_via2_5
* cell instance $15490 r0 *1 95.095,49.91
X$15490 1239 VIA_via2_5
* cell instance $15491 r0 *1 93.385,49.91
X$15491 1239 VIA_via2_5
* cell instance $15492 r0 *1 93.765,53.83
X$15492 1239 VIA_via2_5
* cell instance $15493 r0 *1 82.175,67.69
X$15493 1239 VIA_via2_5
* cell instance $15494 r0 *1 80.465,67.69
X$15494 1239 VIA_via2_5
* cell instance $15495 r0 *1 92.625,65.03
X$15495 1239 VIA_via2_5
* cell instance $15496 r0 *1 94.335,65.03
X$15496 1239 VIA_via2_5
* cell instance $15497 r0 *1 92.625,68.39
X$15497 1239 VIA_via2_5
* cell instance $15498 r0 *1 92.245,67.69
X$15498 1239 VIA_via2_5
* cell instance $15499 r0 *1 92.245,68.39
X$15499 1239 VIA_via2_5
* cell instance $15500 r0 *1 88.445,48.37
X$15500 1239 VIA_via1_4
* cell instance $15501 r0 *1 92.245,67.97
X$15501 1239 VIA_via1_4
* cell instance $15502 r0 *1 94.525,65.17
X$15502 1239 VIA_via1_4
* cell instance $15503 r0 *1 80.465,67.97
X$15503 1239 VIA_via1_4
* cell instance $15504 r0 *1 88.065,56.77
X$15504 1239 VIA_via1_4
* cell instance $15505 r0 *1 94.145,51.17
X$15505 1239 VIA_via1_4
* cell instance $15506 r0 *1 95.095,49.63
X$15506 1239 VIA_via1_4
* cell instance $15507 r0 *1 92.815,53.97
X$15507 1239 VIA_via1_4
* cell instance $15508 r0 *1 92.815,53.83
X$15508 1239 VIA_via2_5
* cell instance $15509 r0 *1 92.775,53.83
X$15509 1239 VIA_via3_2
* cell instance $15510 r0 *1 94.525,59.57
X$15510 1239 VIA_via1_4
* cell instance $15511 r0 *1 93.005,60.83
X$15511 1239 VIA_via1_4
* cell instance $15512 r0 *1 92.775,57.47
X$15512 1239 VIA_via3_2
* cell instance $15513 r0 *1 94.175,57.47
X$15513 1239 VIA_via3_2
* cell instance $15514 r0 *1 94.175,59.57
X$15514 1239 VIA_via3_2
* cell instance $15515 r0 *1 79.325,94.15
X$15515 1240 VIA_via2_5
* cell instance $15516 r0 *1 57.095,50.89
X$15516 1240 VIA_via2_5
* cell instance $15517 r0 *1 86.165,51.31
X$15517 1240 VIA_via2_5
* cell instance $15518 r0 *1 90.345,50.61
X$15518 1240 VIA_via2_5
* cell instance $15519 r0 *1 90.725,50.61
X$15519 1240 VIA_via2_5
* cell instance $15520 r0 *1 86.355,51.31
X$15520 1240 VIA_via2_5
* cell instance $15521 r0 *1 86.165,50.61
X$15521 1240 VIA_via2_5
* cell instance $15522 r0 *1 83.695,51.45
X$15522 1240 VIA_via2_5
* cell instance $15523 r0 *1 83.885,50.61
X$15523 1240 VIA_via2_5
* cell instance $15524 r0 *1 65.835,92.89
X$15524 1240 VIA_via2_5
* cell instance $15525 r0 *1 92.055,49.63
X$15525 1240 VIA_via2_5
* cell instance $15526 r0 *1 79.325,92.89
X$15526 1240 VIA_via2_5
* cell instance $15527 r0 *1 78.375,94.43
X$15527 1240 VIA_via1_4
* cell instance $15528 r0 *1 78.375,94.43
X$15528 1240 VIA_via2_5
* cell instance $15529 r0 *1 85.785,48.37
X$15529 1240 VIA_via1_4
* cell instance $15530 r0 *1 92.055,48.37
X$15530 1240 VIA_via1_4
* cell instance $15531 r0 *1 82.175,78.05
X$15531 1240 VIA_via1_4
* cell instance $15532 r0 *1 82.175,78.05
X$15532 1240 VIA_via2_5
* cell instance $15533 r0 *1 65.835,93.17
X$15533 1240 VIA_via1_4
* cell instance $15534 r0 *1 57.095,52.43
X$15534 1240 VIA_via1_4
* cell instance $15535 r0 *1 91.295,52.43
X$15535 1240 VIA_via1_4
* cell instance $15536 r0 *1 86.355,53.97
X$15536 1240 VIA_via1_4
* cell instance $15537 r0 *1 90.345,49.63
X$15537 1240 VIA_via1_4
* cell instance $15538 r0 *1 90.345,49.63
X$15538 1240 VIA_via2_5
* cell instance $15539 r0 *1 83.885,51.17
X$15539 1240 VIA_via1_4
* cell instance $15540 r0 *1 83.885,51.31
X$15540 1240 VIA_via2_5
* cell instance $15541 r0 *1 83.695,52.43
X$15541 1240 VIA_via1_4
* cell instance $15542 r0 *1 83.815,94.15
X$15542 1240 VIA_via3_2
* cell instance $15543 r0 *1 83.815,78.05
X$15543 1240 VIA_via3_2
* cell instance $15544 r0 *1 83.815,52.15
X$15544 1240 VIA_via3_2
* cell instance $15545 r0 *1 83.695,52.15
X$15545 1240 VIA_via2_5
* cell instance $15546 r0 *1 73.055,65.59
X$15546 1241 VIA_via1_7
* cell instance $15547 r0 *1 73.055,65.59
X$15547 1241 VIA_via2_5
* cell instance $15548 r0 *1 68.495,65.45
X$15548 1241 VIA_via2_5
* cell instance $15549 r0 *1 90.155,49.91
X$15549 1241 VIA_via2_5
* cell instance $15550 r0 *1 85.785,54.25
X$15550 1241 VIA_via2_5
* cell instance $15551 r0 *1 85.595,49.91
X$15551 1241 VIA_via2_5
* cell instance $15552 r0 *1 92.245,57.33
X$15552 1241 VIA_via2_5
* cell instance $15553 r0 *1 92.215,57.33
X$15553 1241 VIA_via3_2
* cell instance $15554 r0 *1 91.865,49.35
X$15554 1241 VIA_via2_5
* cell instance $15555 r0 *1 92.245,54.53
X$15555 1241 VIA_via2_5
* cell instance $15556 r0 *1 89.775,64.33
X$15556 1241 VIA_via2_5
* cell instance $15557 r0 *1 89.775,65.59
X$15557 1241 VIA_via2_5
* cell instance $15558 r0 *1 92.245,64.33
X$15558 1241 VIA_via2_5
* cell instance $15559 r0 *1 92.245,63.35
X$15559 1241 VIA_via2_5
* cell instance $15560 r0 *1 92.215,63.35
X$15560 1241 VIA_via3_2
* cell instance $15561 r0 *1 68.495,67.97
X$15561 1241 VIA_via1_4
* cell instance $15562 r0 *1 85.595,48.37
X$15562 1241 VIA_via1_4
* cell instance $15563 r0 *1 91.865,48.37
X$15563 1241 VIA_via1_4
* cell instance $15564 r0 *1 89.775,65.17
X$15564 1241 VIA_via1_4
* cell instance $15565 r0 *1 92.245,63.63
X$15565 1241 VIA_via1_4
* cell instance $15566 r0 *1 90.155,49.63
X$15566 1241 VIA_via1_4
* cell instance $15567 r0 *1 91.105,52.43
X$15567 1241 VIA_via1_4
* cell instance $15568 r0 *1 91.105,52.57
X$15568 1241 VIA_via2_5
* cell instance $15569 r0 *1 85.785,53.97
X$15569 1241 VIA_via1_4
* cell instance $15570 r0 *1 92.245,56.77
X$15570 1241 VIA_via1_4
* cell instance $15571 r0 *1 92.245,56.63
X$15571 1241 VIA_via2_5
* cell instance $15572 r0 *1 90.915,56.77
X$15572 1241 VIA_via1_4
* cell instance $15573 r0 *1 90.915,56.77
X$15573 1241 VIA_via2_5
* cell instance $15574 r0 *1 91.655,49.35
X$15574 1241 VIA_via3_2
* cell instance $15575 r0 *1 91.655,49.91
X$15575 1241 VIA_via3_2
* cell instance $15576 r0 *1 91.655,54.53
X$15576 1241 VIA_via3_2
* cell instance $15577 r0 *1 91.655,52.57
X$15577 1241 VIA_via3_2
* cell instance $15578 r0 *1 23.275,49.63
X$15578 1242 VIA_via1_4
* cell instance $15579 r0 *1 23.275,49.63
X$15579 1242 VIA_via2_5
* cell instance $15580 r0 *1 22.705,49.63
X$15580 1242 VIA_via1_4
* cell instance $15581 r0 *1 22.705,49.63
X$15581 1242 VIA_via2_5
* cell instance $15582 r0 *1 28.025,50.61
X$15582 1243 VIA_via1_7
* cell instance $15583 r0 *1 28.025,49.63
X$15583 1243 VIA_via2_5
* cell instance $15584 r0 *1 24.985,49.63
X$15584 1243 VIA_via1_4
* cell instance $15585 r0 *1 24.985,49.63
X$15585 1243 VIA_via2_5
* cell instance $15586 r0 *1 27.455,48.37
X$15586 1244 VIA_via1_4
* cell instance $15587 r0 *1 27.455,48.37
X$15587 1244 VIA_via2_5
* cell instance $15588 r0 *1 28.215,48.37
X$15588 1244 VIA_via1_4
* cell instance $15589 r0 *1 28.215,48.37
X$15589 1244 VIA_via2_5
* cell instance $15590 r0 *1 88.255,48.37
X$15590 1245 VIA_via1_4
* cell instance $15591 r0 *1 88.255,48.37
X$15591 1245 VIA_via2_5
* cell instance $15592 r0 *1 87.305,48.37
X$15592 1245 VIA_via1_4
* cell instance $15593 r0 *1 87.305,48.37
X$15593 1245 VIA_via2_5
* cell instance $15594 r0 *1 31.635,49.63
X$15594 1246 VIA_via2_5
* cell instance $15595 r0 *1 30.305,49.63
X$15595 1246 VIA_via1_4
* cell instance $15596 r0 *1 30.305,49.63
X$15596 1246 VIA_via2_5
* cell instance $15597 r0 *1 31.635,48.51
X$15597 1246 VIA_via1_4
* cell instance $15598 r0 *1 86.355,49.07
X$15598 1247 VIA_via2_5
* cell instance $15599 r0 *1 87.115,49.07
X$15599 1247 VIA_via2_5
* cell instance $15600 r0 *1 87.115,48.51
X$15600 1247 VIA_via1_4
* cell instance $15601 r0 *1 86.355,49.63
X$15601 1247 VIA_via1_4
* cell instance $15602 r0 *1 34.865,49.63
X$15602 1248 VIA_via1_4
* cell instance $15603 r0 *1 34.865,49.49
X$15603 1248 VIA_via2_5
* cell instance $15604 r0 *1 36.385,49.49
X$15604 1248 VIA_via1_4
* cell instance $15605 r0 *1 36.385,49.49
X$15605 1248 VIA_via2_5
* cell instance $15606 r0 *1 33.345,50.61
X$15606 1249 VIA_via1_7
* cell instance $15607 r0 *1 33.345,49.63
X$15607 1249 VIA_via2_5
* cell instance $15608 r0 *1 34.675,49.63
X$15608 1249 VIA_via1_4
* cell instance $15609 r0 *1 34.675,49.63
X$15609 1249 VIA_via2_5
* cell instance $15610 r0 *1 81.985,49.49
X$15610 1250 VIA_via2_5
* cell instance $15611 r0 *1 81.985,48.23
X$15611 1250 VIA_via1_4
* cell instance $15612 r0 *1 81.035,49.63
X$15612 1250 VIA_via1_4
* cell instance $15613 r0 *1 81.035,49.49
X$15613 1250 VIA_via2_5
* cell instance $15614 r0 *1 37.145,50.61
X$15614 1251 VIA_via1_7
* cell instance $15615 r0 *1 37.145,49.63
X$15615 1251 VIA_via2_5
* cell instance $15616 r0 *1 35.435,49.7
X$15616 1251 VIA_via1_4
* cell instance $15617 r0 *1 35.435,49.63
X$15617 1251 VIA_via2_5
* cell instance $15618 r0 *1 76.475,48.37
X$15618 1252 VIA_via1_4
* cell instance $15619 r0 *1 76.475,48.37
X$15619 1252 VIA_via2_5
* cell instance $15620 r0 *1 74.955,48.37
X$15620 1252 VIA_via1_4
* cell instance $15621 r0 *1 74.955,48.37
X$15621 1252 VIA_via2_5
* cell instance $15622 r0 *1 44.365,49.91
X$15622 1253 VIA_via1_7
* cell instance $15623 r0 *1 44.365,49.63
X$15623 1253 VIA_via2_5
* cell instance $15624 r0 *1 41.135,49.63
X$15624 1253 VIA_via1_4
* cell instance $15625 r0 *1 41.135,49.63
X$15625 1253 VIA_via2_5
* cell instance $15626 r0 *1 53.295,49.35
X$15626 1254 VIA_via2_5
* cell instance $15627 r0 *1 53.295,48.65
X$15627 1254 VIA_via2_5
* cell instance $15628 r0 *1 49.875,48.65
X$15628 1254 VIA_via2_5
* cell instance $15629 r0 *1 53.295,48.37
X$15629 1254 VIA_via1_4
* cell instance $15630 r0 *1 49.875,48.37
X$15630 1254 VIA_via1_4
* cell instance $15631 r0 *1 53.865,49.35
X$15631 1254 VIA_via1_4
* cell instance $15632 r0 *1 53.865,49.35
X$15632 1254 VIA_via2_5
* cell instance $15633 r0 *1 54.815,48.37
X$15633 1255 VIA_via1_4
* cell instance $15634 r0 *1 54.815,48.37
X$15634 1255 VIA_via2_5
* cell instance $15635 r0 *1 53.675,48.37
X$15635 1255 VIA_via1_4
* cell instance $15636 r0 *1 53.675,48.37
X$15636 1255 VIA_via2_5
* cell instance $15637 r0 *1 57.665,48.79
X$15637 1256 VIA_via2_5
* cell instance $15638 r0 *1 59.185,48.79
X$15638 1256 VIA_via2_5
* cell instance $15639 r0 *1 59.185,48.23
X$15639 1256 VIA_via1_4
* cell instance $15640 r0 *1 57.665,49.63
X$15640 1256 VIA_via1_4
* cell instance $15641 r0 *1 61.275,49.21
X$15641 1257 VIA_via1_7
* cell instance $15642 r0 *1 61.275,48.37
X$15642 1257 VIA_via1_4
* cell instance $15643 r0 *1 3.705,49.91
X$15643 1258 VIA_via1_4
* cell instance $15644 r0 *1 3.705,49.91
X$15644 1258 VIA_via2_5
* cell instance $15645 r0 *1 1.775,49.91
X$15645 1258 VIA_via3_2
* cell instance $15646 r0 *1 1.775,49.91
X$15646 1258 VIA_via4_0
* cell instance $15647 r0 *1 5.605,50.19
X$15647 1259 VIA_via1_7
* cell instance $15648 r0 *1 5.605,50.47
X$15648 1259 VIA_via2_5
* cell instance $15649 r0 *1 5.415,50.47
X$15649 1259 VIA_via4_0
* cell instance $15650 r0 *1 5.415,50.47
X$15650 1259 VIA_via3_2
* cell instance $15651 r0 *1 4.275,50.19
X$15651 1260 VIA_via1_7
* cell instance $15652 r0 *1 4.295,51.03
X$15652 1260 VIA_via3_2
* cell instance $15653 r0 *1 4.275,51.03
X$15653 1260 VIA_via2_5
* cell instance $15654 r0 *1 4.295,51.03
X$15654 1260 VIA_via4_0
* cell instance $15655 r0 *1 20.045,50.61
X$15655 1261 VIA_via1_7
* cell instance $15656 r0 *1 18.905,52.43
X$15656 1261 VIA_via1_4
* cell instance $15657 r0 *1 35.245,50.47
X$15657 1262 VIA_via2_5
* cell instance $15658 r0 *1 30.495,60.83
X$15658 1262 VIA_via2_5
* cell instance $15659 r0 *1 30.685,56.77
X$15659 1262 VIA_via2_5
* cell instance $15660 r0 *1 30.685,52.43
X$15660 1262 VIA_via2_5
* cell instance $15661 r0 *1 31.065,50.19
X$15661 1262 VIA_via2_5
* cell instance $15662 r0 *1 30.495,56.77
X$15662 1262 VIA_via2_5
* cell instance $15663 r0 *1 26.695,52.43
X$15663 1262 VIA_via2_5
* cell instance $15664 r0 *1 32.395,60.83
X$15664 1262 VIA_via2_5
* cell instance $15665 r0 *1 28.595,56.77
X$15665 1262 VIA_via1_4
* cell instance $15666 r0 *1 28.595,56.77
X$15666 1262 VIA_via2_5
* cell instance $15667 r0 *1 31.255,56.77
X$15667 1262 VIA_via1_4
* cell instance $15668 r0 *1 31.255,56.77
X$15668 1262 VIA_via2_5
* cell instance $15669 r0 *1 30.305,60.83
X$15669 1262 VIA_via1_4
* cell instance $15670 r0 *1 31.445,58.03
X$15670 1262 VIA_via1_4
* cell instance $15671 r0 *1 31.255,53.97
X$15671 1262 VIA_via1_4
* cell instance $15672 r0 *1 35.245,51.17
X$15672 1262 VIA_via1_4
* cell instance $15673 r0 *1 31.065,49.63
X$15673 1262 VIA_via1_4
* cell instance $15674 r0 *1 26.695,53.97
X$15674 1262 VIA_via1_4
* cell instance $15675 r0 *1 32.015,65.17
X$15675 1262 VIA_via1_4
* cell instance $15676 r0 *1 31.635,50.61
X$15676 1263 VIA_via1_7
* cell instance $15677 r0 *1 31.825,48.37
X$15677 1263 VIA_via1_4
* cell instance $15678 r0 *1 34.865,49.91
X$15678 1264 VIA_via1_7
* cell instance $15679 r0 *1 34.485,51.17
X$15679 1264 VIA_via1_4
* cell instance $15680 r0 *1 37.905,50.61
X$15680 1265 VIA_via1_7
* cell instance $15681 r0 *1 38.475,49.49
X$15681 1265 VIA_via1_4
* cell instance $15682 r0 *1 54.815,50.89
X$15682 1266 VIA_via1_4
* cell instance $15683 r0 *1 55.195,52.43
X$15683 1266 VIA_via1_4
* cell instance $15684 r0 *1 66.785,50.89
X$15684 1267 VIA_via1_4
* cell instance $15685 r0 *1 65.645,52.43
X$15685 1267 VIA_via1_4
* cell instance $15686 r0 *1 66.405,52.43
X$15686 1267 VIA_via1_4
* cell instance $15687 r0 *1 58.425,51.59
X$15687 1268 VIA_via2_5
* cell instance $15688 r0 *1 58.615,54.11
X$15688 1268 VIA_via2_5
* cell instance $15689 r0 *1 85.975,50.89
X$15689 1268 VIA_via2_5
* cell instance $15690 r0 *1 86.165,52.57
X$15690 1268 VIA_via2_5
* cell instance $15691 r0 *1 86.165,53.69
X$15691 1268 VIA_via2_5
* cell instance $15692 r0 *1 84.075,53.69
X$15692 1268 VIA_via2_5
* cell instance $15693 r0 *1 44.365,53.97
X$15693 1268 VIA_via1_4
* cell instance $15694 r0 *1 44.365,54.11
X$15694 1268 VIA_via2_5
* cell instance $15695 r0 *1 44.365,70.77
X$15695 1268 VIA_via1_4
* cell instance $15696 r0 *1 44.365,70.77
X$15696 1268 VIA_via2_5
* cell instance $15697 r0 *1 89.585,72.03
X$15697 1268 VIA_via1_4
* cell instance $15698 r0 *1 89.585,72.03
X$15698 1268 VIA_via2_5
* cell instance $15699 r0 *1 88.065,72.03
X$15699 1268 VIA_via1_4
* cell instance $15700 r0 *1 88.065,72.03
X$15700 1268 VIA_via2_5
* cell instance $15701 r0 *1 88.015,72.03
X$15701 1268 VIA_via3_2
* cell instance $15702 r0 *1 58.615,52.43
X$15702 1268 VIA_via1_4
* cell instance $15703 r0 *1 85.975,52.43
X$15703 1268 VIA_via1_4
* cell instance $15704 r0 *1 84.075,53.97
X$15704 1268 VIA_via1_4
* cell instance $15705 r0 *1 62.815,51.59
X$15705 1268 VIA_via3_2
* cell instance $15706 r0 *1 63.095,51.31
X$15706 1268 VIA_via3_2
* cell instance $15707 r0 *1 44.895,54.11
X$15707 1268 VIA_via3_2
* cell instance $15708 r0 *1 88.015,52.57
X$15708 1268 VIA_via3_2
* cell instance $15709 r0 *1 44.895,70.77
X$15709 1268 VIA_via3_2
* cell instance $15710 r0 *1 81.035,51.45
X$15710 1269 VIA_via2_5
* cell instance $15711 r0 *1 81.415,51.1
X$15711 1269 VIA_via1_4
* cell instance $15712 r0 *1 80.465,51.45
X$15712 1269 VIA_via1_4
* cell instance $15713 r0 *1 80.465,51.45
X$15713 1269 VIA_via2_5
* cell instance $15714 r0 *1 81.035,52.43
X$15714 1269 VIA_via1_4
* cell instance $15715 r0 *1 89.015,50.19
X$15715 1270 VIA_via1_7
* cell instance $15716 r0 *1 89.395,51.17
X$15716 1270 VIA_via1_4
* cell instance $15717 r0 *1 91.865,50.61
X$15717 1271 VIA_via1_7
* cell instance $15718 r0 *1 91.675,49.63
X$15718 1271 VIA_via1_4
* cell instance $15719 r0 *1 93.765,51.17
X$15719 1272 VIA_via1_4
* cell instance $15720 r0 *1 93.765,51.17
X$15720 1272 VIA_via2_5
* cell instance $15721 r0 *1 93.955,50.05
X$15721 1272 VIA_via1_4
* cell instance $15722 r0 *1 94.525,51.17
X$15722 1272 VIA_via1_4
* cell instance $15723 r0 *1 94.525,51.17
X$15723 1272 VIA_via2_5
* cell instance $15724 r0 *1 93.385,51.17
X$15724 1272 VIA_via1_4
* cell instance $15725 r0 *1 90.155,51.03
X$15725 1273 VIA_via1_4
* cell instance $15726 r0 *1 90.155,51.03
X$15726 1273 VIA_via2_5
* cell instance $15727 r0 *1 95.665,51.17
X$15727 1273 VIA_via1_4
* cell instance $15728 r0 *1 95.665,51.17
X$15728 1273 VIA_via2_5
* cell instance $15729 r0 *1 96.805,50.19
X$15729 1274 VIA_via1_7
* cell instance $15730 r0 *1 96.805,50.19
X$15730 1274 VIA_via2_5
* cell instance $15731 r0 *1 96.975,51.03
X$15731 1274 VIA_via4_0
* cell instance $15732 r0 *1 96.975,50.19
X$15732 1274 VIA_via3_2
* cell instance $15733 r0 *1 96.235,50.61
X$15733 1275 VIA_via1_7
* cell instance $15734 r0 *1 96.235,50.47
X$15734 1275 VIA_via2_5
* cell instance $15735 r0 *1 97.255,50.47
X$15735 1275 VIA_via3_2
* cell instance $15736 r0 *1 97.255,50.47
X$15736 1275 VIA_via4_0
* cell instance $15737 r0 *1 96.995,52.71
X$15737 1276 VIA_via1_4
* cell instance $15738 r0 *1 96.995,52.71
X$15738 1276 VIA_via2_5
* cell instance $15739 r0 *1 97.815,49.91
X$15739 1276 VIA_via4_0
* cell instance $15740 r0 *1 97.815,52.71
X$15740 1276 VIA_via3_2
* cell instance $15741 r0 *1 92.435,50.75
X$15741 1277 VIA_via1_7
* cell instance $15742 r0 *1 92.435,50.61
X$15742 1277 VIA_via2_5
* cell instance $15743 r0 *1 96.995,50.61
X$15743 1277 VIA_via2_5
* cell instance $15744 r0 *1 96.995,51.17
X$15744 1277 VIA_via1_4
* cell instance $15745 r0 *1 84.645,50.61
X$15745 1278 VIA_via1_7
* cell instance $15746 r0 *1 84.645,49.77
X$15746 1278 VIA_via2_5
* cell instance $15747 r0 *1 96.425,49.63
X$15747 1278 VIA_via1_4
* cell instance $15748 r0 *1 96.425,49.77
X$15748 1278 VIA_via2_5
* cell instance $15749 r0 *1 90.725,50.19
X$15749 1279 VIA_via1_7
* cell instance $15750 r0 *1 90.725,50.19
X$15750 1279 VIA_via2_5
* cell instance $15751 r0 *1 91.295,50.19
X$15751 1279 VIA_via2_5
* cell instance $15752 r0 *1 91.295,51.17
X$15752 1279 VIA_via1_4
* cell instance $15753 r0 *1 25.935,49.91
X$15753 1280 VIA_via1_7
* cell instance $15754 r0 *1 25.935,49.91
X$15754 1280 VIA_via2_5
* cell instance $15755 r0 *1 24.415,49.91
X$15755 1280 VIA_via2_5
* cell instance $15756 r0 *1 24.415,49.63
X$15756 1280 VIA_via1_4
* cell instance $15757 r0 *1 27.455,50.61
X$15757 1281 VIA_via1_7
* cell instance $15758 r0 *1 27.455,50.61
X$15758 1281 VIA_via2_5
* cell instance $15759 r0 *1 24.225,50.61
X$15759 1281 VIA_via2_5
* cell instance $15760 r0 *1 24.225,49.63
X$15760 1281 VIA_via1_4
* cell instance $15761 r0 *1 34.295,49.77
X$15761 1282 VIA_via1_4
* cell instance $15762 r0 *1 34.295,49.77
X$15762 1282 VIA_via2_5
* cell instance $15763 r0 *1 27.455,49.63
X$15763 1282 VIA_via1_4
* cell instance $15764 r0 *1 27.455,49.77
X$15764 1282 VIA_via2_5
* cell instance $15765 r0 *1 81.605,50.05
X$15765 1283 VIA_via2_5
* cell instance $15766 r0 *1 81.605,48.37
X$15766 1283 VIA_via1_4
* cell instance $15767 r0 *1 83.315,50.05
X$15767 1283 VIA_via1_4
* cell instance $15768 r0 *1 83.315,50.05
X$15768 1283 VIA_via2_5
* cell instance $15769 r0 *1 81.605,52.43
X$15769 1283 VIA_via1_4
* cell instance $15770 r0 *1 68.115,50.61
X$15770 1284 VIA_via1_7
* cell instance $15771 r0 *1 68.115,50.61
X$15771 1284 VIA_via2_5
* cell instance $15772 r0 *1 65.455,50.61
X$15772 1284 VIA_via2_5
* cell instance $15773 r0 *1 65.455,49.63
X$15773 1284 VIA_via1_4
* cell instance $15774 r0 *1 37.905,49.91
X$15774 1285 VIA_via1_7
* cell instance $15775 r0 *1 37.905,49.91
X$15775 1285 VIA_via2_5
* cell instance $15776 r0 *1 37.895,49.91
X$15776 1285 VIA_via3_2
* cell instance $15777 r0 *1 2.185,52.43
X$15777 1285 VIA_via1_4
* cell instance $15778 r0 *1 2.185,52.43
X$15778 1285 VIA_via2_5
* cell instance $15779 r0 *1 37.895,52.43
X$15779 1285 VIA_via4_0
* cell instance $15780 r0 *1 2.615,52.43
X$15780 1285 VIA_via4_0
* cell instance $15781 r0 *1 2.615,52.43
X$15781 1285 VIA_via3_2
* cell instance $15782 r0 *1 39.235,50.61
X$15782 1286 VIA_via1_7
* cell instance $15783 r0 *1 39.235,50.61
X$15783 1286 VIA_via2_5
* cell instance $15784 r0 *1 37.525,50.61
X$15784 1286 VIA_via2_5
* cell instance $15785 r0 *1 37.525,49.63
X$15785 1286 VIA_via1_4
* cell instance $15786 r0 *1 38.475,50.61
X$15786 1287 VIA_via1_7
* cell instance $15787 r0 *1 38.475,50.47
X$15787 1287 VIA_via2_5
* cell instance $15788 r0 *1 42.085,50.47
X$15788 1287 VIA_via2_5
* cell instance $15789 r0 *1 42.085,49.49
X$15789 1287 VIA_via1_4
* cell instance $15790 r0 *1 60.515,50.47
X$15790 1288 VIA_via2_5
* cell instance $15791 r0 *1 58.615,50.47
X$15791 1288 VIA_via2_5
* cell instance $15792 r0 *1 60.515,48.23
X$15792 1288 VIA_via1_4
* cell instance $15793 r0 *1 58.615,51.17
X$15793 1288 VIA_via1_4
* cell instance $15794 r0 *1 37.525,88.97
X$15794 1289 VIA_via1_7
* cell instance $15795 r0 *1 37.525,88.97
X$15795 1289 VIA_via2_5
* cell instance $15796 r0 *1 28.215,88.97
X$15796 1289 VIA_via1_7
* cell instance $15797 r0 *1 28.215,89.11
X$15797 1289 VIA_via2_5
* cell instance $15798 r0 *1 12.445,53.83
X$15798 1289 VIA_via1_7
* cell instance $15799 r0 *1 11.495,89.25
X$15799 1289 VIA_via2_5
* cell instance $15800 r0 *1 11.495,88.41
X$15800 1289 VIA_via2_5
* cell instance $15801 r0 *1 10.545,88.41
X$15801 1289 VIA_via2_5
* cell instance $15802 r0 *1 10.735,71.47
X$15802 1289 VIA_via2_5
* cell instance $15803 r0 *1 21.185,89.11
X$15803 1289 VIA_via2_5
* cell instance $15804 r0 *1 13.205,65.31
X$15804 1289 VIA_via2_5
* cell instance $15805 r0 *1 45.315,88.27
X$15805 1289 VIA_via2_5
* cell instance $15806 r0 *1 45.315,90.23
X$15806 1289 VIA_via2_5
* cell instance $15807 r0 *1 37.525,88.27
X$15807 1289 VIA_via2_5
* cell instance $15808 r0 *1 12.825,54.39
X$15808 1289 VIA_via2_5
* cell instance $15809 r0 *1 48.355,56.77
X$15809 1289 VIA_via1_4
* cell instance $15810 r0 *1 48.355,56.91
X$15810 1289 VIA_via2_5
* cell instance $15811 r0 *1 21.185,87.57
X$15811 1289 VIA_via1_4
* cell instance $15812 r0 *1 45.695,90.37
X$15812 1289 VIA_via1_4
* cell instance $15813 r0 *1 45.695,90.23
X$15813 1289 VIA_via2_5
* cell instance $15814 r0 *1 48.735,86.03
X$15814 1289 VIA_via1_4
* cell instance $15815 r0 *1 48.735,86.03
X$15815 1289 VIA_via2_5
* cell instance $15816 r0 *1 47.405,50.75
X$15816 1289 VIA_via1_4
* cell instance $15817 r0 *1 47.415,50.75
X$15817 1289 VIA_via3_2
* cell instance $15818 r0 *1 47.405,50.75
X$15818 1289 VIA_via2_5
* cell instance $15819 r0 *1 13.965,65.17
X$15819 1289 VIA_via1_4
* cell instance $15820 r0 *1 10.735,72.03
X$15820 1289 VIA_via1_4
* cell instance $15821 r0 *1 10.545,88.83
X$15821 1289 VIA_via1_4
* cell instance $15822 r0 *1 47.415,54.11
X$15822 1289 VIA_via4_0
* cell instance $15823 r0 *1 49.095,54.11
X$15823 1289 VIA_via4_0
* cell instance $15824 r0 *1 13.815,65.31
X$15824 1289 VIA_via3_2
* cell instance $15825 r0 *1 13.775,65.31
X$15825 1289 VIA_via2_5
* cell instance $15826 r0 *1 13.535,54.39
X$15826 1289 VIA_via3_2
* cell instance $15827 r0 *1 13.395,54.39
X$15827 1289 VIA_via2_5
* cell instance $15828 r0 *1 13.535,54.39
X$15828 1289 VIA_via4_0
* cell instance $15829 r0 *1 13.815,71.47
X$15829 1289 VIA_via3_2
* cell instance $15830 r0 *1 49.095,90.23
X$15830 1289 VIA_via3_2
* cell instance $15831 r0 *1 49.095,56.91
X$15831 1289 VIA_via3_2
* cell instance $15832 r0 *1 49.095,86.03
X$15832 1289 VIA_via3_2
* cell instance $15833 r0 *1 2.565,52.01
X$15833 1290 VIA_via1_7
* cell instance $15834 r0 *1 2.565,51.59
X$15834 1290 VIA_via2_5
* cell instance $15835 r0 *1 0.375,51.59
X$15835 1290 VIA_via4_0
* cell instance $15836 r0 *1 0.375,51.59
X$15836 1290 VIA_via3_2
* cell instance $15837 r0 *1 4.655,53.41
X$15837 1291 VIA_via1_7
* cell instance $15838 r0 *1 4.655,53.41
X$15838 1291 VIA_via2_5
* cell instance $15839 r0 *1 3.515,53.41
X$15839 1291 VIA_via2_5
* cell instance $15840 r0 *1 2.945,51.17
X$15840 1291 VIA_via1_4
* cell instance $15841 r0 *1 3.515,58.87
X$15841 1292 VIA_via2_5
* cell instance $15842 r0 *1 8.835,58.87
X$15842 1292 VIA_via2_5
* cell instance $15843 r0 *1 8.835,59.57
X$15843 1292 VIA_via2_5
* cell instance $15844 r0 *1 6.365,58.87
X$15844 1292 VIA_via2_5
* cell instance $15845 r0 *1 3.895,52.43
X$15845 1292 VIA_via2_5
* cell instance $15846 r0 *1 3.325,56.77
X$15846 1292 VIA_via1_4
* cell instance $15847 r0 *1 6.365,59.57
X$15847 1292 VIA_via1_4
* cell instance $15848 r0 *1 10.735,60.83
X$15848 1292 VIA_via1_4
* cell instance $15849 r0 *1 10.545,59.57
X$15849 1292 VIA_via1_4
* cell instance $15850 r0 *1 10.545,59.57
X$15850 1292 VIA_via2_5
* cell instance $15851 r0 *1 3.705,51.17
X$15851 1292 VIA_via1_4
* cell instance $15852 r0 *1 8.835,58.03
X$15852 1292 VIA_via1_4
* cell instance $15853 r0 *1 5.605,52.43
X$15853 1292 VIA_via1_4
* cell instance $15854 r0 *1 5.605,52.43
X$15854 1292 VIA_via2_5
* cell instance $15855 r0 *1 8.835,59.15
X$15855 1292 VIA_via1_4
* cell instance $15856 r0 *1 9.025,56.77
X$15856 1292 VIA_via1_4
* cell instance $15857 r0 *1 8.455,52.57
X$15857 1293 VIA_via1_4
* cell instance $15858 r0 *1 8.075,51.17
X$15858 1293 VIA_via1_4
* cell instance $15859 r0 *1 8.075,51.45
X$15859 1294 VIA_via2_5
* cell instance $15860 r0 *1 11.305,51.45
X$15860 1294 VIA_via2_5
* cell instance $15861 r0 *1 8.075,52.43
X$15861 1294 VIA_via1_4
* cell instance $15862 r0 *1 10.355,51.45
X$15862 1294 VIA_via1_4
* cell instance $15863 r0 *1 10.355,51.45
X$15863 1294 VIA_via2_5
* cell instance $15864 r0 *1 11.305,51.17
X$15864 1294 VIA_via1_4
* cell instance $15865 r0 *1 12.065,51.59
X$15865 1295 VIA_via1_7
* cell instance $15866 r0 *1 12.445,55.23
X$15866 1295 VIA_via1_4
* cell instance $15867 r0 *1 17.765,53.41
X$15867 1296 VIA_via1_7
* cell instance $15868 r0 *1 18.335,51.17
X$15868 1296 VIA_via1_4
* cell instance $15869 r0 *1 22.325,52.43
X$15869 1297 VIA_via1_4
* cell instance $15870 r0 *1 22.135,51.31
X$15870 1297 VIA_via1_4
* cell instance $15871 r0 *1 47.595,51.31
X$15871 1298 VIA_via2_5
* cell instance $15872 r0 *1 44.175,51.73
X$15872 1298 VIA_via2_5
* cell instance $15873 r0 *1 44.175,59.57
X$15873 1298 VIA_via1_4
* cell instance $15874 r0 *1 38.285,51.17
X$15874 1298 VIA_via1_4
* cell instance $15875 r0 *1 38.285,51.31
X$15875 1298 VIA_via2_5
* cell instance $15876 r0 *1 42.465,51.17
X$15876 1298 VIA_via1_4
* cell instance $15877 r0 *1 42.465,51.31
X$15877 1298 VIA_via2_5
* cell instance $15878 r0 *1 47.595,52.15
X$15878 1298 VIA_via1_4
* cell instance $15879 r0 *1 52.535,53.41
X$15879 1299 VIA_via1_7
* cell instance $15880 r0 *1 52.535,51.17
X$15880 1299 VIA_via2_5
* cell instance $15881 r0 *1 41.895,51.17
X$15881 1299 VIA_via2_5
* cell instance $15882 r0 *1 41.895,56.77
X$15882 1299 VIA_via1_4
* cell instance $15883 r0 *1 45.315,51.17
X$15883 1299 VIA_via1_4
* cell instance $15884 r0 *1 45.315,51.17
X$15884 1299 VIA_via2_5
* cell instance $15885 r0 *1 43.985,51.17
X$15885 1299 VIA_via1_4
* cell instance $15886 r0 *1 43.985,51.17
X$15886 1299 VIA_via2_5
* cell instance $15887 r0 *1 51.395,51.17
X$15887 1299 VIA_via1_4
* cell instance $15888 r0 *1 51.395,51.17
X$15888 1299 VIA_via2_5
* cell instance $15889 r0 *1 77.615,86.31
X$15889 1300 VIA_via2_5
* cell instance $15890 r0 *1 78.375,86.31
X$15890 1300 VIA_via2_5
* cell instance $15891 r0 *1 79.515,88.13
X$15891 1300 VIA_via2_5
* cell instance $15892 r0 *1 70.585,57.05
X$15892 1300 VIA_via2_5
* cell instance $15893 r0 *1 54.625,57.05
X$15893 1300 VIA_via2_5
* cell instance $15894 r0 *1 84.075,88.13
X$15894 1300 VIA_via2_5
* cell instance $15895 r0 *1 71.345,76.09
X$15895 1300 VIA_via2_5
* cell instance $15896 r0 *1 85.975,52.71
X$15896 1300 VIA_via2_5
* cell instance $15897 r0 *1 82.935,51.45
X$15897 1300 VIA_via2_5
* cell instance $15898 r0 *1 79.895,52.85
X$15898 1300 VIA_via2_5
* cell instance $15899 r0 *1 80.655,51.87
X$15899 1300 VIA_via2_5
* cell instance $15900 r0 *1 87.685,88.13
X$15900 1300 VIA_via2_5
* cell instance $15901 r0 *1 87.115,88.13
X$15901 1300 VIA_via2_5
* cell instance $15902 r0 *1 79.895,56.91
X$15902 1300 VIA_via2_5
* cell instance $15903 r0 *1 77.425,76.09
X$15903 1300 VIA_via2_5
* cell instance $15904 r0 *1 70.965,66.43
X$15904 1300 VIA_via1_4
* cell instance $15905 r0 *1 78.375,87.15
X$15905 1300 VIA_via1_4
* cell instance $15906 r0 *1 79.515,87.85
X$15906 1300 VIA_via1_4
* cell instance $15907 r0 *1 84.265,90.37
X$15907 1300 VIA_via1_4
* cell instance $15908 r0 *1 87.115,87.57
X$15908 1300 VIA_via1_4
* cell instance $15909 r0 *1 87.685,88.83
X$15909 1300 VIA_via1_4
* cell instance $15910 r0 *1 54.815,51.17
X$15910 1300 VIA_via1_4
* cell instance $15911 r0 *1 54.625,56.77
X$15911 1300 VIA_via1_4
* cell instance $15912 r0 *1 55.005,51.17
X$15912 1300 VIA_via1_4
* cell instance $15913 r0 *1 85.975,53.97
X$15913 1300 VIA_via1_4
* cell instance $15914 r0 *1 82.935,51.17
X$15914 1300 VIA_via1_4
* cell instance $15915 r0 *1 80.655,52.43
X$15915 1300 VIA_via1_4
* cell instance $15916 r0 *1 80.655,52.57
X$15916 1300 VIA_via2_5
* cell instance $15917 r0 *1 68.115,56.63
X$15917 1301 VIA_via2_5
* cell instance $15918 r0 *1 66.975,54.67
X$15918 1301 VIA_via2_5
* cell instance $15919 r0 *1 56.525,51.17
X$15919 1301 VIA_via2_5
* cell instance $15920 r0 *1 66.785,51.17
X$15920 1301 VIA_via2_5
* cell instance $15921 r0 *1 66.215,51.17
X$15921 1301 VIA_via2_5
* cell instance $15922 r0 *1 68.495,54.67
X$15922 1301 VIA_via2_5
* cell instance $15923 r0 *1 66.215,49.63
X$15923 1301 VIA_via1_4
* cell instance $15924 r0 *1 65.265,51.17
X$15924 1301 VIA_via1_4
* cell instance $15925 r0 *1 65.265,51.17
X$15925 1301 VIA_via2_5
* cell instance $15926 r0 *1 66.975,53.97
X$15926 1301 VIA_via1_4
* cell instance $15927 r0 *1 67.165,56.77
X$15927 1301 VIA_via1_4
* cell instance $15928 r0 *1 67.165,56.63
X$15928 1301 VIA_via2_5
* cell instance $15929 r0 *1 56.335,53.97
X$15929 1301 VIA_via1_4
* cell instance $15930 r0 *1 70.775,59.57
X$15930 1301 VIA_via1_4
* cell instance $15931 r0 *1 71.155,55.23
X$15931 1301 VIA_via1_4
* cell instance $15932 r0 *1 71.155,55.23
X$15932 1301 VIA_via2_5
* cell instance $15933 r0 *1 59.375,51.17
X$15933 1301 VIA_via1_4
* cell instance $15934 r0 *1 59.375,51.17
X$15934 1301 VIA_via2_5
* cell instance $15935 r0 *1 68.495,55.23
X$15935 1301 VIA_via1_4
* cell instance $15936 r0 *1 68.495,55.23
X$15936 1301 VIA_via2_5
* cell instance $15937 r0 *1 68.115,55.65
X$15937 1301 VIA_via1_4
* cell instance $15938 r0 *1 67.735,52.43
X$15938 1302 VIA_via2_5
* cell instance $15939 r0 *1 67.735,50.05
X$15939 1302 VIA_via1_4
* cell instance $15940 r0 *1 67.735,51.17
X$15940 1302 VIA_via1_4
* cell instance $15941 r0 *1 66.975,52.43
X$15941 1302 VIA_via1_4
* cell instance $15942 r0 *1 66.975,52.43
X$15942 1302 VIA_via2_5
* cell instance $15943 r0 *1 83.885,53.41
X$15943 1303 VIA_via1_7
* cell instance $15944 r0 *1 84.645,51.17
X$15944 1303 VIA_via1_4
* cell instance $15945 r0 *1 90.155,59.01
X$15945 1304 VIA_via2_5
* cell instance $15946 r0 *1 90.345,51.45
X$15946 1304 VIA_via2_5
* cell instance $15947 r0 *1 85.785,52.01
X$15947 1304 VIA_via2_5
* cell instance $15948 r0 *1 93.385,58.87
X$15948 1304 VIA_via2_5
* cell instance $15949 r0 *1 94.335,51.45
X$15949 1304 VIA_via2_5
* cell instance $15950 r0 *1 92.625,51.45
X$15950 1304 VIA_via2_5
* cell instance $15951 r0 *1 94.335,54.11
X$15951 1304 VIA_via2_5
* cell instance $15952 r0 *1 93.765,54.11
X$15952 1304 VIA_via2_5
* cell instance $15953 r0 *1 89.965,63.21
X$15953 1304 VIA_via2_5
* cell instance $15954 r0 *1 93.765,63.21
X$15954 1304 VIA_via2_5
* cell instance $15955 r0 *1 85.025,59.01
X$15955 1304 VIA_via2_5
* cell instance $15956 r0 *1 84.835,52.71
X$15956 1304 VIA_via2_5
* cell instance $15957 r0 *1 89.965,63.63
X$15957 1304 VIA_via1_4
* cell instance $15958 r0 *1 93.765,62.37
X$15958 1304 VIA_via1_4
* cell instance $15959 r0 *1 93.765,62.23
X$15959 1304 VIA_via2_5
* cell instance $15960 r0 *1 90.345,52.43
X$15960 1304 VIA_via1_4
* cell instance $15961 r0 *1 96.615,53.97
X$15961 1304 VIA_via1_4
* cell instance $15962 r0 *1 96.615,54.11
X$15962 1304 VIA_via2_5
* cell instance $15963 r0 *1 90.345,51.17
X$15963 1304 VIA_via1_4
* cell instance $15964 r0 *1 90.155,56.77
X$15964 1304 VIA_via1_4
* cell instance $15965 r0 *1 92.625,51.205
X$15965 1304 VIA_via1_4
* cell instance $15966 r0 *1 84.645,59.15
X$15966 1304 VIA_via1_4
* cell instance $15967 r0 *1 93.765,55.23
X$15967 1304 VIA_via1_4
* cell instance $15968 r0 *1 85.595,51.17
X$15968 1304 VIA_via1_4
* cell instance $15969 r0 *1 85.025,53.97
X$15969 1304 VIA_via1_4
* cell instance $15970 r0 *1 93.615,62.23
X$15970 1304 VIA_via3_2
* cell instance $15971 r0 *1 93.615,58.87
X$15971 1304 VIA_via3_2
* cell instance $15972 r0 *1 67.735,66.99
X$15972 1305 VIA_via2_5
* cell instance $15973 r0 *1 90.345,58.45
X$15973 1305 VIA_via2_5
* cell instance $15974 r0 *1 91.295,58.45
X$15974 1305 VIA_via2_5
* cell instance $15975 r0 *1 90.535,51.59
X$15975 1305 VIA_via2_5
* cell instance $15976 r0 *1 85.785,51.45
X$15976 1305 VIA_via2_5
* cell instance $15977 r0 *1 85.025,51.45
X$15977 1305 VIA_via2_5
* cell instance $15978 r0 *1 93.955,58.45
X$15978 1305 VIA_via2_5
* cell instance $15979 r0 *1 92.815,51.59
X$15979 1305 VIA_via2_5
* cell instance $15980 r0 *1 91.295,63.07
X$15980 1305 VIA_via2_5
* cell instance $15981 r0 *1 89.015,63.63
X$15981 1305 VIA_via2_5
* cell instance $15982 r0 *1 89.015,66.99
X$15982 1305 VIA_via2_5
* cell instance $15983 r0 *1 90.155,63.07
X$15983 1305 VIA_via2_5
* cell instance $15984 r0 *1 93.955,63.07
X$15984 1305 VIA_via2_5
* cell instance $15985 r0 *1 67.735,67.97
X$15985 1305 VIA_via1_4
* cell instance $15986 r0 *1 71.915,66.85
X$15986 1305 VIA_via1_4
* cell instance $15987 r0 *1 71.915,66.99
X$15987 1305 VIA_via2_5
* cell instance $15988 r0 *1 90.155,63.63
X$15988 1305 VIA_via1_4
* cell instance $15989 r0 *1 90.155,63.63
X$15989 1305 VIA_via2_5
* cell instance $15990 r0 *1 93.955,62.37
X$15990 1305 VIA_via1_4
* cell instance $15991 r0 *1 85.785,51.17
X$15991 1305 VIA_via1_4
* cell instance $15992 r0 *1 90.535,51.17
X$15992 1305 VIA_via1_4
* cell instance $15993 r0 *1 90.535,51.31
X$15993 1305 VIA_via2_5
* cell instance $15994 r0 *1 90.345,56.77
X$15994 1305 VIA_via1_4
* cell instance $15995 r0 *1 90.535,52.43
X$15995 1305 VIA_via1_4
* cell instance $15996 r0 *1 92.815,51.17
X$15996 1305 VIA_via1_4
* cell instance $15997 r0 *1 93.955,55.23
X$15997 1305 VIA_via1_4
* cell instance $15998 r0 *1 93.955,55.23
X$15998 1305 VIA_via2_5
* cell instance $15999 r0 *1 85.215,53.97
X$15999 1305 VIA_via1_4
* cell instance $16000 r0 *1 93.615,55.23
X$16000 1305 VIA_via3_2
* cell instance $16001 r0 *1 93.615,51.59
X$16001 1305 VIA_via3_2
* cell instance $16002 r0 *1 89.015,52.01
X$16002 1306 VIA_via2_5
* cell instance $16003 r0 *1 94.905,57.19
X$16003 1306 VIA_via2_5
* cell instance $16004 r0 *1 94.905,61.25
X$16004 1306 VIA_via2_5
* cell instance $16005 r0 *1 93.195,57.19
X$16005 1306 VIA_via2_5
* cell instance $16006 r0 *1 96.615,57.19
X$16006 1306 VIA_via2_5
* cell instance $16007 r0 *1 95.285,61.25
X$16007 1306 VIA_via2_5
* cell instance $16008 r0 *1 95.095,52.29
X$16008 1306 VIA_via2_5
* cell instance $16009 r0 *1 95.095,51.73
X$16009 1306 VIA_via2_5
* cell instance $16010 r0 *1 94.905,62.23
X$16010 1306 VIA_via2_5
* cell instance $16011 r0 *1 95.665,62.37
X$16011 1306 VIA_via1_4
* cell instance $16012 r0 *1 95.665,62.23
X$16012 1306 VIA_via2_5
* cell instance $16013 r0 *1 94.905,63.63
X$16013 1306 VIA_via1_4
* cell instance $16014 r0 *1 89.015,53.97
X$16014 1306 VIA_via1_4
* cell instance $16015 r0 *1 89.015,51.17
X$16015 1306 VIA_via1_4
* cell instance $16016 r0 *1 96.615,56.77
X$16016 1306 VIA_via1_4
* cell instance $16017 r0 *1 90.725,61.25
X$16017 1306 VIA_via1_4
* cell instance $16018 r0 *1 90.725,61.25
X$16018 1306 VIA_via2_5
* cell instance $16019 r0 *1 94.905,56.77
X$16019 1306 VIA_via1_4
* cell instance $16020 r0 *1 93.195,56.77
X$16020 1306 VIA_via1_4
* cell instance $16021 r0 *1 95.095,51.17
X$16021 1306 VIA_via1_4
* cell instance $16022 r0 *1 95.095,51.31
X$16022 1306 VIA_via2_5
* cell instance $16023 r0 *1 96.425,51.17
X$16023 1306 VIA_via1_4
* cell instance $16024 r0 *1 96.425,51.31
X$16024 1306 VIA_via2_5
* cell instance $16025 r0 *1 93.195,52.43
X$16025 1306 VIA_via1_4
* cell instance $16026 r0 *1 93.195,52.29
X$16026 1306 VIA_via2_5
* cell instance $16027 r0 *1 91.105,51.17
X$16027 1307 VIA_via1_4
* cell instance $16028 r0 *1 91.105,51.31
X$16028 1307 VIA_via2_5
* cell instance $16029 r0 *1 93.195,51.17
X$16029 1307 VIA_via1_4
* cell instance $16030 r0 *1 93.195,51.17
X$16030 1307 VIA_via2_5
* cell instance $16031 r0 *1 95.855,52.57
X$16031 1308 VIA_via1_4
* cell instance $16032 r0 *1 95.855,52.57
X$16032 1308 VIA_via2_5
* cell instance $16033 r0 *1 95.855,52.57
X$16033 1308 VIA_via3_2
* cell instance $16034 r0 *1 95.855,51.59
X$16034 1308 VIA_via4_0
* cell instance $16035 r0 *1 94.905,51.59
X$16035 1309 VIA_via1_7
* cell instance $16036 r0 *1 94.905,51.59
X$16036 1309 VIA_via2_5
* cell instance $16037 r0 *1 95.475,51.59
X$16037 1309 VIA_via2_5
* cell instance $16038 r0 *1 95.475,51.17
X$16038 1309 VIA_via1_4
* cell instance $16039 r0 *1 95.285,51.45
X$16039 1310 VIA_via1_7
* cell instance $16040 r0 *1 95.285,51.45
X$16040 1310 VIA_via2_5
* cell instance $16041 r0 *1 96.045,51.45
X$16041 1310 VIA_via2_5
* cell instance $16042 r0 *1 96.045,52.43
X$16042 1310 VIA_via1_4
* cell instance $16043 r0 *1 11.875,51.17
X$16043 1311 VIA_via1_4
* cell instance $16044 r0 *1 11.685,51.17
X$16044 1311 VIA_via1_4
* cell instance $16045 r0 *1 17.005,51.17
X$16045 1312 VIA_via1_4
* cell instance $16046 r0 *1 17.005,51.17
X$16046 1312 VIA_via2_5
* cell instance $16047 r0 *1 17.575,51.17
X$16047 1312 VIA_via1_4
* cell instance $16048 r0 *1 17.575,51.17
X$16048 1312 VIA_via2_5
* cell instance $16049 r0 *1 94.145,51.59
X$16049 1313 VIA_via1_7
* cell instance $16050 r0 *1 94.145,51.87
X$16050 1313 VIA_via2_5
* cell instance $16051 r0 *1 91.865,51.87
X$16051 1313 VIA_via2_5
* cell instance $16052 r0 *1 91.865,51.17
X$16052 1313 VIA_via1_4
* cell instance $16053 r0 *1 22.895,51.59
X$16053 1314 VIA_via1_7
* cell instance $16054 r0 *1 22.895,51.73
X$16054 1314 VIA_via2_5
* cell instance $16055 r0 *1 20.425,51.73
X$16055 1314 VIA_via2_5
* cell instance $16056 r0 *1 20.425,52.43
X$16056 1314 VIA_via1_4
* cell instance $16057 r0 *1 24.605,49.91
X$16057 1315 VIA_via1_7
* cell instance $16058 r0 *1 24.605,51.17
X$16058 1315 VIA_via1_4
* cell instance $16059 r0 *1 89.585,51.17
X$16059 1316 VIA_via1_4
* cell instance $16060 r0 *1 89.585,51.17
X$16060 1316 VIA_via2_5
* cell instance $16061 r0 *1 85.405,51.17
X$16061 1316 VIA_via1_4
* cell instance $16062 r0 *1 85.405,51.17
X$16062 1316 VIA_via2_5
* cell instance $16063 r0 *1 83.695,51.17
X$16063 1317 VIA_via1_4
* cell instance $16064 r0 *1 83.695,51.17
X$16064 1317 VIA_via2_5
* cell instance $16065 r0 *1 84.835,51.17
X$16065 1317 VIA_via1_4
* cell instance $16066 r0 *1 84.835,51.17
X$16066 1317 VIA_via2_5
* cell instance $16067 r0 *1 72.295,66.57
X$16067 1318 VIA_via2_5
* cell instance $16068 r0 *1 72.295,65.17
X$16068 1318 VIA_via1_4
* cell instance $16069 r0 *1 54.625,72.03
X$16069 1318 VIA_via1_4
* cell instance $16070 r0 *1 54.625,71.89
X$16070 1318 VIA_via2_5
* cell instance $16071 r0 *1 80.465,76.23
X$16071 1318 VIA_via1_4
* cell instance $16072 r0 *1 80.465,76.23
X$16072 1318 VIA_via2_5
* cell instance $16073 r0 *1 52.915,51.17
X$16073 1318 VIA_via1_4
* cell instance $16074 r0 *1 52.915,51.17
X$16074 1318 VIA_via2_5
* cell instance $16075 r0 *1 53.015,51.17
X$16075 1318 VIA_via3_2
* cell instance $16076 r0 *1 53.015,51.31
X$16076 1318 VIA_via4_0
* cell instance $16077 r0 *1 82.365,51.17
X$16077 1318 VIA_via1_4
* cell instance $16078 r0 *1 82.365,51.31
X$16078 1318 VIA_via2_5
* cell instance $16079 r0 *1 80.085,52.43
X$16079 1318 VIA_via1_4
* cell instance $16080 r0 *1 80.085,52.29
X$16080 1318 VIA_via2_5
* cell instance $16081 r0 *1 61.135,69.51
X$16081 1318 VIA_via4_0
* cell instance $16082 r0 *1 72.895,69.51
X$16082 1318 VIA_via4_0
* cell instance $16083 r0 *1 81.015,51.31
X$16083 1318 VIA_via4_0
* cell instance $16084 r0 *1 81.015,51.31
X$16084 1318 VIA_via3_2
* cell instance $16085 r0 *1 79.895,76.23
X$16085 1318 VIA_via3_2
* cell instance $16086 r0 *1 81.015,52.29
X$16086 1318 VIA_via3_2
* cell instance $16087 r0 *1 61.135,71.89
X$16087 1318 VIA_via3_2
* cell instance $16088 r0 *1 72.895,66.57
X$16088 1318 VIA_via3_2
* cell instance $16089 r0 *1 79.895,66.57
X$16089 1318 VIA_via3_2
* cell instance $16090 r0 *1 81.015,66.57
X$16090 1318 VIA_via3_2
* cell instance $16091 r0 *1 88.445,91.21
X$16091 1319 VIA_via2_5
* cell instance $16092 r0 *1 87.685,91.21
X$16092 1319 VIA_via2_5
* cell instance $16093 r0 *1 81.605,77.77
X$16093 1319 VIA_via2_5
* cell instance $16094 r0 *1 80.465,91.49
X$16094 1319 VIA_via2_5
* cell instance $16095 r0 *1 80.465,90.65
X$16095 1319 VIA_via2_5
* cell instance $16096 r0 *1 84.835,91.07
X$16096 1319 VIA_via2_5
* cell instance $16097 r0 *1 62.605,51.45
X$16097 1319 VIA_via2_5
* cell instance $16098 r0 *1 62.605,51.73
X$16098 1319 VIA_via2_5
* cell instance $16099 r0 *1 55.385,51.45
X$16099 1319 VIA_via2_5
* cell instance $16100 r0 *1 55.385,52.15
X$16100 1319 VIA_via2_5
* cell instance $16101 r0 *1 74.005,85.05
X$16101 1319 VIA_via2_5
* cell instance $16102 r0 *1 81.795,53.83
X$16102 1319 VIA_via2_5
* cell instance $16103 r0 *1 80.655,53.83
X$16103 1319 VIA_via2_5
* cell instance $16104 r0 *1 81.795,51.73
X$16104 1319 VIA_via2_5
* cell instance $16105 r0 *1 70.205,90.65
X$16105 1319 VIA_via2_5
* cell instance $16106 r0 *1 48.355,52.15
X$16106 1319 VIA_via2_5
* cell instance $16107 r0 *1 80.655,95.97
X$16107 1319 VIA_via1_4
* cell instance $16108 r0 *1 74.005,84.77
X$16108 1319 VIA_via1_4
* cell instance $16109 r0 *1 84.835,91.63
X$16109 1319 VIA_via1_4
* cell instance $16110 r0 *1 84.835,91.49
X$16110 1319 VIA_via2_5
* cell instance $16111 r0 *1 88.635,93.17
X$16111 1319 VIA_via1_4
* cell instance $16112 r0 *1 87.495,91.63
X$16112 1319 VIA_via1_4
* cell instance $16113 r0 *1 70.205,90.37
X$16113 1319 VIA_via1_4
* cell instance $16114 r0 *1 80.845,77.77
X$16114 1319 VIA_via1_4
* cell instance $16115 r0 *1 80.845,77.77
X$16115 1319 VIA_via2_5
* cell instance $16116 r0 *1 80.735,77.77
X$16116 1319 VIA_via3_2
* cell instance $16117 r0 *1 48.355,52.43
X$16117 1319 VIA_via1_4
* cell instance $16118 r0 *1 55.385,52.36
X$16118 1319 VIA_via1_4
* cell instance $16119 r0 *1 80.655,56.77
X$16119 1319 VIA_via1_4
* cell instance $16120 r0 *1 82.555,53.97
X$16120 1319 VIA_via1_4
* cell instance $16121 r0 *1 82.555,53.83
X$16121 1319 VIA_via2_5
* cell instance $16122 r0 *1 80.735,85.05
X$16122 1319 VIA_via3_2
* cell instance $16123 r0 *1 80.735,90.65
X$16123 1319 VIA_via3_2
* cell instance $16124 r0 *1 73.735,90.65
X$16124 1319 VIA_via3_2
* cell instance $16125 r0 *1 73.735,85.05
X$16125 1319 VIA_via3_2
* cell instance $16126 r0 *1 78.185,51.17
X$16126 1320 VIA_via1_4
* cell instance $16127 r0 *1 78.185,51.17
X$16127 1320 VIA_via2_5
* cell instance $16128 r0 *1 81.795,51.17
X$16128 1320 VIA_via1_4
* cell instance $16129 r0 *1 81.795,51.17
X$16129 1320 VIA_via2_5
* cell instance $16130 r0 *1 68.305,51.17
X$16130 1321 VIA_via1_4
* cell instance $16131 r0 *1 68.305,51.17
X$16131 1321 VIA_via2_5
* cell instance $16132 r0 *1 70.395,51.17
X$16132 1321 VIA_via1_4
* cell instance $16133 r0 *1 70.395,51.17
X$16133 1321 VIA_via2_5
* cell instance $16134 r0 *1 3.325,52.15
X$16134 1322 VIA_via2_5
* cell instance $16135 r0 *1 3.325,52.43
X$16135 1322 VIA_via1_4
* cell instance $16136 r0 *1 1.775,52.15
X$16136 1322 VIA_via4_0
* cell instance $16137 r0 *1 1.775,52.15
X$16137 1322 VIA_via3_2
* cell instance $16138 r0 *1 3.135,52.71
X$16138 1323 VIA_via1_4
* cell instance $16139 r0 *1 3.135,52.71
X$16139 1323 VIA_via2_5
* cell instance $16140 r0 *1 1.495,52.71
X$16140 1323 VIA_via3_2
* cell instance $16141 r0 *1 1.495,52.71
X$16141 1323 VIA_via4_0
* cell instance $16142 r0 *1 19.095,52.71
X$16142 1324 VIA_via1_7
* cell instance $16143 r0 *1 19.095,52.57
X$16143 1324 VIA_via2_5
* cell instance $16144 r0 *1 2.755,52.43
X$16144 1324 VIA_via1_4
* cell instance $16145 r0 *1 2.755,52.29
X$16145 1324 VIA_via2_5
* cell instance $16146 r0 *1 6.935,57.75
X$16146 1325 VIA_via2_5
* cell instance $16147 r0 *1 9.785,57.75
X$16147 1325 VIA_via2_5
* cell instance $16148 r0 *1 5.985,57.75
X$16148 1325 VIA_via2_5
* cell instance $16149 r0 *1 4.085,57.75
X$16149 1325 VIA_via2_5
* cell instance $16150 r0 *1 4.085,52.85
X$16150 1325 VIA_via2_5
* cell instance $16151 r0 *1 8.835,54.25
X$16151 1325 VIA_via2_5
* cell instance $16152 r0 *1 7.695,54.25
X$16152 1325 VIA_via2_5
* cell instance $16153 r0 *1 6.935,54.25
X$16153 1325 VIA_via2_5
* cell instance $16154 r0 *1 8.835,53.97
X$16154 1325 VIA_via1_4
* cell instance $16155 r0 *1 6.935,55.23
X$16155 1325 VIA_via1_4
* cell instance $16156 r0 *1 7.505,52.43
X$16156 1325 VIA_via1_4
* cell instance $16157 r0 *1 4.085,58.03
X$16157 1325 VIA_via1_4
* cell instance $16158 r0 *1 5.985,58.03
X$16158 1325 VIA_via1_4
* cell instance $16159 r0 *1 3.705,52.85
X$16159 1325 VIA_via1_4
* cell instance $16160 r0 *1 3.705,52.85
X$16160 1325 VIA_via2_5
* cell instance $16161 r0 *1 9.785,58.03
X$16161 1325 VIA_via1_4
* cell instance $16162 r0 *1 22.515,58.03
X$16162 1325 VIA_via1_4
* cell instance $16163 r0 *1 22.515,57.89
X$16163 1325 VIA_via2_5
* cell instance $16164 r0 *1 15.105,55.23
X$16164 1326 VIA_via2_5
* cell instance $16165 r0 *1 17.005,53.55
X$16165 1326 VIA_via2_5
* cell instance $16166 r0 *1 13.965,52.43
X$16166 1326 VIA_via2_5
* cell instance $16167 r0 *1 14.535,53.55
X$16167 1326 VIA_via2_5
* cell instance $16168 r0 *1 25.365,53.55
X$16168 1326 VIA_via2_5
* cell instance $16169 r0 *1 8.835,52.43
X$16169 1326 VIA_via2_5
* cell instance $16170 r0 *1 25.365,51.17
X$16170 1326 VIA_via1_4
* cell instance $16171 r0 *1 16.625,53.97
X$16171 1326 VIA_via1_4
* cell instance $16172 r0 *1 13.965,49.63
X$16172 1326 VIA_via1_4
* cell instance $16173 r0 *1 16.435,53.97
X$16173 1326 VIA_via1_4
* cell instance $16174 r0 *1 14.535,52.43
X$16174 1326 VIA_via1_4
* cell instance $16175 r0 *1 14.535,52.43
X$16175 1326 VIA_via2_5
* cell instance $16176 r0 *1 10.545,52.43
X$16176 1326 VIA_via1_4
* cell instance $16177 r0 *1 10.545,52.43
X$16177 1326 VIA_via2_5
* cell instance $16178 r0 *1 8.835,51.17
X$16178 1326 VIA_via1_4
* cell instance $16179 r0 *1 15.105,59.57
X$16179 1326 VIA_via1_4
* cell instance $16180 r0 *1 17.005,55.23
X$16180 1326 VIA_via1_4
* cell instance $16181 r0 *1 17.005,55.23
X$16181 1326 VIA_via2_5
* cell instance $16182 r0 *1 9.405,52.71
X$16182 1327 VIA_via2_5
* cell instance $16183 r0 *1 10.735,52.71
X$16183 1327 VIA_via2_5
* cell instance $16184 r0 *1 12.065,52.71
X$16184 1327 VIA_via1_4
* cell instance $16185 r0 *1 12.065,52.71
X$16185 1327 VIA_via2_5
* cell instance $16186 r0 *1 10.735,51.17
X$16186 1327 VIA_via1_4
* cell instance $16187 r0 *1 9.405,53.97
X$16187 1327 VIA_via1_4
* cell instance $16188 r0 *1 13.585,53.41
X$16188 1328 VIA_via1_7
* cell instance $16189 r0 *1 13.775,52.43
X$16189 1328 VIA_via1_4
* cell instance $16190 r0 *1 22.135,52.43
X$16190 1329 VIA_via1_4
* cell instance $16191 r0 *1 21.755,52.15
X$16191 1329 VIA_via1_4
* cell instance $16192 r0 *1 22.515,52.15
X$16192 1330 VIA_via2_5
* cell instance $16193 r0 *1 24.035,52.29
X$16193 1330 VIA_via2_5
* cell instance $16194 r0 *1 23.085,52.43
X$16194 1330 VIA_via1_4
* cell instance $16195 r0 *1 23.085,52.29
X$16195 1330 VIA_via2_5
* cell instance $16196 r0 *1 24.035,53.55
X$16196 1330 VIA_via1_4
* cell instance $16197 r0 *1 21.755,52.43
X$16197 1330 VIA_via1_4
* cell instance $16198 r0 *1 21.755,52.43
X$16198 1330 VIA_via2_5
* cell instance $16199 r0 *1 22.515,51.17
X$16199 1330 VIA_via1_4
* cell instance $16200 r0 *1 80.085,74.55
X$16200 1331 VIA_via1_7
* cell instance $16201 r0 *1 84.075,74.55
X$16201 1331 VIA_via1_7
* cell instance $16202 r0 *1 84.075,74.55
X$16202 1331 VIA_via2_5
* cell instance $16203 r0 *1 89.775,62.09
X$16203 1331 VIA_via2_5
* cell instance $16204 r0 *1 37.335,54.39
X$16204 1331 VIA_via2_5
* cell instance $16205 r0 *1 41.515,54.67
X$16205 1331 VIA_via2_5
* cell instance $16206 r0 *1 45.315,69.51
X$16206 1331 VIA_via2_5
* cell instance $16207 r0 *1 41.515,55.23
X$16207 1331 VIA_via1_4
* cell instance $16208 r0 *1 42.275,55.51
X$16208 1331 VIA_via1_4
* cell instance $16209 r0 *1 37.145,52.71
X$16209 1331 VIA_via1_4
* cell instance $16210 r0 *1 45.315,77.63
X$16210 1331 VIA_via1_4
* cell instance $16211 r0 *1 43.225,69.37
X$16211 1331 VIA_via1_4
* cell instance $16212 r0 *1 44.745,69.51
X$16212 1331 VIA_via1_4
* cell instance $16213 r0 *1 44.745,69.51
X$16213 1331 VIA_via2_5
* cell instance $16214 r0 *1 90.155,62.37
X$16214 1331 VIA_via1_4
* cell instance $16215 r0 *1 90.155,62.37
X$16215 1331 VIA_via2_5
* cell instance $16216 r0 *1 89.775,60.83
X$16216 1331 VIA_via1_4
* cell instance $16217 r0 *1 89.415,62.37
X$16217 1331 VIA_via3_2
* cell instance $16218 r0 *1 89.415,74.55
X$16218 1331 VIA_via3_2
* cell instance $16219 r0 *1 45.455,74.27
X$16219 1331 VIA_via3_2
* cell instance $16220 r0 *1 45.315,74.27
X$16220 1331 VIA_via2_5
* cell instance $16221 r0 *1 45.455,74.27
X$16221 1331 VIA_via4_0
* cell instance $16222 r0 *1 80.175,74.27
X$16222 1331 VIA_via3_2
* cell instance $16223 r0 *1 80.085,74.27
X$16223 1331 VIA_via2_5
* cell instance $16224 r0 *1 80.175,74.27
X$16224 1331 VIA_via4_0
* cell instance $16225 r0 *1 71.345,60.55
X$16225 1332 VIA_via1_7
* cell instance $16226 r0 *1 55.005,55.65
X$16226 1332 VIA_via2_5
* cell instance $16227 r0 *1 54.815,52.71
X$16227 1332 VIA_via2_5
* cell instance $16228 r0 *1 54.695,52.71
X$16228 1332 VIA_via3_2
* cell instance $16229 r0 *1 81.985,54.39
X$16229 1332 VIA_via2_5
* cell instance $16230 r0 *1 80.085,57.19
X$16230 1332 VIA_via2_5
* cell instance $16231 r0 *1 36.195,52.57
X$16231 1332 VIA_via2_5
* cell instance $16232 r0 *1 90.155,73.57
X$16232 1332 VIA_via1_4
* cell instance $16233 r0 *1 90.155,73.57
X$16233 1332 VIA_via2_5
* cell instance $16234 r0 *1 90.255,73.57
X$16234 1332 VIA_via3_2
* cell instance $16235 r0 *1 36.195,53.97
X$16235 1332 VIA_via1_4
* cell instance $16236 r0 *1 47.785,52.43
X$16236 1332 VIA_via1_4
* cell instance $16237 r0 *1 47.785,52.57
X$16237 1332 VIA_via2_5
* cell instance $16238 r0 *1 54.815,52.43
X$16238 1332 VIA_via1_4
* cell instance $16239 r0 *1 80.085,56.77
X$16239 1332 VIA_via1_4
* cell instance $16240 r0 *1 81.985,53.97
X$16240 1332 VIA_via1_4
* cell instance $16241 r0 *1 48.255,52.43
X$16241 1332 VIA_via4_0
* cell instance $16242 r0 *1 48.255,52.43
X$16242 1332 VIA_via3_2
* cell instance $16243 r0 *1 79.895,56.91
X$16243 1332 VIA_via4_0
* cell instance $16244 r0 *1 54.695,52.43
X$16244 1332 VIA_via4_0
* cell instance $16245 r0 *1 90.255,57.19
X$16245 1332 VIA_via3_2
* cell instance $16246 r0 *1 79.895,57.19
X$16246 1332 VIA_via3_2
* cell instance $16247 r0 *1 82.135,57.19
X$16247 1332 VIA_via3_2
* cell instance $16248 r0 *1 71.215,56.91
X$16248 1332 VIA_via3_2
* cell instance $16249 r0 *1 71.215,56.91
X$16249 1332 VIA_via4_0
* cell instance $16250 r0 *1 71.345,56.91
X$16250 1332 VIA_via2_5
* cell instance $16251 r0 *1 82.135,54.39
X$16251 1332 VIA_via3_2
* cell instance $16252 r0 *1 71.215,55.65
X$16252 1332 VIA_via3_2
* cell instance $16253 r0 *1 54.625,52.43
X$16253 1333 VIA_via1_4
* cell instance $16254 r0 *1 54.625,52.43
X$16254 1333 VIA_via2_5
* cell instance $16255 r0 *1 57.665,52.43
X$16255 1333 VIA_via1_4
* cell instance $16256 r0 *1 57.665,52.29
X$16256 1333 VIA_via2_5
* cell instance $16257 r0 *1 57.855,53.55
X$16257 1333 VIA_via1_4
* cell instance $16258 r0 *1 58.235,52.43
X$16258 1333 VIA_via1_4
* cell instance $16259 r0 *1 58.235,52.29
X$16259 1333 VIA_via2_5
* cell instance $16260 r0 *1 54.625,52.15
X$16260 1334 VIA_via1_4
* cell instance $16261 r0 *1 55.005,52.43
X$16261 1334 VIA_via1_4
* cell instance $16262 r0 *1 66.025,58.03
X$16262 1335 VIA_via2_5
* cell instance $16263 r0 *1 66.595,58.03
X$16263 1335 VIA_via2_5
* cell instance $16264 r0 *1 65.265,52.57
X$16264 1335 VIA_via2_5
* cell instance $16265 r0 *1 65.265,54.53
X$16265 1335 VIA_via2_5
* cell instance $16266 r0 *1 66.595,54.53
X$16266 1335 VIA_via2_5
* cell instance $16267 r0 *1 67.165,52.57
X$16267 1335 VIA_via2_5
* cell instance $16268 r0 *1 65.265,67.97
X$16268 1335 VIA_via2_5
* cell instance $16269 r0 *1 66.025,62.93
X$16269 1335 VIA_via2_5
* cell instance $16270 r0 *1 65.265,62.93
X$16270 1335 VIA_via2_5
* cell instance $16271 r0 *1 70.395,72.31
X$16271 1335 VIA_via2_5
* cell instance $16272 r0 *1 69.635,54.39
X$16272 1335 VIA_via2_5
* cell instance $16273 r0 *1 66.215,67.97
X$16273 1335 VIA_via1_4
* cell instance $16274 r0 *1 66.215,67.97
X$16274 1335 VIA_via2_5
* cell instance $16275 r0 *1 67.165,72.03
X$16275 1335 VIA_via1_4
* cell instance $16276 r0 *1 67.165,71.89
X$16276 1335 VIA_via2_5
* cell instance $16277 r0 *1 70.585,70.77
X$16277 1335 VIA_via1_4
* cell instance $16278 r0 *1 94.525,72.45
X$16278 1335 VIA_via1_4
* cell instance $16279 r0 *1 94.525,72.31
X$16279 1335 VIA_via2_5
* cell instance $16280 r0 *1 67.165,51.17
X$16280 1335 VIA_via1_4
* cell instance $16281 r0 *1 69.825,53.97
X$16281 1335 VIA_via1_4
* cell instance $16282 r0 *1 65.075,52.43
X$16282 1335 VIA_via1_4
* cell instance $16283 r0 *1 66.595,55.23
X$16283 1335 VIA_via1_4
* cell instance $16284 r0 *1 66.735,71.89
X$16284 1335 VIA_via3_2
* cell instance $16285 r0 *1 66.735,67.97
X$16285 1335 VIA_via3_2
* cell instance $16286 r0 *1 76.665,60.83
X$16286 1336 VIA_via2_5
* cell instance $16287 r0 *1 76.665,59.57
X$16287 1336 VIA_via2_5
* cell instance $16288 r0 *1 73.625,56.21
X$16288 1336 VIA_via2_5
* cell instance $16289 r0 *1 74.765,59.57
X$16289 1336 VIA_via2_5
* cell instance $16290 r0 *1 74.955,56.21
X$16290 1336 VIA_via2_5
* cell instance $16291 r0 *1 74.765,56.21
X$16291 1336 VIA_via2_5
* cell instance $16292 r0 *1 78.185,65.17
X$16292 1336 VIA_via2_5
* cell instance $16293 r0 *1 77.045,65.17
X$16293 1336 VIA_via2_5
* cell instance $16294 r0 *1 77.045,63.63
X$16294 1336 VIA_via2_5
* cell instance $16295 r0 *1 76.475,65.17
X$16295 1336 VIA_via1_4
* cell instance $16296 r0 *1 76.475,65.17
X$16296 1336 VIA_via2_5
* cell instance $16297 r0 *1 78.185,66.43
X$16297 1336 VIA_via1_4
* cell instance $16298 r0 *1 76.665,60.55
X$16298 1336 VIA_via1_4
* cell instance $16299 r0 *1 77.045,61.25
X$16299 1336 VIA_via1_4
* cell instance $16300 r0 *1 76.095,59.57
X$16300 1336 VIA_via1_4
* cell instance $16301 r0 *1 76.095,59.57
X$16301 1336 VIA_via2_5
* cell instance $16302 r0 *1 73.625,56.77
X$16302 1336 VIA_via1_4
* cell instance $16303 r0 *1 75.145,52.43
X$16303 1336 VIA_via1_4
* cell instance $16304 r0 *1 73.815,63.63
X$16304 1336 VIA_via1_4
* cell instance $16305 r0 *1 73.815,63.63
X$16305 1336 VIA_via2_5
* cell instance $16306 r0 *1 80.845,60.83
X$16306 1336 VIA_via1_4
* cell instance $16307 r0 *1 80.845,60.83
X$16307 1336 VIA_via2_5
* cell instance $16308 r0 *1 74.955,55.23
X$16308 1336 VIA_via1_4
* cell instance $16309 r0 *1 76.665,52.43
X$16309 1337 VIA_via1_4
* cell instance $16310 r0 *1 76.665,52.43
X$16310 1337 VIA_via2_5
* cell instance $16311 r0 *1 77.615,52.43
X$16311 1337 VIA_via1_4
* cell instance $16312 r0 *1 77.615,52.43
X$16312 1337 VIA_via2_5
* cell instance $16313 r0 *1 77.805,53.97
X$16313 1337 VIA_via1_4
* cell instance $16314 r0 *1 85.785,52.29
X$16314 1338 VIA_via1_4
* cell instance $16315 r0 *1 85.215,52.43
X$16315 1338 VIA_via1_4
* cell instance $16316 r0 *1 95.475,52.71
X$16316 1339 VIA_via2_5
* cell instance $16317 r0 *1 95.475,52.43
X$16317 1339 VIA_via1_4
* cell instance $16318 r0 *1 84.455,52.85
X$16318 1339 VIA_via1_4
* cell instance $16319 r0 *1 84.455,52.85
X$16319 1339 VIA_via2_5
* cell instance $16320 r0 *1 85.215,52.99
X$16320 1340 VIA_via1_7
* cell instance $16321 r0 *1 85.215,52.99
X$16321 1340 VIA_via2_5
* cell instance $16322 r0 *1 95.665,52.99
X$16322 1340 VIA_via2_5
* cell instance $16323 r0 *1 95.855,51.17
X$16323 1340 VIA_via1_4
* cell instance $16324 r0 *1 96.425,52.57
X$16324 1341 VIA_via1_4
* cell instance $16325 r0 *1 96.425,52.57
X$16325 1341 VIA_via2_5
* cell instance $16326 r0 *1 97.255,52.15
X$16326 1341 VIA_via4_0
* cell instance $16327 r0 *1 97.255,52.57
X$16327 1341 VIA_via3_2
* cell instance $16328 r0 *1 96.425,53.41
X$16328 1342 VIA_via1_7
* cell instance $16329 r0 *1 96.425,53.41
X$16329 1342 VIA_via2_5
* cell instance $16330 r0 *1 97.535,52.71
X$16330 1342 VIA_via4_0
* cell instance $16331 r0 *1 97.535,53.41
X$16331 1342 VIA_via3_2
* cell instance $16332 r0 *1 17.385,50.89
X$16332 1343 VIA_via1_7
* cell instance $16333 r0 *1 1.425,52.01
X$16333 1343 VIA_via2_5
* cell instance $16334 r0 *1 17.385,52.01
X$16334 1343 VIA_via2_5
* cell instance $16335 r0 *1 1.425,52.43
X$16335 1343 VIA_via1_4
* cell instance $16336 r0 *1 96.615,51.45
X$16336 1344 VIA_via1_7
* cell instance $16337 r0 *1 96.615,52.43
X$16337 1344 VIA_via1_4
* cell instance $16338 r0 *1 5.985,53.41
X$16338 1345 VIA_via1_7
* cell instance $16339 r0 *1 5.985,52.57
X$16339 1345 VIA_via2_5
* cell instance $16340 r0 *1 4.845,52.43
X$16340 1345 VIA_via1_4
* cell instance $16341 r0 *1 4.845,52.57
X$16341 1345 VIA_via2_5
* cell instance $16342 r0 *1 50.255,94.57
X$16342 1346 VIA_via1_7
* cell instance $16343 r0 *1 50.255,94.57
X$16343 1346 VIA_via2_5
* cell instance $16344 r0 *1 36.955,95.83
X$16344 1346 VIA_via1_7
* cell instance $16345 r0 *1 36.955,95.83
X$16345 1346 VIA_via2_5
* cell instance $16346 r0 *1 4.655,65.45
X$16346 1346 VIA_via2_5
* cell instance $16347 r0 *1 32.965,94.15
X$16347 1346 VIA_via2_5
* cell instance $16348 r0 *1 4.845,82.53
X$16348 1346 VIA_via2_5
* cell instance $16349 r0 *1 3.705,82.53
X$16349 1346 VIA_via2_5
* cell instance $16350 r0 *1 6.745,82.53
X$16350 1346 VIA_via2_5
* cell instance $16351 r0 *1 5.035,65.45
X$16351 1346 VIA_via2_5
* cell instance $16352 r0 *1 6.555,94.15
X$16352 1346 VIA_via2_5
* cell instance $16353 r0 *1 14.725,94.15
X$16353 1346 VIA_via2_5
* cell instance $16354 r0 *1 50.635,94.57
X$16354 1346 VIA_via2_5
* cell instance $16355 r0 *1 50.635,95.83
X$16355 1346 VIA_via2_5
* cell instance $16356 r0 *1 54.245,86.17
X$16356 1346 VIA_via2_5
* cell instance $16357 r0 *1 54.245,84.91
X$16357 1346 VIA_via2_5
* cell instance $16358 r0 *1 36.955,94.15
X$16358 1346 VIA_via2_5
* cell instance $16359 r0 *1 57.475,84.77
X$16359 1346 VIA_via1_4
* cell instance $16360 r0 *1 57.495,84.91
X$16360 1346 VIA_via3_2
* cell instance $16361 r0 *1 57.475,84.91
X$16361 1346 VIA_via2_5
* cell instance $16362 r0 *1 14.725,93.17
X$16362 1346 VIA_via1_4
* cell instance $16363 r0 *1 32.965,94.43
X$16363 1346 VIA_via1_4
* cell instance $16364 r0 *1 7.315,52.43
X$16364 1346 VIA_via1_4
* cell instance $16365 r0 *1 7.315,52.43
X$16365 1346 VIA_via2_5
* cell instance $16366 r0 *1 7.375,52.43
X$16366 1346 VIA_via3_2
* cell instance $16367 r0 *1 5.035,65.17
X$16367 1346 VIA_via1_4
* cell instance $16368 r0 *1 3.705,83.23
X$16368 1346 VIA_via1_4
* cell instance $16369 r0 *1 6.555,94.43
X$16369 1346 VIA_via1_4
* cell instance $16370 r0 *1 57.475,58.45
X$16370 1346 VIA_via1_4
* cell instance $16371 r0 *1 57.495,58.45
X$16371 1346 VIA_via3_2
* cell instance $16372 r0 *1 57.475,58.45
X$16372 1346 VIA_via2_5
* cell instance $16373 r0 *1 55.385,60.83
X$16373 1346 VIA_via1_4
* cell instance $16374 r0 *1 55.385,60.83
X$16374 1346 VIA_via2_5
* cell instance $16375 r0 *1 7.375,65.45
X$16375 1346 VIA_via3_2
* cell instance $16376 r0 *1 57.495,60.83
X$16376 1346 VIA_via3_2
* cell instance $16377 r0 *1 51.055,94.57
X$16377 1346 VIA_via3_2
* cell instance $16378 r0 *1 51.055,86.17
X$16378 1346 VIA_via3_2
* cell instance $16379 r0 *1 95.285,52.57
X$16379 1347 VIA_via2_5
* cell instance $16380 r0 *1 95.285,53.97
X$16380 1347 VIA_via1_4
* cell instance $16381 r0 *1 93.385,52.57
X$16381 1347 VIA_via1_4
* cell instance $16382 r0 *1 93.385,52.57
X$16382 1347 VIA_via2_5
* cell instance $16383 r0 *1 90.155,52.43
X$16383 1348 VIA_via1_4
* cell instance $16384 r0 *1 90.155,52.43
X$16384 1348 VIA_via2_5
* cell instance $16385 r0 *1 93.765,52.43
X$16385 1348 VIA_via1_4
* cell instance $16386 r0 *1 93.765,52.43
X$16386 1348 VIA_via2_5
* cell instance $16387 r0 *1 23.275,52.43
X$16387 1349 VIA_via1_4
* cell instance $16388 r0 *1 23.275,52.43
X$16388 1349 VIA_via2_5
* cell instance $16389 r0 *1 22.895,52.43
X$16389 1349 VIA_via1_4
* cell instance $16390 r0 *1 22.895,52.43
X$16390 1349 VIA_via2_5
* cell instance $16391 r0 *1 85.405,52.43
X$16391 1350 VIA_via1_4
* cell instance $16392 r0 *1 85.405,52.43
X$16392 1350 VIA_via2_5
* cell instance $16393 r0 *1 83.505,52.43
X$16393 1350 VIA_via1_4
* cell instance $16394 r0 *1 83.505,52.43
X$16394 1350 VIA_via2_5
* cell instance $16395 r0 *1 58.615,52.15
X$16395 1351 VIA_via2_5
* cell instance $16396 r0 *1 58.615,52.15
X$16396 1351 VIA_via3_2
* cell instance $16397 r0 *1 58.615,52.15
X$16397 1351 VIA_via4_0
* cell instance $16398 r0 *1 58.615,52.15
X$16398 1351 VIA_via1_4
* cell instance $16399 r0 *1 84.455,52.43
X$16399 1351 VIA_via1_4
* cell instance $16400 r0 *1 84.455,52.57
X$16400 1351 VIA_via2_5
* cell instance $16401 r0 *1 84.375,52.57
X$16401 1351 VIA_via3_2
* cell instance $16402 r0 *1 84.375,52.15
X$16402 1351 VIA_via4_0
* cell instance $16403 r0 *1 57.475,52.57
X$16403 1352 VIA_via1_4
* cell instance $16404 r0 *1 57.475,52.71
X$16404 1352 VIA_via2_5
* cell instance $16405 r0 *1 84.645,52.43
X$16405 1352 VIA_via1_4
* cell instance $16406 r0 *1 84.645,52.29
X$16406 1352 VIA_via2_5
* cell instance $16407 r0 *1 82.135,52.71
X$16407 1352 VIA_via4_0
* cell instance $16408 r0 *1 58.615,52.71
X$16408 1352 VIA_via4_0
* cell instance $16409 r0 *1 58.615,52.71
X$16409 1352 VIA_via3_2
* cell instance $16410 r0 *1 82.135,52.29
X$16410 1352 VIA_via3_2
* cell instance $16411 r0 *1 42.465,51.59
X$16411 1353 VIA_via1_7
* cell instance $16412 r0 *1 42.465,52.43
X$16412 1353 VIA_via2_5
* cell instance $16413 r0 *1 47.975,52.43
X$16413 1353 VIA_via1_4
* cell instance $16414 r0 *1 47.975,52.43
X$16414 1353 VIA_via2_5
* cell instance $16415 r0 *1 74.385,52.43
X$16415 1354 VIA_via1_4
* cell instance $16416 r0 *1 74.385,52.57
X$16416 1354 VIA_via2_5
* cell instance $16417 r0 *1 77.995,52.57
X$16417 1354 VIA_via1_4
* cell instance $16418 r0 *1 77.995,52.57
X$16418 1354 VIA_via2_5
* cell instance $16419 r0 *1 71.535,52.29
X$16419 1355 VIA_via2_5
* cell instance $16420 r0 *1 70.585,52.29
X$16420 1355 VIA_via2_5
* cell instance $16421 r0 *1 71.725,75.95
X$16421 1355 VIA_via1_4
* cell instance $16422 r0 *1 71.725,75.95
X$16422 1355 VIA_via2_5
* cell instance $16423 r0 *1 71.775,75.95
X$16423 1355 VIA_via3_2
* cell instance $16424 r0 *1 69.825,52.43
X$16424 1355 VIA_via1_4
* cell instance $16425 r0 *1 69.825,52.29
X$16425 1355 VIA_via2_5
* cell instance $16426 r0 *1 70.585,51.17
X$16426 1355 VIA_via1_4
* cell instance $16427 r0 *1 71.535,49.63
X$16427 1355 VIA_via1_4
* cell instance $16428 r0 *1 71.775,52.29
X$16428 1355 VIA_via3_2
* cell instance $16429 r0 *1 69.065,52.43
X$16429 1356 VIA_via1_4
* cell instance $16430 r0 *1 69.065,52.43
X$16430 1356 VIA_via2_5
* cell instance $16431 r0 *1 70.395,52.43
X$16431 1356 VIA_via1_4
* cell instance $16432 r0 *1 70.395,52.43
X$16432 1356 VIA_via2_5
* cell instance $16433 r0 *1 55.765,52.43
X$16433 1357 VIA_via1_4
* cell instance $16434 r0 *1 55.765,52.43
X$16434 1357 VIA_via2_5
* cell instance $16435 r0 *1 57.855,52.43
X$16435 1357 VIA_via1_4
* cell instance $16436 r0 *1 57.855,52.43
X$16436 1357 VIA_via2_5
* cell instance $16437 r0 *1 17.385,93.03
X$16437 1358 VIA_via1_7
* cell instance $16438 r0 *1 54.435,63.77
X$16438 1358 VIA_via1_7
* cell instance $16439 r0 *1 54.435,63.77
X$16439 1358 VIA_via2_5
* cell instance $16440 r0 *1 32.015,93.03
X$16440 1358 VIA_via1_7
* cell instance $16441 r0 *1 32.015,92.89
X$16441 1358 VIA_via2_5
* cell instance $16442 r0 *1 56.525,86.17
X$16442 1358 VIA_via1_7
* cell instance $16443 r0 *1 56.525,86.17
X$16443 1358 VIA_via2_5
* cell instance $16444 r0 *1 56.655,86.17
X$16444 1358 VIA_via3_2
* cell instance $16445 r0 *1 56.655,86.31
X$16445 1358 VIA_via4_0
* cell instance $16446 r0 *1 56.655,86.31
X$16446 1358 VIA_via5_0
* cell instance $16447 r0 *1 8.455,64.05
X$16447 1358 VIA_via2_5
* cell instance $16448 r0 *1 8.455,65.31
X$16448 1358 VIA_via2_5
* cell instance $16449 r0 *1 9.025,82.25
X$16449 1358 VIA_via2_5
* cell instance $16450 r0 *1 9.025,94.29
X$16450 1358 VIA_via2_5
* cell instance $16451 r0 *1 17.385,92.61
X$16451 1358 VIA_via2_5
* cell instance $16452 r0 *1 23.655,92.47
X$16452 1358 VIA_via2_5
* cell instance $16453 r0 *1 23.655,92.89
X$16453 1358 VIA_via2_5
* cell instance $16454 r0 *1 50.445,92.75
X$16454 1358 VIA_via2_5
* cell instance $16455 r0 *1 50.445,93.73
X$16455 1358 VIA_via2_5
* cell instance $16456 r0 *1 39.045,93.73
X$16456 1358 VIA_via2_5
* cell instance $16457 r0 *1 38.475,92.89
X$16457 1358 VIA_via2_5
* cell instance $16458 r0 *1 38.475,94.29
X$16458 1358 VIA_via2_5
* cell instance $16459 r0 *1 50.445,93.17
X$16459 1358 VIA_via1_4
* cell instance $16460 r0 *1 42.655,53.69
X$16460 1358 VIA_via1_4
* cell instance $16461 r0 *1 42.655,53.69
X$16461 1358 VIA_via2_5
* cell instance $16462 r0 *1 42.275,54.25
X$16462 1358 VIA_via1_4
* cell instance $16463 r0 *1 42.275,54.25
X$16463 1358 VIA_via2_5
* cell instance $16464 r0 *1 42.375,54.25
X$16464 1358 VIA_via3_2
* cell instance $16465 r0 *1 6.555,65.17
X$16465 1358 VIA_via1_4
* cell instance $16466 r0 *1 6.555,65.31
X$16466 1358 VIA_via2_5
* cell instance $16467 r0 *1 5.415,81.97
X$16467 1358 VIA_via1_4
* cell instance $16468 r0 *1 5.415,81.97
X$16468 1358 VIA_via2_5
* cell instance $16469 r0 *1 8.455,94.43
X$16469 1358 VIA_via1_4
* cell instance $16470 r0 *1 8.455,94.29
X$16470 1358 VIA_via2_5
* cell instance $16471 r0 *1 66.215,52.43
X$16471 1358 VIA_via1_4
* cell instance $16472 r0 *1 66.215,52.43
X$16472 1358 VIA_via2_5
* cell instance $16473 r0 *1 39.045,94.43
X$16473 1358 VIA_via1_4
* cell instance $16474 r0 *1 39.045,94.29
X$16474 1358 VIA_via2_5
* cell instance $16475 r0 *1 17.175,94.43
X$16475 1358 VIA_via4_0
* cell instance $16476 r0 *1 56.655,63.91
X$16476 1358 VIA_via4_0
* cell instance $16477 r0 *1 56.655,63.77
X$16477 1358 VIA_via3_2
* cell instance $16478 r0 *1 56.655,63.91
X$16478 1358 VIA_via5_0
* cell instance $16479 r0 *1 65.335,53.55
X$16479 1358 VIA_via4_0
* cell instance $16480 r0 *1 9.335,94.29
X$16480 1358 VIA_via3_2
* cell instance $16481 r0 *1 9.335,94.43
X$16481 1358 VIA_via4_0
* cell instance $16482 r0 *1 65.335,52.43
X$16482 1358 VIA_via3_2
* cell instance $16483 r0 *1 17.175,92.61
X$16483 1358 VIA_via3_2
* cell instance $16484 r0 *1 56.375,92.75
X$16484 1358 VIA_via3_2
* cell instance $16485 r0 *1 55.535,63.77
X$16485 1358 VIA_via3_2
* cell instance $16486 r0 *1 42.375,64.05
X$16486 1358 VIA_via3_2
* cell instance $16487 r0 *1 55.535,53.69
X$16487 1358 VIA_via3_2
* cell instance $16488 r0 *1 55.535,53.55
X$16488 1358 VIA_via4_0
* cell instance $16489 r0 *1 66.025,52.01
X$16489 1359 VIA_via1_7
* cell instance $16490 r0 *1 66.025,52.01
X$16490 1359 VIA_via2_5
* cell instance $16491 r0 *1 64.505,52.01
X$16491 1359 VIA_via2_5
* cell instance $16492 r0 *1 64.505,51.17
X$16492 1359 VIA_via1_4
* cell instance $16493 r0 *1 1.805,52.99
X$16493 1360 VIA_via1_7
* cell instance $16494 r0 *1 1.805,52.99
X$16494 1360 VIA_via2_5
* cell instance $16495 r0 *1 1.775,52.99
X$16495 1360 VIA_via3_2
* cell instance $16496 r0 *1 1.775,53.27
X$16496 1360 VIA_via4_0
* cell instance $16497 r0 *1 7.695,55.65
X$16497 1361 VIA_via2_5
* cell instance $16498 r0 *1 13.205,55.65
X$16498 1361 VIA_via2_5
* cell instance $16499 r0 *1 14.915,55.65
X$16499 1361 VIA_via2_5
* cell instance $16500 r0 *1 5.605,54.67
X$16500 1361 VIA_via2_5
* cell instance $16501 r0 *1 24.795,55.65
X$16501 1361 VIA_via2_5
* cell instance $16502 r0 *1 26.505,55.65
X$16502 1361 VIA_via2_5
* cell instance $16503 r0 *1 4.465,54.67
X$16503 1361 VIA_via2_5
* cell instance $16504 r0 *1 5.605,55.65
X$16504 1361 VIA_via2_5
* cell instance $16505 r0 *1 29.165,56.35
X$16505 1361 VIA_via2_5
* cell instance $16506 r0 *1 29.165,55.65
X$16506 1361 VIA_via2_5
* cell instance $16507 r0 *1 33.915,56.49
X$16507 1361 VIA_via2_5
* cell instance $16508 r0 *1 24.795,58.03
X$16508 1361 VIA_via1_4
* cell instance $16509 r0 *1 29.165,53.97
X$16509 1361 VIA_via1_4
* cell instance $16510 r0 *1 33.915,56.77
X$16510 1361 VIA_via1_4
* cell instance $16511 r0 *1 13.205,53.97
X$16511 1361 VIA_via1_4
* cell instance $16512 r0 *1 14.915,55.23
X$16512 1361 VIA_via1_4
* cell instance $16513 r0 *1 7.315,55.65
X$16513 1361 VIA_via1_4
* cell instance $16514 r0 *1 7.315,55.65
X$16514 1361 VIA_via2_5
* cell instance $16515 r0 *1 4.275,53.97
X$16515 1361 VIA_via1_4
* cell instance $16516 r0 *1 7.695,58.03
X$16516 1361 VIA_via1_4
* cell instance $16517 r0 *1 5.605,53.97
X$16517 1361 VIA_via1_4
* cell instance $16518 r0 *1 33.915,58.03
X$16518 1361 VIA_via1_4
* cell instance $16519 r0 *1 26.505,55.23
X$16519 1361 VIA_via1_4
* cell instance $16520 r0 *1 5.225,53.83
X$16520 1362 VIA_via2_5
* cell instance $16521 r0 *1 6.935,53.97
X$16521 1362 VIA_via1_4
* cell instance $16522 r0 *1 6.935,53.83
X$16522 1362 VIA_via2_5
* cell instance $16523 r0 *1 3.705,53.97
X$16523 1362 VIA_via1_4
* cell instance $16524 r0 *1 3.705,53.97
X$16524 1362 VIA_via2_5
* cell instance $16525 r0 *1 5.225,51.45
X$16525 1362 VIA_via1_4
* cell instance $16526 r0 *1 11.305,53.55
X$16526 1363 VIA_via1_4
* cell instance $16527 r0 *1 11.875,55.23
X$16527 1363 VIA_via1_4
* cell instance $16528 r0 *1 22.705,53.97
X$16528 1364 VIA_via2_5
* cell instance $16529 r0 *1 22.705,54.95
X$16529 1364 VIA_via1_4
* cell instance $16530 r0 *1 18.525,53.97
X$16530 1364 VIA_via1_4
* cell instance $16531 r0 *1 18.525,53.97
X$16531 1364 VIA_via2_5
* cell instance $16532 r0 *1 17.575,53.97
X$16532 1364 VIA_via1_4
* cell instance $16533 r0 *1 17.575,53.97
X$16533 1364 VIA_via2_5
* cell instance $16534 r0 *1 22.895,55.23
X$16534 1364 VIA_via1_4
* cell instance $16535 r0 *1 19.475,53.41
X$16535 1365 VIA_via2_5
* cell instance $16536 r0 *1 20.995,53.41
X$16536 1365 VIA_via2_5
* cell instance $16537 r0 *1 20.805,53.69
X$16537 1365 VIA_via1_4
* cell instance $16538 r0 *1 19.095,53.97
X$16538 1365 VIA_via1_4
* cell instance $16539 r0 *1 28.025,53.97
X$16539 1366 VIA_via2_5
* cell instance $16540 r0 *1 32.775,53.97
X$16540 1366 VIA_via1_4
* cell instance $16541 r0 *1 32.775,53.97
X$16541 1366 VIA_via2_5
* cell instance $16542 r0 *1 28.595,53.97
X$16542 1366 VIA_via1_4
* cell instance $16543 r0 *1 28.595,53.97
X$16543 1366 VIA_via2_5
* cell instance $16544 r0 *1 28.025,55.23
X$16544 1366 VIA_via1_4
* cell instance $16545 r0 *1 36.575,54.81
X$16545 1367 VIA_via1_7
* cell instance $16546 r0 *1 37.145,53.97
X$16546 1367 VIA_via1_4
* cell instance $16547 r0 *1 37.715,54.53
X$16547 1368 VIA_via2_5
* cell instance $16548 r0 *1 38.095,54.53
X$16548 1368 VIA_via2_5
* cell instance $16549 r0 *1 37.715,53.55
X$16549 1368 VIA_via2_5
* cell instance $16550 r0 *1 36.195,54.67
X$16550 1368 VIA_via2_5
* cell instance $16551 r0 *1 40.375,53.55
X$16551 1368 VIA_via1_4
* cell instance $16552 r0 *1 40.375,53.55
X$16552 1368 VIA_via2_5
* cell instance $16553 r0 *1 37.715,51.17
X$16553 1368 VIA_via1_4
* cell instance $16554 r0 *1 38.475,56.77
X$16554 1368 VIA_via1_4
* cell instance $16555 r0 *1 36.195,55.23
X$16555 1368 VIA_via1_4
* cell instance $16556 r0 *1 16.055,87.43
X$16556 1369 VIA_via1_7
* cell instance $16557 r0 *1 16.055,87.43
X$16557 1369 VIA_via2_5
* cell instance $16558 r0 *1 49.115,90.23
X$16558 1369 VIA_via1_7
* cell instance $16559 r0 *1 7.125,70.63
X$16559 1369 VIA_via1_7
* cell instance $16560 r0 *1 7.125,67.27
X$16560 1369 VIA_via2_5
* cell instance $16561 r0 *1 26.505,87.43
X$16561 1369 VIA_via2_5
* cell instance $16562 r0 *1 12.445,68.25
X$16562 1369 VIA_via2_5
* cell instance $16563 r0 *1 12.445,67.55
X$16563 1369 VIA_via2_5
* cell instance $16564 r0 *1 49.115,88.13
X$16564 1369 VIA_via2_5
* cell instance $16565 r0 *1 7.125,68.25
X$16565 1369 VIA_via2_5
* cell instance $16566 r0 *1 10.735,68.25
X$16566 1369 VIA_via2_5
* cell instance $16567 r0 *1 16.055,86.03
X$16567 1369 VIA_via2_5
* cell instance $16568 r0 *1 51.395,60.97
X$16568 1369 VIA_via2_5
* cell instance $16569 r0 *1 41.515,87.99
X$16569 1369 VIA_via2_5
* cell instance $16570 r0 *1 40.945,64.75
X$16570 1369 VIA_via2_5
* cell instance $16571 r0 *1 25.745,64.75
X$16571 1369 VIA_via2_5
* cell instance $16572 r0 *1 25.745,67.55
X$16572 1369 VIA_via2_5
* cell instance $16573 r0 *1 51.775,83.23
X$16573 1369 VIA_via1_4
* cell instance $16574 r0 *1 51.775,83.23
X$16574 1369 VIA_via2_5
* cell instance $16575 r0 *1 26.885,88.83
X$16575 1369 VIA_via1_4
* cell instance $16576 r0 *1 41.515,87.57
X$16576 1369 VIA_via1_4
* cell instance $16577 r0 *1 41.515,87.43
X$16577 1369 VIA_via2_5
* cell instance $16578 r0 *1 4.845,53.97
X$16578 1369 VIA_via1_4
* cell instance $16579 r0 *1 4.845,53.97
X$16579 1369 VIA_via2_5
* cell instance $16580 r0 *1 10.735,67.97
X$16580 1369 VIA_via1_4
* cell instance $16581 r0 *1 5.035,86.03
X$16581 1369 VIA_via1_4
* cell instance $16582 r0 *1 5.035,86.03
X$16582 1369 VIA_via2_5
* cell instance $16583 r0 *1 40.945,62.37
X$16583 1369 VIA_via1_4
* cell instance $16584 r0 *1 51.205,52.85
X$16584 1369 VIA_via1_4
* cell instance $16585 r0 *1 50.775,62.79
X$16585 1369 VIA_via4_0
* cell instance $16586 r0 *1 6.535,67.27
X$16586 1369 VIA_via3_2
* cell instance $16587 r0 *1 6.535,53.97
X$16587 1369 VIA_via3_2
* cell instance $16588 r0 *1 50.775,88.13
X$16588 1369 VIA_via3_2
* cell instance $16589 r0 *1 50.775,83.23
X$16589 1369 VIA_via3_2
* cell instance $16590 r0 *1 40.975,62.79
X$16590 1369 VIA_via3_2
* cell instance $16591 r0 *1 40.945,62.79
X$16591 1369 VIA_via2_5
* cell instance $16592 r0 *1 40.975,62.79
X$16592 1369 VIA_via4_0
* cell instance $16593 r0 *1 50.775,60.97
X$16593 1369 VIA_via3_2
* cell instance $16594 r0 *1 60.515,66.71
X$16594 1370 VIA_via2_5
* cell instance $16595 r0 *1 51.965,66.71
X$16595 1370 VIA_via2_5
* cell instance $16596 r0 *1 60.515,90.65
X$16596 1370 VIA_via2_5
* cell instance $16597 r0 *1 64.315,90.65
X$16597 1370 VIA_via1_4
* cell instance $16598 r0 *1 64.315,90.65
X$16598 1370 VIA_via2_5
* cell instance $16599 r0 *1 52.155,53.97
X$16599 1370 VIA_via1_4
* cell instance $16600 r0 *1 67.355,52.99
X$16600 1371 VIA_via1_7
* cell instance $16601 r0 *1 67.165,59.57
X$16601 1371 VIA_via1_4
* cell instance $16602 r0 *1 70.205,54.67
X$16602 1372 VIA_via2_5
* cell instance $16603 r0 *1 69.635,54.67
X$16603 1372 VIA_via2_5
* cell instance $16604 r0 *1 72.675,54.67
X$16604 1372 VIA_via2_5
* cell instance $16605 r0 *1 70.395,53.97
X$16605 1372 VIA_via1_4
* cell instance $16606 r0 *1 72.675,54.95
X$16606 1372 VIA_via1_4
* cell instance $16607 r0 *1 69.635,56.77
X$16607 1372 VIA_via1_4
* cell instance $16608 r0 *1 11.875,91.77
X$16608 1373 VIA_via1_7
* cell instance $16609 r0 *1 11.875,91.77
X$16609 1373 VIA_via2_5
* cell instance $16610 r0 *1 68.875,56.63
X$16610 1373 VIA_via1_7
* cell instance $16611 r0 *1 80.845,52.57
X$16611 1373 VIA_via1_7
* cell instance $16612 r0 *1 80.845,52.71
X$16612 1373 VIA_via2_5
* cell instance $16613 r0 *1 56.335,90.23
X$16613 1373 VIA_via1_7
* cell instance $16614 r0 *1 56.335,90.23
X$16614 1373 VIA_via2_5
* cell instance $16615 r0 *1 58.425,56.07
X$16615 1373 VIA_via2_5
* cell instance $16616 r0 *1 57.855,56.07
X$16616 1373 VIA_via2_5
* cell instance $16617 r0 *1 68.875,56.07
X$16617 1373 VIA_via2_5
* cell instance $16618 r0 *1 58.425,53.55
X$16618 1373 VIA_via2_5
* cell instance $16619 r0 *1 42.275,92.89
X$16619 1373 VIA_via2_5
* cell instance $16620 r0 *1 42.275,94.15
X$16620 1373 VIA_via2_5
* cell instance $16621 r0 *1 37.905,93.03
X$16621 1373 VIA_via2_5
* cell instance $16622 r0 *1 37.905,91.77
X$16622 1373 VIA_via2_5
* cell instance $16623 r0 *1 68.875,54.81
X$16623 1373 VIA_via2_5
* cell instance $16624 r0 *1 77.425,52.99
X$16624 1373 VIA_via2_5
* cell instance $16625 r0 *1 77.045,54.67
X$16625 1373 VIA_via2_5
* cell instance $16626 r0 *1 58.235,65.17
X$16626 1373 VIA_via1_4
* cell instance $16627 r0 *1 58.235,65.31
X$16627 1373 VIA_via2_5
* cell instance $16628 r0 *1 58.335,65.31
X$16628 1373 VIA_via3_2
* cell instance $16629 r0 *1 56.145,94.43
X$16629 1373 VIA_via1_4
* cell instance $16630 r0 *1 56.145,94.43
X$16630 1373 VIA_via2_5
* cell instance $16631 r0 *1 20.615,91.63
X$16631 1373 VIA_via1_4
* cell instance $16632 r0 *1 20.615,91.49
X$16632 1373 VIA_via2_5
* cell instance $16633 r0 *1 20.615,91.77
X$16633 1373 VIA_via2_5
* cell instance $16634 r0 *1 28.025,91.63
X$16634 1373 VIA_via1_4
* cell instance $16635 r0 *1 28.025,91.49
X$16635 1373 VIA_via2_5
* cell instance $16636 r0 *1 43.985,53.55
X$16636 1373 VIA_via1_4
* cell instance $16637 r0 *1 43.985,53.55
X$16637 1373 VIA_via2_5
* cell instance $16638 r0 *1 42.275,93.17
X$16638 1373 VIA_via1_4
* cell instance $16639 r0 *1 77.045,53.97
X$16639 1373 VIA_via1_4
* cell instance $16640 r0 *1 58.335,90.23
X$16640 1373 VIA_via3_2
* cell instance $16641 r0 *1 77.425,55.51
X$16641 1374 VIA_via2_5
* cell instance $16642 r0 *1 77.235,53.97
X$16642 1374 VIA_via1_4
* cell instance $16643 r0 *1 76.475,55.51
X$16643 1374 VIA_via1_4
* cell instance $16644 r0 *1 76.475,55.51
X$16644 1374 VIA_via2_5
* cell instance $16645 r0 *1 77.425,55.23
X$16645 1374 VIA_via1_4
* cell instance $16646 r0 *1 80.655,52.99
X$16646 1375 VIA_via1_7
* cell instance $16647 r0 *1 80.845,56.63
X$16647 1375 VIA_via2_5
* cell instance $16648 r0 *1 80.465,56.77
X$16648 1375 VIA_via1_4
* cell instance $16649 r0 *1 80.465,56.77
X$16649 1375 VIA_via2_5
* cell instance $16650 r0 *1 82.745,51.31
X$16650 1376 VIA_via1_4
* cell instance $16651 r0 *1 82.365,53.97
X$16651 1376 VIA_via1_4
* cell instance $16652 r0 *1 85.595,53.55
X$16652 1377 VIA_via2_5
* cell instance $16653 r0 *1 84.455,53.55
X$16653 1377 VIA_via2_5
* cell instance $16654 r0 *1 84.265,54.95
X$16654 1377 VIA_via2_5
* cell instance $16655 r0 *1 81.605,56.77
X$16655 1377 VIA_via1_4
* cell instance $16656 r0 *1 81.795,56.77
X$16656 1377 VIA_via1_4
* cell instance $16657 r0 *1 81.985,54.95
X$16657 1377 VIA_via1_4
* cell instance $16658 r0 *1 81.985,54.95
X$16658 1377 VIA_via2_5
* cell instance $16659 r0 *1 85.595,52.5
X$16659 1377 VIA_via1_4
* cell instance $16660 r0 *1 91.105,53.69
X$16660 1378 VIA_via1_7
* cell instance $16661 r0 *1 90.535,55.23
X$16661 1378 VIA_via1_4
* cell instance $16662 r0 *1 91.675,52.99
X$16662 1379 VIA_via1_7
* cell instance $16663 r0 *1 91.485,54.11
X$16663 1379 VIA_via2_5
* cell instance $16664 r0 *1 91.105,53.97
X$16664 1379 VIA_via1_4
* cell instance $16665 r0 *1 91.105,54.11
X$16665 1379 VIA_via2_5
* cell instance $16666 r0 *1 93.195,53.41
X$16666 1380 VIA_via1_7
* cell instance $16667 r0 *1 93.575,52.43
X$16667 1380 VIA_via1_4
* cell instance $16668 r0 *1 94.525,53.97
X$16668 1381 VIA_via1_4
* cell instance $16669 r0 *1 94.525,53.83
X$16669 1381 VIA_via2_5
* cell instance $16670 r0 *1 96.415,53.83
X$16670 1381 VIA_via4_0
* cell instance $16671 r0 *1 96.415,53.83
X$16671 1381 VIA_via3_2
* cell instance $16672 r0 *1 95.665,53.41
X$16672 1382 VIA_via1_7
* cell instance $16673 r0 *1 95.665,53.27
X$16673 1382 VIA_via2_5
* cell instance $16674 r0 *1 96.975,53.27
X$16674 1382 VIA_via4_0
* cell instance $16675 r0 *1 96.975,53.27
X$16675 1382 VIA_via3_2
* cell instance $16676 r0 *1 13.775,88.97
X$16676 1383 VIA_via1_7
* cell instance $16677 r0 *1 13.775,89.11
X$16677 1383 VIA_via2_5
* cell instance $16678 r0 *1 13.815,89.11
X$16678 1383 VIA_via3_2
* cell instance $16679 r0 *1 5.795,88.97
X$16679 1383 VIA_via1_7
* cell instance $16680 r0 *1 39.805,87.43
X$16680 1383 VIA_via1_7
* cell instance $16681 r0 *1 39.805,87.29
X$16681 1383 VIA_via2_5
* cell instance $16682 r0 *1 50.065,84.63
X$16682 1383 VIA_via1_7
* cell instance $16683 r0 *1 50.065,84.63
X$16683 1383 VIA_via2_5
* cell instance $16684 r0 *1 3.515,53.83
X$16684 1383 VIA_via1_7
* cell instance $16685 r0 *1 3.515,53.83
X$16685 1383 VIA_via2_5
* cell instance $16686 r0 *1 4.845,77.91
X$16686 1383 VIA_via2_5
* cell instance $16687 r0 *1 4.275,77.91
X$16687 1383 VIA_via2_5
* cell instance $16688 r0 *1 4.465,88.27
X$16688 1383 VIA_via2_5
* cell instance $16689 r0 *1 5.795,88.27
X$16689 1383 VIA_via2_5
* cell instance $16690 r0 *1 5.795,89.53
X$16690 1383 VIA_via2_5
* cell instance $16691 r0 *1 13.775,89.53
X$16691 1383 VIA_via2_5
* cell instance $16692 r0 *1 50.065,87.29
X$16692 1383 VIA_via2_5
* cell instance $16693 r0 *1 49.495,87.85
X$16693 1383 VIA_via2_5
* cell instance $16694 r0 *1 49.495,88.83
X$16694 1383 VIA_via1_4
* cell instance $16695 r0 *1 42.085,60.83
X$16695 1383 VIA_via1_4
* cell instance $16696 r0 *1 26.125,86.03
X$16696 1383 VIA_via1_4
* cell instance $16697 r0 *1 26.125,86.03
X$16697 1383 VIA_via2_5
* cell instance $16698 r0 *1 5.225,69.23
X$16698 1383 VIA_via1_4
* cell instance $16699 r0 *1 5.225,69.23
X$16699 1383 VIA_via2_5
* cell instance $16700 r0 *1 7.695,69.23
X$16700 1383 VIA_via1_4
* cell instance $16701 r0 *1 7.695,69.09
X$16701 1383 VIA_via2_5
* cell instance $16702 r0 *1 49.495,52.85
X$16702 1383 VIA_via1_4
* cell instance $16703 r0 *1 49.495,52.85
X$16703 1383 VIA_via2_5
* cell instance $16704 r0 *1 43.495,53.83
X$16704 1383 VIA_via4_0
* cell instance $16705 r0 *1 42.095,53.83
X$16705 1383 VIA_via4_0
* cell instance $16706 r0 *1 13.815,88.83
X$16706 1383 VIA_via4_0
* cell instance $16707 r0 *1 43.495,54.39
X$16707 1383 VIA_via4_0
* cell instance $16708 r0 *1 49.655,54.39
X$16708 1383 VIA_via4_0
* cell instance $16709 r0 *1 25.855,88.83
X$16709 1383 VIA_via4_0
* cell instance $16710 r0 *1 49.655,84.63
X$16710 1383 VIA_via3_2
* cell instance $16711 r0 *1 25.855,86.03
X$16711 1383 VIA_via3_2
* cell instance $16712 r0 *1 25.855,87.01
X$16712 1383 VIA_via3_2
* cell instance $16713 r0 *1 42.095,60.27
X$16713 1383 VIA_via3_2
* cell instance $16714 r0 *1 42.085,60.27
X$16714 1383 VIA_via2_5
* cell instance $16715 r0 *1 49.655,52.85
X$16715 1383 VIA_via3_2
* cell instance $16716 r0 *1 4.015,53.83
X$16716 1383 VIA_via3_2
* cell instance $16717 r0 *1 4.015,53.83
X$16717 1383 VIA_via4_0
* cell instance $16718 r0 *1 89.205,51.45
X$16718 1384 VIA_via1_7
* cell instance $16719 r0 *1 89.205,52.85
X$16719 1384 VIA_via2_5
* cell instance $16720 r0 *1 96.045,52.85
X$16720 1384 VIA_via2_5
* cell instance $16721 r0 *1 96.045,53.97
X$16721 1384 VIA_via1_4
* cell instance $16722 r0 *1 9.785,53.41
X$16722 1385 VIA_via1_7
* cell instance $16723 r0 *1 9.785,52.43
X$16723 1385 VIA_via1_4
* cell instance $16724 r0 *1 93.955,53.69
X$16724 1386 VIA_via2_5
* cell instance $16725 r0 *1 93.955,53.97
X$16725 1386 VIA_via1_4
* cell instance $16726 r0 *1 89.395,53.69
X$16726 1386 VIA_via1_4
* cell instance $16727 r0 *1 89.395,53.69
X$16727 1386 VIA_via2_5
* cell instance $16728 r0 *1 15.105,52.85
X$16728 1387 VIA_via2_5
* cell instance $16729 r0 *1 12.635,53.97
X$16729 1387 VIA_via1_4
* cell instance $16730 r0 *1 12.635,53.83
X$16730 1387 VIA_via2_5
* cell instance $16731 r0 *1 16.055,52.85
X$16731 1387 VIA_via1_4
* cell instance $16732 r0 *1 16.055,52.85
X$16732 1387 VIA_via2_5
* cell instance $16733 r0 *1 15.105,53.97
X$16733 1387 VIA_via1_4
* cell instance $16734 r0 *1 15.105,53.83
X$16734 1387 VIA_via2_5
* cell instance $16735 r0 *1 89.585,53.97
X$16735 1388 VIA_via1_4
* cell instance $16736 r0 *1 89.585,53.83
X$16736 1388 VIA_via2_5
* cell instance $16737 r0 *1 84.835,53.83
X$16737 1388 VIA_via1_4
* cell instance $16738 r0 *1 84.835,53.83
X$16738 1388 VIA_via2_5
* cell instance $16739 r0 *1 19.095,53.69
X$16739 1389 VIA_via1_7
* cell instance $16740 r0 *1 19.095,53.69
X$16740 1389 VIA_via2_5
* cell instance $16741 r0 *1 20.615,53.69
X$16741 1389 VIA_via2_5
* cell instance $16742 r0 *1 20.425,55.23
X$16742 1389 VIA_via1_4
* cell instance $16743 r0 *1 79.325,53.69
X$16743 1390 VIA_via2_5
* cell instance $16744 r0 *1 79.325,53.97
X$16744 1390 VIA_via1_4
* cell instance $16745 r0 *1 82.935,53.69
X$16745 1390 VIA_via1_4
* cell instance $16746 r0 *1 82.935,53.69
X$16746 1390 VIA_via2_5
* cell instance $16747 r0 *1 81.985,52.99
X$16747 1391 VIA_via1_7
* cell instance $16748 r0 *1 81.985,52.99
X$16748 1391 VIA_via2_5
* cell instance $16749 r0 *1 85.215,54.39
X$16749 1391 VIA_via2_5
* cell instance $16750 r0 *1 83.315,54.39
X$16750 1391 VIA_via2_5
* cell instance $16751 r0 *1 83.315,52.99
X$16751 1391 VIA_via2_5
* cell instance $16752 r0 *1 85.215,55.23
X$16752 1391 VIA_via1_4
* cell instance $16753 r0 *1 75.905,66.01
X$16753 1392 VIA_via1_7
* cell instance $16754 r0 *1 75.905,66.01
X$16754 1392 VIA_via2_5
* cell instance $16755 r0 *1 75.905,66.85
X$16755 1392 VIA_via1_4
* cell instance $16756 r0 *1 75.905,66.85
X$16756 1392 VIA_via2_5
* cell instance $16757 r0 *1 73.245,66.01
X$16757 1392 VIA_via2_5
* cell instance $16758 r0 *1 67.735,59.99
X$16758 1392 VIA_via2_5
* cell instance $16759 r0 *1 62.605,66.43
X$16759 1392 VIA_via2_5
* cell instance $16760 r0 *1 68.875,66.43
X$16760 1392 VIA_via2_5
* cell instance $16761 r0 *1 82.175,53.55
X$16761 1392 VIA_via2_5
* cell instance $16762 r0 *1 80.275,67.97
X$16762 1392 VIA_via2_5
* cell instance $16763 r0 *1 76.285,60.55
X$16763 1392 VIA_via2_5
* cell instance $16764 r0 *1 76.285,59.99
X$16764 1392 VIA_via2_5
* cell instance $16765 r0 *1 82.745,59.99
X$16765 1392 VIA_via2_5
* cell instance $16766 r0 *1 82.745,53.55
X$16766 1392 VIA_via2_5
* cell instance $16767 r0 *1 80.085,66.85
X$16767 1392 VIA_via2_5
* cell instance $16768 r0 *1 52.535,66.43
X$16768 1392 VIA_via1_4
* cell instance $16769 r0 *1 52.535,66.43
X$16769 1392 VIA_via2_5
* cell instance $16770 r0 *1 69.065,65.17
X$16770 1392 VIA_via1_4
* cell instance $16771 r0 *1 62.605,67.97
X$16771 1392 VIA_via1_4
* cell instance $16772 r0 *1 73.245,66.43
X$16772 1392 VIA_via1_4
* cell instance $16773 r0 *1 73.245,66.43
X$16773 1392 VIA_via2_5
* cell instance $16774 r0 *1 89.015,67.97
X$16774 1392 VIA_via1_4
* cell instance $16775 r0 *1 89.015,67.97
X$16775 1392 VIA_via2_5
* cell instance $16776 r0 *1 80.085,69.23
X$16776 1392 VIA_via1_4
* cell instance $16777 r0 *1 67.735,55.23
X$16777 1392 VIA_via1_4
* cell instance $16778 r0 *1 91.105,58.03
X$16778 1392 VIA_via1_4
* cell instance $16779 r0 *1 91.105,58.03
X$16779 1392 VIA_via2_5
* cell instance $16780 r0 *1 76.285,60.83
X$16780 1392 VIA_via1_4
* cell instance $16781 r0 *1 82.175,52.43
X$16781 1392 VIA_via1_4
* cell instance $16782 r0 *1 90.535,67.97
X$16782 1392 VIA_via3_2
* cell instance $16783 r0 *1 90.535,58.03
X$16783 1392 VIA_via3_2
* cell instance $16784 r0 *1 38.095,53.69
X$16784 1393 VIA_via2_5
* cell instance $16785 r0 *1 37.145,53.69
X$16785 1393 VIA_via1_4
* cell instance $16786 r0 *1 37.145,53.69
X$16786 1393 VIA_via2_5
* cell instance $16787 r0 *1 38.095,53.97
X$16787 1393 VIA_via1_4
* cell instance $16788 r0 *1 48.355,52.71
X$16788 1394 VIA_via1_7
* cell instance $16789 r0 *1 48.355,52.71
X$16789 1394 VIA_via2_5
* cell instance $16790 r0 *1 45.315,52.71
X$16790 1394 VIA_via2_5
* cell instance $16791 r0 *1 45.315,52.43
X$16791 1394 VIA_via1_4
* cell instance $16792 r0 *1 4.275,54.81
X$16792 1395 VIA_via1_7
* cell instance $16793 r0 *1 4.295,54.39
X$16793 1395 VIA_via3_2
* cell instance $16794 r0 *1 4.275,54.39
X$16794 1395 VIA_via2_5
* cell instance $16795 r0 *1 4.295,54.39
X$16795 1395 VIA_via4_0
* cell instance $16796 r0 *1 14.535,53.97
X$16796 1396 VIA_via1_4
* cell instance $16797 r0 *1 18.525,55.37
X$16797 1396 VIA_via1_4
* cell instance $16798 r0 *1 18.525,55.37
X$16798 1396 VIA_via2_5
* cell instance $16799 r0 *1 14.345,55.23
X$16799 1396 VIA_via1_4
* cell instance $16800 r0 *1 14.345,55.37
X$16800 1396 VIA_via2_5
* cell instance $16801 r0 *1 29.735,55.51
X$16801 1397 VIA_via1_7
* cell instance $16802 r0 *1 29.735,55.37
X$16802 1397 VIA_via2_5
* cell instance $16803 r0 *1 3.895,55.23
X$16803 1397 VIA_via1_4
* cell instance $16804 r0 *1 3.895,55.37
X$16804 1397 VIA_via2_5
* cell instance $16805 r0 *1 18.905,53.97
X$16805 1398 VIA_via1_4
* cell instance $16806 r0 *1 18.525,54.25
X$16806 1398 VIA_via1_4
* cell instance $16807 r0 *1 23.845,59.57
X$16807 1399 VIA_via2_5
* cell instance $16808 r0 *1 21.565,59.57
X$16808 1399 VIA_via2_5
* cell instance $16809 r0 *1 21.565,60.83
X$16809 1399 VIA_via2_5
* cell instance $16810 r0 *1 17.765,60.83
X$16810 1399 VIA_via2_5
* cell instance $16811 r0 *1 17.005,60.83
X$16811 1399 VIA_via2_5
* cell instance $16812 r0 *1 25.935,59.57
X$16812 1399 VIA_via1_4
* cell instance $16813 r0 *1 25.935,59.57
X$16813 1399 VIA_via2_5
* cell instance $16814 r0 *1 22.515,53.97
X$16814 1399 VIA_via1_4
* cell instance $16815 r0 *1 17.005,62.37
X$16815 1399 VIA_via1_4
* cell instance $16816 r0 *1 22.135,59.57
X$16816 1399 VIA_via1_4
* cell instance $16817 r0 *1 22.135,59.57
X$16817 1399 VIA_via2_5
* cell instance $16818 r0 *1 24.415,56.77
X$16818 1399 VIA_via1_4
* cell instance $16819 r0 *1 17.955,58.03
X$16819 1399 VIA_via1_4
* cell instance $16820 r0 *1 21.185,55.23
X$16820 1399 VIA_via1_4
* cell instance $16821 r0 *1 18.715,60.83
X$16821 1399 VIA_via1_4
* cell instance $16822 r0 *1 18.715,60.83
X$16822 1399 VIA_via2_5
* cell instance $16823 r0 *1 21.565,59.85
X$16823 1399 VIA_via1_4
* cell instance $16824 r0 *1 22.325,52.71
X$16824 1400 VIA_via1_7
* cell instance $16825 r0 *1 21.755,53.97
X$16825 1400 VIA_via1_4
* cell instance $16826 r0 *1 28.215,55.23
X$16826 1401 VIA_via2_5
* cell instance $16827 r0 *1 28.215,54.25
X$16827 1401 VIA_via1_4
* cell instance $16828 r0 *1 27.455,55.23
X$16828 1401 VIA_via1_4
* cell instance $16829 r0 *1 27.455,55.23
X$16829 1401 VIA_via2_5
* cell instance $16830 r0 *1 25.935,55.23
X$16830 1401 VIA_via1_4
* cell instance $16831 r0 *1 25.935,55.23
X$16831 1401 VIA_via2_5
* cell instance $16832 r0 *1 29.545,56.21
X$16832 1402 VIA_via1_7
* cell instance $16833 r0 *1 29.355,55.23
X$16833 1402 VIA_via1_4
* cell instance $16834 r0 *1 18.905,88.97
X$16834 1403 VIA_via1_7
* cell instance $16835 r0 *1 9.405,87.43
X$16835 1403 VIA_via1_7
* cell instance $16836 r0 *1 9.975,74.97
X$16836 1403 VIA_via1_7
* cell instance $16837 r0 *1 9.975,74.97
X$16837 1403 VIA_via2_5
* cell instance $16838 r0 *1 35.625,90.23
X$16838 1403 VIA_via1_7
* cell instance $16839 r0 *1 12.635,67.83
X$16839 1403 VIA_via1_7
* cell instance $16840 r0 *1 12.635,67.83
X$16840 1403 VIA_via2_5
* cell instance $16841 r0 *1 14.155,55.37
X$16841 1403 VIA_via1_7
* cell instance $16842 r0 *1 29.925,88.27
X$16842 1403 VIA_via2_5
* cell instance $16843 r0 *1 29.925,89.53
X$16843 1403 VIA_via2_5
* cell instance $16844 r0 *1 31.255,88.27
X$16844 1403 VIA_via2_5
* cell instance $16845 r0 *1 31.255,89.39
X$16845 1403 VIA_via2_5
* cell instance $16846 r0 *1 35.815,89.11
X$16846 1403 VIA_via2_5
* cell instance $16847 r0 *1 47.025,89.11
X$16847 1403 VIA_via2_5
* cell instance $16848 r0 *1 9.405,74.97
X$16848 1403 VIA_via2_5
* cell instance $16849 r0 *1 9.405,87.15
X$16849 1403 VIA_via2_5
* cell instance $16850 r0 *1 18.905,89.53
X$16850 1403 VIA_via2_5
* cell instance $16851 r0 *1 18.905,87.15
X$16851 1403 VIA_via2_5
* cell instance $16852 r0 *1 47.025,55.51
X$16852 1403 VIA_via2_5
* cell instance $16853 r0 *1 14.155,56.49
X$16853 1403 VIA_via2_5
* cell instance $16854 r0 *1 14.095,56.49
X$16854 1403 VIA_via3_2
* cell instance $16855 r0 *1 47.025,56.77
X$16855 1403 VIA_via1_4
* cell instance $16856 r0 *1 47.025,56.63
X$16856 1403 VIA_via2_5
* cell instance $16857 r0 *1 47.595,84.77
X$16857 1403 VIA_via1_4
* cell instance $16858 r0 *1 47.595,84.77
X$16858 1403 VIA_via2_5
* cell instance $16859 r0 *1 47.695,84.77
X$16859 1403 VIA_via3_2
* cell instance $16860 r0 *1 29.545,86.03
X$16860 1403 VIA_via1_4
* cell instance $16861 r0 *1 47.405,88.83
X$16861 1403 VIA_via1_4
* cell instance $16862 r0 *1 47.215,54.25
X$16862 1403 VIA_via1_4
* cell instance $16863 r0 *1 14.095,55.51
X$16863 1403 VIA_via4_0
* cell instance $16864 r0 *1 46.855,55.51
X$16864 1403 VIA_via3_2
* cell instance $16865 r0 *1 46.855,55.51
X$16865 1403 VIA_via4_0
* cell instance $16866 r0 *1 47.695,56.63
X$16866 1403 VIA_via3_2
* cell instance $16867 r0 *1 14.095,67.83
X$16867 1403 VIA_via3_2
* cell instance $16868 r0 *1 49.685,54.95
X$16868 1404 VIA_via2_5
* cell instance $16869 r0 *1 51.015,54.95
X$16869 1404 VIA_via2_5
* cell instance $16870 r0 *1 51.015,60.41
X$16870 1404 VIA_via2_5
* cell instance $16871 r0 *1 45.315,60.83
X$16871 1404 VIA_via2_5
* cell instance $16872 r0 *1 42.465,60.83
X$16872 1404 VIA_via2_5
* cell instance $16873 r0 *1 46.075,60.83
X$16873 1404 VIA_via2_5
* cell instance $16874 r0 *1 45.125,56.77
X$16874 1404 VIA_via1_4
* cell instance $16875 r0 *1 40.375,60.83
X$16875 1404 VIA_via1_4
* cell instance $16876 r0 *1 40.375,60.83
X$16876 1404 VIA_via2_5
* cell instance $16877 r0 *1 46.265,59.57
X$16877 1404 VIA_via1_4
* cell instance $16878 r0 *1 47.215,60.83
X$16878 1404 VIA_via1_4
* cell instance $16879 r0 *1 47.215,60.83
X$16879 1404 VIA_via2_5
* cell instance $16880 r0 *1 47.595,60.41
X$16880 1404 VIA_via1_7
* cell instance $16881 r0 *1 47.595,60.41
X$16881 1404 VIA_via2_5
* cell instance $16882 r0 *1 42.275,63.63
X$16882 1404 VIA_via1_4
* cell instance $16883 r0 *1 46.265,62.37
X$16883 1404 VIA_via1_4
* cell instance $16884 r0 *1 51.015,59.57
X$16884 1404 VIA_via1_4
* cell instance $16885 r0 *1 51.205,55.23
X$16885 1404 VIA_via1_4
* cell instance $16886 r0 *1 49.685,53.97
X$16886 1404 VIA_via1_4
* cell instance $16887 r0 *1 51.205,54.67
X$16887 1405 VIA_via2_5
* cell instance $16888 r0 *1 53.105,54.67
X$16888 1405 VIA_via2_5
* cell instance $16889 r0 *1 47.215,54.67
X$16889 1405 VIA_via2_5
* cell instance $16890 r0 *1 47.215,56.77
X$16890 1405 VIA_via1_4
* cell instance $16891 r0 *1 51.205,54.25
X$16891 1405 VIA_via1_4
* cell instance $16892 r0 *1 53.105,55.23
X$16892 1405 VIA_via1_4
* cell instance $16893 r0 *1 52.345,63.77
X$16893 1406 VIA_via1_7
* cell instance $16894 r0 *1 2.375,83.37
X$16894 1406 VIA_via1_7
* cell instance $16895 r0 *1 38.855,93.03
X$16895 1406 VIA_via1_7
* cell instance $16896 r0 *1 29.545,93.03
X$16896 1406 VIA_via1_7
* cell instance $16897 r0 *1 48.735,93.03
X$16897 1406 VIA_via1_7
* cell instance $16898 r0 *1 48.735,92.89
X$16898 1406 VIA_via2_5
* cell instance $16899 r0 *1 48.815,92.89
X$16899 1406 VIA_via3_2
* cell instance $16900 r0 *1 55.955,87.43
X$16900 1406 VIA_via1_7
* cell instance $16901 r0 *1 55.955,87.43
X$16901 1406 VIA_via2_5
* cell instance $16902 r0 *1 56.095,87.43
X$16902 1406 VIA_via3_2
* cell instance $16903 r0 *1 56.095,87.43
X$16903 1406 VIA_via4_0
* cell instance $16904 r0 *1 56.935,87.43
X$16904 1406 VIA_via5_0
* cell instance $16905 r0 *1 56.935,64.19
X$16905 1406 VIA_via5_0
* cell instance $16906 r0 *1 29.545,92.75
X$16906 1406 VIA_via2_5
* cell instance $16907 r0 *1 8.455,63.63
X$16907 1406 VIA_via2_5
* cell instance $16908 r0 *1 2.375,83.79
X$16908 1406 VIA_via2_5
* cell instance $16909 r0 *1 9.975,83.79
X$16909 1406 VIA_via2_5
* cell instance $16910 r0 *1 9.975,91.35
X$16910 1406 VIA_via2_5
* cell instance $16911 r0 *1 10.165,91.77
X$16911 1406 VIA_via2_5
* cell instance $16912 r0 *1 8.455,91.35
X$16912 1406 VIA_via2_5
* cell instance $16913 r0 *1 16.055,91.91
X$16913 1406 VIA_via2_5
* cell instance $16914 r0 *1 56.335,64.19
X$16914 1406 VIA_via2_5
* cell instance $16915 r0 *1 52.535,64.19
X$16915 1406 VIA_via2_5
* cell instance $16916 r0 *1 56.335,54.95
X$16916 1406 VIA_via2_5
* cell instance $16917 r0 *1 55.955,88.13
X$16917 1406 VIA_via2_5
* cell instance $16918 r0 *1 38.855,92.75
X$16918 1406 VIA_via2_5
* cell instance $16919 r0 *1 16.055,93.17
X$16919 1406 VIA_via1_4
* cell instance $16920 r0 *1 16.055,93.31
X$16920 1406 VIA_via2_5
* cell instance $16921 r0 *1 8.645,53.97
X$16921 1406 VIA_via1_4
* cell instance $16922 r0 *1 3.325,63.63
X$16922 1406 VIA_via1_4
* cell instance $16923 r0 *1 3.325,63.63
X$16923 1406 VIA_via2_5
* cell instance $16924 r0 *1 8.455,91.63
X$16924 1406 VIA_via1_4
* cell instance $16925 r0 *1 54.975,64.19
X$16925 1406 VIA_via4_0
* cell instance $16926 r0 *1 54.975,64.19
X$16926 1406 VIA_via3_2
* cell instance $16927 r0 *1 54.695,54.95
X$16927 1406 VIA_via4_0
* cell instance $16928 r0 *1 54.695,54.95
X$16928 1406 VIA_via3_2
* cell instance $16929 r0 *1 54.815,54.95
X$16929 1406 VIA_via2_5
* cell instance $16930 r0 *1 54.815,54.95
X$16930 1406 VIA_via1_4
* cell instance $16931 r0 *1 8.775,54.95
X$16931 1406 VIA_via3_2
* cell instance $16932 r0 *1 8.645,54.95
X$16932 1406 VIA_via2_5
* cell instance $16933 r0 *1 8.775,54.95
X$16933 1406 VIA_via4_0
* cell instance $16934 r0 *1 48.815,88.27
X$16934 1406 VIA_via3_2
* cell instance $16935 r0 *1 58.615,56.35
X$16935 1407 VIA_via1_4
* cell instance $16936 r0 *1 58.615,57.19
X$16936 1407 VIA_via1_7
* cell instance $16937 r0 *1 57.665,55.23
X$16937 1407 VIA_via1_4
* cell instance $16938 r0 *1 58.235,58.03
X$16938 1407 VIA_via1_4
* cell instance $16939 r0 *1 60.325,59.01
X$16939 1408 VIA_via1_7
* cell instance $16940 r0 *1 58.995,55.23
X$16940 1408 VIA_via1_4
* cell instance $16941 r0 *1 60.325,54.81
X$16941 1409 VIA_via1_7
* cell instance $16942 r0 *1 59.945,53.97
X$16942 1409 VIA_via1_4
* cell instance $16943 r0 *1 61.275,57.61
X$16943 1410 VIA_via1_7
* cell instance $16944 r0 *1 60.325,55.79
X$16944 1410 VIA_via2_5
* cell instance $16945 r0 *1 61.275,55.79
X$16945 1410 VIA_via2_5
* cell instance $16946 r0 *1 60.515,55.23
X$16946 1410 VIA_via1_4
* cell instance $16947 r0 *1 66.405,78.61
X$16947 1411 VIA_via1_7
* cell instance $16948 r0 *1 64.315,55.23
X$16948 1411 VIA_via2_5
* cell instance $16949 r0 *1 63.935,55.23
X$16949 1411 VIA_via2_5
* cell instance $16950 r0 *1 65.265,56.77
X$16950 1411 VIA_via2_5
* cell instance $16951 r0 *1 66.405,72.45
X$16951 1411 VIA_via2_5
* cell instance $16952 r0 *1 63.935,53.97
X$16952 1411 VIA_via1_4
* cell instance $16953 r0 *1 64.315,56.77
X$16953 1411 VIA_via1_4
* cell instance $16954 r0 *1 64.315,56.77
X$16954 1411 VIA_via2_5
* cell instance $16955 r0 *1 62.035,53.97
X$16955 1411 VIA_via1_4
* cell instance $16956 r0 *1 62.225,55.23
X$16956 1411 VIA_via1_4
* cell instance $16957 r0 *1 62.225,55.23
X$16957 1411 VIA_via2_5
* cell instance $16958 r0 *1 65.335,72.45
X$16958 1411 VIA_via3_2
* cell instance $16959 r0 *1 65.335,61.39
X$16959 1411 VIA_via3_2
* cell instance $16960 r0 *1 65.265,61.39
X$16960 1411 VIA_via2_5
* cell instance $16961 r0 *1 63.555,57.61
X$16961 1412 VIA_via1_7
* cell instance $16962 r0 *1 62.985,55.23
X$16962 1412 VIA_via1_4
* cell instance $16963 r0 *1 66.785,56.77
X$16963 1413 VIA_via2_5
* cell instance $16964 r0 *1 69.065,56.77
X$16964 1413 VIA_via1_4
* cell instance $16965 r0 *1 69.065,56.77
X$16965 1413 VIA_via2_5
* cell instance $16966 r0 *1 68.685,56.77
X$16966 1413 VIA_via1_4
* cell instance $16967 r0 *1 68.685,56.77
X$16967 1413 VIA_via2_5
* cell instance $16968 r0 *1 67.165,55.23
X$16968 1413 VIA_via1_4
* cell instance $16969 r0 *1 70.775,54.39
X$16969 1414 VIA_via1_7
* cell instance $16970 r0 *1 70.395,55.23
X$16970 1414 VIA_via1_4
* cell instance $16971 r0 *1 82.365,55.09
X$16971 1415 VIA_via1_4
* cell instance $16972 r0 *1 82.175,53.97
X$16972 1415 VIA_via1_4
* cell instance $16973 r0 *1 82.555,54.25
X$16973 1416 VIA_via2_5
* cell instance $16974 r0 *1 83.695,54.25
X$16974 1416 VIA_via2_5
* cell instance $16975 r0 *1 82.555,55.23
X$16975 1416 VIA_via1_4
* cell instance $16976 r0 *1 82.555,55.23
X$16976 1416 VIA_via2_5
* cell instance $16977 r0 *1 82.935,55.23
X$16977 1416 VIA_via1_4
* cell instance $16978 r0 *1 82.935,55.23
X$16978 1416 VIA_via2_5
* cell instance $16979 r0 *1 81.605,54.25
X$16979 1416 VIA_via1_4
* cell instance $16980 r0 *1 81.605,54.25
X$16980 1416 VIA_via2_5
* cell instance $16981 r0 *1 83.695,53.97
X$16981 1416 VIA_via1_4
* cell instance $16982 r0 *1 82.935,53.97
X$16982 1417 VIA_via1_4
* cell instance $16983 r0 *1 83.125,55.09
X$16983 1417 VIA_via1_4
* cell instance $16984 r0 *1 86.165,54.11
X$16984 1418 VIA_via1_4
* cell instance $16985 r0 *1 86.355,56.77
X$16985 1418 VIA_via1_4
* cell instance $16986 r0 *1 87.495,55.65
X$16986 1419 VIA_via2_5
* cell instance $16987 r0 *1 88.825,55.65
X$16987 1419 VIA_via1_4
* cell instance $16988 r0 *1 88.825,55.65
X$16988 1419 VIA_via2_5
* cell instance $16989 r0 *1 87.495,56.77
X$16989 1419 VIA_via1_4
* cell instance $16990 r0 *1 87.685,56.77
X$16990 1419 VIA_via1_4
* cell instance $16991 r0 *1 89.015,55.23
X$16991 1419 VIA_via1_4
* cell instance $16992 r0 *1 92.815,54.95
X$16992 1420 VIA_via1_4
* cell instance $16993 r0 *1 93.005,53.97
X$16993 1420 VIA_via1_4
* cell instance $16994 r0 *1 93.005,53.97
X$16994 1420 VIA_via2_5
* cell instance $16995 r0 *1 92.245,53.97
X$16995 1420 VIA_via1_4
* cell instance $16996 r0 *1 92.435,53.97
X$16996 1420 VIA_via1_4
* cell instance $16997 r0 *1 92.435,53.97
X$16997 1420 VIA_via2_5
* cell instance $16998 r0 *1 96.995,54.39
X$16998 1421 VIA_via1_7
* cell instance $16999 r0 *1 96.995,54.39
X$16999 1421 VIA_via2_5
* cell instance $17000 r0 *1 97.255,54.95
X$17000 1421 VIA_via4_0
* cell instance $17001 r0 *1 97.255,54.39
X$17001 1421 VIA_via3_2
* cell instance $17002 r0 *1 94.335,54.39
X$17002 1422 VIA_via1_7
* cell instance $17003 r0 *1 94.335,54.39
X$17003 1422 VIA_via2_5
* cell instance $17004 r0 *1 94.735,54.39
X$17004 1422 VIA_via4_0
* cell instance $17005 r0 *1 94.735,54.39
X$17005 1422 VIA_via3_2
* cell instance $17006 r0 *1 7.125,54.11
X$17006 1423 VIA_via2_5
* cell instance $17007 r0 *1 7.125,52.85
X$17007 1423 VIA_via1_4
* cell instance $17008 r0 *1 7.505,53.97
X$17008 1423 VIA_via1_4
* cell instance $17009 r0 *1 7.505,54.11
X$17009 1423 VIA_via2_5
* cell instance $17010 r0 *1 5.035,53.97
X$17010 1423 VIA_via1_4
* cell instance $17011 r0 *1 5.035,54.11
X$17011 1423 VIA_via2_5
* cell instance $17012 r0 *1 7.885,53.97
X$17012 1424 VIA_via1_4
* cell instance $17013 r0 *1 7.885,53.97
X$17013 1424 VIA_via2_5
* cell instance $17014 r0 *1 10.925,53.97
X$17014 1424 VIA_via1_4
* cell instance $17015 r0 *1 10.925,53.97
X$17015 1424 VIA_via2_5
* cell instance $17016 r0 *1 57.215,76.79
X$17016 1425 VIA_via5_0
* cell instance $17017 r0 *1 57.215,65.31
X$17017 1425 VIA_via5_0
* cell instance $17018 r0 *1 32.395,90.65
X$17018 1425 VIA_via2_5
* cell instance $17019 r0 *1 12.065,91.07
X$17019 1425 VIA_via2_5
* cell instance $17020 r0 *1 11.305,90.37
X$17020 1425 VIA_via2_5
* cell instance $17021 r0 *1 11.875,90.37
X$17021 1425 VIA_via2_5
* cell instance $17022 r0 *1 19.665,91.07
X$17022 1425 VIA_via2_5
* cell instance $17023 r0 *1 19.665,90.65
X$17023 1425 VIA_via2_5
* cell instance $17024 r0 *1 53.865,54.67
X$17024 1425 VIA_via2_5
* cell instance $17025 r0 *1 53.855,54.67
X$17025 1425 VIA_via3_2
* cell instance $17026 r0 *1 50.445,91.07
X$17026 1425 VIA_via2_5
* cell instance $17027 r0 *1 55.005,86.03
X$17027 1425 VIA_via1_4
* cell instance $17028 r0 *1 55.005,85.89
X$17028 1425 VIA_via2_5
* cell instance $17029 r0 *1 50.445,91.63
X$17029 1425 VIA_via1_4
* cell instance $17030 r0 *1 19.475,90.37
X$17030 1425 VIA_via1_4
* cell instance $17031 r0 *1 40.375,90.37
X$17031 1425 VIA_via1_4
* cell instance $17032 r0 *1 40.375,90.37
X$17032 1425 VIA_via2_5
* cell instance $17033 r0 *1 40.415,90.37
X$17033 1425 VIA_via3_2
* cell instance $17034 r0 *1 32.395,88.83
X$17034 1425 VIA_via1_4
* cell instance $17035 r0 *1 11.495,55.23
X$17035 1425 VIA_via1_4
* cell instance $17036 r0 *1 11.495,55.09
X$17036 1425 VIA_via2_5
* cell instance $17037 r0 *1 11.115,65.17
X$17037 1425 VIA_via1_4
* cell instance $17038 r0 *1 12.065,90.37
X$17038 1425 VIA_via1_4
* cell instance $17039 r0 *1 11.875,74.83
X$17039 1425 VIA_via1_4
* cell instance $17040 r0 *1 53.865,54.25
X$17040 1425 VIA_via1_4
* cell instance $17041 r0 *1 56.375,76.79
X$17041 1425 VIA_via4_0
* cell instance $17042 r0 *1 53.855,55.23
X$17042 1425 VIA_via4_0
* cell instance $17043 r0 *1 54.695,65.31
X$17043 1425 VIA_via4_0
* cell instance $17044 r0 *1 54.695,65.31
X$17044 1425 VIA_via3_2
* cell instance $17045 r0 *1 54.815,65.31
X$17045 1425 VIA_via2_5
* cell instance $17046 r0 *1 54.815,65.17
X$17046 1425 VIA_via1_4
* cell instance $17047 r0 *1 54.135,65.31
X$17047 1425 VIA_via4_0
* cell instance $17048 r0 *1 40.415,91.63
X$17048 1425 VIA_via4_0
* cell instance $17049 r0 *1 54.695,91.07
X$17049 1425 VIA_via4_0
* cell instance $17050 r0 *1 51.615,91.07
X$17050 1425 VIA_via4_0
* cell instance $17051 r0 *1 51.615,91.07
X$17051 1425 VIA_via3_2
* cell instance $17052 r0 *1 51.615,91.63
X$17052 1425 VIA_via4_0
* cell instance $17053 r0 *1 12.415,55.09
X$17053 1425 VIA_via3_2
* cell instance $17054 r0 *1 12.415,55.23
X$17054 1425 VIA_via4_0
* cell instance $17055 r0 *1 54.695,85.89
X$17055 1425 VIA_via3_2
* cell instance $17056 r0 *1 56.375,85.61
X$17056 1425 VIA_via3_2
* cell instance $17057 r0 *1 29.545,57.05
X$17057 1426 VIA_via2_5
* cell instance $17058 r0 *1 29.495,57.05
X$17058 1426 VIA_via3_2
* cell instance $17059 r0 *1 29.545,59.57
X$17059 1426 VIA_via1_4
* cell instance $17060 r0 *1 29.545,59.57
X$17060 1426 VIA_via2_5
* cell instance $17061 r0 *1 29.495,59.57
X$17061 1426 VIA_via3_2
* cell instance $17062 r0 *1 29.545,56.77
X$17062 1426 VIA_via1_4
* cell instance $17063 r0 *1 12.065,55.09
X$17063 1426 VIA_via1_4
* cell instance $17064 r0 *1 12.065,54.95
X$17064 1426 VIA_via2_5
* cell instance $17065 r0 *1 29.495,54.95
X$17065 1426 VIA_via3_2
* cell instance $17066 r0 *1 13.965,54.39
X$17066 1427 VIA_via1_7
* cell instance $17067 r0 *1 13.965,54.81
X$17067 1427 VIA_via2_5
* cell instance $17068 r0 *1 11.685,54.81
X$17068 1427 VIA_via2_5
* cell instance $17069 r0 *1 11.685,55.23
X$17069 1427 VIA_via1_4
* cell instance $17070 r0 *1 15.485,53.97
X$17070 1428 VIA_via1_4
* cell instance $17071 r0 *1 15.485,53.97
X$17071 1428 VIA_via2_5
* cell instance $17072 r0 *1 13.775,53.97
X$17072 1428 VIA_via1_4
* cell instance $17073 r0 *1 13.775,53.97
X$17073 1428 VIA_via2_5
* cell instance $17074 r0 *1 91.675,54.25
X$17074 1429 VIA_via2_5
* cell instance $17075 r0 *1 91.675,53.97
X$17075 1429 VIA_via1_4
* cell instance $17076 r0 *1 92.815,54.25
X$17076 1429 VIA_via1_4
* cell instance $17077 r0 *1 92.815,54.25
X$17077 1429 VIA_via2_5
* cell instance $17078 r0 *1 15.295,55.09
X$17078 1430 VIA_via1_4
* cell instance $17079 r0 *1 15.295,55.09
X$17079 1430 VIA_via2_5
* cell instance $17080 r0 *1 16.245,55.23
X$17080 1430 VIA_via1_4
* cell instance $17081 r0 *1 16.245,55.09
X$17081 1430 VIA_via2_5
* cell instance $17082 r0 *1 23.275,54.81
X$17082 1431 VIA_via1_7
* cell instance $17083 r0 *1 23.275,54.81
X$17083 1431 VIA_via2_5
* cell instance $17084 r0 *1 19.665,54.81
X$17084 1431 VIA_via2_5
* cell instance $17085 r0 *1 19.665,53.97
X$17085 1431 VIA_via1_4
* cell instance $17086 r0 *1 26.885,54.81
X$17086 1432 VIA_via1_7
* cell instance $17087 r0 *1 26.885,54.81
X$17087 1432 VIA_via2_5
* cell instance $17088 r0 *1 25.935,54.81
X$17088 1432 VIA_via2_5
* cell instance $17089 r0 *1 25.935,53.97
X$17089 1432 VIA_via1_4
* cell instance $17090 r0 *1 90.915,54.81
X$17090 1433 VIA_via2_5
* cell instance $17091 r0 *1 92.055,54.81
X$17091 1433 VIA_via2_5
* cell instance $17092 r0 *1 90.915,54.04
X$17092 1433 VIA_via1_4
* cell instance $17093 r0 *1 92.055,54.11
X$17093 1433 VIA_via1_4
* cell instance $17094 r0 *1 36.385,66.57
X$17094 1434 VIA_via1_7
* cell instance $17095 r0 *1 36.385,66.57
X$17095 1434 VIA_via2_5
* cell instance $17096 r0 *1 48.165,67.83
X$17096 1434 VIA_via1_7
* cell instance $17097 r0 *1 23.845,74.97
X$17097 1434 VIA_via1_7
* cell instance $17098 r0 *1 23.845,74.97
X$17098 1434 VIA_via2_5
* cell instance $17099 r0 *1 25.935,66.57
X$17099 1434 VIA_via1_7
* cell instance $17100 r0 *1 25.935,66.71
X$17100 1434 VIA_via2_5
* cell instance $17101 r0 *1 44.935,58.17
X$17101 1434 VIA_via1_7
* cell instance $17102 r0 *1 44.935,58.17
X$17102 1434 VIA_via2_5
* cell instance $17103 r0 *1 17.385,69.09
X$17103 1434 VIA_via2_5
* cell instance $17104 r0 *1 17.385,66.71
X$17104 1434 VIA_via2_5
* cell instance $17105 r0 *1 17.385,74.97
X$17105 1434 VIA_via2_5
* cell instance $17106 r0 *1 18.715,66.71
X$17106 1434 VIA_via2_5
* cell instance $17107 r0 *1 36.385,67.41
X$17107 1434 VIA_via2_5
* cell instance $17108 r0 *1 48.165,67.41
X$17108 1434 VIA_via2_5
* cell instance $17109 r0 *1 43.795,67.41
X$17109 1434 VIA_via2_5
* cell instance $17110 r0 *1 27.075,54.11
X$17110 1434 VIA_via2_5
* cell instance $17111 r0 *1 26.885,66.71
X$17111 1434 VIA_via2_5
* cell instance $17112 r0 *1 43.605,74.83
X$17112 1434 VIA_via1_4
* cell instance $17113 r0 *1 28.405,53.97
X$17113 1434 VIA_via1_4
* cell instance $17114 r0 *1 28.405,54.11
X$17114 1434 VIA_via2_5
* cell instance $17115 r0 *1 45.885,54.25
X$17115 1434 VIA_via1_4
* cell instance $17116 r0 *1 18.715,62.37
X$17116 1434 VIA_via1_4
* cell instance $17117 r0 *1 16.055,69.23
X$17117 1434 VIA_via1_4
* cell instance $17118 r0 *1 16.055,69.09
X$17118 1434 VIA_via2_5
* cell instance $17119 r0 *1 17.955,77.63
X$17119 1434 VIA_via1_4
* cell instance $17120 r0 *1 46.015,67.41
X$17120 1434 VIA_via3_2
* cell instance $17121 r0 *1 46.015,58.17
X$17121 1434 VIA_via3_2
* cell instance $17122 r0 *1 45.885,58.17
X$17122 1434 VIA_via2_5
* cell instance $17123 r0 *1 89.395,54.81
X$17123 1435 VIA_via1_7
* cell instance $17124 r0 *1 89.395,53.97
X$17124 1435 VIA_via1_4
* cell instance $17125 r0 *1 29.545,54.11
X$17125 1436 VIA_via1_4
* cell instance $17126 r0 *1 29.545,54.11
X$17126 1436 VIA_via2_5
* cell instance $17127 r0 *1 30.495,53.97
X$17127 1436 VIA_via1_4
* cell instance $17128 r0 *1 30.495,54.11
X$17128 1436 VIA_via2_5
* cell instance $17129 r0 *1 38.285,56.21
X$17129 1437 VIA_via1_7
* cell instance $17130 r0 *1 38.285,54.11
X$17130 1437 VIA_via2_5
* cell instance $17131 r0 *1 36.385,53.97
X$17131 1437 VIA_via1_4
* cell instance $17132 r0 *1 36.385,54.11
X$17132 1437 VIA_via2_5
* cell instance $17133 r0 *1 41.325,53.97
X$17133 1438 VIA_via1_4
* cell instance $17134 r0 *1 41.325,53.97
X$17134 1438 VIA_via2_5
* cell instance $17135 r0 *1 36.575,53.97
X$17135 1438 VIA_via1_4
* cell instance $17136 r0 *1 36.575,53.97
X$17136 1438 VIA_via2_5
* cell instance $17137 r0 *1 48.165,56.21
X$17137 1439 VIA_via1_7
* cell instance $17138 r0 *1 48.165,53.97
X$17138 1439 VIA_via2_5
* cell instance $17139 r0 *1 48.925,53.97
X$17139 1439 VIA_via1_4
* cell instance $17140 r0 *1 48.925,53.97
X$17140 1439 VIA_via2_5
* cell instance $17141 r0 *1 55.575,52.71
X$17141 1440 VIA_via1_4
* cell instance $17142 r0 *1 55.575,53.97
X$17142 1440 VIA_via1_4
* cell instance $17143 r0 *1 64.725,53.97
X$17143 1441 VIA_via1_4
* cell instance $17144 r0 *1 64.505,53.97
X$17144 1441 VIA_via1_4
* cell instance $17145 r0 *1 59.945,55.51
X$17145 1442 VIA_via2_5
* cell instance $17146 r0 *1 61.655,59.71
X$17146 1442 VIA_via2_5
* cell instance $17147 r0 *1 64.125,54.67
X$17147 1442 VIA_via2_5
* cell instance $17148 r0 *1 62.415,54.67
X$17148 1442 VIA_via2_5
* cell instance $17149 r0 *1 62.225,55.51
X$17149 1442 VIA_via2_5
* cell instance $17150 r0 *1 64.505,82.95
X$17150 1442 VIA_via1_4
* cell instance $17151 r0 *1 64.505,82.95
X$17151 1442 VIA_via2_5
* cell instance $17152 r0 *1 59.945,55.23
X$17152 1442 VIA_via1_4
* cell instance $17153 r0 *1 59.945,59.57
X$17153 1442 VIA_via1_4
* cell instance $17154 r0 *1 59.945,59.71
X$17154 1442 VIA_via2_5
* cell instance $17155 r0 *1 61.655,58.03
X$17155 1442 VIA_via1_4
* cell instance $17156 r0 *1 64.125,53.97
X$17156 1442 VIA_via1_4
* cell instance $17157 r0 *1 61.415,59.71
X$17157 1442 VIA_via3_2
* cell instance $17158 r0 *1 61.415,82.95
X$17158 1442 VIA_via3_2
* cell instance $17159 r0 *1 62.825,53.97
X$17159 1443 VIA_via1_4
* cell instance $17160 r0 *1 62.605,53.97
X$17160 1443 VIA_via1_4
* cell instance $17161 r0 *1 61.085,58.03
X$17161 1444 VIA_via2_5
* cell instance $17162 r0 *1 61.085,57.75
X$17162 1444 VIA_via2_5
* cell instance $17163 r0 *1 61.845,53.97
X$17163 1444 VIA_via2_5
* cell instance $17164 r0 *1 61.655,57.75
X$17164 1444 VIA_via2_5
* cell instance $17165 r0 *1 63.175,68.95
X$17165 1444 VIA_via2_5
* cell instance $17166 r0 *1 63.745,68.95
X$17166 1444 VIA_via2_5
* cell instance $17167 r0 *1 63.745,76.23
X$17167 1444 VIA_via2_5
* cell instance $17168 r0 *1 63.365,76.23
X$17168 1444 VIA_via2_5
* cell instance $17169 r0 *1 63.365,82.95
X$17169 1444 VIA_via1_4
* cell instance $17170 r0 *1 60.895,58.03
X$17170 1444 VIA_via1_4
* cell instance $17171 r0 *1 63.175,58.03
X$17171 1444 VIA_via1_4
* cell instance $17172 r0 *1 63.175,58.03
X$17172 1444 VIA_via2_5
* cell instance $17173 r0 *1 61.655,56.77
X$17173 1444 VIA_via1_4
* cell instance $17174 r0 *1 62.225,53.97
X$17174 1444 VIA_via1_4
* cell instance $17175 r0 *1 62.225,53.97
X$17175 1444 VIA_via2_5
* cell instance $17176 r0 *1 23.465,57.61
X$17176 1445 VIA_via1_7
* cell instance $17177 r0 *1 23.655,56.77
X$17177 1445 VIA_via1_4
* cell instance $17178 r0 *1 25.745,55.37
X$17178 1446 VIA_via1_7
* cell instance $17179 r0 *1 47.975,65.03
X$17179 1446 VIA_via1_7
* cell instance $17180 r0 *1 22.705,76.23
X$17180 1446 VIA_via1_7
* cell instance $17181 r0 *1 22.705,76.23
X$17181 1446 VIA_via2_5
* cell instance $17182 r0 *1 15.295,74.97
X$17182 1446 VIA_via1_7
* cell instance $17183 r0 *1 46.265,58.17
X$17183 1446 VIA_via1_7
* cell instance $17184 r0 *1 16.435,63.77
X$17184 1446 VIA_via1_7
* cell instance $17185 r0 *1 16.435,63.91
X$17185 1446 VIA_via2_5
* cell instance $17186 r0 *1 15.295,76.23
X$17186 1446 VIA_via2_5
* cell instance $17187 r0 *1 15.295,63.91
X$17187 1446 VIA_via2_5
* cell instance $17188 r0 *1 46.265,58.45
X$17188 1446 VIA_via2_5
* cell instance $17189 r0 *1 47.405,58.45
X$17189 1446 VIA_via2_5
* cell instance $17190 r0 *1 47.975,66.29
X$17190 1446 VIA_via2_5
* cell instance $17191 r0 *1 42.085,66.29
X$17191 1446 VIA_via2_5
* cell instance $17192 r0 *1 27.455,64.89
X$17192 1446 VIA_via2_5
* cell instance $17193 r0 *1 27.455,66.15
X$17193 1446 VIA_via2_5
* cell instance $17194 r0 *1 25.555,64.89
X$17194 1446 VIA_via2_5
* cell instance $17195 r0 *1 25.555,63.91
X$17195 1446 VIA_via2_5
* cell instance $17196 r0 *1 48.165,58.45
X$17196 1446 VIA_via1_4
* cell instance $17197 r0 *1 48.165,58.45
X$17197 1446 VIA_via2_5
* cell instance $17198 r0 *1 27.455,66.43
X$17198 1446 VIA_via1_4
* cell instance $17199 r0 *1 41.895,72.03
X$17199 1446 VIA_via1_4
* cell instance $17200 r0 *1 37.715,66.43
X$17200 1446 VIA_via1_4
* cell instance $17201 r0 *1 37.715,66.29
X$17201 1446 VIA_via2_5
* cell instance $17202 r0 *1 16.055,73.57
X$17202 1446 VIA_via1_4
* cell instance $17203 r0 *1 28.405,55.79
X$17203 1447 VIA_via1_7
* cell instance $17204 r0 *1 27.455,56.77
X$17204 1447 VIA_via1_4
* cell instance $17205 r0 *1 27.835,56.35
X$17205 1448 VIA_via1_4
* cell instance $17206 r0 *1 28.975,58.03
X$17206 1448 VIA_via1_4
* cell instance $17207 r0 *1 28.025,56.77
X$17207 1449 VIA_via1_4
* cell instance $17208 r0 *1 28.025,56.77
X$17208 1449 VIA_via2_5
* cell instance $17209 r0 *1 32.965,56.49
X$17209 1449 VIA_via1_4
* cell instance $17210 r0 *1 32.965,56.49
X$17210 1449 VIA_via2_5
* cell instance $17211 r0 *1 30.685,60.55
X$17211 1450 VIA_via2_5
* cell instance $17212 r0 *1 30.685,61.95
X$17212 1450 VIA_via2_5
* cell instance $17213 r0 *1 31.825,60.55
X$17213 1450 VIA_via1_4
* cell instance $17214 r0 *1 31.825,60.55
X$17214 1450 VIA_via2_5
* cell instance $17215 r0 *1 29.545,62.3
X$17215 1450 VIA_via1_4
* cell instance $17216 r0 *1 29.545,62.23
X$17216 1450 VIA_via2_5
* cell instance $17217 r0 *1 31.445,55.23
X$17217 1450 VIA_via1_4
* cell instance $17218 r0 *1 30.875,62.37
X$17218 1450 VIA_via1_4
* cell instance $17219 r0 *1 33.345,58.03
X$17219 1451 VIA_via1_4
* cell instance $17220 r0 *1 32.585,56.77
X$17220 1451 VIA_via1_4
* cell instance $17221 r0 *1 32.965,57.75
X$17221 1451 VIA_via1_4
* cell instance $17222 r0 *1 33.345,55.65
X$17222 1452 VIA_via2_5
* cell instance $17223 r0 *1 33.345,56.77
X$17223 1452 VIA_via1_4
* cell instance $17224 r0 *1 33.345,56.63
X$17224 1452 VIA_via2_5
* cell instance $17225 r0 *1 32.015,56.77
X$17225 1452 VIA_via1_4
* cell instance $17226 r0 *1 32.015,56.63
X$17226 1452 VIA_via2_5
* cell instance $17227 r0 *1 36.005,55.51
X$17227 1452 VIA_via1_4
* cell instance $17228 r0 *1 36.005,55.51
X$17228 1452 VIA_via2_5
* cell instance $17229 r0 *1 34.295,56.21
X$17229 1453 VIA_via1_7
* cell instance $17230 r0 *1 33.725,55.23
X$17230 1453 VIA_via1_4
* cell instance $17231 r0 *1 46.265,66.57
X$17231 1454 VIA_via1_7
* cell instance $17232 r0 *1 46.265,66.57
X$17232 1454 VIA_via2_5
* cell instance $17233 r0 *1 42.085,59.43
X$17233 1454 VIA_via1_7
* cell instance $17234 r0 *1 42.085,59.43
X$17234 1454 VIA_via2_5
* cell instance $17235 r0 *1 74.765,70.63
X$17235 1454 VIA_via1_7
* cell instance $17236 r0 *1 20.615,71.05
X$17236 1454 VIA_via2_5
* cell instance $17237 r0 *1 53.295,72.03
X$17237 1454 VIA_via2_5
* cell instance $17238 r0 *1 53.295,71.05
X$17238 1454 VIA_via2_5
* cell instance $17239 r0 *1 64.505,70.07
X$17239 1454 VIA_via2_5
* cell instance $17240 r0 *1 64.505,71.89
X$17240 1454 VIA_via2_5
* cell instance $17241 r0 *1 74.765,70.07
X$17241 1454 VIA_via2_5
* cell instance $17242 r0 *1 43.035,59.43
X$17242 1454 VIA_via2_5
* cell instance $17243 r0 *1 35.625,71.05
X$17243 1454 VIA_via2_5
* cell instance $17244 r0 *1 40.565,71.05
X$17244 1454 VIA_via2_5
* cell instance $17245 r0 *1 25.175,71.05
X$17245 1454 VIA_via2_5
* cell instance $17246 r0 *1 62.795,72.03
X$17246 1454 VIA_via1_4
* cell instance $17247 r0 *1 62.795,71.89
X$17247 1454 VIA_via2_5
* cell instance $17248 r0 *1 52.725,72.03
X$17248 1454 VIA_via1_4
* cell instance $17249 r0 *1 52.725,72.03
X$17249 1454 VIA_via2_5
* cell instance $17250 r0 *1 43.225,51.45
X$17250 1454 VIA_via1_4
* cell instance $17251 r0 *1 20.615,72.03
X$17251 1454 VIA_via1_4
* cell instance $17252 r0 *1 25.175,72.03
X$17252 1454 VIA_via1_4
* cell instance $17253 r0 *1 40.565,70.77
X$17253 1454 VIA_via1_4
* cell instance $17254 r0 *1 35.625,70.77
X$17254 1454 VIA_via1_4
* cell instance $17255 r0 *1 74.575,62.37
X$17255 1454 VIA_via1_4
* cell instance $17256 r0 *1 43.495,66.57
X$17256 1454 VIA_via3_2
* cell instance $17257 r0 *1 44.055,66.57
X$17257 1454 VIA_via3_2
* cell instance $17258 r0 *1 44.055,71.05
X$17258 1454 VIA_via3_2
* cell instance $17259 r0 *1 43.495,59.43
X$17259 1454 VIA_via3_2
* cell instance $17260 r0 *1 52.535,56.77
X$17260 1455 VIA_via2_5
* cell instance $17261 r0 *1 53.675,56.77
X$17261 1455 VIA_via2_5
* cell instance $17262 r0 *1 48.545,56.77
X$17262 1455 VIA_via1_4
* cell instance $17263 r0 *1 48.545,56.77
X$17263 1455 VIA_via2_5
* cell instance $17264 r0 *1 52.725,55.65
X$17264 1455 VIA_via1_4
* cell instance $17265 r0 *1 53.675,55.23
X$17265 1455 VIA_via1_4
* cell instance $17266 r0 *1 65.455,77.21
X$17266 1456 VIA_via1_7
* cell instance $17267 r0 *1 59.755,58.31
X$17267 1456 VIA_via2_5
* cell instance $17268 r0 *1 62.985,58.31
X$17268 1456 VIA_via2_5
* cell instance $17269 r0 *1 63.175,58.45
X$17269 1456 VIA_via2_5
* cell instance $17270 r0 *1 65.645,58.45
X$17270 1456 VIA_via2_5
* cell instance $17271 r0 *1 59.755,56.77
X$17271 1456 VIA_via1_4
* cell instance $17272 r0 *1 59.755,55.23
X$17272 1456 VIA_via1_4
* cell instance $17273 r0 *1 62.985,58.03
X$17273 1456 VIA_via1_4
* cell instance $17274 r0 *1 65.645,58.03
X$17274 1456 VIA_via1_4
* cell instance $17275 r0 *1 59.945,56.91
X$17275 1457 VIA_via2_5
* cell instance $17276 r0 *1 61.655,56.49
X$17276 1457 VIA_via2_5
* cell instance $17277 r0 *1 61.465,63.49
X$17277 1457 VIA_via2_5
* cell instance $17278 r0 *1 61.845,63.49
X$17278 1457 VIA_via2_5
* cell instance $17279 r0 *1 61.275,58.17
X$17279 1457 VIA_via2_5
* cell instance $17280 r0 *1 62.605,82.95
X$17280 1457 VIA_via1_4
* cell instance $17281 r0 *1 59.945,58.17
X$17281 1457 VIA_via1_4
* cell instance $17282 r0 *1 59.945,58.17
X$17282 1457 VIA_via2_5
* cell instance $17283 r0 *1 59.185,56.77
X$17283 1457 VIA_via1_4
* cell instance $17284 r0 *1 59.185,56.91
X$17284 1457 VIA_via2_5
* cell instance $17285 r0 *1 62.605,56.77
X$17285 1457 VIA_via1_4
* cell instance $17286 r0 *1 62.605,56.91
X$17286 1457 VIA_via2_5
* cell instance $17287 r0 *1 61.655,55.23
X$17287 1457 VIA_via1_4
* cell instance $17288 r0 *1 63.175,81.97
X$17288 1458 VIA_via1_4
* cell instance $17289 r0 *1 63.175,81.97
X$17289 1458 VIA_via2_5
* cell instance $17290 r0 *1 63.175,84.35
X$17290 1458 VIA_via1_4
* cell instance $17291 r0 *1 63.745,56.77
X$17291 1458 VIA_via1_4
* cell instance $17292 r0 *1 65.075,58.03
X$17292 1458 VIA_via1_4
* cell instance $17293 r0 *1 65.075,58.17
X$17293 1458 VIA_via2_5
* cell instance $17294 r0 *1 63.935,58.17
X$17294 1458 VIA_via1_4
* cell instance $17295 r0 *1 63.935,58.17
X$17295 1458 VIA_via3_2
* cell instance $17296 r0 *1 63.935,58.17
X$17296 1458 VIA_via2_5
* cell instance $17297 r0 *1 63.935,81.97
X$17297 1458 VIA_via3_2
* cell instance $17298 r0 *1 74.955,58.03
X$17298 1459 VIA_via2_5
* cell instance $17299 r0 *1 73.625,58.03
X$17299 1459 VIA_via1_4
* cell instance $17300 r0 *1 73.625,58.03
X$17300 1459 VIA_via2_5
* cell instance $17301 r0 *1 75.145,56.77
X$17301 1459 VIA_via1_4
* cell instance $17302 r0 *1 75.525,58.03
X$17302 1459 VIA_via1_4
* cell instance $17303 r0 *1 75.525,58.03
X$17303 1459 VIA_via2_5
* cell instance $17304 r0 *1 76.095,57.19
X$17304 1460 VIA_via1_7
* cell instance $17305 r0 *1 88.255,81.83
X$17305 1460 VIA_via2_5
* cell instance $17306 r0 *1 87.115,77.63
X$17306 1460 VIA_via2_5
* cell instance $17307 r0 *1 88.635,77.49
X$17307 1460 VIA_via2_5
* cell instance $17308 r0 *1 81.605,82.25
X$17308 1460 VIA_via2_5
* cell instance $17309 r0 *1 83.125,80.15
X$17309 1460 VIA_via2_5
* cell instance $17310 r0 *1 83.885,80.15
X$17310 1460 VIA_via2_5
* cell instance $17311 r0 *1 70.205,83.65
X$17311 1460 VIA_via2_5
* cell instance $17312 r0 *1 69.445,83.65
X$17312 1460 VIA_via2_5
* cell instance $17313 r0 *1 83.885,82.25
X$17313 1460 VIA_via2_5
* cell instance $17314 r0 *1 81.605,87.85
X$17314 1460 VIA_via2_5
* cell instance $17315 r0 *1 81.605,83.65
X$17315 1460 VIA_via2_5
* cell instance $17316 r0 *1 88.635,87.85
X$17316 1460 VIA_via2_5
* cell instance $17317 r0 *1 76.095,57.61
X$17317 1460 VIA_via2_5
* cell instance $17318 r0 *1 82.935,58.59
X$17318 1460 VIA_via2_5
* cell instance $17319 r0 *1 81.225,58.59
X$17319 1460 VIA_via2_5
* cell instance $17320 r0 *1 81.225,57.61
X$17320 1460 VIA_via2_5
* cell instance $17321 r0 *1 82.365,58.59
X$17321 1460 VIA_via2_5
* cell instance $17322 r0 *1 69.445,81.97
X$17322 1460 VIA_via1_4
* cell instance $17323 r0 *1 83.885,80.43
X$17323 1460 VIA_via1_4
* cell instance $17324 r0 *1 81.605,88.83
X$17324 1460 VIA_via1_4
* cell instance $17325 r0 *1 89.395,88.83
X$17325 1460 VIA_via1_4
* cell instance $17326 r0 *1 70.585,87.57
X$17326 1460 VIA_via1_4
* cell instance $17327 r0 *1 88.635,76.37
X$17327 1460 VIA_via1_4
* cell instance $17328 r0 *1 88.635,83.23
X$17328 1460 VIA_via1_4
* cell instance $17329 r0 *1 86.925,77.63
X$17329 1460 VIA_via1_4
* cell instance $17330 r0 *1 81.225,56.77
X$17330 1460 VIA_via1_4
* cell instance $17331 r0 *1 82.175,55.23
X$17331 1460 VIA_via1_4
* cell instance $17332 r0 *1 88.015,77.63
X$17332 1460 VIA_via3_2
* cell instance $17333 r0 *1 88.015,81.83
X$17333 1460 VIA_via3_2
* cell instance $17334 r0 *1 91.485,60.13
X$17334 1461 VIA_via2_5
* cell instance $17335 r0 *1 91.865,60.13
X$17335 1461 VIA_via2_5
* cell instance $17336 r0 *1 91.485,56.35
X$17336 1461 VIA_via1_4
* cell instance $17337 r0 *1 91.865,60.83
X$17337 1461 VIA_via1_4
* cell instance $17338 r0 *1 92.815,56.49
X$17338 1462 VIA_via1_4
* cell instance $17339 r0 *1 92.815,59.57
X$17339 1462 VIA_via1_4
* cell instance $17340 r0 *1 93.575,55.65
X$17340 1463 VIA_via1_7
* cell instance $17341 r0 *1 93.765,56.77
X$17341 1463 VIA_via1_4
* cell instance $17342 r0 *1 95.665,55.79
X$17342 1464 VIA_via1_7
* cell instance $17343 r0 *1 95.665,55.79
X$17343 1464 VIA_via2_5
* cell instance $17344 r0 *1 95.855,56.63
X$17344 1464 VIA_via4_0
* cell instance $17345 r0 *1 95.855,55.79
X$17345 1464 VIA_via3_2
* cell instance $17346 r0 *1 96.995,56.21
X$17346 1465 VIA_via1_7
* cell instance $17347 r0 *1 96.995,55.51
X$17347 1465 VIA_via2_5
* cell instance $17348 r0 *1 97.815,55.51
X$17348 1465 VIA_via3_2
* cell instance $17349 r0 *1 97.815,55.51
X$17349 1465 VIA_via4_0
* cell instance $17350 r0 *1 96.045,56.21
X$17350 1466 VIA_via1_7
* cell instance $17351 r0 *1 96.045,56.07
X$17351 1466 VIA_via2_5
* cell instance $17352 r0 *1 97.255,56.07
X$17352 1466 VIA_via4_0
* cell instance $17353 r0 *1 97.255,56.07
X$17353 1466 VIA_via3_2
* cell instance $17354 r0 *1 11.115,56.21
X$17354 1467 VIA_via1_7
* cell instance $17355 r0 *1 11.115,55.23
X$17355 1467 VIA_via2_5
* cell instance $17356 r0 *1 12.635,55.23
X$17356 1467 VIA_via1_4
* cell instance $17357 r0 *1 12.635,55.23
X$17357 1467 VIA_via2_5
* cell instance $17358 r0 *1 6.745,56.63
X$17358 1468 VIA_via1_4
* cell instance $17359 r0 *1 6.745,56.63
X$17359 1468 VIA_via2_5
* cell instance $17360 r0 *1 10.735,56.77
X$17360 1468 VIA_via1_4
* cell instance $17361 r0 *1 10.735,56.63
X$17361 1468 VIA_via2_5
* cell instance $17362 r0 *1 95.665,56.49
X$17362 1469 VIA_via2_5
* cell instance $17363 r0 *1 93.575,56.49
X$17363 1469 VIA_via1_4
* cell instance $17364 r0 *1 93.575,56.49
X$17364 1469 VIA_via2_5
* cell instance $17365 r0 *1 95.665,56.77
X$17365 1469 VIA_via1_4
* cell instance $17366 r0 *1 95.285,56.21
X$17366 1470 VIA_via1_7
* cell instance $17367 r0 *1 95.285,55.23
X$17367 1470 VIA_via1_4
* cell instance $17368 r0 *1 89.395,56.35
X$17368 1471 VIA_via2_5
* cell instance $17369 r0 *1 89.585,60.83
X$17369 1471 VIA_via1_4
* cell instance $17370 r0 *1 78.565,56.35
X$17370 1471 VIA_via1_4
* cell instance $17371 r0 *1 78.565,56.35
X$17371 1471 VIA_via2_5
* cell instance $17372 r0 *1 86.545,56.49
X$17372 1472 VIA_via1_7
* cell instance $17373 r0 *1 86.545,55.23
X$17373 1472 VIA_via1_4
* cell instance $17374 r0 *1 80.465,56.49
X$17374 1473 VIA_via1_7
* cell instance $17375 r0 *1 80.465,56.49
X$17375 1473 VIA_via2_5
* cell instance $17376 r0 *1 79.705,56.49
X$17376 1473 VIA_via2_5
* cell instance $17377 r0 *1 79.705,55.23
X$17377 1473 VIA_via1_4
* cell instance $17378 r0 *1 31.635,55.23
X$17378 1474 VIA_via1_4
* cell instance $17379 r0 *1 31.635,55.23
X$17379 1474 VIA_via2_5
* cell instance $17380 r0 *1 30.875,55.23
X$17380 1474 VIA_via1_4
* cell instance $17381 r0 *1 30.875,55.23
X$17381 1474 VIA_via2_5
* cell instance $17382 r0 *1 77.805,55.23
X$17382 1475 VIA_via1_4
* cell instance $17383 r0 *1 77.805,55.23
X$17383 1475 VIA_via2_5
* cell instance $17384 r0 *1 74.195,55.23
X$17384 1475 VIA_via1_4
* cell instance $17385 r0 *1 74.195,55.23
X$17385 1475 VIA_via2_5
* cell instance $17386 r0 *1 67.545,55.79
X$17386 1476 VIA_via1_7
* cell instance $17387 r0 *1 67.545,55.93
X$17387 1476 VIA_via2_5
* cell instance $17388 r0 *1 66.405,55.93
X$17388 1476 VIA_via2_5
* cell instance $17389 r0 *1 66.405,56.77
X$17389 1476 VIA_via1_4
* cell instance $17390 r0 *1 49.495,56.21
X$17390 1477 VIA_via1_7
* cell instance $17391 r0 *1 49.495,55.23
X$17391 1477 VIA_via2_5
* cell instance $17392 r0 *1 50.445,55.23
X$17392 1477 VIA_via1_4
* cell instance $17393 r0 *1 50.445,55.23
X$17393 1477 VIA_via2_5
* cell instance $17394 r0 *1 59.565,72.03
X$17394 1478 VIA_via2_5
* cell instance $17395 r0 *1 77.235,80.15
X$17395 1478 VIA_via2_5
* cell instance $17396 r0 *1 72.295,82.95
X$17396 1478 VIA_via2_5
* cell instance $17397 r0 *1 59.565,77.91
X$17397 1478 VIA_via2_5
* cell instance $17398 r0 *1 77.235,82.95
X$17398 1478 VIA_via2_5
* cell instance $17399 r0 *1 68.875,77.91
X$17399 1478 VIA_via2_5
* cell instance $17400 r0 *1 68.685,92.75
X$17400 1478 VIA_via2_5
* cell instance $17401 r0 *1 69.255,92.75
X$17401 1478 VIA_via2_5
* cell instance $17402 r0 *1 79.325,76.23
X$17402 1478 VIA_via2_5
* cell instance $17403 r0 *1 79.135,92.75
X$17403 1478 VIA_via2_5
* cell instance $17404 r0 *1 75.335,57.33
X$17404 1478 VIA_via2_5
* cell instance $17405 r0 *1 72.295,83.23
X$17405 1478 VIA_via1_4
* cell instance $17406 r0 *1 55.575,72.03
X$17406 1478 VIA_via1_4
* cell instance $17407 r0 *1 55.575,72.03
X$17407 1478 VIA_via2_5
* cell instance $17408 r0 *1 79.135,93.17
X$17408 1478 VIA_via1_4
* cell instance $17409 r0 *1 79.135,93.17
X$17409 1478 VIA_via2_5
* cell instance $17410 r0 *1 79.325,80.43
X$17410 1478 VIA_via1_4
* cell instance $17411 r0 *1 79.335,80.43
X$17411 1478 VIA_via3_2
* cell instance $17412 r0 *1 79.325,80.43
X$17412 1478 VIA_via2_5
* cell instance $17413 r0 *1 77.235,80.43
X$17413 1478 VIA_via1_4
* cell instance $17414 r0 *1 78.565,76.37
X$17414 1478 VIA_via1_4
* cell instance $17415 r0 *1 78.565,76.23
X$17415 1478 VIA_via2_5
* cell instance $17416 r0 *1 68.685,95.55
X$17416 1478 VIA_via1_4
* cell instance $17417 r0 *1 55.575,55.23
X$17417 1478 VIA_via1_4
* cell instance $17418 r0 *1 55.575,55.23
X$17418 1478 VIA_via2_5
* cell instance $17419 r0 *1 75.335,56.77
X$17419 1478 VIA_via1_4
* cell instance $17420 r0 *1 79.895,66.43
X$17420 1478 VIA_via1_4
* cell instance $17421 r0 *1 79.895,66.43
X$17421 1478 VIA_via2_5
* cell instance $17422 r0 *1 79.615,66.43
X$17422 1478 VIA_via3_2
* cell instance $17423 r0 *1 79.335,93.17
X$17423 1478 VIA_via3_2
* cell instance $17424 r0 *1 79.615,76.23
X$17424 1478 VIA_via3_2
* cell instance $17425 r0 *1 55.815,55.23
X$17425 1478 VIA_via3_2
* cell instance $17426 r0 *1 55.815,72.03
X$17426 1478 VIA_via3_2
* cell instance $17427 r0 *1 79.615,57.33
X$17427 1478 VIA_via3_2
* cell instance $17428 r0 *1 5.795,57.05
X$17428 1479 VIA_via2_5
* cell instance $17429 r0 *1 5.795,56.77
X$17429 1479 VIA_via1_4
* cell instance $17430 r0 *1 4.655,58.03
X$17430 1479 VIA_via1_4
* cell instance $17431 r0 *1 4.845,57.05
X$17431 1479 VIA_via1_4
* cell instance $17432 r0 *1 4.845,57.05
X$17432 1479 VIA_via2_5
* cell instance $17433 r0 *1 56.095,58.47
X$17433 1480 VIA_via6_0
* cell instance $17434 r0 *1 5.975,58.47
X$17434 1480 VIA_via6_0
* cell instance $17435 r0 *1 58.425,94.57
X$17435 1480 VIA_via1_7
* cell instance $17436 r0 *1 19.285,91.77
X$17436 1480 VIA_via1_7
* cell instance $17437 r0 *1 19.285,91.91
X$17437 1480 VIA_via2_5
* cell instance $17438 r0 *1 12.825,93.03
X$17438 1480 VIA_via1_7
* cell instance $17439 r0 *1 5.605,76.23
X$17439 1480 VIA_via1_7
* cell instance $17440 r0 *1 5.605,76.23
X$17440 1480 VIA_via2_5
* cell instance $17441 r0 *1 26.315,91.77
X$17441 1480 VIA_via1_7
* cell instance $17442 r0 *1 5.415,62.23
X$17442 1480 VIA_via1_7
* cell instance $17443 r0 *1 5.415,62.37
X$17443 1480 VIA_via2_5
* cell instance $17444 r0 *1 5.415,62.37
X$17444 1480 VIA_via3_2
* cell instance $17445 r0 *1 5.795,58.17
X$17445 1480 VIA_via1_7
* cell instance $17446 r0 *1 5.795,58.17
X$17446 1480 VIA_via2_5
* cell instance $17447 r0 *1 57.495,65.59
X$17447 1480 VIA_via5_0
* cell instance $17448 r0 *1 57.495,58.31
X$17448 1480 VIA_via5_0
* cell instance $17449 r0 *1 26.315,92.05
X$17449 1480 VIA_via2_5
* cell instance $17450 r0 *1 13.015,92.75
X$17450 1480 VIA_via2_5
* cell instance $17451 r0 *1 19.285,92.75
X$17451 1480 VIA_via2_5
* cell instance $17452 r0 *1 56.715,65.59
X$17452 1480 VIA_via2_5
* cell instance $17453 r0 *1 58.425,90.37
X$17453 1480 VIA_via2_5
* cell instance $17454 r0 *1 40.375,94.01
X$17454 1480 VIA_via2_5
* cell instance $17455 r0 *1 40.375,91.91
X$17455 1480 VIA_via2_5
* cell instance $17456 r0 *1 58.425,94.15
X$17456 1480 VIA_via2_5
* cell instance $17457 r0 *1 5.415,58.17
X$17457 1480 VIA_via2_5
* cell instance $17458 r0 *1 58.045,90.37
X$17458 1480 VIA_via1_4
* cell instance $17459 r0 *1 58.055,90.37
X$17459 1480 VIA_via3_2
* cell instance $17460 r0 *1 58.045,90.37
X$17460 1480 VIA_via2_5
* cell instance $17461 r0 *1 58.055,90.51
X$17461 1480 VIA_via4_0
* cell instance $17462 r0 *1 58.055,90.51
X$17462 1480 VIA_via5_0
* cell instance $17463 r0 *1 56.715,65.17
X$17463 1480 VIA_via1_4
* cell instance $17464 r0 *1 40.375,94.43
X$17464 1480 VIA_via1_4
* cell instance $17465 r0 *1 56.095,58.31
X$17465 1480 VIA_via4_0
* cell instance $17466 r0 *1 56.095,58.31
X$17466 1480 VIA_via5_0
* cell instance $17467 r0 *1 56.095,58.31
X$17467 1480 VIA_via3_2
* cell instance $17468 r0 *1 56.145,58.31
X$17468 1480 VIA_via2_5
* cell instance $17469 r0 *1 56.145,58.31
X$17469 1480 VIA_via1_4
* cell instance $17470 r0 *1 56.935,65.59
X$17470 1480 VIA_via4_0
* cell instance $17471 r0 *1 56.935,65.59
X$17471 1480 VIA_via3_2
* cell instance $17472 r0 *1 5.975,58.31
X$17472 1480 VIA_via4_0
* cell instance $17473 r0 *1 5.975,58.17
X$17473 1480 VIA_via3_2
* cell instance $17474 r0 *1 5.975,58.31
X$17474 1480 VIA_via5_0
* cell instance $17475 r0 *1 5.415,76.23
X$17475 1480 VIA_via3_2
* cell instance $17476 r0 *1 6.365,56.77
X$17476 1481 VIA_via1_4
* cell instance $17477 r0 *1 7.885,59.15
X$17477 1481 VIA_via1_4
* cell instance $17478 r0 *1 6.555,58.03
X$17478 1481 VIA_via1_4
* cell instance $17479 r0 *1 48.735,63.77
X$17479 1482 VIA_via1_7
* cell instance $17480 r0 *1 48.735,63.91
X$17480 1482 VIA_via2_5
* cell instance $17481 r0 *1 20.805,84.63
X$17481 1482 VIA_via1_7
* cell instance $17482 r0 *1 10.165,80.57
X$17482 1482 VIA_via1_7
* cell instance $17483 r0 *1 9.405,83.37
X$17483 1482 VIA_via1_7
* cell instance $17484 r0 *1 9.405,83.37
X$17484 1482 VIA_via2_5
* cell instance $17485 r0 *1 32.585,83.37
X$17485 1482 VIA_via1_7
* cell instance $17486 r0 *1 32.585,83.37
X$17486 1482 VIA_via2_5
* cell instance $17487 r0 *1 41.135,84.63
X$17487 1482 VIA_via1_7
* cell instance $17488 r0 *1 48.165,83.37
X$17488 1482 VIA_via1_7
* cell instance $17489 r0 *1 48.165,83.37
X$17489 1482 VIA_via2_5
* cell instance $17490 r0 *1 9.595,58.17
X$17490 1482 VIA_via1_7
* cell instance $17491 r0 *1 9.595,58.17
X$17491 1482 VIA_via2_5
* cell instance $17492 r0 *1 32.585,82.95
X$17492 1482 VIA_via2_5
* cell instance $17493 r0 *1 9.975,83.37
X$17493 1482 VIA_via2_5
* cell instance $17494 r0 *1 9.975,82.95
X$17494 1482 VIA_via2_5
* cell instance $17495 r0 *1 21.185,83.37
X$17495 1482 VIA_via2_5
* cell instance $17496 r0 *1 21.185,82.81
X$17496 1482 VIA_via2_5
* cell instance $17497 r0 *1 41.135,82.95
X$17497 1482 VIA_via2_5
* cell instance $17498 r0 *1 41.135,83.37
X$17498 1482 VIA_via2_5
* cell instance $17499 r0 *1 55.195,61.25
X$17499 1482 VIA_via2_5
* cell instance $17500 r0 *1 49.685,64.47
X$17500 1482 VIA_via2_5
* cell instance $17501 r0 *1 49.685,83.37
X$17501 1482 VIA_via2_5
* cell instance $17502 r0 *1 55.195,83.37
X$17502 1482 VIA_via2_5
* cell instance $17503 r0 *1 48.735,64.47
X$17503 1482 VIA_via2_5
* cell instance $17504 r0 *1 55.195,81.97
X$17504 1482 VIA_via1_4
* cell instance $17505 r0 *1 11.305,62.37
X$17505 1482 VIA_via1_4
* cell instance $17506 r0 *1 11.305,62.37
X$17506 1482 VIA_via2_5
* cell instance $17507 r0 *1 54.815,58.45
X$17507 1482 VIA_via1_4
* cell instance $17508 r0 *1 48.535,62.51
X$17508 1482 VIA_via4_0
* cell instance $17509 r0 *1 11.575,62.37
X$17509 1482 VIA_via3_2
* cell instance $17510 r0 *1 11.575,62.51
X$17510 1482 VIA_via4_0
* cell instance $17511 r0 *1 48.535,63.91
X$17511 1482 VIA_via3_2
* cell instance $17512 r0 *1 11.575,58.31
X$17512 1482 VIA_via3_2
* cell instance $17513 r0 *1 48.535,61.25
X$17513 1482 VIA_via3_2
* cell instance $17514 r0 *1 31.635,90.37
X$17514 1483 VIA_via2_5
* cell instance $17515 r0 *1 11.685,75.11
X$17515 1483 VIA_via2_5
* cell instance $17516 r0 *1 21.375,90.79
X$17516 1483 VIA_via2_5
* cell instance $17517 r0 *1 55.765,66.15
X$17517 1483 VIA_via2_5
* cell instance $17518 r0 *1 55.765,66.99
X$17518 1483 VIA_via2_5
* cell instance $17519 r0 *1 56.525,66.99
X$17519 1483 VIA_via2_5
* cell instance $17520 r0 *1 56.145,91.49
X$17520 1483 VIA_via2_5
* cell instance $17521 r0 *1 42.085,91.49
X$17521 1483 VIA_via2_5
* cell instance $17522 r0 *1 43.985,60.97
X$17522 1483 VIA_via2_5
* cell instance $17523 r0 *1 43.985,66.01
X$17523 1483 VIA_via2_5
* cell instance $17524 r0 *1 35.435,60.97
X$17524 1483 VIA_via2_5
* cell instance $17525 r0 *1 53.485,91.63
X$17525 1483 VIA_via1_4
* cell instance $17526 r0 *1 53.485,91.49
X$17526 1483 VIA_via2_5
* cell instance $17527 r0 *1 56.335,88.83
X$17527 1483 VIA_via1_4
* cell instance $17528 r0 *1 56.335,88.69
X$17528 1483 VIA_via2_5
* cell instance $17529 r0 *1 13.585,91.63
X$17529 1483 VIA_via1_4
* cell instance $17530 r0 *1 13.585,91.49
X$17530 1483 VIA_via2_5
* cell instance $17531 r0 *1 21.375,90.37
X$17531 1483 VIA_via1_4
* cell instance $17532 r0 *1 21.375,90.37
X$17532 1483 VIA_via2_5
* cell instance $17533 r0 *1 42.085,90.37
X$17533 1483 VIA_via1_4
* cell instance $17534 r0 *1 31.635,91.63
X$17534 1483 VIA_via1_4
* cell instance $17535 r0 *1 11.115,63.63
X$17535 1483 VIA_via1_4
* cell instance $17536 r0 *1 11.115,63.63
X$17536 1483 VIA_via2_5
* cell instance $17537 r0 *1 11.115,56.77
X$17537 1483 VIA_via1_4
* cell instance $17538 r0 *1 11.115,56.77
X$17538 1483 VIA_via2_5
* cell instance $17539 r0 *1 35.435,57.05
X$17539 1483 VIA_via1_4
* cell instance $17540 r0 *1 35.435,57.19
X$17540 1483 VIA_via2_5
* cell instance $17541 r0 *1 35.375,57.19
X$17541 1483 VIA_via3_2
* cell instance $17542 r0 *1 11.685,74.83
X$17542 1483 VIA_via1_4
* cell instance $17543 r0 *1 56.525,65.17
X$17543 1483 VIA_via1_4
* cell instance $17544 r0 *1 35.375,56.91
X$17544 1483 VIA_via4_0
* cell instance $17545 r0 *1 14.095,91.49
X$17545 1483 VIA_via3_2
* cell instance $17546 r0 *1 14.095,90.79
X$17546 1483 VIA_via3_2
* cell instance $17547 r0 *1 11.295,63.63
X$17547 1483 VIA_via3_2
* cell instance $17548 r0 *1 56.935,66.99
X$17548 1483 VIA_via3_2
* cell instance $17549 r0 *1 11.295,56.77
X$17549 1483 VIA_via3_2
* cell instance $17550 r0 *1 11.295,56.91
X$17550 1483 VIA_via4_0
* cell instance $17551 r0 *1 14.095,75.11
X$17551 1483 VIA_via3_2
* cell instance $17552 r0 *1 11.295,75.11
X$17552 1483 VIA_via3_2
* cell instance $17553 r0 *1 56.935,88.69
X$17553 1483 VIA_via3_2
* cell instance $17554 r0 *1 23.275,57.05
X$17554 1484 VIA_via2_5
* cell instance $17555 r0 *1 26.885,57.05
X$17555 1484 VIA_via2_5
* cell instance $17556 r0 *1 26.885,58.03
X$17556 1484 VIA_via1_4
* cell instance $17557 r0 *1 25.935,57.05
X$17557 1484 VIA_via1_4
* cell instance $17558 r0 *1 25.935,57.05
X$17558 1484 VIA_via2_5
* cell instance $17559 r0 *1 23.085,58.03
X$17559 1484 VIA_via1_4
* cell instance $17560 r0 *1 52.345,52.29
X$17560 1485 VIA_via1_7
* cell instance $17561 r0 *1 26.125,76.65
X$17561 1485 VIA_via2_5
* cell instance $17562 r0 *1 19.855,76.51
X$17562 1485 VIA_via2_5
* cell instance $17563 r0 *1 47.975,75.39
X$17563 1485 VIA_via2_5
* cell instance $17564 r0 *1 52.345,58.17
X$17564 1485 VIA_via2_5
* cell instance $17565 r0 *1 52.915,58.87
X$17565 1485 VIA_via2_5
* cell instance $17566 r0 *1 52.915,60.55
X$17566 1485 VIA_via2_5
* cell instance $17567 r0 *1 52.345,58.87
X$17567 1485 VIA_via2_5
* cell instance $17568 r0 *1 53.485,75.39
X$17568 1485 VIA_via2_5
* cell instance $17569 r0 *1 21.185,61.25
X$17569 1485 VIA_via2_5
* cell instance $17570 r0 *1 53.865,74.83
X$17570 1485 VIA_via1_4
* cell instance $17571 r0 *1 39.805,76.37
X$17571 1485 VIA_via1_4
* cell instance $17572 r0 *1 39.805,76.23
X$17572 1485 VIA_via2_5
* cell instance $17573 r0 *1 39.855,76.23
X$17573 1485 VIA_via3_2
* cell instance $17574 r0 *1 39.855,76.23
X$17574 1485 VIA_via4_0
* cell instance $17575 r0 *1 34.105,76.37
X$17575 1485 VIA_via1_4
* cell instance $17576 r0 *1 34.105,76.23
X$17576 1485 VIA_via2_5
* cell instance $17577 r0 *1 28.595,58.03
X$17577 1485 VIA_via1_4
* cell instance $17578 r0 *1 28.595,58.17
X$17578 1485 VIA_via2_5
* cell instance $17579 r0 *1 26.125,76.37
X$17579 1485 VIA_via1_4
* cell instance $17580 r0 *1 21.185,62.37
X$17580 1485 VIA_via1_4
* cell instance $17581 r0 *1 20.615,76.37
X$17581 1485 VIA_via1_4
* cell instance $17582 r0 *1 20.615,76.51
X$17582 1485 VIA_via2_5
* cell instance $17583 r0 *1 53.865,60.9
X$17583 1485 VIA_via1_4
* cell instance $17584 r0 *1 53.865,60.97
X$17584 1485 VIA_via2_5
* cell instance $17585 r0 *1 19.855,73.57
X$17585 1485 VIA_via1_4
* cell instance $17586 r0 *1 28.375,58.03
X$17586 1485 VIA_via4_0
* cell instance $17587 r0 *1 28.375,58.17
X$17587 1485 VIA_via3_2
* cell instance $17588 r0 *1 53.015,75.39
X$17588 1485 VIA_via3_2
* cell instance $17589 r0 *1 47.975,76.23
X$17589 1485 VIA_via3_2
* cell instance $17590 r0 *1 47.975,76.23
X$17590 1485 VIA_via4_0
* cell instance $17591 r0 *1 47.975,76.23
X$17591 1485 VIA_via2_5
* cell instance $17592 r0 *1 47.975,76.37
X$17592 1485 VIA_via1_4
* cell instance $17593 r0 *1 28.375,61.25
X$17593 1485 VIA_via3_2
* cell instance $17594 r0 *1 53.015,60.69
X$17594 1485 VIA_via3_2
* cell instance $17595 r0 *1 51.895,58.17
X$17595 1485 VIA_via3_2
* cell instance $17596 r0 *1 51.895,58.03
X$17596 1485 VIA_via4_0
* cell instance $17597 r0 *1 8.075,66.29
X$17597 1486 VIA_via2_5
* cell instance $17598 r0 *1 14.155,66.57
X$17598 1486 VIA_via2_5
* cell instance $17599 r0 *1 22.515,66.57
X$17599 1486 VIA_via2_5
* cell instance $17600 r0 *1 23.465,66.57
X$17600 1486 VIA_via2_5
* cell instance $17601 r0 *1 46.835,58.73
X$17601 1486 VIA_via2_5
* cell instance $17602 r0 *1 37.715,56.91
X$17602 1486 VIA_via2_5
* cell instance $17603 r0 *1 37.715,58.73
X$17603 1486 VIA_via2_5
* cell instance $17604 r0 *1 21.185,56.91
X$17604 1486 VIA_via2_5
* cell instance $17605 r0 *1 22.515,58.73
X$17605 1486 VIA_via2_5
* cell instance $17606 r0 *1 21.185,58.73
X$17606 1486 VIA_via2_5
* cell instance $17607 r0 *1 15.675,58.73
X$17607 1486 VIA_via2_5
* cell instance $17608 r0 *1 37.715,55.23
X$17608 1486 VIA_via1_4
* cell instance $17609 r0 *1 46.835,60.83
X$17609 1486 VIA_via1_4
* cell instance $17610 r0 *1 30.875,56.77
X$17610 1486 VIA_via1_4
* cell instance $17611 r0 *1 30.875,56.91
X$17611 1486 VIA_via2_5
* cell instance $17612 r0 *1 15.675,53.97
X$17612 1486 VIA_via1_4
* cell instance $17613 r0 *1 24.605,66.43
X$17613 1486 VIA_via1_4
* cell instance $17614 r0 *1 24.605,66.57
X$17614 1486 VIA_via2_5
* cell instance $17615 r0 *1 24.065,67.97
X$17615 1486 VIA_via1_4
* cell instance $17616 r0 *1 23.465,67.55
X$17616 1486 VIA_via1_4
* cell instance $17617 r0 *1 23.845,67.97
X$17617 1486 VIA_via1_4
* cell instance $17618 r0 *1 14.155,69.23
X$17618 1486 VIA_via1_4
* cell instance $17619 r0 *1 8.075,59.57
X$17619 1486 VIA_via1_4
* cell instance $17620 r0 *1 21.185,59.57
X$17620 1486 VIA_via1_4
* cell instance $17621 r0 *1 5.985,66.43
X$17621 1486 VIA_via1_4
* cell instance $17622 r0 *1 5.985,66.29
X$17622 1486 VIA_via2_5
* cell instance $17623 r0 *1 40.565,67.97
X$17623 1486 VIA_via1_4
* cell instance $17624 r0 *1 40.565,67.97
X$17624 1486 VIA_via2_5
* cell instance $17625 r0 *1 40.415,58.73
X$17625 1486 VIA_via3_2
* cell instance $17626 r0 *1 40.415,67.97
X$17626 1486 VIA_via3_2
* cell instance $17627 r0 *1 39.235,70.63
X$17627 1487 VIA_via1_7
* cell instance $17628 r0 *1 41.515,67.83
X$17628 1487 VIA_via1_7
* cell instance $17629 r0 *1 41.515,67.69
X$17629 1487 VIA_via2_5
* cell instance $17630 r0 *1 33.155,67.83
X$17630 1487 VIA_via1_7
* cell instance $17631 r0 *1 33.155,67.83
X$17631 1487 VIA_via2_5
* cell instance $17632 r0 *1 39.805,59.43
X$17632 1487 VIA_via1_7
* cell instance $17633 r0 *1 39.805,59.43
X$17633 1487 VIA_via2_5
* cell instance $17634 r0 *1 24.225,69.09
X$17634 1487 VIA_via2_5
* cell instance $17635 r0 *1 19.285,67.97
X$17635 1487 VIA_via2_5
* cell instance $17636 r0 *1 19.285,69.09
X$17636 1487 VIA_via2_5
* cell instance $17637 r0 *1 23.465,62.37
X$17637 1487 VIA_via2_5
* cell instance $17638 r0 *1 25.745,67.83
X$17638 1487 VIA_via2_5
* cell instance $17639 r0 *1 48.545,67.69
X$17639 1487 VIA_via2_5
* cell instance $17640 r0 *1 39.235,67.69
X$17640 1487 VIA_via2_5
* cell instance $17641 r0 *1 33.535,59.43
X$17641 1487 VIA_via2_5
* cell instance $17642 r0 *1 32.965,59.43
X$17642 1487 VIA_via2_5
* cell instance $17643 r0 *1 48.735,59.85
X$17643 1487 VIA_via1_4
* cell instance $17644 r0 *1 33.155,56.77
X$17644 1487 VIA_via1_4
* cell instance $17645 r0 *1 22.895,62.37
X$17645 1487 VIA_via1_4
* cell instance $17646 r0 *1 22.895,62.37
X$17646 1487 VIA_via2_5
* cell instance $17647 r0 *1 19.285,72.03
X$17647 1487 VIA_via1_4
* cell instance $17648 r0 *1 19.855,67.97
X$17648 1487 VIA_via1_4
* cell instance $17649 r0 *1 19.855,67.97
X$17649 1487 VIA_via2_5
* cell instance $17650 r0 *1 48.165,72.03
X$17650 1487 VIA_via1_4
* cell instance $17651 r0 *1 25.745,69.23
X$17651 1487 VIA_via1_4
* cell instance $17652 r0 *1 25.745,69.09
X$17652 1487 VIA_via2_5
* cell instance $17653 r0 *1 33.155,58.17
X$17653 1488 VIA_via1_7
* cell instance $17654 r0 *1 33.155,58.17
X$17654 1488 VIA_via2_5
* cell instance $17655 r0 *1 51.585,70.63
X$17655 1488 VIA_via1_7
* cell instance $17656 r0 *1 51.585,70.63
X$17656 1488 VIA_via2_5
* cell instance $17657 r0 *1 32.775,70.63
X$17657 1488 VIA_via1_7
* cell instance $17658 r0 *1 32.775,70.63
X$17658 1488 VIA_via2_5
* cell instance $17659 r0 *1 25.745,70.63
X$17659 1488 VIA_via1_7
* cell instance $17660 r0 *1 25.745,70.63
X$17660 1488 VIA_via2_5
* cell instance $17661 r0 *1 42.085,58.17
X$17661 1488 VIA_via1_7
* cell instance $17662 r0 *1 42.085,58.17
X$17662 1488 VIA_via2_5
* cell instance $17663 r0 *1 17.955,70.63
X$17663 1488 VIA_via1_7
* cell instance $17664 r0 *1 23.275,63.77
X$17664 1488 VIA_via1_7
* cell instance $17665 r0 *1 18.145,66.57
X$17665 1488 VIA_via1_7
* cell instance $17666 r0 *1 18.145,69.37
X$17666 1488 VIA_via2_5
* cell instance $17667 r0 *1 23.655,69.37
X$17667 1488 VIA_via2_5
* cell instance $17668 r0 *1 23.655,70.63
X$17668 1488 VIA_via2_5
* cell instance $17669 r0 *1 50.635,57.61
X$17669 1488 VIA_via2_5
* cell instance $17670 r0 *1 43.795,58.17
X$17670 1488 VIA_via2_5
* cell instance $17671 r0 *1 43.795,57.61
X$17671 1488 VIA_via2_5
* cell instance $17672 r0 *1 43.415,67.97
X$17672 1488 VIA_via2_5
* cell instance $17673 r0 *1 40.375,70.63
X$17673 1488 VIA_via2_5
* cell instance $17674 r0 *1 42.845,69.51
X$17674 1488 VIA_via2_5
* cell instance $17675 r0 *1 42.845,70.63
X$17675 1488 VIA_via2_5
* cell instance $17676 r0 *1 40.375,69.51
X$17676 1488 VIA_via2_5
* cell instance $17677 r0 *1 42.845,67.97
X$17677 1488 VIA_via1_4
* cell instance $17678 r0 *1 42.845,67.97
X$17678 1488 VIA_via2_5
* cell instance $17679 r0 *1 40.755,69.23
X$17679 1488 VIA_via1_4
* cell instance $17680 r0 *1 50.635,57.05
X$17680 1488 VIA_via1_4
* cell instance $17681 r0 *1 42.275,58.31
X$17681 1489 VIA_via2_5
* cell instance $17682 r0 *1 42.845,58.31
X$17682 1489 VIA_via2_5
* cell instance $17683 r0 *1 41.705,58.31
X$17683 1489 VIA_via2_5
* cell instance $17684 r0 *1 42.845,59.57
X$17684 1489 VIA_via1_4
* cell instance $17685 r0 *1 42.275,58.03
X$17685 1489 VIA_via1_4
* cell instance $17686 r0 *1 41.705,57.05
X$17686 1489 VIA_via1_4
* cell instance $17687 r0 *1 49.115,58.03
X$17687 1490 VIA_via2_5
* cell instance $17688 r0 *1 49.115,57.05
X$17688 1490 VIA_via2_5
* cell instance $17689 r0 *1 45.695,60.41
X$17689 1490 VIA_via2_5
* cell instance $17690 r0 *1 41.705,60.41
X$17690 1490 VIA_via2_5
* cell instance $17691 r0 *1 40.565,60.41
X$17691 1490 VIA_via2_5
* cell instance $17692 r0 *1 42.845,60.41
X$17692 1490 VIA_via2_5
* cell instance $17693 r0 *1 47.025,57.05
X$17693 1490 VIA_via2_5
* cell instance $17694 r0 *1 47.785,57.05
X$17694 1490 VIA_via2_5
* cell instance $17695 r0 *1 49.115,56.77
X$17695 1490 VIA_via1_4
* cell instance $17696 r0 *1 45.695,58.03
X$17696 1490 VIA_via1_4
* cell instance $17697 r0 *1 45.695,58.03
X$17697 1490 VIA_via2_5
* cell instance $17698 r0 *1 40.565,59.57
X$17698 1490 VIA_via1_4
* cell instance $17699 r0 *1 47.025,58.03
X$17699 1490 VIA_via1_4
* cell instance $17700 r0 *1 47.025,58.03
X$17700 1490 VIA_via2_5
* cell instance $17701 r0 *1 47.785,56.77
X$17701 1490 VIA_via1_4
* cell instance $17702 r0 *1 45.695,60.83
X$17702 1490 VIA_via1_4
* cell instance $17703 r0 *1 42.845,60.83
X$17703 1490 VIA_via1_4
* cell instance $17704 r0 *1 42.845,58.03
X$17704 1490 VIA_via1_4
* cell instance $17705 r0 *1 42.845,58.03
X$17705 1490 VIA_via2_5
* cell instance $17706 r0 *1 41.705,62.37
X$17706 1490 VIA_via1_4
* cell instance $17707 r0 *1 49.685,60.55
X$17707 1490 VIA_via1_4
* cell instance $17708 r0 *1 49.875,58.03
X$17708 1490 VIA_via1_4
* cell instance $17709 r0 *1 49.875,58.03
X$17709 1490 VIA_via2_5
* cell instance $17710 r0 *1 46.455,59.85
X$17710 1491 VIA_via2_5
* cell instance $17711 r0 *1 48.165,59.85
X$17711 1491 VIA_via2_5
* cell instance $17712 r0 *1 46.455,58.03
X$17712 1491 VIA_via1_4
* cell instance $17713 r0 *1 46.645,57.05
X$17713 1491 VIA_via1_4
* cell instance $17714 r0 *1 48.165,60.83
X$17714 1491 VIA_via1_4
* cell instance $17715 r0 *1 16.625,77.77
X$17715 1492 VIA_via1_7
* cell instance $17716 r0 *1 56.905,76.23
X$17716 1492 VIA_via1_7
* cell instance $17717 r0 *1 16.815,59.43
X$17717 1492 VIA_via1_7
* cell instance $17718 r0 *1 24.605,58.17
X$17718 1492 VIA_via1_7
* cell instance $17719 r0 *1 24.605,58.17
X$17719 1492 VIA_via2_5
* cell instance $17720 r0 *1 24.735,58.17
X$17720 1492 VIA_via3_2
* cell instance $17721 r0 *1 24.735,58.31
X$17721 1492 VIA_via4_0
* cell instance $17722 r0 *1 28.215,80.15
X$17722 1492 VIA_via2_5
* cell instance $17723 r0 *1 17.005,80.29
X$17723 1492 VIA_via2_5
* cell instance $17724 r0 *1 23.465,80.15
X$17724 1492 VIA_via2_5
* cell instance $17725 r0 *1 49.685,58.31
X$17725 1492 VIA_via2_5
* cell instance $17726 r0 *1 49.685,57.05
X$17726 1492 VIA_via2_5
* cell instance $17727 r0 *1 56.905,75.67
X$17727 1492 VIA_via2_5
* cell instance $17728 r0 *1 36.955,80.15
X$17728 1492 VIA_via2_5
* cell instance $17729 r0 *1 24.605,58.87
X$17729 1492 VIA_via2_5
* cell instance $17730 r0 *1 16.815,58.87
X$17730 1492 VIA_via2_5
* cell instance $17731 r0 *1 36.955,81.97
X$17731 1492 VIA_via1_4
* cell instance $17732 r0 *1 47.405,74.83
X$17732 1492 VIA_via1_4
* cell instance $17733 r0 *1 47.405,74.83
X$17733 1492 VIA_via2_5
* cell instance $17734 r0 *1 28.215,80.43
X$17734 1492 VIA_via1_4
* cell instance $17735 r0 *1 23.465,80.43
X$17735 1492 VIA_via1_4
* cell instance $17736 r0 *1 15.295,80.43
X$17736 1492 VIA_via1_4
* cell instance $17737 r0 *1 15.295,80.29
X$17737 1492 VIA_via2_5
* cell instance $17738 r0 *1 49.685,58.03
X$17738 1492 VIA_via1_4
* cell instance $17739 r0 *1 52.725,57.05
X$17739 1492 VIA_via1_4
* cell instance $17740 r0 *1 52.725,57.05
X$17740 1492 VIA_via2_5
* cell instance $17741 r0 *1 46.855,75.67
X$17741 1492 VIA_via4_0
* cell instance $17742 r0 *1 46.855,74.83
X$17742 1492 VIA_via3_2
* cell instance $17743 r0 *1 56.375,75.67
X$17743 1492 VIA_via3_2
* cell instance $17744 r0 *1 56.375,75.67
X$17744 1492 VIA_via4_0
* cell instance $17745 r0 *1 47.135,80.01
X$17745 1492 VIA_via3_2
* cell instance $17746 r0 *1 46.855,58.31
X$17746 1492 VIA_via3_2
* cell instance $17747 r0 *1 46.295,58.31
X$17747 1492 VIA_via3_2
* cell instance $17748 r0 *1 46.295,58.31
X$17748 1492 VIA_via4_0
* cell instance $17749 r0 *1 10.355,91.77
X$17749 1493 VIA_via1_7
* cell instance $17750 r0 *1 21.945,93.03
X$17750 1493 VIA_via1_7
* cell instance $17751 r0 *1 21.945,92.89
X$17751 1493 VIA_via2_5
* cell instance $17752 r0 *1 55.005,93.03
X$17752 1493 VIA_via1_7
* cell instance $17753 r0 *1 55.005,93.03
X$17753 1493 VIA_via2_5
* cell instance $17754 r0 *1 53.105,93.03
X$17754 1493 VIA_via1_7
* cell instance $17755 r0 *1 53.105,93.03
X$17755 1493 VIA_via2_5
* cell instance $17756 r0 *1 2.945,74.97
X$17756 1493 VIA_via1_7
* cell instance $17757 r0 *1 2.945,74.97
X$17757 1493 VIA_via2_5
* cell instance $17758 r0 *1 40.945,93.03
X$17758 1493 VIA_via1_7
* cell instance $17759 r0 *1 40.945,93.03
X$17759 1493 VIA_via2_5
* cell instance $17760 r0 *1 28.215,93.03
X$17760 1493 VIA_via1_7
* cell instance $17761 r0 *1 28.215,93.03
X$17761 1493 VIA_via2_5
* cell instance $17762 r0 *1 3.895,58.17
X$17762 1493 VIA_via1_7
* cell instance $17763 r0 *1 56.375,93.03
X$17763 1493 VIA_via5_0
* cell instance $17764 r0 *1 56.375,93.03
X$17764 1493 VIA_via4_0
* cell instance $17765 r0 *1 56.375,93.03
X$17765 1493 VIA_via3_2
* cell instance $17766 r0 *1 28.785,92.61
X$17766 1493 VIA_via2_5
* cell instance $17767 r0 *1 28.785,93.03
X$17767 1493 VIA_via2_5
* cell instance $17768 r0 *1 7.315,74.97
X$17768 1493 VIA_via2_5
* cell instance $17769 r0 *1 4.465,74.97
X$17769 1493 VIA_via2_5
* cell instance $17770 r0 *1 10.925,86.17
X$17770 1493 VIA_via2_5
* cell instance $17771 r0 *1 7.315,86.17
X$17771 1493 VIA_via2_5
* cell instance $17772 r0 *1 10.545,92.89
X$17772 1493 VIA_via2_5
* cell instance $17773 r0 *1 56.145,66.15
X$17773 1493 VIA_via2_5
* cell instance $17774 r0 *1 57.095,66.15
X$17774 1493 VIA_via2_5
* cell instance $17775 r0 *1 40.945,92.61
X$17775 1493 VIA_via2_5
* cell instance $17776 r0 *1 4.085,62.37
X$17776 1493 VIA_via1_4
* cell instance $17777 r0 *1 56.145,66.43
X$17777 1493 VIA_via1_4
* cell instance $17778 r0 *1 57.665,57.05
X$17778 1493 VIA_via1_4
* cell instance $17779 r0 *1 56.375,66.15
X$17779 1493 VIA_via4_0
* cell instance $17780 r0 *1 56.375,66.15
X$17780 1493 VIA_via5_0
* cell instance $17781 r0 *1 56.375,66.15
X$17781 1493 VIA_via3_2
* cell instance $17782 r0 *1 58.045,59.43
X$17782 1494 VIA_via2_5
* cell instance $17783 r0 *1 62.415,61.25
X$17783 1494 VIA_via2_5
* cell instance $17784 r0 *1 67.165,77.77
X$17784 1494 VIA_via1_4
* cell instance $17785 r0 *1 67.165,77.77
X$17785 1494 VIA_via2_5
* cell instance $17786 r0 *1 57.095,59.57
X$17786 1494 VIA_via1_4
* cell instance $17787 r0 *1 57.095,59.43
X$17787 1494 VIA_via2_5
* cell instance $17788 r0 *1 58.425,56.77
X$17788 1494 VIA_via1_4
* cell instance $17789 r0 *1 62.225,59.57
X$17789 1494 VIA_via1_4
* cell instance $17790 r0 *1 62.225,59.43
X$17790 1494 VIA_via2_5
* cell instance $17791 r0 *1 66.175,77.77
X$17791 1494 VIA_via3_2
* cell instance $17792 r0 *1 66.175,61.25
X$17792 1494 VIA_via3_2
* cell instance $17793 r0 *1 65.075,59.01
X$17793 1495 VIA_via1_7
* cell instance $17794 r0 *1 65.075,59.01
X$17794 1495 VIA_via2_5
* cell instance $17795 r0 *1 60.705,59.01
X$17795 1495 VIA_via2_5
* cell instance $17796 r0 *1 60.705,59.57
X$17796 1495 VIA_via2_5
* cell instance $17797 r0 *1 64.125,59.01
X$17797 1495 VIA_via2_5
* cell instance $17798 r0 *1 60.705,58.03
X$17798 1495 VIA_via1_4
* cell instance $17799 r0 *1 60.135,58.03
X$17799 1495 VIA_via1_4
* cell instance $17800 r0 *1 59.755,59.57
X$17800 1495 VIA_via1_4
* cell instance $17801 r0 *1 59.755,59.57
X$17801 1495 VIA_via2_5
* cell instance $17802 r0 *1 64.125,58.03
X$17802 1495 VIA_via1_4
* cell instance $17803 r0 *1 62.795,57.33
X$17803 1496 VIA_via2_5
* cell instance $17804 r0 *1 61.465,57.33
X$17804 1496 VIA_via2_5
* cell instance $17805 r0 *1 63.745,63.49
X$17805 1496 VIA_via2_5
* cell instance $17806 r0 *1 62.605,63.49
X$17806 1496 VIA_via2_5
* cell instance $17807 r0 *1 63.935,86.03
X$17807 1496 VIA_via2_5
* cell instance $17808 r0 *1 64.315,86.03
X$17808 1496 VIA_via2_5
* cell instance $17809 r0 *1 63.745,81.97
X$17809 1496 VIA_via1_4
* cell instance $17810 r0 *1 65.265,86.03
X$17810 1496 VIA_via1_4
* cell instance $17811 r0 *1 65.265,86.03
X$17811 1496 VIA_via2_5
* cell instance $17812 r0 *1 64.315,87.57
X$17812 1496 VIA_via1_4
* cell instance $17813 r0 *1 61.465,58.03
X$17813 1496 VIA_via1_4
* cell instance $17814 r0 *1 61.465,56.77
X$17814 1496 VIA_via1_4
* cell instance $17815 r0 *1 62.795,56.77
X$17815 1496 VIA_via1_4
* cell instance $17816 r0 *1 73.245,61.11
X$17816 1497 VIA_via2_5
* cell instance $17817 r0 *1 86.165,63.07
X$17817 1497 VIA_via2_5
* cell instance $17818 r0 *1 74.005,61.11
X$17818 1497 VIA_via2_5
* cell instance $17819 r0 *1 85.595,60.55
X$17819 1497 VIA_via2_5
* cell instance $17820 r0 *1 84.645,60.55
X$17820 1497 VIA_via2_5
* cell instance $17821 r0 *1 83.505,60.55
X$17821 1497 VIA_via2_5
* cell instance $17822 r0 *1 83.505,63.07
X$17822 1497 VIA_via2_5
* cell instance $17823 r0 *1 78.945,63.07
X$17823 1497 VIA_via2_5
* cell instance $17824 r0 *1 74.005,62.93
X$17824 1497 VIA_via2_5
* cell instance $17825 r0 *1 76.285,62.93
X$17825 1497 VIA_via2_5
* cell instance $17826 r0 *1 76.285,63.21
X$17826 1497 VIA_via2_5
* cell instance $17827 r0 *1 86.165,63.63
X$17827 1497 VIA_via1_4
* cell instance $17828 r0 *1 76.285,63.63
X$17828 1497 VIA_via1_4
* cell instance $17829 r0 *1 73.245,59.57
X$17829 1497 VIA_via1_4
* cell instance $17830 r0 *1 73.245,60.83
X$17830 1497 VIA_via1_4
* cell instance $17831 r0 *1 73.055,58.03
X$17831 1497 VIA_via1_4
* cell instance $17832 r0 *1 83.315,60.83
X$17832 1497 VIA_via1_4
* cell instance $17833 r0 *1 85.595,59.57
X$17833 1497 VIA_via1_4
* cell instance $17834 r0 *1 83.315,58.45
X$17834 1497 VIA_via1_4
* cell instance $17835 r0 *1 78.945,63.63
X$17835 1497 VIA_via1_4
* cell instance $17836 r0 *1 74.005,62.37
X$17836 1497 VIA_via1_4
* cell instance $17837 r0 *1 84.645,60.83
X$17837 1497 VIA_via1_4
* cell instance $17838 r0 *1 77.615,59.15
X$17838 1498 VIA_via1_4
* cell instance $17839 r0 *1 76.095,58.03
X$17839 1498 VIA_via1_4
* cell instance $17840 r0 *1 76.095,58.03
X$17840 1498 VIA_via2_5
* cell instance $17841 r0 *1 77.425,58.03
X$17841 1498 VIA_via1_4
* cell instance $17842 r0 *1 77.425,58.03
X$17842 1498 VIA_via2_5
* cell instance $17843 r0 *1 76.475,58.17
X$17843 1499 VIA_via1_4
* cell instance $17844 r0 *1 76.475,58.17
X$17844 1499 VIA_via2_5
* cell instance $17845 r0 *1 77.995,58.03
X$17845 1499 VIA_via1_4
* cell instance $17846 r0 *1 77.995,58.03
X$17846 1499 VIA_via2_5
* cell instance $17847 r0 *1 95.475,57.05
X$17847 1500 VIA_via2_5
* cell instance $17848 r0 *1 95.475,56.77
X$17848 1500 VIA_via1_4
* cell instance $17849 r0 *1 89.965,56.91
X$17849 1500 VIA_via1_4
* cell instance $17850 r0 *1 89.965,57.05
X$17850 1500 VIA_via2_5
* cell instance $17851 r0 *1 5.035,57.61
X$17851 1501 VIA_via1_7
* cell instance $17852 r0 *1 5.035,56.77
X$17852 1501 VIA_via2_5
* cell instance $17853 r0 *1 2.565,56.77
X$17853 1501 VIA_via1_4
* cell instance $17854 r0 *1 2.565,56.77
X$17854 1501 VIA_via2_5
* cell instance $17855 r0 *1 94.145,57.75
X$17855 1502 VIA_via2_5
* cell instance $17856 r0 *1 95.095,56.77
X$17856 1502 VIA_via2_5
* cell instance $17857 r0 *1 95.095,57.75
X$17857 1502 VIA_via1_4
* cell instance $17858 r0 *1 95.095,57.75
X$17858 1502 VIA_via2_5
* cell instance $17859 r0 *1 94.145,59.57
X$17859 1502 VIA_via1_4
* cell instance $17860 r0 *1 93.955,59.57
X$17860 1502 VIA_via1_4
* cell instance $17861 r0 *1 94.145,56.77
X$17861 1502 VIA_via1_4
* cell instance $17862 r0 *1 94.145,56.77
X$17862 1502 VIA_via2_5
* cell instance $17863 r0 *1 93.575,56.77
X$17863 1503 VIA_via1_4
* cell instance $17864 r0 *1 93.575,56.91
X$17864 1503 VIA_via2_5
* cell instance $17865 r0 *1 94.335,56.91
X$17865 1503 VIA_via1_4
* cell instance $17866 r0 *1 94.335,56.91
X$17866 1503 VIA_via2_5
* cell instance $17867 r0 *1 8.645,57.61
X$17867 1504 VIA_via1_7
* cell instance $17868 r0 *1 8.645,57.61
X$17868 1504 VIA_via2_5
* cell instance $17869 r0 *1 8.265,57.61
X$17869 1504 VIA_via2_5
* cell instance $17870 r0 *1 8.265,56.77
X$17870 1504 VIA_via1_4
* cell instance $17871 r0 *1 11.875,57.05
X$17871 1505 VIA_via2_5
* cell instance $17872 r0 *1 10.545,57.89
X$17872 1505 VIA_via2_5
* cell instance $17873 r0 *1 11.875,58.03
X$17873 1505 VIA_via1_4
* cell instance $17874 r0 *1 10.545,57.05
X$17874 1505 VIA_via1_4
* cell instance $17875 r0 *1 10.545,57.05
X$17875 1505 VIA_via2_5
* cell instance $17876 r0 *1 8.265,58.03
X$17876 1505 VIA_via1_4
* cell instance $17877 r0 *1 8.265,57.89
X$17877 1505 VIA_via2_5
* cell instance $17878 r0 *1 36.385,77.35
X$17878 1506 VIA_via2_5
* cell instance $17879 r0 *1 41.705,77.63
X$17879 1506 VIA_via2_5
* cell instance $17880 r0 *1 55.005,67.83
X$17880 1506 VIA_via2_5
* cell instance $17881 r0 *1 55.575,77.35
X$17881 1506 VIA_via2_5
* cell instance $17882 r0 *1 54.815,77.91
X$17882 1506 VIA_via2_5
* cell instance $17883 r0 *1 54.815,77.35
X$17883 1506 VIA_via2_5
* cell instance $17884 r0 *1 51.015,77.91
X$17884 1506 VIA_via2_5
* cell instance $17885 r0 *1 68.685,68.25
X$17885 1506 VIA_via2_5
* cell instance $17886 r0 *1 68.685,67.69
X$17886 1506 VIA_via2_5
* cell instance $17887 r0 *1 91.105,57.19
X$17887 1506 VIA_via2_5
* cell instance $17888 r0 *1 89.965,64.05
X$17888 1506 VIA_via2_5
* cell instance $17889 r0 *1 85.025,67.55
X$17889 1506 VIA_via2_5
* cell instance $17890 r0 *1 85.025,68.25
X$17890 1506 VIA_via2_5
* cell instance $17891 r0 *1 89.965,67.55
X$17891 1506 VIA_via2_5
* cell instance $17892 r0 *1 51.585,76.37
X$17892 1506 VIA_via1_4
* cell instance $17893 r0 *1 55.005,66.43
X$17893 1506 VIA_via1_4
* cell instance $17894 r0 *1 55.575,76.37
X$17894 1506 VIA_via1_4
* cell instance $17895 r0 *1 55.575,76.37
X$17895 1506 VIA_via2_5
* cell instance $17896 r0 *1 68.685,67.97
X$17896 1506 VIA_via1_4
* cell instance $17897 r0 *1 85.025,74.55
X$17897 1506 VIA_via1_4
* cell instance $17898 r0 *1 41.705,76.37
X$17898 1506 VIA_via1_4
* cell instance $17899 r0 *1 36.385,76.37
X$17899 1506 VIA_via1_4
* cell instance $17900 r0 *1 89.965,65.17
X$17900 1506 VIA_via1_4
* cell instance $17901 r0 *1 92.435,63.63
X$17901 1506 VIA_via1_4
* cell instance $17902 r0 *1 92.435,56.77
X$17902 1506 VIA_via1_4
* cell instance $17903 r0 *1 91.105,56.77
X$17903 1506 VIA_via1_4
* cell instance $17904 r0 *1 56.655,76.37
X$17904 1506 VIA_via3_2
* cell instance $17905 r0 *1 92.495,63.91
X$17905 1506 VIA_via3_2
* cell instance $17906 r0 *1 92.435,63.91
X$17906 1506 VIA_via2_5
* cell instance $17907 r0 *1 92.495,57.19
X$17907 1506 VIA_via3_2
* cell instance $17908 r0 *1 92.435,57.19
X$17908 1506 VIA_via2_5
* cell instance $17909 r0 *1 56.655,67.83
X$17909 1506 VIA_via3_2
* cell instance $17910 r0 *1 12.065,58.03
X$17910 1507 VIA_via2_5
* cell instance $17911 r0 *1 10.355,58.03
X$17911 1507 VIA_via1_4
* cell instance $17912 r0 *1 10.355,58.03
X$17912 1507 VIA_via2_5
* cell instance $17913 r0 *1 12.065,59.15
X$17913 1507 VIA_via1_4
* cell instance $17914 r0 *1 12.445,58.03
X$17914 1507 VIA_via1_4
* cell instance $17915 r0 *1 12.445,58.03
X$17915 1507 VIA_via2_5
* cell instance $17916 r0 *1 12.825,58.03
X$17916 1508 VIA_via1_4
* cell instance $17917 r0 *1 12.825,58.03
X$17917 1508 VIA_via2_5
* cell instance $17918 r0 *1 24.035,58.03
X$17918 1508 VIA_via1_4
* cell instance $17919 r0 *1 24.035,58.03
X$17919 1508 VIA_via2_5
* cell instance $17920 r0 *1 27.265,58.03
X$17920 1509 VIA_via1_4
* cell instance $17921 r0 *1 27.645,58.03
X$17921 1509 VIA_via1_4
* cell instance $17922 r0 *1 28.215,57.19
X$17922 1510 VIA_via1_7
* cell instance $17923 r0 *1 28.215,57.33
X$17923 1510 VIA_via2_5
* cell instance $17924 r0 *1 28.785,57.33
X$17924 1510 VIA_via2_5
* cell instance $17925 r0 *1 28.785,58.03
X$17925 1510 VIA_via1_4
* cell instance $17926 r0 *1 31.825,66.57
X$17926 1511 VIA_via1_7
* cell instance $17927 r0 *1 55.575,57.19
X$17927 1511 VIA_via1_7
* cell instance $17928 r0 *1 55.575,57.33
X$17928 1511 VIA_via2_5
* cell instance $17929 r0 *1 36.765,77.21
X$17929 1511 VIA_via2_5
* cell instance $17930 r0 *1 29.925,77.21
X$17930 1511 VIA_via2_5
* cell instance $17931 r0 *1 41.895,77.35
X$17931 1511 VIA_via2_5
* cell instance $17932 r0 *1 52.915,67.41
X$17932 1511 VIA_via2_5
* cell instance $17933 r0 *1 54.245,67.55
X$17933 1511 VIA_via2_5
* cell instance $17934 r0 *1 52.725,57.33
X$17934 1511 VIA_via2_5
* cell instance $17935 r0 *1 32.015,57.33
X$17935 1511 VIA_via2_5
* cell instance $17936 r0 *1 29.925,57.33
X$17936 1511 VIA_via2_5
* cell instance $17937 r0 *1 51.205,77.63
X$17937 1511 VIA_via1_4
* cell instance $17938 r0 *1 51.205,77.49
X$17938 1511 VIA_via2_5
* cell instance $17939 r0 *1 55.765,77.63
X$17939 1511 VIA_via1_4
* cell instance $17940 r0 *1 55.765,77.49
X$17940 1511 VIA_via2_5
* cell instance $17941 r0 *1 54.245,67.97
X$17941 1511 VIA_via1_4
* cell instance $17942 r0 *1 41.895,77.63
X$17942 1511 VIA_via1_4
* cell instance $17943 r0 *1 29.925,56.77
X$17943 1511 VIA_via1_4
* cell instance $17944 r0 *1 29.925,77.63
X$17944 1511 VIA_via1_4
* cell instance $17945 r0 *1 36.765,77.63
X$17945 1511 VIA_via1_4
* cell instance $17946 r0 *1 36.775,77.63
X$17946 1511 VIA_via3_2
* cell instance $17947 r0 *1 36.765,77.63
X$17947 1511 VIA_via2_5
* cell instance $17948 r0 *1 29.735,76.37
X$17948 1511 VIA_via1_4
* cell instance $17949 r0 *1 29.735,76.37
X$17949 1511 VIA_via2_5
* cell instance $17950 r0 *1 29.775,76.37
X$17950 1511 VIA_via3_2
* cell instance $17951 r0 *1 29.735,73.57
X$17951 1511 VIA_via1_4
* cell instance $17952 r0 *1 29.735,73.71
X$17952 1511 VIA_via2_5
* cell instance $17953 r0 *1 29.775,73.71
X$17953 1511 VIA_via3_2
* cell instance $17954 r0 *1 42.095,77.07
X$17954 1511 VIA_via4_0
* cell instance $17955 r0 *1 36.775,77.07
X$17955 1511 VIA_via4_0
* cell instance $17956 r0 *1 51.055,77.07
X$17956 1511 VIA_via4_0
* cell instance $17957 r0 *1 42.095,77.35
X$17957 1511 VIA_via3_2
* cell instance $17958 r0 *1 53.295,67.41
X$17958 1511 VIA_via3_2
* cell instance $17959 r0 *1 51.055,77.49
X$17959 1511 VIA_via3_2
* cell instance $17960 r0 *1 53.295,77.49
X$17960 1511 VIA_via3_2
* cell instance $17961 r0 *1 27.835,58.03
X$17961 1512 VIA_via1_4
* cell instance $17962 r0 *1 27.835,58.03
X$17962 1512 VIA_via2_5
* cell instance $17963 r0 *1 29.735,58.03
X$17963 1512 VIA_via1_4
* cell instance $17964 r0 *1 29.735,58.03
X$17964 1512 VIA_via2_5
* cell instance $17965 r0 *1 29.735,56.63
X$17965 1513 VIA_via1_7
* cell instance $17966 r0 *1 29.355,59.57
X$17966 1513 VIA_via1_4
* cell instance $17967 r0 *1 29.735,57.75
X$17967 1513 VIA_via1_4
* cell instance $17968 r0 *1 29.165,58.31
X$17968 1513 VIA_via1_4
* cell instance $17969 r0 *1 29.545,58.03
X$17969 1514 VIA_via1_4
* cell instance $17970 r0 *1 29.545,57.89
X$17970 1514 VIA_via2_5
* cell instance $17971 r0 *1 24.225,57.89
X$17971 1514 VIA_via1_4
* cell instance $17972 r0 *1 24.225,57.89
X$17972 1514 VIA_via2_5
* cell instance $17973 r0 *1 89.965,57.33
X$17973 1515 VIA_via2_5
* cell instance $17974 r0 *1 85.405,57.33
X$17974 1515 VIA_via2_5
* cell instance $17975 r0 *1 89.965,62.37
X$17975 1515 VIA_via1_4
* cell instance $17976 r0 *1 85.405,55.51
X$17976 1515 VIA_via1_4
* cell instance $17977 r0 *1 86.925,56.77
X$17977 1516 VIA_via1_4
* cell instance $17978 r0 *1 86.925,56.91
X$17978 1516 VIA_via2_5
* cell instance $17979 r0 *1 87.875,56.91
X$17979 1516 VIA_via1_4
* cell instance $17980 r0 *1 87.875,56.91
X$17980 1516 VIA_via2_5
* cell instance $17981 r0 *1 30.685,58.03
X$17981 1517 VIA_via1_4
* cell instance $17982 r0 *1 30.685,58.03
X$17982 1517 VIA_via2_5
* cell instance $17983 r0 *1 34.295,58.03
X$17983 1517 VIA_via1_4
* cell instance $17984 r0 *1 34.295,58.03
X$17984 1517 VIA_via2_5
* cell instance $17985 r0 *1 86.165,56.77
X$17985 1518 VIA_via1_4
* cell instance $17986 r0 *1 86.165,56.77
X$17986 1518 VIA_via2_5
* cell instance $17987 r0 *1 87.305,56.77
X$17987 1518 VIA_via1_4
* cell instance $17988 r0 *1 87.305,56.77
X$17988 1518 VIA_via2_5
* cell instance $17989 r0 *1 80.655,76.37
X$17989 1519 VIA_via1_7
* cell instance $17990 r0 *1 80.655,78.61
X$17990 1519 VIA_via1_7
* cell instance $17991 r0 *1 80.655,77.21
X$17991 1519 VIA_via2_5
* cell instance $17992 r0 *1 56.715,58.73
X$17992 1519 VIA_via2_5
* cell instance $17993 r0 *1 56.905,77.35
X$17993 1519 VIA_via2_5
* cell instance $17994 r0 *1 83.315,56.91
X$17994 1519 VIA_via2_5
* cell instance $17995 r0 *1 80.655,65.17
X$17995 1519 VIA_via2_5
* cell instance $17996 r0 *1 81.795,65.17
X$17996 1519 VIA_via2_5
* cell instance $17997 r0 *1 56.905,77.63
X$17997 1519 VIA_via1_4
* cell instance $17998 r0 *1 56.715,55.23
X$17998 1519 VIA_via1_4
* cell instance $17999 r0 *1 81.415,65.17
X$17999 1519 VIA_via1_4
* cell instance $18000 r0 *1 81.415,65.17
X$18000 1519 VIA_via2_5
* cell instance $18001 r0 *1 82.175,56.77
X$18001 1519 VIA_via1_4
* cell instance $18002 r0 *1 82.175,56.91
X$18002 1519 VIA_via2_5
* cell instance $18003 r0 *1 83.315,55.23
X$18003 1519 VIA_via1_4
* cell instance $18004 r0 *1 57.215,77.35
X$18004 1519 VIA_via3_2
* cell instance $18005 r0 *1 57.215,58.73
X$18005 1519 VIA_via3_2
* cell instance $18006 r0 *1 81.605,57.19
X$18006 1520 VIA_via1_7
* cell instance $18007 r0 *1 81.605,57.33
X$18007 1520 VIA_via2_5
* cell instance $18008 r0 *1 80.275,57.33
X$18008 1520 VIA_via2_5
* cell instance $18009 r0 *1 80.275,56.77
X$18009 1520 VIA_via1_4
* cell instance $18010 r0 *1 81.985,56.77
X$18010 1521 VIA_via1_4
* cell instance $18011 r0 *1 81.985,56.77
X$18011 1521 VIA_via2_5
* cell instance $18012 r0 *1 81.035,56.77
X$18012 1521 VIA_via1_4
* cell instance $18013 r0 *1 81.035,56.77
X$18013 1521 VIA_via2_5
* cell instance $18014 r0 *1 43.225,57.61
X$18014 1522 VIA_via1_7
* cell instance $18015 r0 *1 43.225,56.77
X$18015 1522 VIA_via2_5
* cell instance $18016 r0 *1 39.425,56.77
X$18016 1522 VIA_via1_4
* cell instance $18017 r0 *1 39.425,56.77
X$18017 1522 VIA_via2_5
* cell instance $18018 r0 *1 47.405,57.61
X$18018 1523 VIA_via1_7
* cell instance $18019 r0 *1 47.405,56.77
X$18019 1523 VIA_via2_5
* cell instance $18020 r0 *1 44.365,56.77
X$18020 1523 VIA_via1_4
* cell instance $18021 r0 *1 44.365,56.77
X$18021 1523 VIA_via2_5
* cell instance $18022 r0 *1 78.185,54.39
X$18022 1524 VIA_via1_7
* cell instance $18023 r0 *1 78.185,56.77
X$18023 1524 VIA_via1_4
* cell instance $18024 r0 *1 52.535,58.03
X$18024 1525 VIA_via2_5
* cell instance $18025 r0 *1 52.535,60.83
X$18025 1525 VIA_via1_4
* cell instance $18026 r0 *1 52.535,59.15
X$18026 1525 VIA_via1_4
* cell instance $18027 r0 *1 50.445,58.03
X$18027 1525 VIA_via1_4
* cell instance $18028 r0 *1 50.445,58.03
X$18028 1525 VIA_via2_5
* cell instance $18029 r0 *1 74.005,57.61
X$18029 1526 VIA_via1_7
* cell instance $18030 r0 *1 74.005,57.61
X$18030 1526 VIA_via2_5
* cell instance $18031 r0 *1 72.865,57.61
X$18031 1526 VIA_via2_5
* cell instance $18032 r0 *1 72.865,56.77
X$18032 1526 VIA_via1_4
* cell instance $18033 r0 *1 70.205,56.77
X$18033 1527 VIA_via1_4
* cell instance $18034 r0 *1 70.015,56.77
X$18034 1527 VIA_via1_4
* cell instance $18035 r0 *1 60.705,56.77
X$18035 1528 VIA_via1_4
* cell instance $18036 r0 *1 60.705,56.77
X$18036 1528 VIA_via2_5
* cell instance $18037 r0 *1 62.035,56.77
X$18037 1528 VIA_via1_4
* cell instance $18038 r0 *1 62.035,56.77
X$18038 1528 VIA_via2_5
* cell instance $18039 r0 *1 62.035,58.03
X$18039 1529 VIA_via1_4
* cell instance $18040 r0 *1 62.225,58.03
X$18040 1529 VIA_via1_4
* cell instance $18041 r0 *1 22.325,84.63
X$18041 1530 VIA_via1_7
* cell instance $18042 r0 *1 50.255,60.97
X$18042 1530 VIA_via1_7
* cell instance $18043 r0 *1 37.525,84.63
X$18043 1530 VIA_via1_7
* cell instance $18044 r0 *1 48.165,80.57
X$18044 1530 VIA_via1_7
* cell instance $18045 r0 *1 48.165,80.57
X$18045 1530 VIA_via2_5
* cell instance $18046 r0 *1 22.325,58.17
X$18046 1530 VIA_via1_7
* cell instance $18047 r0 *1 57.665,81.83
X$18047 1530 VIA_via1_7
* cell instance $18048 r0 *1 12.255,59.43
X$18048 1530 VIA_via1_7
* cell instance $18049 r0 *1 12.255,59.15
X$18049 1530 VIA_via2_5
* cell instance $18050 r0 *1 11.875,77.35
X$18050 1530 VIA_via2_5
* cell instance $18051 r0 *1 13.205,77.35
X$18051 1530 VIA_via2_5
* cell instance $18052 r0 *1 22.325,83.23
X$18052 1530 VIA_via2_5
* cell instance $18053 r0 *1 22.325,82.11
X$18053 1530 VIA_via2_5
* cell instance $18054 r0 *1 10.925,77.35
X$18054 1530 VIA_via2_5
* cell instance $18055 r0 *1 11.115,70.91
X$18055 1530 VIA_via2_5
* cell instance $18056 r0 *1 12.255,70.91
X$18056 1530 VIA_via2_5
* cell instance $18057 r0 *1 37.335,83.37
X$18057 1530 VIA_via2_5
* cell instance $18058 r0 *1 48.545,80.57
X$18058 1530 VIA_via2_5
* cell instance $18059 r0 *1 37.335,82.11
X$18059 1530 VIA_via2_5
* cell instance $18060 r0 *1 48.545,82.39
X$18060 1530 VIA_via2_5
* cell instance $18061 r0 *1 50.445,61.11
X$18061 1530 VIA_via2_5
* cell instance $18062 r0 *1 57.665,80.57
X$18062 1530 VIA_via2_5
* cell instance $18063 r0 *1 22.325,59.01
X$18063 1530 VIA_via2_5
* cell instance $18064 r0 *1 57.665,80.85
X$18064 1530 VIA_via1_4
* cell instance $18065 r0 *1 27.835,83.23
X$18065 1530 VIA_via1_4
* cell instance $18066 r0 *1 27.835,83.23
X$18066 1530 VIA_via2_5
* cell instance $18067 r0 *1 11.875,77.63
X$18067 1530 VIA_via1_4
* cell instance $18068 r0 *1 13.015,81.97
X$18068 1530 VIA_via1_4
* cell instance $18069 r0 *1 13.015,82.11
X$18069 1530 VIA_via2_5
* cell instance $18070 r0 *1 51.615,80.57
X$18070 1530 VIA_via3_2
* cell instance $18071 r0 *1 51.615,61.11
X$18071 1530 VIA_via3_2
* cell instance $18072 r0 *1 13.015,59.57
X$18072 1531 VIA_via1_4
* cell instance $18073 r0 *1 13.015,59.57
X$18073 1531 VIA_via2_5
* cell instance $18074 r0 *1 16.625,59.57
X$18074 1531 VIA_via1_4
* cell instance $18075 r0 *1 16.625,59.57
X$18075 1531 VIA_via2_5
* cell instance $18076 r0 *1 18.905,59.57
X$18076 1531 VIA_via1_4
* cell instance $18077 r0 *1 18.905,59.57
X$18077 1531 VIA_via2_5
* cell instance $18078 r0 *1 9.025,62.79
X$18078 1532 VIA_via1_7
* cell instance $18079 r0 *1 9.025,62.37
X$18079 1532 VIA_via2_5
* cell instance $18080 r0 *1 14.725,68.11
X$18080 1532 VIA_via2_5
* cell instance $18081 r0 *1 8.455,68.11
X$18081 1532 VIA_via2_5
* cell instance $18082 r0 *1 17.195,62.37
X$18082 1532 VIA_via2_5
* cell instance $18083 r0 *1 14.725,63.77
X$18083 1532 VIA_via2_5
* cell instance $18084 r0 *1 23.655,62.65
X$18084 1532 VIA_via2_5
* cell instance $18085 r0 *1 23.655,62.37
X$18085 1532 VIA_via1_4
* cell instance $18086 r0 *1 24.035,63.63
X$18086 1532 VIA_via1_4
* cell instance $18087 r0 *1 19.475,62.37
X$18087 1532 VIA_via1_4
* cell instance $18088 r0 *1 19.475,62.37
X$18088 1532 VIA_via2_5
* cell instance $18089 r0 *1 13.395,67.97
X$18089 1532 VIA_via1_4
* cell instance $18090 r0 *1 13.395,68.11
X$18090 1532 VIA_via2_5
* cell instance $18091 r0 *1 14.725,65.17
X$18091 1532 VIA_via1_4
* cell instance $18092 r0 *1 17.195,63.63
X$18092 1532 VIA_via1_4
* cell instance $18093 r0 *1 17.195,63.77
X$18093 1532 VIA_via2_5
* cell instance $18094 r0 *1 10.165,62.37
X$18094 1532 VIA_via1_4
* cell instance $18095 r0 *1 10.165,62.37
X$18095 1532 VIA_via2_5
* cell instance $18096 r0 *1 17.005,59.57
X$18096 1532 VIA_via1_4
* cell instance $18097 r0 *1 11.495,67.97
X$18097 1532 VIA_via1_4
* cell instance $18098 r0 *1 11.495,68.11
X$18098 1532 VIA_via2_5
* cell instance $18099 r0 *1 8.455,69.23
X$18099 1532 VIA_via1_4
* cell instance $18100 r0 *1 19.475,59.43
X$18100 1533 VIA_via2_5
* cell instance $18101 r0 *1 18.335,59.57
X$18101 1533 VIA_via1_4
* cell instance $18102 r0 *1 18.335,59.43
X$18102 1533 VIA_via2_5
* cell instance $18103 r0 *1 17.575,59.57
X$18103 1533 VIA_via1_4
* cell instance $18104 r0 *1 17.575,59.43
X$18104 1533 VIA_via2_5
* cell instance $18105 r0 *1 19.475,58.45
X$18105 1533 VIA_via1_4
* cell instance $18106 r0 *1 25.365,59.15
X$18106 1534 VIA_via2_5
* cell instance $18107 r0 *1 26.315,59.15
X$18107 1534 VIA_via2_5
* cell instance $18108 r0 *1 27.455,59.15
X$18108 1534 VIA_via1_4
* cell instance $18109 r0 *1 27.455,59.15
X$18109 1534 VIA_via2_5
* cell instance $18110 r0 *1 26.315,58.03
X$18110 1534 VIA_via1_4
* cell instance $18111 r0 *1 25.365,58.03
X$18111 1534 VIA_via1_4
* cell instance $18112 r0 *1 10.925,65.73
X$18112 1535 VIA_via2_5
* cell instance $18113 r0 *1 33.345,91.35
X$18113 1535 VIA_via2_5
* cell instance $18114 r0 *1 15.485,64.61
X$18114 1535 VIA_via2_5
* cell instance $18115 r0 *1 11.115,90.65
X$18115 1535 VIA_via2_5
* cell instance $18116 r0 *1 15.485,65.73
X$18116 1535 VIA_via2_5
* cell instance $18117 r0 *1 18.715,90.65
X$18117 1535 VIA_via2_5
* cell instance $18118 r0 *1 55.955,59.43
X$18118 1535 VIA_via2_5
* cell instance $18119 r0 *1 52.155,91.35
X$18119 1535 VIA_via2_5
* cell instance $18120 r0 *1 67.545,59.29
X$18120 1535 VIA_via2_5
* cell instance $18121 r0 *1 57.285,84.35
X$18121 1535 VIA_via2_5
* cell instance $18122 r0 *1 39.995,91.35
X$18122 1535 VIA_via2_5
* cell instance $18123 r0 *1 57.285,84.77
X$18123 1535 VIA_via1_4
* cell instance $18124 r0 *1 52.155,91.63
X$18124 1535 VIA_via1_4
* cell instance $18125 r0 *1 39.425,59.57
X$18125 1535 VIA_via1_4
* cell instance $18126 r0 *1 39.425,59.57
X$18126 1535 VIA_via2_5
* cell instance $18127 r0 *1 18.905,90.37
X$18127 1535 VIA_via1_4
* cell instance $18128 r0 *1 39.995,90.37
X$18128 1535 VIA_via1_4
* cell instance $18129 r0 *1 33.345,91.63
X$18129 1535 VIA_via1_4
* cell instance $18130 r0 *1 10.925,65.17
X$18130 1535 VIA_via1_4
* cell instance $18131 r0 *1 11.115,90.37
X$18131 1535 VIA_via1_4
* cell instance $18132 r0 *1 12.825,81.97
X$18132 1535 VIA_via1_4
* cell instance $18133 r0 *1 12.825,81.97
X$18133 1535 VIA_via2_5
* cell instance $18134 r0 *1 67.545,59.57
X$18134 1535 VIA_via1_4
* cell instance $18135 r0 *1 56.095,84.35
X$18135 1535 VIA_via4_0
* cell instance $18136 r0 *1 56.095,84.35
X$18136 1535 VIA_via3_2
* cell instance $18137 r0 *1 56.095,84.35
X$18137 1535 VIA_via5_0
* cell instance $18138 r0 *1 55.815,91.35
X$18138 1535 VIA_via3_2
* cell instance $18139 r0 *1 14.655,90.65
X$18139 1535 VIA_via3_2
* cell instance $18140 r0 *1 14.655,81.97
X$18140 1535 VIA_via3_2
* cell instance $18141 r0 *1 56.095,63.63
X$18141 1535 VIA_via3_2
* cell instance $18142 r0 *1 56.095,63.63
X$18142 1535 VIA_via4_0
* cell instance $18143 r0 *1 56.095,63.63
X$18143 1535 VIA_via5_0
* cell instance $18144 r0 *1 56.145,63.63
X$18144 1535 VIA_via2_5
* cell instance $18145 r0 *1 56.145,63.63
X$18145 1535 VIA_via1_4
* cell instance $18146 r0 *1 55.535,59.43
X$18146 1535 VIA_via3_2
* cell instance $18147 r0 *1 55.535,59.43
X$18147 1535 VIA_via4_0
* cell instance $18148 r0 *1 39.575,59.57
X$18148 1535 VIA_via3_2
* cell instance $18149 r0 *1 39.575,59.43
X$18149 1535 VIA_via4_0
* cell instance $18150 r0 *1 39.015,64.61
X$18150 1535 VIA_via3_2
* cell instance $18151 r0 *1 39.015,59.57
X$18151 1535 VIA_via3_2
* cell instance $18152 r0 *1 50.775,91.21
X$18152 1535 VIA_via3_2
* cell instance $18153 r0 *1 50.775,91.35
X$18153 1535 VIA_via4_0
* cell instance $18154 r0 *1 41.815,91.35
X$18154 1535 VIA_via3_2
* cell instance $18155 r0 *1 41.815,91.35
X$18155 1535 VIA_via4_0
* cell instance $18156 r0 *1 14.655,65.73
X$18156 1535 VIA_via3_2
* cell instance $18157 r0 *1 45.125,59.15
X$18157 1536 VIA_via2_5
* cell instance $18158 r0 *1 48.925,59.15
X$18158 1536 VIA_via2_5
* cell instance $18159 r0 *1 45.125,58.03
X$18159 1536 VIA_via1_4
* cell instance $18160 r0 *1 47.785,59.15
X$18160 1536 VIA_via1_4
* cell instance $18161 r0 *1 47.785,59.15
X$18161 1536 VIA_via2_5
* cell instance $18162 r0 *1 48.735,60.83
X$18162 1536 VIA_via1_4
* cell instance $18163 r0 *1 38.455,76.07
X$18163 1537 VIA_via6_0
* cell instance $18164 r0 *1 49.375,76.07
X$18164 1537 VIA_via6_0
* cell instance $18165 r0 *1 38.455,77.35
X$18165 1537 VIA_via5_0
* cell instance $18166 r0 *1 38.455,77.35
X$18166 1537 VIA_via4_0
* cell instance $18167 r0 *1 38.455,77.49
X$18167 1537 VIA_via3_2
* cell instance $18168 r0 *1 19.665,77.49
X$18168 1537 VIA_via2_5
* cell instance $18169 r0 *1 60.325,67.13
X$18169 1537 VIA_via2_5
* cell instance $18170 r0 *1 60.325,59.85
X$18170 1537 VIA_via2_5
* cell instance $18171 r0 *1 54.625,59.85
X$18171 1537 VIA_via2_5
* cell instance $18172 r0 *1 54.435,59.15
X$18172 1537 VIA_via2_5
* cell instance $18173 r0 *1 70.015,67.13
X$18173 1537 VIA_via2_5
* cell instance $18174 r0 *1 70.015,68.53
X$18174 1537 VIA_via2_5
* cell instance $18175 r0 *1 78.945,68.81
X$18175 1537 VIA_via2_5
* cell instance $18176 r0 *1 49.685,76.37
X$18176 1537 VIA_via1_4
* cell instance $18177 r0 *1 49.685,76.23
X$18177 1537 VIA_via2_5
* cell instance $18178 r0 *1 70.015,67.97
X$18178 1537 VIA_via1_4
* cell instance $18179 r0 *1 38.285,77.63
X$18179 1537 VIA_via1_4
* cell instance $18180 r0 *1 38.285,77.49
X$18180 1537 VIA_via2_5
* cell instance $18181 r0 *1 35.055,59.15
X$18181 1537 VIA_via1_4
* cell instance $18182 r0 *1 35.055,59.15
X$18182 1537 VIA_via2_5
* cell instance $18183 r0 *1 35.095,59.15
X$18183 1537 VIA_via3_2
* cell instance $18184 r0 *1 35.095,59.15
X$18184 1537 VIA_via4_0
* cell instance $18185 r0 *1 35.055,77.63
X$18185 1537 VIA_via1_4
* cell instance $18186 r0 *1 35.055,77.63
X$18186 1537 VIA_via2_5
* cell instance $18187 r0 *1 27.265,77.63
X$18187 1537 VIA_via1_4
* cell instance $18188 r0 *1 27.265,77.63
X$18188 1537 VIA_via2_5
* cell instance $18189 r0 *1 27.255,77.63
X$18189 1537 VIA_via3_2
* cell instance $18190 r0 *1 20.235,77.63
X$18190 1537 VIA_via1_4
* cell instance $18191 r0 *1 20.235,77.49
X$18191 1537 VIA_via2_5
* cell instance $18192 r0 *1 19.665,79.17
X$18192 1537 VIA_via1_4
* cell instance $18193 r0 *1 78.945,69.23
X$18193 1537 VIA_via1_4
* cell instance $18194 r0 *1 54.625,59.57
X$18194 1537 VIA_via1_4
* cell instance $18195 r0 *1 34.535,76.79
X$18195 1537 VIA_via4_0
* cell instance $18196 r0 *1 36.495,77.35
X$18196 1537 VIA_via4_0
* cell instance $18197 r0 *1 49.375,76.23
X$18197 1537 VIA_via4_0
* cell instance $18198 r0 *1 49.375,76.23
X$18198 1537 VIA_via5_0
* cell instance $18199 r0 *1 49.375,76.23
X$18199 1537 VIA_via3_2
* cell instance $18200 r0 *1 54.695,76.23
X$18200 1537 VIA_via4_0
* cell instance $18201 r0 *1 54.695,76.37
X$18201 1537 VIA_via3_2
* cell instance $18202 r0 *1 54.815,76.37
X$18202 1537 VIA_via2_5
* cell instance $18203 r0 *1 54.815,76.37
X$18203 1537 VIA_via1_4
* cell instance $18204 r0 *1 27.255,76.79
X$18204 1537 VIA_via4_0
* cell instance $18205 r0 *1 36.215,77.63
X$18205 1537 VIA_via3_2
* cell instance $18206 r0 *1 34.535,77.63
X$18206 1537 VIA_via3_2
* cell instance $18207 r0 *1 54.135,59.15
X$18207 1537 VIA_via3_2
* cell instance $18208 r0 *1 54.135,59.15
X$18208 1537 VIA_via4_0
* cell instance $18209 r0 *1 74.005,59.71
X$18209 1538 VIA_via2_5
* cell instance $18210 r0 *1 72.295,59.29
X$18210 1538 VIA_via1_4
* cell instance $18211 r0 *1 72.675,59.57
X$18211 1538 VIA_via1_4
* cell instance $18212 r0 *1 72.675,59.71
X$18212 1538 VIA_via2_5
* cell instance $18213 r0 *1 74.005,60.83
X$18213 1538 VIA_via1_4
* cell instance $18214 r0 *1 78.375,58.59
X$18214 1539 VIA_via1_7
* cell instance $18215 r0 *1 78.755,62.37
X$18215 1539 VIA_via1_4
* cell instance $18216 r0 *1 79.895,60.69
X$18216 1540 VIA_via2_5
* cell instance $18217 r0 *1 82.365,60.69
X$18217 1540 VIA_via1_4
* cell instance $18218 r0 *1 82.365,60.69
X$18218 1540 VIA_via2_5
* cell instance $18219 r0 *1 80.085,59.57
X$18219 1540 VIA_via1_4
* cell instance $18220 r0 *1 79.895,62.37
X$18220 1540 VIA_via1_4
* cell instance $18221 r0 *1 92.625,59.29
X$18221 1541 VIA_via2_5
* cell instance $18222 r0 *1 92.815,58.03
X$18222 1541 VIA_via1_4
* cell instance $18223 r0 *1 93.195,59.29
X$18223 1541 VIA_via1_4
* cell instance $18224 r0 *1 93.195,59.29
X$18224 1541 VIA_via2_5
* cell instance $18225 r0 *1 94.905,59.01
X$18225 1542 VIA_via1_7
* cell instance $18226 r0 *1 94.905,59.01
X$18226 1542 VIA_via2_5
* cell instance $18227 r0 *1 95.285,59.01
X$18227 1542 VIA_via2_5
* cell instance $18228 r0 *1 95.285,56.77
X$18228 1542 VIA_via1_4
* cell instance $18229 r0 *1 93.385,59.15
X$18229 1543 VIA_via2_5
* cell instance $18230 r0 *1 93.385,59.57
X$18230 1543 VIA_via1_4
* cell instance $18231 r0 *1 94.335,59.15
X$18231 1543 VIA_via1_4
* cell instance $18232 r0 *1 94.335,59.15
X$18232 1543 VIA_via2_5
* cell instance $18233 r0 *1 18.525,80.57
X$18233 1544 VIA_via1_7
* cell instance $18234 r0 *1 18.525,80.71
X$18234 1544 VIA_via2_5
* cell instance $18235 r0 *1 45.125,79.03
X$18235 1544 VIA_via1_7
* cell instance $18236 r0 *1 9.975,62.23
X$18236 1544 VIA_via1_7
* cell instance $18237 r0 *1 7.505,58.17
X$18237 1544 VIA_via1_7
* cell instance $18238 r0 *1 45.125,80.15
X$18238 1544 VIA_via2_5
* cell instance $18239 r0 *1 7.505,58.73
X$18239 1544 VIA_via2_5
* cell instance $18240 r0 *1 9.595,58.73
X$18240 1544 VIA_via2_5
* cell instance $18241 r0 *1 34.105,80.71
X$18241 1544 VIA_via2_5
* cell instance $18242 r0 *1 7.505,80.71
X$18242 1544 VIA_via2_5
* cell instance $18243 r0 *1 9.595,61.39
X$18243 1544 VIA_via2_5
* cell instance $18244 r0 *1 40.565,80.15
X$18244 1544 VIA_via2_5
* cell instance $18245 r0 *1 40.565,80.71
X$18245 1544 VIA_via2_5
* cell instance $18246 r0 *1 51.395,80.15
X$18246 1544 VIA_via2_5
* cell instance $18247 r0 *1 45.885,61.11
X$18247 1544 VIA_via2_5
* cell instance $18248 r0 *1 45.505,61.11
X$18248 1544 VIA_via2_5
* cell instance $18249 r0 *1 51.395,80.43
X$18249 1544 VIA_via1_4
* cell instance $18250 r0 *1 45.505,60.83
X$18250 1544 VIA_via1_4
* cell instance $18251 r0 *1 45.505,60.69
X$18251 1544 VIA_via2_5
* cell instance $18252 r0 *1 40.565,80.43
X$18252 1544 VIA_via1_4
* cell instance $18253 r0 *1 34.105,83.23
X$18253 1544 VIA_via1_4
* cell instance $18254 r0 *1 7.505,81.97
X$18254 1544 VIA_via1_4
* cell instance $18255 r0 *1 7.695,76.37
X$18255 1544 VIA_via1_4
* cell instance $18256 r0 *1 52.155,58.45
X$18256 1544 VIA_via1_4
* cell instance $18257 r0 *1 52.155,58.45
X$18257 1544 VIA_via2_5
* cell instance $18258 r0 *1 50.495,60.83
X$18258 1544 VIA_via4_0
* cell instance $18259 r0 *1 45.735,60.69
X$18259 1544 VIA_via3_2
* cell instance $18260 r0 *1 45.735,60.83
X$18260 1544 VIA_via4_0
* cell instance $18261 r0 *1 50.495,58.45
X$18261 1544 VIA_via3_2
* cell instance $18262 r0 *1 10.735,58.59
X$18262 1545 VIA_via1_7
* cell instance $18263 r0 *1 9.785,59.15
X$18263 1545 VIA_via2_5
* cell instance $18264 r0 *1 10.735,59.15
X$18264 1545 VIA_via2_5
* cell instance $18265 r0 *1 9.785,59.57
X$18265 1545 VIA_via1_4
* cell instance $18266 r0 *1 17.955,59.01
X$18266 1546 VIA_via1_7
* cell instance $18267 r0 *1 17.955,59.01
X$18267 1546 VIA_via2_5
* cell instance $18268 r0 *1 17.195,59.01
X$18268 1546 VIA_via2_5
* cell instance $18269 r0 *1 17.195,58.03
X$18269 1546 VIA_via1_4
* cell instance $18270 r0 *1 25.745,58.59
X$18270 1547 VIA_via1_7
* cell instance $18271 r0 *1 25.175,59.29
X$18271 1547 VIA_via2_5
* cell instance $18272 r0 *1 25.745,59.29
X$18272 1547 VIA_via2_5
* cell instance $18273 r0 *1 25.175,59.57
X$18273 1547 VIA_via1_4
* cell instance $18274 r0 *1 77.805,58.59
X$18274 1548 VIA_via1_7
* cell instance $18275 r0 *1 77.805,58.59
X$18275 1548 VIA_via2_5
* cell instance $18276 r0 *1 75.335,58.59
X$18276 1548 VIA_via2_5
* cell instance $18277 r0 *1 75.335,59.57
X$18277 1548 VIA_via1_4
* cell instance $18278 r0 *1 40.945,59.01
X$18278 1549 VIA_via1_7
* cell instance $18279 r0 *1 40.945,59.01
X$18279 1549 VIA_via2_5
* cell instance $18280 r0 *1 39.615,59.01
X$18280 1549 VIA_via2_5
* cell instance $18281 r0 *1 39.615,58.03
X$18281 1549 VIA_via1_4
* cell instance $18282 r0 *1 53.105,59.29
X$18282 1550 VIA_via2_5
* cell instance $18283 r0 *1 53.295,60.69
X$18283 1550 VIA_via2_5
* cell instance $18284 r0 *1 43.985,59.15
X$18284 1550 VIA_via1_4
* cell instance $18285 r0 *1 43.985,59.29
X$18285 1550 VIA_via2_5
* cell instance $18286 r0 *1 54.055,60.83
X$18286 1550 VIA_via1_4
* cell instance $18287 r0 *1 54.055,60.83
X$18287 1550 VIA_via2_5
* cell instance $18288 r0 *1 49.115,60.41
X$18288 1551 VIA_via1_7
* cell instance $18289 r0 *1 53.295,59.15
X$18289 1551 VIA_via2_5
* cell instance $18290 r0 *1 49.305,59.15
X$18290 1551 VIA_via2_5
* cell instance $18291 r0 *1 53.295,59.57
X$18291 1551 VIA_via1_4
* cell instance $18292 r0 *1 44.365,59.01
X$18292 1552 VIA_via1_7
* cell instance $18293 r0 *1 44.365,58.87
X$18293 1552 VIA_via2_5
* cell instance $18294 r0 *1 48.735,58.87
X$18294 1552 VIA_via2_5
* cell instance $18295 r0 *1 48.735,52.43
X$18295 1552 VIA_via1_4
* cell instance $18296 r0 *1 50.825,58.59
X$18296 1553 VIA_via1_7
* cell instance $18297 r0 *1 50.825,58.59
X$18297 1553 VIA_via2_5
* cell instance $18298 r0 *1 50.255,58.59
X$18298 1553 VIA_via2_5
* cell instance $18299 r0 *1 50.255,59.57
X$18299 1553 VIA_via1_4
* cell instance $18300 r0 *1 46.075,58.59
X$18300 1554 VIA_via1_7
* cell instance $18301 r0 *1 46.075,58.59
X$18301 1554 VIA_via2_5
* cell instance $18302 r0 *1 45.505,58.59
X$18302 1554 VIA_via2_5
* cell instance $18303 r0 *1 45.505,59.57
X$18303 1554 VIA_via1_4
* cell instance $18304 r0 *1 2.755,61.11
X$18304 1555 VIA_via2_5
* cell instance $18305 r0 *1 2.755,60.83
X$18305 1555 VIA_via1_4
* cell instance $18306 r0 *1 1.495,61.11
X$18306 1555 VIA_via3_2
* cell instance $18307 r0 *1 1.495,61.11
X$18307 1555 VIA_via4_0
* cell instance $18308 r0 *1 4.275,65.17
X$18308 1556 VIA_via2_5
* cell instance $18309 r0 *1 5.035,63.49
X$18309 1556 VIA_via2_5
* cell instance $18310 r0 *1 6.365,66.43
X$18310 1556 VIA_via2_5
* cell instance $18311 r0 *1 8.835,67.97
X$18311 1556 VIA_via1_4
* cell instance $18312 r0 *1 8.645,66.43
X$18312 1556 VIA_via1_4
* cell instance $18313 r0 *1 8.645,66.43
X$18313 1556 VIA_via2_5
* cell instance $18314 r0 *1 6.555,63.63
X$18314 1556 VIA_via1_4
* cell instance $18315 r0 *1 6.555,63.49
X$18315 1556 VIA_via2_5
* cell instance $18316 r0 *1 4.845,60.83
X$18316 1556 VIA_via1_4
* cell instance $18317 r0 *1 3.515,69.23
X$18317 1556 VIA_via1_4
* cell instance $18318 r0 *1 4.085,70.77
X$18318 1556 VIA_via1_4
* cell instance $18319 r0 *1 6.365,66.15
X$18319 1556 VIA_via1_4
* cell instance $18320 r0 *1 4.275,66.43
X$18320 1556 VIA_via1_4
* cell instance $18321 r0 *1 4.275,66.43
X$18321 1556 VIA_via2_5
* cell instance $18322 r0 *1 3.325,65.17
X$18322 1556 VIA_via1_4
* cell instance $18323 r0 *1 3.325,65.17
X$18323 1556 VIA_via2_5
* cell instance $18324 r0 *1 43.035,60.55
X$18324 1557 VIA_via2_5
* cell instance $18325 r0 *1 42.275,60.55
X$18325 1557 VIA_via2_5
* cell instance $18326 r0 *1 42.275,60.83
X$18326 1557 VIA_via1_4
* cell instance $18327 r0 *1 41.895,60.55
X$18327 1557 VIA_via1_4
* cell instance $18328 r0 *1 41.895,60.55
X$18328 1557 VIA_via2_5
* cell instance $18329 r0 *1 43.225,62.37
X$18329 1557 VIA_via1_4
* cell instance $18330 r0 *1 48.165,61.95
X$18330 1558 VIA_via2_5
* cell instance $18331 r0 *1 46.455,61.95
X$18331 1558 VIA_via2_5
* cell instance $18332 r0 *1 46.265,60.83
X$18332 1558 VIA_via1_4
* cell instance $18333 r0 *1 47.785,61.95
X$18333 1558 VIA_via1_4
* cell instance $18334 r0 *1 47.785,61.95
X$18334 1558 VIA_via2_5
* cell instance $18335 r0 *1 48.165,62.37
X$18335 1558 VIA_via1_4
* cell instance $18336 r0 *1 52.915,60.83
X$18336 1559 VIA_via2_5
* cell instance $18337 r0 *1 52.535,61.39
X$18337 1559 VIA_via2_5
* cell instance $18338 r0 *1 53.105,61.39
X$18338 1559 VIA_via2_5
* cell instance $18339 r0 *1 52.535,61.95
X$18339 1559 VIA_via1_4
* cell instance $18340 r0 *1 53.105,60.83
X$18340 1559 VIA_via1_4
* cell instance $18341 r0 *1 51.015,60.83
X$18341 1559 VIA_via1_4
* cell instance $18342 r0 *1 51.015,60.83
X$18342 1559 VIA_via2_5
* cell instance $18343 r0 *1 53.485,59.99
X$18343 1560 VIA_via1_7
* cell instance $18344 r0 *1 54.245,60.55
X$18344 1560 VIA_via2_5
* cell instance $18345 r0 *1 53.675,60.55
X$18345 1560 VIA_via2_5
* cell instance $18346 r0 *1 54.245,60.83
X$18346 1560 VIA_via1_4
* cell instance $18347 r0 *1 67.545,67.27
X$18347 1561 VIA_via2_5
* cell instance $18348 r0 *1 67.355,61.11
X$18348 1561 VIA_via2_5
* cell instance $18349 r0 *1 63.935,68.25
X$18349 1561 VIA_via2_5
* cell instance $18350 r0 *1 62.795,68.25
X$18350 1561 VIA_via2_5
* cell instance $18351 r0 *1 63.935,70.49
X$18351 1561 VIA_via2_5
* cell instance $18352 r0 *1 62.035,68.25
X$18352 1561 VIA_via2_5
* cell instance $18353 r0 *1 66.595,67.27
X$18353 1561 VIA_via2_5
* cell instance $18354 r0 *1 62.035,70.49
X$18354 1561 VIA_via2_5
* cell instance $18355 r0 *1 68.115,68.25
X$18355 1561 VIA_via2_5
* cell instance $18356 r0 *1 67.355,63.63
X$18356 1561 VIA_via1_4
* cell instance $18357 r0 *1 62.795,63.63
X$18357 1561 VIA_via1_4
* cell instance $18358 r0 *1 62.035,67.97
X$18358 1561 VIA_via1_4
* cell instance $18359 r0 *1 63.935,70.77
X$18359 1561 VIA_via1_4
* cell instance $18360 r0 *1 64.315,72.03
X$18360 1561 VIA_via1_4
* cell instance $18361 r0 *1 68.305,70.77
X$18361 1561 VIA_via1_4
* cell instance $18362 r0 *1 64.125,65.17
X$18362 1561 VIA_via1_4
* cell instance $18363 r0 *1 66.595,68.25
X$18363 1561 VIA_via1_4
* cell instance $18364 r0 *1 66.595,68.25
X$18364 1561 VIA_via2_5
* cell instance $18365 r0 *1 67.735,65.17
X$18365 1561 VIA_via1_4
* cell instance $18366 r0 *1 62.035,73.57
X$18366 1561 VIA_via1_4
* cell instance $18367 r0 *1 65.455,60.83
X$18367 1561 VIA_via1_4
* cell instance $18368 r0 *1 65.455,60.83
X$18368 1561 VIA_via2_5
* cell instance $18369 r0 *1 70.395,60.69
X$18369 1562 VIA_via2_5
* cell instance $18370 r0 *1 70.395,56.63
X$18370 1562 VIA_via1_4
* cell instance $18371 r0 *1 67.545,60.83
X$18371 1562 VIA_via1_4
* cell instance $18372 r0 *1 67.545,60.97
X$18372 1562 VIA_via2_5
* cell instance $18373 r0 *1 67.925,67.83
X$18373 1563 VIA_via2_5
* cell instance $18374 r0 *1 68.305,67.97
X$18374 1563 VIA_via1_4
* cell instance $18375 r0 *1 68.305,67.83
X$18375 1563 VIA_via2_5
* cell instance $18376 r0 *1 67.165,67.97
X$18376 1563 VIA_via1_4
* cell instance $18377 r0 *1 67.165,67.83
X$18377 1563 VIA_via2_5
* cell instance $18378 r0 *1 67.545,60.55
X$18378 1563 VIA_via1_4
* cell instance $18379 r0 *1 71.725,60.83
X$18379 1564 VIA_via2_5
* cell instance $18380 r0 *1 71.725,61.95
X$18380 1564 VIA_via1_4
* cell instance $18381 r0 *1 72.675,60.83
X$18381 1564 VIA_via1_4
* cell instance $18382 r0 *1 72.675,60.83
X$18382 1564 VIA_via2_5
* cell instance $18383 r0 *1 74.575,60.83
X$18383 1564 VIA_via1_4
* cell instance $18384 r0 *1 74.575,60.69
X$18384 1564 VIA_via2_5
* cell instance $18385 r0 *1 80.465,59.99
X$18385 1565 VIA_via1_7
* cell instance $18386 r0 *1 80.085,60.83
X$18386 1565 VIA_via1_4
* cell instance $18387 r0 *1 89.015,60.41
X$18387 1566 VIA_via2_5
* cell instance $18388 r0 *1 92.055,61.11
X$18388 1566 VIA_via2_5
* cell instance $18389 r0 *1 93.385,60.69
X$18389 1566 VIA_via2_5
* cell instance $18390 r0 *1 93.385,62.37
X$18390 1566 VIA_via1_4
* cell instance $18391 r0 *1 92.055,63.63
X$18391 1566 VIA_via1_4
* cell instance $18392 r0 *1 89.015,60.69
X$18392 1566 VIA_via1_4
* cell instance $18393 r0 *1 91.675,60.83
X$18393 1567 VIA_via1_4
* cell instance $18394 r0 *1 92.055,59.71
X$18394 1567 VIA_via1_4
* cell instance $18395 r0 *1 92.815,60.69
X$18395 1568 VIA_via1_4
* cell instance $18396 r0 *1 92.435,60.83
X$18396 1568 VIA_via1_4
* cell instance $18397 r0 *1 96.805,61.81
X$18397 1569 VIA_via1_7
* cell instance $18398 r0 *1 96.805,61.11
X$18398 1569 VIA_via2_5
* cell instance $18399 r0 *1 97.535,61.11
X$18399 1569 VIA_via3_2
* cell instance $18400 r0 *1 97.535,61.11
X$18400 1569 VIA_via4_0
* cell instance $18401 r0 *1 92.245,60.27
X$18401 1570 VIA_via2_5
* cell instance $18402 r0 *1 94.715,60.55
X$18402 1570 VIA_via2_5
* cell instance $18403 r0 *1 92.625,60.27
X$18403 1570 VIA_via2_5
* cell instance $18404 r0 *1 94.715,60.27
X$18404 1570 VIA_via2_5
* cell instance $18405 r0 *1 94.715,59.57
X$18405 1570 VIA_via1_4
* cell instance $18406 r0 *1 92.245,59.57
X$18406 1570 VIA_via1_4
* cell instance $18407 r0 *1 92.625,60.83
X$18407 1570 VIA_via1_4
* cell instance $18408 r0 *1 96.425,60.55
X$18408 1570 VIA_via1_4
* cell instance $18409 r0 *1 96.425,60.55
X$18409 1570 VIA_via2_5
* cell instance $18410 r0 *1 6.935,58.59
X$18410 1571 VIA_via1_7
* cell instance $18411 r0 *1 6.935,59.57
X$18411 1571 VIA_via2_5
* cell instance $18412 r0 *1 5.605,59.57
X$18412 1571 VIA_via1_4
* cell instance $18413 r0 *1 5.605,59.57
X$18413 1571 VIA_via2_5
* cell instance $18414 r0 *1 92.245,60.83
X$18414 1572 VIA_via1_4
* cell instance $18415 r0 *1 92.245,60.83
X$18415 1572 VIA_via2_5
* cell instance $18416 r0 *1 94.145,60.83
X$18416 1572 VIA_via1_4
* cell instance $18417 r0 *1 94.145,60.83
X$18417 1572 VIA_via2_5
* cell instance $18418 r0 *1 92.625,59.57
X$18418 1573 VIA_via1_4
* cell instance $18419 r0 *1 92.625,59.57
X$18419 1573 VIA_via2_5
* cell instance $18420 r0 *1 93.765,59.57
X$18420 1573 VIA_via1_4
* cell instance $18421 r0 *1 93.765,59.57
X$18421 1573 VIA_via2_5
* cell instance $18422 r0 *1 14.345,59.57
X$18422 1574 VIA_via1_4
* cell instance $18423 r0 *1 14.345,59.71
X$18423 1574 VIA_via2_5
* cell instance $18424 r0 *1 13.395,59.71
X$18424 1574 VIA_via1_4
* cell instance $18425 r0 *1 13.395,59.71
X$18425 1574 VIA_via2_5
* cell instance $18426 r0 *1 19.285,59.71
X$18426 1575 VIA_via1_4
* cell instance $18427 r0 *1 19.285,59.71
X$18427 1575 VIA_via2_5
* cell instance $18428 r0 *1 22.705,59.57
X$18428 1575 VIA_via1_4
* cell instance $18429 r0 *1 22.705,59.71
X$18429 1575 VIA_via2_5
* cell instance $18430 r0 *1 21.945,60.83
X$18430 1576 VIA_via1_4
* cell instance $18431 r0 *1 21.945,60.97
X$18431 1576 VIA_via2_5
* cell instance $18432 r0 *1 24.605,60.97
X$18432 1576 VIA_via1_4
* cell instance $18433 r0 *1 24.605,60.97
X$18433 1576 VIA_via2_5
* cell instance $18434 r0 *1 86.355,59.71
X$18434 1577 VIA_via2_5
* cell instance $18435 r0 *1 87.115,62.37
X$18435 1577 VIA_via1_4
* cell instance $18436 r0 *1 89.205,59.71
X$18436 1577 VIA_via1_4
* cell instance $18437 r0 *1 89.205,59.71
X$18437 1577 VIA_via2_5
* cell instance $18438 r0 *1 85.025,59.57
X$18438 1577 VIA_via1_4
* cell instance $18439 r0 *1 85.025,59.71
X$18439 1577 VIA_via2_5
* cell instance $18440 r0 *1 86.545,61.81
X$18440 1578 VIA_via1_7
* cell instance $18441 r0 *1 86.545,60.83
X$18441 1578 VIA_via2_5
* cell instance $18442 r0 *1 88.825,60.83
X$18442 1578 VIA_via1_4
* cell instance $18443 r0 *1 88.825,60.83
X$18443 1578 VIA_via2_5
* cell instance $18444 r0 *1 54.625,62.93
X$18444 1579 VIA_via2_5
* cell instance $18445 r0 *1 54.625,62.65
X$18445 1579 VIA_via2_5
* cell instance $18446 r0 *1 50.255,90.51
X$18446 1579 VIA_via2_5
* cell instance $18447 r0 *1 50.255,90.93
X$18447 1579 VIA_via2_5
* cell instance $18448 r0 *1 66.785,62.79
X$18448 1579 VIA_via2_5
* cell instance $18449 r0 *1 38.665,88.69
X$18449 1579 VIA_via2_5
* cell instance $18450 r0 *1 38.665,90.93
X$18450 1579 VIA_via2_5
* cell instance $18451 r0 *1 88.635,62.79
X$18451 1579 VIA_via2_5
* cell instance $18452 r0 *1 37.905,59.85
X$18452 1579 VIA_via2_5
* cell instance $18453 r0 *1 37.905,62.51
X$18453 1579 VIA_via2_5
* cell instance $18454 r0 *1 54.625,62.37
X$18454 1579 VIA_via1_4
* cell instance $18455 r0 *1 66.785,62.37
X$18455 1579 VIA_via1_4
* cell instance $18456 r0 *1 50.445,87.57
X$18456 1579 VIA_via1_4
* cell instance $18457 r0 *1 50.445,87.57
X$18457 1579 VIA_via2_5
* cell instance $18458 r0 *1 50.495,87.57
X$18458 1579 VIA_via3_2
* cell instance $18459 r0 *1 50.255,91.63
X$18459 1579 VIA_via1_4
* cell instance $18460 r0 *1 13.015,88.83
X$18460 1579 VIA_via1_4
* cell instance $18461 r0 *1 13.015,88.69
X$18461 1579 VIA_via2_5
* cell instance $18462 r0 *1 20.615,88.83
X$18462 1579 VIA_via1_4
* cell instance $18463 r0 *1 20.615,88.97
X$18463 1579 VIA_via2_5
* cell instance $18464 r0 *1 36.765,59.85
X$18464 1579 VIA_via1_4
* cell instance $18465 r0 *1 36.765,59.85
X$18465 1579 VIA_via2_5
* cell instance $18466 r0 *1 38.665,90.37
X$18466 1579 VIA_via1_4
* cell instance $18467 r0 *1 32.015,88.83
X$18467 1579 VIA_via1_4
* cell instance $18468 r0 *1 32.015,88.69
X$18468 1579 VIA_via2_5
* cell instance $18469 r0 *1 32.015,88.97
X$18469 1579 VIA_via2_5
* cell instance $18470 r0 *1 88.825,65.17
X$18470 1579 VIA_via1_4
* cell instance $18471 r0 *1 88.635,62.37
X$18471 1579 VIA_via1_4
* cell instance $18472 r0 *1 50.495,90.51
X$18472 1579 VIA_via3_2
* cell instance $18473 r0 *1 50.495,62.93
X$18473 1579 VIA_via3_2
* cell instance $18474 r0 *1 43.225,60.69
X$18474 1580 VIA_via1_4
* cell instance $18475 r0 *1 43.225,60.69
X$18475 1580 VIA_via2_5
* cell instance $18476 r0 *1 39.615,60.83
X$18476 1580 VIA_via1_4
* cell instance $18477 r0 *1 39.615,60.69
X$18477 1580 VIA_via2_5
* cell instance $18478 r0 *1 86.925,59.57
X$18478 1581 VIA_via1_4
* cell instance $18479 r0 *1 86.925,59.57
X$18479 1581 VIA_via2_5
* cell instance $18480 r0 *1 85.975,59.57
X$18480 1581 VIA_via1_4
* cell instance $18481 r0 *1 85.975,59.57
X$18481 1581 VIA_via2_5
* cell instance $18482 r0 *1 87.875,60.69
X$18482 1582 VIA_via2_5
* cell instance $18483 r0 *1 87.685,62.37
X$18483 1582 VIA_via1_4
* cell instance $18484 r0 *1 88.255,60.69
X$18484 1582 VIA_via1_4
* cell instance $18485 r0 *1 88.255,60.69
X$18485 1582 VIA_via2_5
* cell instance $18486 r0 *1 84.075,60.83
X$18486 1582 VIA_via1_4
* cell instance $18487 r0 *1 84.075,60.69
X$18487 1582 VIA_via2_5
* cell instance $18488 r0 *1 41.895,59.57
X$18488 1583 VIA_via2_5
* cell instance $18489 r0 *1 41.895,58.45
X$18489 1583 VIA_via1_4
* cell instance $18490 r0 *1 42.275,59.57
X$18490 1583 VIA_via1_4
* cell instance $18491 r0 *1 42.275,59.57
X$18491 1583 VIA_via2_5
* cell instance $18492 r0 *1 39.995,59.57
X$18492 1583 VIA_via1_4
* cell instance $18493 r0 *1 39.995,59.57
X$18493 1583 VIA_via2_5
* cell instance $18494 r0 *1 85.975,60.83
X$18494 1584 VIA_via1_4
* cell instance $18495 r0 *1 85.025,60.83
X$18495 1584 VIA_via1_4
* cell instance $18496 r0 *1 43.225,59.57
X$18496 1585 VIA_via1_4
* cell instance $18497 r0 *1 43.605,59.57
X$18497 1585 VIA_via1_4
* cell instance $18498 r0 *1 84.455,60.83
X$18498 1586 VIA_via2_5
* cell instance $18499 r0 *1 84.645,61.95
X$18499 1586 VIA_via1_4
* cell instance $18500 r0 *1 82.745,60.83
X$18500 1586 VIA_via1_4
* cell instance $18501 r0 *1 82.745,60.83
X$18501 1586 VIA_via2_5
* cell instance $18502 r0 *1 85.025,62.37
X$18502 1586 VIA_via1_4
* cell instance $18503 r0 *1 56.335,66.01
X$18503 1587 VIA_via2_5
* cell instance $18504 r0 *1 56.335,65.31
X$18504 1587 VIA_via2_5
* cell instance $18505 r0 *1 55.575,59.99
X$18505 1587 VIA_via2_5
* cell instance $18506 r0 *1 52.725,66.01
X$18506 1587 VIA_via2_5
* cell instance $18507 r0 *1 49.685,63.77
X$18507 1587 VIA_via2_5
* cell instance $18508 r0 *1 50.445,59.99
X$18508 1587 VIA_via2_5
* cell instance $18509 r0 *1 46.645,63.77
X$18509 1587 VIA_via2_5
* cell instance $18510 r0 *1 52.535,63.63
X$18510 1587 VIA_via1_4
* cell instance $18511 r0 *1 52.535,63.63
X$18511 1587 VIA_via2_5
* cell instance $18512 r0 *1 48.925,63.63
X$18512 1587 VIA_via1_4
* cell instance $18513 r0 *1 48.925,63.77
X$18513 1587 VIA_via2_5
* cell instance $18514 r0 *1 50.445,60.83
X$18514 1587 VIA_via1_4
* cell instance $18515 r0 *1 50.445,60.83
X$18515 1587 VIA_via2_5
* cell instance $18516 r0 *1 49.305,60.83
X$18516 1587 VIA_via1_4
* cell instance $18517 r0 *1 49.305,60.83
X$18517 1587 VIA_via2_5
* cell instance $18518 r0 *1 56.335,66.43
X$18518 1587 VIA_via1_4
* cell instance $18519 r0 *1 56.905,65.17
X$18519 1587 VIA_via1_4
* cell instance $18520 r0 *1 56.905,65.31
X$18520 1587 VIA_via2_5
* cell instance $18521 r0 *1 55.575,60.83
X$18521 1587 VIA_via1_4
* cell instance $18522 r0 *1 46.835,94.43
X$18522 1587 VIA_via1_4
* cell instance $18523 r0 *1 77.235,60.83
X$18523 1588 VIA_via1_4
* cell instance $18524 r0 *1 77.235,60.97
X$18524 1588 VIA_via2_5
* cell instance $18525 r0 *1 74.955,60.97
X$18525 1588 VIA_via1_4
* cell instance $18526 r0 *1 74.955,60.97
X$18526 1588 VIA_via2_5
* cell instance $18527 r0 *1 53.485,60.41
X$18527 1589 VIA_via1_7
* cell instance $18528 r0 *1 53.485,60.27
X$18528 1589 VIA_via2_5
* cell instance $18529 r0 *1 54.245,60.27
X$18529 1589 VIA_via2_5
* cell instance $18530 r0 *1 54.245,59.57
X$18530 1589 VIA_via1_4
* cell instance $18531 r0 *1 54.435,59.99
X$18531 1590 VIA_via1_7
* cell instance $18532 r0 *1 54.435,60.83
X$18532 1590 VIA_via2_5
* cell instance $18533 r0 *1 55.005,60.83
X$18533 1590 VIA_via1_4
* cell instance $18534 r0 *1 55.005,60.83
X$18534 1590 VIA_via2_5
* cell instance $18535 r0 *1 54.055,55.79
X$18535 1591 VIA_via1_7
* cell instance $18536 r0 *1 54.055,59.71
X$18536 1591 VIA_via2_5
* cell instance $18537 r0 *1 54.245,62.37
X$18537 1591 VIA_via1_4
* cell instance $18538 r0 *1 54.245,62.37
X$18538 1591 VIA_via2_5
* cell instance $18539 r0 *1 54.695,59.71
X$18539 1591 VIA_via3_2
* cell instance $18540 r0 *1 54.695,62.37
X$18540 1591 VIA_via3_2
* cell instance $18541 r0 *1 70.015,59.57
X$18541 1592 VIA_via1_4
* cell instance $18542 r0 *1 70.015,59.57
X$18542 1592 VIA_via2_5
* cell instance $18543 r0 *1 73.625,59.57
X$18543 1592 VIA_via1_4
* cell instance $18544 r0 *1 73.625,59.57
X$18544 1592 VIA_via2_5
* cell instance $18545 r0 *1 68.495,63.21
X$18545 1593 VIA_via1_7
* cell instance $18546 r0 *1 68.495,60.55
X$18546 1593 VIA_via2_5
* cell instance $18547 r0 *1 66.785,60.55
X$18547 1593 VIA_via2_5
* cell instance $18548 r0 *1 66.785,60.83
X$18548 1593 VIA_via1_4
* cell instance $18549 r0 *1 70.205,74.83
X$18549 1594 VIA_via1_4
* cell instance $18550 r0 *1 70.205,74.83
X$18550 1594 VIA_via2_5
* cell instance $18551 r0 *1 70.095,74.83
X$18551 1594 VIA_via3_2
* cell instance $18552 r0 *1 73.815,74.69
X$18552 1594 VIA_via1_4
* cell instance $18553 r0 *1 73.815,74.69
X$18553 1594 VIA_via2_5
* cell instance $18554 r0 *1 76.475,74.83
X$18554 1594 VIA_via1_4
* cell instance $18555 r0 *1 76.475,74.69
X$18555 1594 VIA_via2_5
* cell instance $18556 r0 *1 67.735,60.83
X$18556 1594 VIA_via1_4
* cell instance $18557 r0 *1 67.735,60.83
X$18557 1594 VIA_via2_5
* cell instance $18558 r0 *1 70.095,60.83
X$18558 1594 VIA_via3_2
* cell instance $18559 r0 *1 62.225,60.83
X$18559 1595 VIA_via1_4
* cell instance $18560 r0 *1 62.225,60.97
X$18560 1595 VIA_via2_5
* cell instance $18561 r0 *1 65.835,60.97
X$18561 1595 VIA_via1_4
* cell instance $18562 r0 *1 65.835,60.97
X$18562 1595 VIA_via2_5
* cell instance $18563 r0 *1 67.355,59.99
X$18563 1596 VIA_via1_7
* cell instance $18564 r0 *1 67.355,60.83
X$18564 1596 VIA_via1_4
* cell instance $18565 r0 *1 66.405,81.97
X$18565 1597 VIA_via1_4
* cell instance $18566 r0 *1 66.405,81.97
X$18566 1597 VIA_via2_5
* cell instance $18567 r0 *1 66.455,81.97
X$18567 1597 VIA_via3_2
* cell instance $18568 r0 *1 64.695,59.57
X$18568 1597 VIA_via1_4
* cell instance $18569 r0 *1 64.695,59.57
X$18569 1597 VIA_via2_5
* cell instance $18570 r0 *1 66.455,59.57
X$18570 1597 VIA_via3_2
* cell instance $18571 r0 *1 3.135,61.39
X$18571 1598 VIA_via1_7
* cell instance $18572 r0 *1 12.445,62.23
X$18572 1598 VIA_via2_5
* cell instance $18573 r0 *1 3.135,62.37
X$18573 1598 VIA_via2_5
* cell instance $18574 r0 *1 5.225,62.23
X$18574 1598 VIA_via2_5
* cell instance $18575 r0 *1 3.515,62.37
X$18575 1598 VIA_via2_5
* cell instance $18576 r0 *1 11.495,62.37
X$18576 1598 VIA_via1_4
* cell instance $18577 r0 *1 11.495,62.23
X$18577 1598 VIA_via2_5
* cell instance $18578 r0 *1 8.645,62.37
X$18578 1598 VIA_via1_4
* cell instance $18579 r0 *1 8.645,62.23
X$18579 1598 VIA_via2_5
* cell instance $18580 r0 *1 12.445,59.57
X$18580 1598 VIA_via1_4
* cell instance $18581 r0 *1 3.515,63.63
X$18581 1598 VIA_via1_4
* cell instance $18582 r0 *1 5.605,62.37
X$18582 1598 VIA_via1_4
* cell instance $18583 r0 *1 5.605,62.23
X$18583 1598 VIA_via2_5
* cell instance $18584 r0 *1 5.225,65.17
X$18584 1598 VIA_via1_4
* cell instance $18585 r0 *1 4.275,62.37
X$18585 1598 VIA_via1_4
* cell instance $18586 r0 *1 4.275,62.37
X$18586 1598 VIA_via2_5
* cell instance $18587 r0 *1 10.735,61.25
X$18587 1599 VIA_via2_5
* cell instance $18588 r0 *1 13.775,61.25
X$18588 1599 VIA_via2_5
* cell instance $18589 r0 *1 13.775,62.37
X$18589 1599 VIA_via1_4
* cell instance $18590 r0 *1 10.735,62.37
X$18590 1599 VIA_via1_4
* cell instance $18591 r0 *1 12.255,61.25
X$18591 1599 VIA_via1_4
* cell instance $18592 r0 *1 12.255,61.25
X$18592 1599 VIA_via2_5
* cell instance $18593 r0 *1 18.905,61.25
X$18593 1600 VIA_via2_5
* cell instance $18594 r0 *1 19.095,63.63
X$18594 1600 VIA_via1_4
* cell instance $18595 r0 *1 18.905,62.37
X$18595 1600 VIA_via1_4
* cell instance $18596 r0 *1 20.235,61.25
X$18596 1600 VIA_via1_4
* cell instance $18597 r0 *1 20.235,61.25
X$18597 1600 VIA_via2_5
* cell instance $18598 r0 *1 23.085,63.35
X$18598 1601 VIA_via1_4
* cell instance $18599 r0 *1 23.085,62.37
X$18599 1601 VIA_via1_4
* cell instance $18600 r0 *1 23.655,60.83
X$18600 1601 VIA_via1_4
* cell instance $18601 r0 *1 29.545,62.65
X$18601 1602 VIA_via1_4
* cell instance $18602 r0 *1 29.545,62.65
X$18602 1602 VIA_via2_5
* cell instance $18603 r0 *1 29.925,62.37
X$18603 1602 VIA_via1_4
* cell instance $18604 r0 *1 29.925,62.37
X$18604 1602 VIA_via2_5
* cell instance $18605 r0 *1 30.115,62.09
X$18605 1603 VIA_via1_7
* cell instance $18606 r0 *1 29.545,60.83
X$18606 1603 VIA_via1_4
* cell instance $18607 r0 *1 30.115,59.71
X$18607 1604 VIA_via1_4
* cell instance $18608 r0 *1 30.115,62.37
X$18608 1604 VIA_via1_4
* cell instance $18609 r0 *1 39.425,62.37
X$18609 1605 VIA_via1_7
* cell instance $18610 r0 *1 39.615,61.95
X$18610 1605 VIA_via1_4
* cell instance $18611 r0 *1 39.615,78.05
X$18611 1605 VIA_via2_5
* cell instance $18612 r0 *1 53.295,61.53
X$18612 1605 VIA_via2_5
* cell instance $18613 r0 *1 50.255,75.95
X$18613 1605 VIA_via2_5
* cell instance $18614 r0 *1 50.215,75.95
X$18614 1605 VIA_via3_2
* cell instance $18615 r0 *1 65.835,72.17
X$18615 1605 VIA_via2_5
* cell instance $18616 r0 *1 65.835,77.63
X$18616 1605 VIA_via2_5
* cell instance $18617 r0 *1 78.185,71.33
X$18617 1605 VIA_via2_5
* cell instance $18618 r0 *1 39.615,61.53
X$18618 1605 VIA_via2_5
* cell instance $18619 r0 *1 50.255,76.3
X$18619 1605 VIA_via1_4
* cell instance $18620 r0 *1 53.105,62.37
X$18620 1605 VIA_via1_4
* cell instance $18621 r0 *1 58.235,77.7
X$18621 1605 VIA_via1_4
* cell instance $18622 r0 *1 58.235,77.77
X$18622 1605 VIA_via2_5
* cell instance $18623 r0 *1 66.785,72.03
X$18623 1605 VIA_via1_4
* cell instance $18624 r0 *1 66.785,72.17
X$18624 1605 VIA_via2_5
* cell instance $18625 r0 *1 42.465,79.17
X$18625 1605 VIA_via1_4
* cell instance $18626 r0 *1 26.315,77.63
X$18626 1605 VIA_via1_4
* cell instance $18627 r0 *1 26.315,77.63
X$18627 1605 VIA_via2_5
* cell instance $18628 r0 *1 26.415,77.63
X$18628 1605 VIA_via3_2
* cell instance $18629 r0 *1 35.815,77.63
X$18629 1605 VIA_via1_4
* cell instance $18630 r0 *1 21.565,77.63
X$18630 1605 VIA_via1_4
* cell instance $18631 r0 *1 21.565,77.63
X$18631 1605 VIA_via2_5
* cell instance $18632 r0 *1 20.805,77.63
X$18632 1605 VIA_via1_4
* cell instance $18633 r0 *1 20.805,77.63
X$18633 1605 VIA_via2_5
* cell instance $18634 r0 *1 78.185,70.77
X$18634 1605 VIA_via1_4
* cell instance $18635 r0 *1 35.935,77.35
X$18635 1605 VIA_via4_0
* cell instance $18636 r0 *1 50.215,77.35
X$18636 1605 VIA_via4_0
* cell instance $18637 r0 *1 42.655,77.35
X$18637 1605 VIA_via4_0
* cell instance $18638 r0 *1 26.415,77.35
X$18638 1605 VIA_via4_0
* cell instance $18639 r0 *1 67.295,71.33
X$18639 1605 VIA_via3_2
* cell instance $18640 r0 *1 67.295,72.17
X$18640 1605 VIA_via3_2
* cell instance $18641 r0 *1 35.935,78.05
X$18641 1605 VIA_via3_2
* cell instance $18642 r0 *1 35.815,78.05
X$18642 1605 VIA_via2_5
* cell instance $18643 r0 *1 58.055,77.49
X$18643 1605 VIA_via3_2
* cell instance $18644 r0 *1 58.055,77.35
X$18644 1605 VIA_via4_0
* cell instance $18645 r0 *1 42.655,78.05
X$18645 1605 VIA_via3_2
* cell instance $18646 r0 *1 42.655,78.05
X$18646 1605 VIA_via2_5
* cell instance $18647 r0 *1 56.145,61.81
X$18647 1606 VIA_via2_5
* cell instance $18648 r0 *1 55.195,61.81
X$18648 1606 VIA_via2_5
* cell instance $18649 r0 *1 55.195,63.63
X$18649 1606 VIA_via1_4
* cell instance $18650 r0 *1 58.805,61.95
X$18650 1606 VIA_via1_4
* cell instance $18651 r0 *1 58.805,61.81
X$18651 1606 VIA_via2_5
* cell instance $18652 r0 *1 56.145,60.83
X$18652 1606 VIA_via1_4
* cell instance $18653 r0 *1 63.175,63.21
X$18653 1607 VIA_via1_7
* cell instance $18654 r0 *1 63.175,63.21
X$18654 1607 VIA_via2_5
* cell instance $18655 r0 *1 61.845,63.21
X$18655 1607 VIA_via2_5
* cell instance $18656 r0 *1 61.655,62.37
X$18656 1607 VIA_via1_4
* cell instance $18657 r0 *1 64.885,62.37
X$18657 1608 VIA_via1_4
* cell instance $18658 r0 *1 64.505,61.25
X$18658 1608 VIA_via1_4
* cell instance $18659 r0 *1 64.885,60.83
X$18659 1608 VIA_via1_4
* cell instance $18660 r0 *1 73.055,63.07
X$18660 1609 VIA_via2_5
* cell instance $18661 r0 *1 74.195,63.07
X$18661 1609 VIA_via2_5
* cell instance $18662 r0 *1 73.055,63.63
X$18662 1609 VIA_via1_4
* cell instance $18663 r0 *1 74.385,62.09
X$18663 1609 VIA_via1_4
* cell instance $18664 r0 *1 75.715,63.91
X$18664 1610 VIA_via2_5
* cell instance $18665 r0 *1 77.995,63.91
X$18665 1610 VIA_via2_5
* cell instance $18666 r0 *1 77.995,64.75
X$18666 1610 VIA_via1_4
* cell instance $18667 r0 *1 75.335,62.37
X$18667 1610 VIA_via1_4
* cell instance $18668 r0 *1 75.715,63.63
X$18668 1610 VIA_via1_4
* cell instance $18669 r0 *1 81.225,63.63
X$18669 1611 VIA_via2_5
* cell instance $18670 r0 *1 81.225,64.75
X$18670 1611 VIA_via1_4
* cell instance $18671 r0 *1 79.325,62.37
X$18671 1611 VIA_via1_4
* cell instance $18672 r0 *1 79.515,63.63
X$18672 1611 VIA_via1_4
* cell instance $18673 r0 *1 79.515,63.63
X$18673 1611 VIA_via2_5
* cell instance $18674 r0 *1 95.855,64.61
X$18674 1612 VIA_via1_7
* cell instance $18675 r0 *1 96.045,62.37
X$18675 1612 VIA_via1_4
* cell instance $18676 r0 *1 96.045,62.09
X$18676 1613 VIA_via1_4
* cell instance $18677 r0 *1 96.425,62.37
X$18677 1613 VIA_via1_4
* cell instance $18678 r0 *1 5.225,61.81
X$18678 1614 VIA_via1_7
* cell instance $18679 r0 *1 5.225,61.81
X$18679 1614 VIA_via2_5
* cell instance $18680 r0 *1 4.085,61.81
X$18680 1614 VIA_via2_5
* cell instance $18681 r0 *1 4.085,60.83
X$18681 1614 VIA_via1_4
* cell instance $18682 r0 *1 91.865,62.09
X$18682 1615 VIA_via2_5
* cell instance $18683 r0 *1 93.195,62.09
X$18683 1615 VIA_via2_5
* cell instance $18684 r0 *1 91.865,62.65
X$18684 1615 VIA_via2_5
* cell instance $18685 r0 *1 91.865,63.63
X$18685 1615 VIA_via1_4
* cell instance $18686 r0 *1 93.195,62.37
X$18686 1615 VIA_via1_4
* cell instance $18687 r0 *1 78.945,62.65
X$18687 1615 VIA_via1_4
* cell instance $18688 r0 *1 78.945,62.65
X$18688 1615 VIA_via2_5
* cell instance $18689 r0 *1 88.635,61.81
X$18689 1616 VIA_via1_7
* cell instance $18690 r0 *1 88.635,60.83
X$18690 1616 VIA_via1_4
* cell instance $18691 r0 *1 10.545,62.09
X$18691 1617 VIA_via2_5
* cell instance $18692 r0 *1 10.735,63.63
X$18692 1617 VIA_via1_4
* cell instance $18693 r0 *1 8.265,62.09
X$18693 1617 VIA_via1_4
* cell instance $18694 r0 *1 8.265,62.09
X$18694 1617 VIA_via2_5
* cell instance $18695 r0 *1 11.115,61.81
X$18695 1618 VIA_via1_7
* cell instance $18696 r0 *1 11.115,61.81
X$18696 1618 VIA_via2_5
* cell instance $18697 r0 *1 9.975,61.81
X$18697 1618 VIA_via2_5
* cell instance $18698 r0 *1 9.975,60.83
X$18698 1618 VIA_via1_4
* cell instance $18699 r0 *1 83.695,61.39
X$18699 1619 VIA_via1_7
* cell instance $18700 r0 *1 83.695,61.39
X$18700 1619 VIA_via2_5
* cell instance $18701 r0 *1 82.365,61.39
X$18701 1619 VIA_via2_5
* cell instance $18702 r0 *1 82.365,62.37
X$18702 1619 VIA_via1_4
* cell instance $18703 r0 *1 80.275,61.81
X$18703 1620 VIA_via1_7
* cell instance $18704 r0 *1 80.275,61.81
X$18704 1620 VIA_via2_5
* cell instance $18705 r0 *1 78.755,61.81
X$18705 1620 VIA_via2_5
* cell instance $18706 r0 *1 78.755,60.83
X$18706 1620 VIA_via1_4
* cell instance $18707 r0 *1 77.615,61.39
X$18707 1621 VIA_via1_7
* cell instance $18708 r0 *1 77.615,61.39
X$18708 1621 VIA_via2_5
* cell instance $18709 r0 *1 78.185,61.39
X$18709 1621 VIA_via2_5
* cell instance $18710 r0 *1 78.185,62.37
X$18710 1621 VIA_via1_4
* cell instance $18711 r0 *1 19.855,61.81
X$18711 1622 VIA_via1_7
* cell instance $18712 r0 *1 19.855,61.81
X$18712 1622 VIA_via2_5
* cell instance $18713 r0 *1 17.955,61.81
X$18713 1622 VIA_via2_5
* cell instance $18714 r0 *1 17.955,60.83
X$18714 1622 VIA_via1_4
* cell instance $18715 r0 *1 14.725,62.23
X$18715 1623 VIA_via1_4
* cell instance $18716 r0 *1 14.725,62.23
X$18716 1623 VIA_via2_5
* cell instance $18717 r0 *1 20.615,62.37
X$18717 1623 VIA_via1_4
* cell instance $18718 r0 *1 20.615,62.23
X$18718 1623 VIA_via2_5
* cell instance $18719 r0 *1 73.625,61.39
X$18719 1624 VIA_via1_7
* cell instance $18720 r0 *1 73.625,61.39
X$18720 1624 VIA_via2_5
* cell instance $18721 r0 *1 69.445,61.39
X$18721 1624 VIA_via2_5
* cell instance $18722 r0 *1 69.445,62.37
X$18722 1624 VIA_via1_4
* cell instance $18723 r0 *1 22.895,59.99
X$18723 1625 VIA_via1_7
* cell instance $18724 r0 *1 22.325,61.11
X$18724 1625 VIA_via2_5
* cell instance $18725 r0 *1 22.895,61.11
X$18725 1625 VIA_via2_5
* cell instance $18726 r0 *1 22.325,62.37
X$18726 1625 VIA_via1_4
* cell instance $18727 r0 *1 22.135,61.53
X$18727 1626 VIA_via2_5
* cell instance $18728 r0 *1 21.375,61.53
X$18728 1626 VIA_via2_5
* cell instance $18729 r0 *1 21.375,62.37
X$18729 1626 VIA_via1_4
* cell instance $18730 r0 *1 22.135,61.11
X$18730 1626 VIA_via1_4
* cell instance $18731 r0 *1 66.595,62.09
X$18731 1627 VIA_via1_4
* cell instance $18732 r0 *1 66.595,60.83
X$18732 1627 VIA_via1_4
* cell instance $18733 r0 *1 53.105,61.81
X$18733 1628 VIA_via1_7
* cell instance $18734 r0 *1 53.105,61.81
X$18734 1628 VIA_via2_5
* cell instance $18735 r0 *1 54.815,61.81
X$18735 1628 VIA_via2_5
* cell instance $18736 r0 *1 54.815,60.83
X$18736 1628 VIA_via1_4
* cell instance $18737 r0 *1 30.305,74.13
X$18737 1629 VIA_via2_5
* cell instance $18738 r0 *1 36.195,74.27
X$18738 1629 VIA_via2_5
* cell instance $18739 r0 *1 32.205,74.27
X$18739 1629 VIA_via2_5
* cell instance $18740 r0 *1 36.195,76.79
X$18740 1629 VIA_via2_5
* cell instance $18741 r0 *1 32.205,73.85
X$18741 1629 VIA_via2_5
* cell instance $18742 r0 *1 30.875,74.13
X$18742 1629 VIA_via2_5
* cell instance $18743 r0 *1 31.065,73.85
X$18743 1629 VIA_via2_5
* cell instance $18744 r0 *1 28.215,74.27
X$18744 1629 VIA_via2_5
* cell instance $18745 r0 *1 29.165,74.27
X$18745 1629 VIA_via2_5
* cell instance $18746 r0 *1 41.515,76.79
X$18746 1629 VIA_via2_5
* cell instance $18747 r0 *1 55.385,76.79
X$18747 1629 VIA_via2_5
* cell instance $18748 r0 *1 50.635,76.79
X$18748 1629 VIA_via2_5
* cell instance $18749 r0 *1 50.635,75.95
X$18749 1629 VIA_via2_5
* cell instance $18750 r0 *1 51.395,75.95
X$18750 1629 VIA_via2_5
* cell instance $18751 r0 *1 30.305,71.89
X$18751 1629 VIA_via2_5
* cell instance $18752 r0 *1 29.545,71.89
X$18752 1629 VIA_via2_5
* cell instance $18753 r0 *1 51.395,76.37
X$18753 1629 VIA_via1_4
* cell instance $18754 r0 *1 54.815,66.43
X$18754 1629 VIA_via1_4
* cell instance $18755 r0 *1 55.385,76.37
X$18755 1629 VIA_via1_4
* cell instance $18756 r0 *1 55.005,71.75
X$18756 1629 VIA_via1_4
* cell instance $18757 r0 *1 55.385,72.45
X$18757 1629 VIA_via1_4
* cell instance $18758 r0 *1 41.515,76.37
X$18758 1629 VIA_via1_4
* cell instance $18759 r0 *1 36.195,76.37
X$18759 1629 VIA_via1_4
* cell instance $18760 r0 *1 29.735,59.57
X$18760 1629 VIA_via1_4
* cell instance $18761 r0 *1 29.165,74.83
X$18761 1629 VIA_via1_4
* cell instance $18762 r0 *1 28.215,76.37
X$18762 1629 VIA_via1_4
* cell instance $18763 r0 *1 29.735,66.43
X$18763 1629 VIA_via1_4
* cell instance $18764 r0 *1 31.065,73.57
X$18764 1629 VIA_via1_4
* cell instance $18765 r0 *1 54.415,75.95
X$18765 1629 VIA_via3_2
* cell instance $18766 r0 *1 54.415,76.79
X$18766 1629 VIA_via3_2
* cell instance $18767 r0 *1 29.775,61.53
X$18767 1629 VIA_via3_2
* cell instance $18768 r0 *1 29.735,61.53
X$18768 1629 VIA_via2_5
* cell instance $18769 r0 *1 29.775,62.79
X$18769 1629 VIA_via3_2
* cell instance $18770 r0 *1 29.735,62.79
X$18770 1629 VIA_via2_5
* cell instance $18771 r0 *1 30.685,62.37
X$18771 1630 VIA_via1_4
* cell instance $18772 r0 *1 30.685,62.23
X$18772 1630 VIA_via2_5
* cell instance $18773 r0 *1 31.065,62.23
X$18773 1630 VIA_via1_4
* cell instance $18774 r0 *1 31.065,62.23
X$18774 1630 VIA_via2_5
* cell instance $18775 r0 *1 51.395,61.39
X$18775 1631 VIA_via1_7
* cell instance $18776 r0 *1 51.395,61.39
X$18776 1631 VIA_via2_5
* cell instance $18777 r0 *1 50.255,61.39
X$18777 1631 VIA_via2_5
* cell instance $18778 r0 *1 50.255,62.37
X$18778 1631 VIA_via1_4
* cell instance $18779 r0 *1 46.645,61.39
X$18779 1632 VIA_via1_7
* cell instance $18780 r0 *1 46.645,61.39
X$18780 1632 VIA_via2_5
* cell instance $18781 r0 *1 45.505,61.39
X$18781 1632 VIA_via2_5
* cell instance $18782 r0 *1 45.505,62.37
X$18782 1632 VIA_via1_4
* cell instance $18783 r0 *1 8.075,63.35
X$18783 1633 VIA_via1_4
* cell instance $18784 r0 *1 7.885,62.37
X$18784 1633 VIA_via1_4
* cell instance $18785 r0 *1 7.885,62.37
X$18785 1633 VIA_via2_5
* cell instance $18786 r0 *1 6.175,62.37
X$18786 1633 VIA_via1_4
* cell instance $18787 r0 *1 6.175,62.37
X$18787 1633 VIA_via2_5
* cell instance $18788 r0 *1 12.445,62.79
X$18788 1634 VIA_via1_7
* cell instance $18789 r0 *1 12.065,63.63
X$18789 1634 VIA_via1_4
* cell instance $18790 r0 *1 15.675,72.03
X$18790 1635 VIA_via2_5
* cell instance $18791 r0 *1 15.675,69.23
X$18791 1635 VIA_via2_5
* cell instance $18792 r0 *1 15.105,72.03
X$18792 1635 VIA_via2_5
* cell instance $18793 r0 *1 13.015,66.43
X$18793 1635 VIA_via2_5
* cell instance $18794 r0 *1 15.675,66.43
X$18794 1635 VIA_via1_4
* cell instance $18795 r0 *1 15.675,66.43
X$18795 1635 VIA_via2_5
* cell instance $18796 r0 *1 9.025,72.03
X$18796 1635 VIA_via1_4
* cell instance $18797 r0 *1 9.025,72.03
X$18797 1635 VIA_via2_5
* cell instance $18798 r0 *1 12.825,63.63
X$18798 1635 VIA_via1_4
* cell instance $18799 r0 *1 19.665,69.23
X$18799 1635 VIA_via1_4
* cell instance $18800 r0 *1 19.665,69.23
X$18800 1635 VIA_via2_5
* cell instance $18801 r0 *1 14.915,69.65
X$18801 1635 VIA_via1_4
* cell instance $18802 r0 *1 14.345,72.03
X$18802 1635 VIA_via1_4
* cell instance $18803 r0 *1 14.345,72.03
X$18803 1635 VIA_via2_5
* cell instance $18804 r0 *1 15.675,70.77
X$18804 1635 VIA_via1_4
* cell instance $18805 r0 *1 15.105,69.23
X$18805 1635 VIA_via1_4
* cell instance $18806 r0 *1 15.105,69.23
X$18806 1635 VIA_via2_5
* cell instance $18807 r0 *1 11.875,66.43
X$18807 1635 VIA_via1_4
* cell instance $18808 r0 *1 11.875,66.43
X$18808 1635 VIA_via2_5
* cell instance $18809 r0 *1 29.925,75.25
X$18809 1636 VIA_via2_5
* cell instance $18810 r0 *1 29.545,75.25
X$18810 1636 VIA_via2_5
* cell instance $18811 r0 *1 42.465,75.11
X$18811 1636 VIA_via2_5
* cell instance $18812 r0 *1 37.525,75.25
X$18812 1636 VIA_via2_5
* cell instance $18813 r0 *1 53.295,72.45
X$18813 1636 VIA_via2_5
* cell instance $18814 r0 *1 53.675,72.45
X$18814 1636 VIA_via2_5
* cell instance $18815 r0 *1 53.105,75.25
X$18815 1636 VIA_via2_5
* cell instance $18816 r0 *1 56.145,76.65
X$18816 1636 VIA_via2_5
* cell instance $18817 r0 *1 53.105,76.93
X$18817 1636 VIA_via2_5
* cell instance $18818 r0 *1 30.685,70.21
X$18818 1636 VIA_via2_5
* cell instance $18819 r0 *1 29.165,63.49
X$18819 1636 VIA_via2_5
* cell instance $18820 r0 *1 30.115,70.21
X$18820 1636 VIA_via2_5
* cell instance $18821 r0 *1 31.065,64.89
X$18821 1636 VIA_via2_5
* cell instance $18822 r0 *1 32.205,64.89
X$18822 1636 VIA_via2_5
* cell instance $18823 r0 *1 56.145,76.37
X$18823 1636 VIA_via1_4
* cell instance $18824 r0 *1 53.105,76.37
X$18824 1636 VIA_via1_4
* cell instance $18825 r0 *1 54.245,69.23
X$18825 1636 VIA_via1_4
* cell instance $18826 r0 *1 55.955,72.45
X$18826 1636 VIA_via1_4
* cell instance $18827 r0 *1 55.955,72.45
X$18827 1636 VIA_via2_5
* cell instance $18828 r0 *1 42.465,74.83
X$18828 1636 VIA_via1_4
* cell instance $18829 r0 *1 37.525,74.83
X$18829 1636 VIA_via1_4
* cell instance $18830 r0 *1 30.115,79.17
X$18830 1636 VIA_via1_4
* cell instance $18831 r0 *1 29.925,74.83
X$18831 1636 VIA_via1_4
* cell instance $18832 r0 *1 29.165,62.37
X$18832 1636 VIA_via1_4
* cell instance $18833 r0 *1 32.205,63.63
X$18833 1636 VIA_via1_4
* cell instance $18834 r0 *1 32.205,63.49
X$18834 1636 VIA_via2_5
* cell instance $18835 r0 *1 31.445,70.77
X$18835 1636 VIA_via1_4
* cell instance $18836 r0 *1 32.775,63.49
X$18836 1637 VIA_via2_5
* cell instance $18837 r0 *1 33.535,66.43
X$18837 1637 VIA_via1_4
* cell instance $18838 r0 *1 32.585,63.63
X$18838 1637 VIA_via1_4
* cell instance $18839 r0 *1 33.155,63.63
X$18839 1637 VIA_via1_4
* cell instance $18840 r0 *1 33.155,63.49
X$18840 1637 VIA_via2_5
* cell instance $18841 r0 *1 33.535,65.45
X$18841 1637 VIA_via1_4
* cell instance $18842 r0 *1 35.245,76.09
X$18842 1638 VIA_via2_5
* cell instance $18843 r0 *1 33.725,77.35
X$18843 1638 VIA_via2_5
* cell instance $18844 r0 *1 34.105,75.95
X$18844 1638 VIA_via2_5
* cell instance $18845 r0 *1 43.605,75.81
X$18845 1638 VIA_via2_5
* cell instance $18846 r0 *1 39.045,76.09
X$18846 1638 VIA_via2_5
* cell instance $18847 r0 *1 39.045,75.81
X$18847 1638 VIA_via2_5
* cell instance $18848 r0 *1 38.475,76.09
X$18848 1638 VIA_via2_5
* cell instance $18849 r0 *1 57.285,76.23
X$18849 1638 VIA_via2_5
* cell instance $18850 r0 *1 54.055,75.81
X$18850 1638 VIA_via2_5
* cell instance $18851 r0 *1 35.245,71.19
X$18851 1638 VIA_via2_5
* cell instance $18852 r0 *1 32.585,71.19
X$18852 1638 VIA_via2_5
* cell instance $18853 r0 *1 33.535,63.91
X$18853 1638 VIA_via2_5
* cell instance $18854 r0 *1 32.775,63.91
X$18854 1638 VIA_via2_5
* cell instance $18855 r0 *1 33.535,62.37
X$18855 1638 VIA_via2_5
* cell instance $18856 r0 *1 54.055,76.37
X$18856 1638 VIA_via1_4
* cell instance $18857 r0 *1 54.055,76.23
X$18857 1638 VIA_via2_5
* cell instance $18858 r0 *1 57.285,74.83
X$18858 1638 VIA_via1_4
* cell instance $18859 r0 *1 57.285,77.35
X$18859 1638 VIA_via1_4
* cell instance $18860 r0 *1 56.905,70.77
X$18860 1638 VIA_via1_4
* cell instance $18861 r0 *1 38.475,76.37
X$18861 1638 VIA_via1_4
* cell instance $18862 r0 *1 34.105,74.83
X$18862 1638 VIA_via1_4
* cell instance $18863 r0 *1 33.725,79.17
X$18863 1638 VIA_via1_4
* cell instance $18864 r0 *1 43.415,74.83
X$18864 1638 VIA_via1_4
* cell instance $18865 r0 *1 33.535,63.63
X$18865 1638 VIA_via1_4
* cell instance $18866 r0 *1 32.585,70.77
X$18866 1638 VIA_via1_4
* cell instance $18867 r0 *1 31.255,62.37
X$18867 1638 VIA_via1_4
* cell instance $18868 r0 *1 31.255,62.37
X$18868 1638 VIA_via2_5
* cell instance $18869 r0 *1 34.255,77.35
X$18869 1638 VIA_via3_2
* cell instance $18870 r0 *1 34.255,76.09
X$18870 1638 VIA_via3_2
* cell instance $18871 r0 *1 49.115,67.55
X$18871 1639 VIA_via2_5
* cell instance $18872 r0 *1 43.605,67.55
X$18872 1639 VIA_via2_5
* cell instance $18873 r0 *1 45.695,67.55
X$18873 1639 VIA_via2_5
* cell instance $18874 r0 *1 40.185,68.25
X$18874 1639 VIA_via2_5
* cell instance $18875 r0 *1 46.835,67.55
X$18875 1639 VIA_via2_5
* cell instance $18876 r0 *1 39.045,68.25
X$18876 1639 VIA_via2_5
* cell instance $18877 r0 *1 49.305,66.43
X$18877 1639 VIA_via1_4
* cell instance $18878 r0 *1 45.695,67.97
X$18878 1639 VIA_via1_4
* cell instance $18879 r0 *1 39.995,65.17
X$18879 1639 VIA_via1_4
* cell instance $18880 r0 *1 39.235,72.03
X$18880 1639 VIA_via1_4
* cell instance $18881 r0 *1 41.325,67.55
X$18881 1639 VIA_via1_4
* cell instance $18882 r0 *1 41.325,67.55
X$18882 1639 VIA_via2_5
* cell instance $18883 r0 *1 40.945,68.25
X$18883 1639 VIA_via1_4
* cell instance $18884 r0 *1 40.945,68.25
X$18884 1639 VIA_via2_5
* cell instance $18885 r0 *1 39.045,69.23
X$18885 1639 VIA_via1_4
* cell instance $18886 r0 *1 43.795,66.43
X$18886 1639 VIA_via1_4
* cell instance $18887 r0 *1 47.025,63.63
X$18887 1639 VIA_via1_4
* cell instance $18888 r0 *1 43.605,65.17
X$18888 1639 VIA_via1_4
* cell instance $18889 r0 *1 49.495,63.63
X$18889 1640 VIA_via1_4
* cell instance $18890 r0 *1 48.545,63.35
X$18890 1640 VIA_via1_4
* cell instance $18891 r0 *1 48.735,62.37
X$18891 1640 VIA_via1_4
* cell instance $18892 r0 *1 54.055,67.83
X$18892 1641 VIA_via1_7
* cell instance $18893 r0 *1 54.435,62.51
X$18893 1641 VIA_via2_5
* cell instance $18894 r0 *1 54.245,62.65
X$18894 1641 VIA_via2_5
* cell instance $18895 r0 *1 54.435,66.43
X$18895 1641 VIA_via1_4
* cell instance $18896 r0 *1 54.435,61.11
X$18896 1641 VIA_via1_4
* cell instance $18897 r0 *1 57.855,64.61
X$18897 1642 VIA_via1_7
* cell instance $18898 r0 *1 57.665,63.63
X$18898 1642 VIA_via1_4
* cell instance $18899 r0 *1 63.935,63.35
X$18899 1643 VIA_via2_5
* cell instance $18900 r0 *1 62.225,63.35
X$18900 1643 VIA_via2_5
* cell instance $18901 r0 *1 64.315,62.37
X$18901 1643 VIA_via1_4
* cell instance $18902 r0 *1 62.225,63.63
X$18902 1643 VIA_via1_4
* cell instance $18903 r0 *1 63.935,62.65
X$18903 1643 VIA_via1_4
* cell instance $18904 r0 *1 69.445,63.63
X$18904 1644 VIA_via2_5
* cell instance $18905 r0 *1 67.545,63.63
X$18905 1644 VIA_via2_5
* cell instance $18906 r0 *1 70.205,63.63
X$18906 1644 VIA_via2_5
* cell instance $18907 r0 *1 62.985,63.63
X$18907 1644 VIA_via2_5
* cell instance $18908 r0 *1 72.485,67.97
X$18908 1644 VIA_via2_5
* cell instance $18909 r0 *1 69.825,67.97
X$18909 1644 VIA_via2_5
* cell instance $18910 r0 *1 64.885,63.63
X$18910 1644 VIA_via1_4
* cell instance $18911 r0 *1 64.885,63.63
X$18911 1644 VIA_via2_5
* cell instance $18912 r0 *1 67.545,66.43
X$18912 1644 VIA_via1_4
* cell instance $18913 r0 *1 70.205,62.37
X$18913 1644 VIA_via1_4
* cell instance $18914 r0 *1 72.485,69.23
X$18914 1644 VIA_via1_4
* cell instance $18915 r0 *1 69.445,64.75
X$18915 1644 VIA_via1_4
* cell instance $18916 r0 *1 69.825,65.59
X$18916 1644 VIA_via1_7
* cell instance $18917 r0 *1 70.015,65.17
X$18917 1644 VIA_via1_4
* cell instance $18918 r0 *1 75.335,67.97
X$18918 1644 VIA_via1_4
* cell instance $18919 r0 *1 75.335,67.97
X$18919 1644 VIA_via2_5
* cell instance $18920 r0 *1 62.985,60.83
X$18920 1644 VIA_via1_4
* cell instance $18921 r0 *1 67.735,63.21
X$18921 1645 VIA_via2_5
* cell instance $18922 r0 *1 66.785,63.21
X$18922 1645 VIA_via2_5
* cell instance $18923 r0 *1 66.785,63.63
X$18923 1645 VIA_via1_4
* cell instance $18924 r0 *1 66.405,63.35
X$18924 1645 VIA_via1_4
* cell instance $18925 r0 *1 66.405,63.21
X$18925 1645 VIA_via2_5
* cell instance $18926 r0 *1 67.735,62.37
X$18926 1645 VIA_via1_4
* cell instance $18927 r0 *1 68.115,62.79
X$18927 1646 VIA_via1_7
* cell instance $18928 r0 *1 68.305,63.63
X$18928 1646 VIA_via1_4
* cell instance $18929 r0 *1 73.435,62.65
X$18929 1647 VIA_via2_5
* cell instance $18930 r0 *1 74.765,62.65
X$18930 1647 VIA_via2_5
* cell instance $18931 r0 *1 75.335,62.65
X$18931 1647 VIA_via2_5
* cell instance $18932 r0 *1 73.435,62.37
X$18932 1647 VIA_via1_4
* cell instance $18933 r0 *1 74.765,62.37
X$18933 1647 VIA_via1_4
* cell instance $18934 r0 *1 75.335,63.35
X$18934 1647 VIA_via1_4
* cell instance $18935 r0 *1 82.745,69.23
X$18935 1648 VIA_via2_5
* cell instance $18936 r0 *1 74.575,69.23
X$18936 1648 VIA_via2_5
* cell instance $18937 r0 *1 80.845,67.27
X$18937 1648 VIA_via2_5
* cell instance $18938 r0 *1 79.705,67.27
X$18938 1648 VIA_via2_5
* cell instance $18939 r0 *1 73.815,73.57
X$18939 1648 VIA_via1_4
* cell instance $18940 r0 *1 74.005,72.03
X$18940 1648 VIA_via1_4
* cell instance $18941 r0 *1 82.555,70.77
X$18941 1648 VIA_via1_4
* cell instance $18942 r0 *1 81.035,69.23
X$18942 1648 VIA_via1_4
* cell instance $18943 r0 *1 81.035,69.23
X$18943 1648 VIA_via2_5
* cell instance $18944 r0 *1 83.315,69.23
X$18944 1648 VIA_via1_4
* cell instance $18945 r0 *1 83.315,69.23
X$18945 1648 VIA_via2_5
* cell instance $18946 r0 *1 80.845,69.23
X$18946 1648 VIA_via1_4
* cell instance $18947 r0 *1 79.705,65.17
X$18947 1648 VIA_via1_4
* cell instance $18948 r0 *1 83.695,63.63
X$18948 1648 VIA_via1_4
* cell instance $18949 r0 *1 83.505,66.43
X$18949 1648 VIA_via1_4
* cell instance $18950 r0 *1 85.595,63.63
X$18950 1649 VIA_via1_4
* cell instance $18951 r0 *1 85.595,62.37
X$18951 1649 VIA_via1_4
* cell instance $18952 r0 *1 85.215,63.35
X$18952 1649 VIA_via1_4
* cell instance $18953 r0 *1 55.535,63.91
X$18953 1650 VIA_via5_0
* cell instance $18954 r0 *1 36.385,87.57
X$18954 1650 VIA_via2_5
* cell instance $18955 r0 *1 30.875,88.41
X$18955 1650 VIA_via2_5
* cell instance $18956 r0 *1 30.875,89.39
X$18956 1650 VIA_via2_5
* cell instance $18957 r0 *1 32.015,88.41
X$18957 1650 VIA_via2_5
* cell instance $18958 r0 *1 17.385,89.39
X$18958 1650 VIA_via2_5
* cell instance $18959 r0 *1 54.055,63.91
X$18959 1650 VIA_via2_5
* cell instance $18960 r0 *1 68.685,63.91
X$18960 1650 VIA_via2_5
* cell instance $18961 r0 *1 55.385,90.79
X$18961 1650 VIA_via2_5
* cell instance $18962 r0 *1 86.355,64.33
X$18962 1650 VIA_via2_5
* cell instance $18963 r0 *1 36.955,64.19
X$18963 1650 VIA_via2_5
* cell instance $18964 r0 *1 54.055,63.63
X$18964 1650 VIA_via1_4
* cell instance $18965 r0 *1 68.685,63.63
X$18965 1650 VIA_via1_4
* cell instance $18966 r0 *1 55.385,90.37
X$18966 1650 VIA_via1_4
* cell instance $18967 r0 *1 55.385,90.37
X$18967 1650 VIA_via2_5
* cell instance $18968 r0 *1 55.255,90.37
X$18968 1650 VIA_via3_2
* cell instance $18969 r0 *1 17.195,88.83
X$18969 1650 VIA_via1_4
* cell instance $18970 r0 *1 17.195,88.97
X$18970 1650 VIA_via2_5
* cell instance $18971 r0 *1 43.795,90.37
X$18971 1650 VIA_via1_4
* cell instance $18972 r0 *1 43.795,90.37
X$18972 1650 VIA_via2_5
* cell instance $18973 r0 *1 32.205,87.57
X$18973 1650 VIA_via1_4
* cell instance $18974 r0 *1 32.205,87.57
X$18974 1650 VIA_via2_5
* cell instance $18975 r0 *1 12.255,88.83
X$18975 1650 VIA_via1_4
* cell instance $18976 r0 *1 12.255,88.97
X$18976 1650 VIA_via2_5
* cell instance $18977 r0 *1 36.955,62.65
X$18977 1650 VIA_via1_4
* cell instance $18978 r0 *1 86.545,62.37
X$18978 1650 VIA_via1_4
* cell instance $18979 r0 *1 86.355,65.17
X$18979 1650 VIA_via1_4
* cell instance $18980 r0 *1 55.255,63.91
X$18980 1650 VIA_via4_0
* cell instance $18981 r0 *1 55.255,63.91
X$18981 1650 VIA_via3_2
* cell instance $18982 r0 *1 55.535,84.63
X$18982 1650 VIA_via4_0
* cell instance $18983 r0 *1 55.535,84.63
X$18983 1650 VIA_via5_0
* cell instance $18984 r0 *1 55.535,84.77
X$18984 1650 VIA_via3_2
* cell instance $18985 r0 *1 55.575,84.77
X$18985 1650 VIA_via2_5
* cell instance $18986 r0 *1 55.575,84.77
X$18986 1650 VIA_via1_4
* cell instance $18987 r0 *1 88.825,64.61
X$18987 1651 VIA_via1_7
* cell instance $18988 r0 *1 89.015,62.37
X$18988 1651 VIA_via1_4
* cell instance $18989 r0 *1 89.585,63.63
X$18989 1652 VIA_via1_4
* cell instance $18990 r0 *1 89.395,62.51
X$18990 1652 VIA_via1_4
* cell instance $18991 r0 *1 89.585,65.17
X$18991 1652 VIA_via1_4
* cell instance $18992 r0 *1 96.995,63.35
X$18992 1653 VIA_via1_4
* cell instance $18993 r0 *1 96.995,63.35
X$18993 1653 VIA_via2_5
* cell instance $18994 r0 *1 97.535,63.35
X$18994 1653 VIA_via3_2
* cell instance $18995 r0 *1 97.535,63.35
X$18995 1653 VIA_via4_0
* cell instance $18996 r0 *1 6.365,62.51
X$18996 1654 VIA_via2_5
* cell instance $18997 r0 *1 7.315,62.37
X$18997 1654 VIA_via1_4
* cell instance $18998 r0 *1 7.315,62.51
X$18998 1654 VIA_via2_5
* cell instance $18999 r0 *1 6.365,61.25
X$18999 1654 VIA_via1_4
* cell instance $19000 r0 *1 4.845,62.37
X$19000 1654 VIA_via1_4
* cell instance $19001 r0 *1 4.845,62.51
X$19001 1654 VIA_via2_5
* cell instance $19002 r0 *1 6.555,62.79
X$19002 1655 VIA_via1_7
* cell instance $19003 r0 *1 6.555,63.07
X$19003 1655 VIA_via2_5
* cell instance $19004 r0 *1 5.795,63.07
X$19004 1655 VIA_via2_5
* cell instance $19005 r0 *1 5.795,63.63
X$19005 1655 VIA_via1_4
* cell instance $19006 r0 *1 89.775,63.49
X$19006 1656 VIA_via1_4
* cell instance $19007 r0 *1 89.775,63.49
X$19007 1656 VIA_via2_5
* cell instance $19008 r0 *1 95.475,63.63
X$19008 1656 VIA_via1_4
* cell instance $19009 r0 *1 95.475,63.49
X$19009 1656 VIA_via2_5
* cell instance $19010 r0 *1 95.095,63.63
X$19010 1657 VIA_via1_4
* cell instance $19011 r0 *1 95.095,63.63
X$19011 1657 VIA_via2_5
* cell instance $19012 r0 *1 96.615,63.63
X$19012 1657 VIA_via1_4
* cell instance $19013 r0 *1 96.615,63.63
X$19013 1657 VIA_via2_5
* cell instance $19014 r0 *1 93.575,62.37
X$19014 1658 VIA_via1_4
* cell instance $19015 r0 *1 93.575,62.37
X$19015 1658 VIA_via2_5
* cell instance $19016 r0 *1 96.235,62.37
X$19016 1658 VIA_via1_4
* cell instance $19017 r0 *1 96.235,62.37
X$19017 1658 VIA_via2_5
* cell instance $19018 r0 *1 14.345,62.37
X$19018 1659 VIA_via1_4
* cell instance $19019 r0 *1 14.345,62.37
X$19019 1659 VIA_via2_5
* cell instance $19020 r0 *1 14.345,63.35
X$19020 1659 VIA_via1_4
* cell instance $19021 r0 *1 12.065,62.37
X$19021 1659 VIA_via1_4
* cell instance $19022 r0 *1 12.065,62.37
X$19022 1659 VIA_via2_5
* cell instance $19023 r0 *1 17.575,63.21
X$19023 1660 VIA_via1_7
* cell instance $19024 r0 *1 17.575,63.21
X$19024 1660 VIA_via2_5
* cell instance $19025 r0 *1 16.245,63.21
X$19025 1660 VIA_via2_5
* cell instance $19026 r0 *1 16.245,62.37
X$19026 1660 VIA_via1_4
* cell instance $19027 r0 *1 16.625,63.63
X$19027 1661 VIA_via1_4
* cell instance $19028 r0 *1 16.625,63.63
X$19028 1661 VIA_via2_5
* cell instance $19029 r0 *1 18.525,63.63
X$19029 1661 VIA_via1_4
* cell instance $19030 r0 *1 18.525,63.63
X$19030 1661 VIA_via2_5
* cell instance $19031 r0 *1 18.525,62.65
X$19031 1661 VIA_via1_4
* cell instance $19032 r0 *1 19.475,63.21
X$19032 1662 VIA_via1_7
* cell instance $19033 r0 *1 19.475,63.21
X$19033 1662 VIA_via2_5
* cell instance $19034 r0 *1 20.045,63.21
X$19034 1662 VIA_via2_5
* cell instance $19035 r0 *1 20.045,62.37
X$19035 1662 VIA_via1_4
* cell instance $19036 r0 *1 21.565,62.37
X$19036 1663 VIA_via1_4
* cell instance $19037 r0 *1 21.565,62.51
X$19037 1663 VIA_via2_5
* cell instance $19038 r0 *1 20.235,62.51
X$19038 1663 VIA_via1_4
* cell instance $19039 r0 *1 20.235,62.51
X$19039 1663 VIA_via2_5
* cell instance $19040 r0 *1 20.805,62.37
X$19040 1664 VIA_via1_4
* cell instance $19041 r0 *1 20.805,62.37
X$19041 1664 VIA_via2_5
* cell instance $19042 r0 *1 22.135,62.37
X$19042 1664 VIA_via1_4
* cell instance $19043 r0 *1 22.135,62.37
X$19043 1664 VIA_via2_5
* cell instance $19044 r0 *1 24.035,62.79
X$19044 1665 VIA_via1_7
* cell instance $19045 r0 *1 24.035,63.35
X$19045 1665 VIA_via2_5
* cell instance $19046 r0 *1 20.805,63.35
X$19046 1665 VIA_via2_5
* cell instance $19047 r0 *1 20.805,63.63
X$19047 1665 VIA_via1_4
* cell instance $19048 r0 *1 24.225,63.63
X$19048 1666 VIA_via2_5
* cell instance $19049 r0 *1 23.465,65.17
X$19049 1666 VIA_via2_5
* cell instance $19050 r0 *1 23.465,63.63
X$19050 1666 VIA_via1_4
* cell instance $19051 r0 *1 23.465,63.63
X$19051 1666 VIA_via2_5
* cell instance $19052 r0 *1 24.225,60.83
X$19052 1666 VIA_via1_4
* cell instance $19053 r0 *1 25.365,65.17
X$19053 1666 VIA_via1_4
* cell instance $19054 r0 *1 25.365,65.17
X$19054 1666 VIA_via2_5
* cell instance $19055 r0 *1 31.255,63.35
X$19055 1667 VIA_via2_5
* cell instance $19056 r0 *1 31.255,63.63
X$19056 1667 VIA_via1_4
* cell instance $19057 r0 *1 32.585,63.35
X$19057 1667 VIA_via1_4
* cell instance $19058 r0 *1 32.585,63.35
X$19058 1667 VIA_via2_5
* cell instance $19059 r0 *1 33.345,63.63
X$19059 1668 VIA_via1_4
* cell instance $19060 r0 *1 33.345,63.63
X$19060 1668 VIA_via2_5
* cell instance $19061 r0 *1 32.015,63.63
X$19061 1668 VIA_via1_4
* cell instance $19062 r0 *1 32.015,63.63
X$19062 1668 VIA_via2_5
* cell instance $19063 r0 *1 88.255,62.37
X$19063 1669 VIA_via1_4
* cell instance $19064 r0 *1 88.065,62.37
X$19064 1669 VIA_via1_4
* cell instance $19065 r0 *1 42.085,62.79
X$19065 1670 VIA_via1_7
* cell instance $19066 r0 *1 42.085,62.79
X$19066 1670 VIA_via2_5
* cell instance $19067 r0 *1 41.515,62.79
X$19067 1670 VIA_via2_5
* cell instance $19068 r0 *1 41.515,63.63
X$19068 1670 VIA_via1_4
* cell instance $19069 r0 *1 41.135,62.37
X$19069 1671 VIA_via1_4
* cell instance $19070 r0 *1 41.135,62.37
X$19070 1671 VIA_via2_5
* cell instance $19071 r0 *1 43.795,62.37
X$19071 1671 VIA_via1_4
* cell instance $19072 r0 *1 43.795,62.37
X$19072 1671 VIA_via2_5
* cell instance $19073 r0 *1 43.795,63.35
X$19073 1671 VIA_via1_4
* cell instance $19074 r0 *1 86.545,63.63
X$19074 1672 VIA_via1_4
* cell instance $19075 r0 *1 86.545,63.63
X$19075 1672 VIA_via2_5
* cell instance $19076 r0 *1 82.935,63.63
X$19076 1672 VIA_via1_4
* cell instance $19077 r0 *1 82.935,63.63
X$19077 1672 VIA_via2_5
* cell instance $19078 r0 *1 44.175,62.79
X$19078 1673 VIA_via1_7
* cell instance $19079 r0 *1 53.675,63.07
X$19079 1673 VIA_via2_5
* cell instance $19080 r0 *1 44.175,63.07
X$19080 1673 VIA_via2_5
* cell instance $19081 r0 *1 53.675,63.63
X$19081 1673 VIA_via1_4
* cell instance $19082 r0 *1 86.165,62.37
X$19082 1674 VIA_via1_4
* cell instance $19083 r0 *1 85.975,62.37
X$19083 1674 VIA_via1_4
* cell instance $19084 r0 *1 49.875,63.63
X$19084 1675 VIA_via1_4
* cell instance $19085 r0 *1 49.875,63.63
X$19085 1675 VIA_via2_5
* cell instance $19086 r0 *1 46.265,63.63
X$19086 1675 VIA_via1_4
* cell instance $19087 r0 *1 46.265,63.63
X$19087 1675 VIA_via2_5
* cell instance $19088 r0 *1 52.725,62.37
X$19088 1676 VIA_via1_4
* cell instance $19089 r0 *1 52.725,62.37
X$19089 1676 VIA_via2_5
* cell instance $19090 r0 *1 49.115,62.37
X$19090 1676 VIA_via1_4
* cell instance $19091 r0 *1 49.115,62.37
X$19091 1676 VIA_via2_5
* cell instance $19092 r0 *1 54.625,64.75
X$19092 1677 VIA_via1_4
* cell instance $19093 r0 *1 53.105,63.63
X$19093 1677 VIA_via1_4
* cell instance $19094 r0 *1 53.105,63.63
X$19094 1677 VIA_via2_5
* cell instance $19095 r0 *1 54.625,63.63
X$19095 1677 VIA_via1_4
* cell instance $19096 r0 *1 54.625,63.63
X$19096 1677 VIA_via2_5
* cell instance $19097 r0 *1 78.945,61.11
X$19097 1678 VIA_via1_4
* cell instance $19098 r0 *1 78.945,62.37
X$19098 1678 VIA_via1_4
* cell instance $19099 r0 *1 54.435,62.79
X$19099 1679 VIA_via1_7
* cell instance $19100 r0 *1 54.435,62.79
X$19100 1679 VIA_via2_5
* cell instance $19101 r0 *1 55.005,62.79
X$19101 1679 VIA_via2_5
* cell instance $19102 r0 *1 55.005,65.17
X$19102 1679 VIA_via1_4
* cell instance $19103 r0 *1 55.575,63.63
X$19103 1680 VIA_via1_4
* cell instance $19104 r0 *1 55.765,63.63
X$19104 1680 VIA_via1_4
* cell instance $19105 r0 *1 76.285,62.51
X$19105 1681 VIA_via1_4
* cell instance $19106 r0 *1 76.285,62.51
X$19106 1681 VIA_via2_5
* cell instance $19107 r0 *1 77.995,62.37
X$19107 1681 VIA_via1_4
* cell instance $19108 r0 *1 77.995,62.51
X$19108 1681 VIA_via2_5
* cell instance $19109 r0 *1 56.525,61.39
X$19109 1682 VIA_via1_7
* cell instance $19110 r0 *1 56.525,62.37
X$19110 1682 VIA_via1_4
* cell instance $19111 r0 *1 76.095,62.37
X$19111 1683 VIA_via1_4
* cell instance $19112 r0 *1 76.095,62.37
X$19112 1683 VIA_via2_5
* cell instance $19113 r0 *1 75.715,62.37
X$19113 1683 VIA_via1_4
* cell instance $19114 r0 *1 75.715,62.37
X$19114 1683 VIA_via2_5
* cell instance $19115 r0 *1 63.365,68.39
X$19115 1684 VIA_via1_7
* cell instance $19116 r0 *1 63.365,68.39
X$19116 1684 VIA_via2_5
* cell instance $19117 r0 *1 66.405,68.39
X$19117 1684 VIA_via2_5
* cell instance $19118 r0 *1 61.655,68.39
X$19118 1684 VIA_via2_5
* cell instance $19119 r0 *1 63.555,68.39
X$19119 1684 VIA_via2_5
* cell instance $19120 r0 *1 61.655,63.63
X$19120 1684 VIA_via2_5
* cell instance $19121 r0 *1 61.655,63.07
X$19121 1684 VIA_via2_5
* cell instance $19122 r0 *1 62.415,63.07
X$19122 1684 VIA_via2_5
* cell instance $19123 r0 *1 62.415,62.37
X$19123 1684 VIA_via1_4
* cell instance $19124 r0 *1 63.555,67.97
X$19124 1684 VIA_via1_4
* cell instance $19125 r0 *1 66.405,70.77
X$19125 1684 VIA_via1_4
* cell instance $19126 r0 *1 61.465,70.77
X$19126 1684 VIA_via1_4
* cell instance $19127 r0 *1 61.655,65.17
X$19127 1684 VIA_via1_4
* cell instance $19128 r0 *1 61.465,66.43
X$19128 1684 VIA_via1_4
* cell instance $19129 r0 *1 61.085,72.03
X$19129 1684 VIA_via1_4
* cell instance $19130 r0 *1 58.425,63.63
X$19130 1684 VIA_via1_4
* cell instance $19131 r0 *1 58.425,63.63
X$19131 1684 VIA_via2_5
* cell instance $19132 r0 *1 64.125,63.63
X$19132 1685 VIA_via1_4
* cell instance $19133 r0 *1 64.125,63.49
X$19133 1685 VIA_via2_5
* cell instance $19134 r0 *1 67.735,63.49
X$19134 1685 VIA_via1_4
* cell instance $19135 r0 *1 67.735,63.49
X$19135 1685 VIA_via2_5
* cell instance $19136 r0 *1 80.845,78.75
X$19136 1686 VIA_via2_5
* cell instance $19137 r0 *1 91.295,85.33
X$19137 1686 VIA_via2_5
* cell instance $19138 r0 *1 67.355,74.55
X$19138 1686 VIA_via2_5
* cell instance $19139 r0 *1 67.355,78.75
X$19139 1686 VIA_via2_5
* cell instance $19140 r0 *1 80.845,85.33
X$19140 1686 VIA_via2_5
* cell instance $19141 r0 *1 66.215,74.55
X$19141 1686 VIA_via2_5
* cell instance $19142 r0 *1 82.935,85.33
X$19142 1686 VIA_via2_5
* cell instance $19143 r0 *1 91.675,64.89
X$19143 1686 VIA_via2_5
* cell instance $19144 r0 *1 90.345,64.89
X$19144 1686 VIA_via2_5
* cell instance $19145 r0 *1 65.455,62.385
X$19145 1686 VIA_via1_4
* cell instance $19146 r0 *1 65.455,62.37
X$19146 1686 VIA_via2_5
* cell instance $19147 r0 *1 66.215,74.83
X$19147 1686 VIA_via1_4
* cell instance $19148 r0 *1 80.275,90.37
X$19148 1686 VIA_via1_4
* cell instance $19149 r0 *1 80.275,90.37
X$19149 1686 VIA_via2_5
* cell instance $19150 r0 *1 80.845,87.15
X$19150 1686 VIA_via1_4
* cell instance $19151 r0 *1 80.465,87.85
X$19151 1686 VIA_via1_4
* cell instance $19152 r0 *1 82.745,86.03
X$19152 1686 VIA_via1_4
* cell instance $19153 r0 *1 91.295,86.03
X$19153 1686 VIA_via1_4
* cell instance $19154 r0 *1 88.825,90.37
X$19154 1686 VIA_via1_4
* cell instance $19155 r0 *1 88.825,90.37
X$19155 1686 VIA_via2_5
* cell instance $19156 r0 *1 90.535,83.23
X$19156 1686 VIA_via1_4
* cell instance $19157 r0 *1 90.535,83.23
X$19157 1686 VIA_via2_5
* cell instance $19158 r0 *1 90.535,83.23
X$19158 1686 VIA_via3_2
* cell instance $19159 r0 *1 90.725,80.43
X$19159 1686 VIA_via1_4
* cell instance $19160 r0 *1 91.485,79.17
X$19160 1686 VIA_via1_4
* cell instance $19161 r0 *1 90.345,63.63
X$19161 1686 VIA_via1_4
* cell instance $19162 r0 *1 81.855,90.51
X$19162 1686 VIA_via4_0
* cell instance $19163 r0 *1 81.855,90.37
X$19163 1686 VIA_via3_2
* cell instance $19164 r0 *1 90.535,85.33
X$19164 1686 VIA_via3_2
* cell instance $19165 r0 *1 65.615,74.55
X$19165 1686 VIA_via3_2
* cell instance $19166 r0 *1 65.615,62.37
X$19166 1686 VIA_via3_2
* cell instance $19167 r0 *1 88.575,90.37
X$19167 1686 VIA_via3_2
* cell instance $19168 r0 *1 88.575,90.51
X$19168 1686 VIA_via4_0
* cell instance $19169 r0 *1 66.405,62.37
X$19169 1687 VIA_via1_4
* cell instance $19170 r0 *1 66.405,62.51
X$19170 1687 VIA_via2_5
* cell instance $19171 r0 *1 65.265,62.51
X$19171 1687 VIA_via1_4
* cell instance $19172 r0 *1 65.265,62.51
X$19172 1687 VIA_via2_5
* cell instance $19173 r0 *1 8.265,64.61
X$19173 1688 VIA_via1_7
* cell instance $19174 r0 *1 8.265,64.47
X$19174 1688 VIA_via2_5
* cell instance $19175 r0 *1 4.295,64.47
X$19175 1688 VIA_via3_2
* cell instance $19176 r0 *1 4.295,64.47
X$19176 1688 VIA_via4_0
* cell instance $19177 r0 *1 4.845,64.89
X$19177 1689 VIA_via2_5
* cell instance $19178 r0 *1 6.745,64.89
X$19178 1689 VIA_via2_5
* cell instance $19179 r0 *1 4.085,64.89
X$19179 1689 VIA_via2_5
* cell instance $19180 r0 *1 6.745,65.17
X$19180 1689 VIA_via1_4
* cell instance $19181 r0 *1 4.085,63.63
X$19181 1689 VIA_via1_4
* cell instance $19182 r0 *1 4.845,65.17
X$19182 1689 VIA_via1_4
* cell instance $19183 r0 *1 11.115,64.19
X$19183 1690 VIA_via1_7
* cell instance $19184 r0 *1 12.255,65.17
X$19184 1690 VIA_via1_4
* cell instance $19185 r0 *1 10.925,64.61
X$19185 1691 VIA_via1_7
* cell instance $19186 r0 *1 12.065,65.17
X$19186 1691 VIA_via1_4
* cell instance $19187 r0 *1 17.195,65.17
X$19187 1692 VIA_via2_5
* cell instance $19188 r0 *1 13.395,65.17
X$19188 1692 VIA_via1_4
* cell instance $19189 r0 *1 13.395,65.17
X$19189 1692 VIA_via2_5
* cell instance $19190 r0 *1 17.195,66.15
X$19190 1692 VIA_via1_4
* cell instance $19191 r0 *1 14.155,65.17
X$19191 1692 VIA_via1_4
* cell instance $19192 r0 *1 14.155,65.17
X$19192 1692 VIA_via2_5
* cell instance $19193 r0 *1 23.845,66.43
X$19193 1693 VIA_via2_5
* cell instance $19194 r0 *1 21.565,65.17
X$19194 1693 VIA_via2_5
* cell instance $19195 r0 *1 23.845,67.13
X$19195 1693 VIA_via2_5
* cell instance $19196 r0 *1 21.565,66.43
X$19196 1693 VIA_via2_5
* cell instance $19197 r0 *1 27.265,67.13
X$19197 1693 VIA_via2_5
* cell instance $19198 r0 *1 27.455,67.13
X$19198 1693 VIA_via2_5
* cell instance $19199 r0 *1 24.985,67.13
X$19199 1693 VIA_via2_5
* cell instance $19200 r0 *1 21.565,63.63
X$19200 1693 VIA_via1_4
* cell instance $19201 r0 *1 23.845,65.17
X$19201 1693 VIA_via1_4
* cell instance $19202 r0 *1 22.895,66.43
X$19202 1693 VIA_via1_4
* cell instance $19203 r0 *1 22.895,66.43
X$19203 1693 VIA_via2_5
* cell instance $19204 r0 *1 19.665,65.17
X$19204 1693 VIA_via1_4
* cell instance $19205 r0 *1 19.665,65.17
X$19205 1693 VIA_via2_5
* cell instance $19206 r0 *1 24.985,66.85
X$19206 1693 VIA_via1_4
* cell instance $19207 r0 *1 27.075,65.17
X$19207 1693 VIA_via1_4
* cell instance $19208 r0 *1 28.595,69.23
X$19208 1693 VIA_via1_4
* cell instance $19209 r0 *1 24.985,67.97
X$19209 1693 VIA_via1_4
* cell instance $19210 r0 *1 27.455,67.97
X$19210 1693 VIA_via1_4
* cell instance $19211 r0 *1 28.785,66.71
X$19211 1694 VIA_via2_5
* cell instance $19212 r0 *1 29.355,66.71
X$19212 1694 VIA_via2_5
* cell instance $19213 r0 *1 27.645,66.71
X$19213 1694 VIA_via2_5
* cell instance $19214 r0 *1 28.595,64.89
X$19214 1694 VIA_via1_4
* cell instance $19215 r0 *1 27.645,66.43
X$19215 1694 VIA_via1_4
* cell instance $19216 r0 *1 29.355,67.97
X$19216 1694 VIA_via1_4
* cell instance $19217 r0 *1 30.685,66.71
X$19217 1695 VIA_via2_5
* cell instance $19218 r0 *1 30.305,66.71
X$19218 1695 VIA_via1_4
* cell instance $19219 r0 *1 30.305,66.71
X$19219 1695 VIA_via2_5
* cell instance $19220 r0 *1 31.445,63.63
X$19220 1695 VIA_via1_4
* cell instance $19221 r0 *1 31.635,63.91
X$19221 1696 VIA_via1_7
* cell instance $19222 r0 *1 31.255,65.17
X$19222 1696 VIA_via1_4
* cell instance $19223 r0 *1 38.855,66.01
X$19223 1697 VIA_via1_7
* cell instance $19224 r0 *1 39.235,65.17
X$19224 1697 VIA_via1_4
* cell instance $19225 r0 *1 49.115,64.89
X$19225 1698 VIA_via1_4
* cell instance $19226 r0 *1 48.545,66.43
X$19226 1698 VIA_via1_4
* cell instance $19227 r0 *1 55.955,63.91
X$19227 1699 VIA_via1_4
* cell instance $19228 r0 *1 55.765,65.17
X$19228 1699 VIA_via1_4
* cell instance $19229 r0 *1 55.955,65.17
X$19229 1700 VIA_via1_4
* cell instance $19230 r0 *1 56.335,64.89
X$19230 1700 VIA_via1_4
* cell instance $19231 r0 *1 59.375,65.03
X$19231 1701 VIA_via1_4
* cell instance $19232 r0 *1 59.375,65.03
X$19232 1701 VIA_via2_5
* cell instance $19233 r0 *1 56.145,65.17
X$19233 1701 VIA_via1_4
* cell instance $19234 r0 *1 56.145,65.17
X$19234 1701 VIA_via2_5
* cell instance $19235 r0 *1 59.945,65.17
X$19235 1702 VIA_via2_5
* cell instance $19236 r0 *1 57.475,65.17
X$19236 1702 VIA_via1_4
* cell instance $19237 r0 *1 57.475,65.17
X$19237 1702 VIA_via2_5
* cell instance $19238 r0 *1 58.995,65.17
X$19238 1702 VIA_via1_4
* cell instance $19239 r0 *1 58.995,65.17
X$19239 1702 VIA_via2_5
* cell instance $19240 r0 *1 59.945,64.05
X$19240 1702 VIA_via1_4
* cell instance $19241 r0 *1 61.085,65.03
X$19241 1703 VIA_via2_5
* cell instance $19242 r0 *1 60.895,65.17
X$19242 1703 VIA_via1_4
* cell instance $19243 r0 *1 64.505,65.03
X$19243 1703 VIA_via1_4
* cell instance $19244 r0 *1 64.505,65.03
X$19244 1703 VIA_via2_5
* cell instance $19245 r0 *1 67.165,66.15
X$19245 1704 VIA_via2_5
* cell instance $19246 r0 *1 67.165,62.37
X$19246 1704 VIA_via1_4
* cell instance $19247 r0 *1 69.065,66.15
X$19247 1704 VIA_via1_4
* cell instance $19248 r0 *1 69.065,66.15
X$19248 1704 VIA_via2_5
* cell instance $19249 r0 *1 67.165,65.17
X$19249 1704 VIA_via1_4
* cell instance $19250 r0 *1 88.635,66.01
X$19250 1705 VIA_via1_7
* cell instance $19251 r0 *1 88.445,65.17
X$19251 1705 VIA_via1_4
* cell instance $19252 r0 *1 78.565,65.31
X$19252 1706 VIA_via2_5
* cell instance $19253 r0 *1 89.395,63.63
X$19253 1706 VIA_via1_4
* cell instance $19254 r0 *1 89.395,65.17
X$19254 1706 VIA_via1_4
* cell instance $19255 r0 *1 89.395,65.31
X$19255 1706 VIA_via2_5
* cell instance $19256 r0 *1 78.375,68.95
X$19256 1706 VIA_via1_4
* cell instance $19257 r0 *1 92.815,64.19
X$19257 1707 VIA_via1_7
* cell instance $19258 r0 *1 93.385,66.43
X$19258 1707 VIA_via1_4
* cell instance $19259 r0 *1 94.905,64.61
X$19259 1708 VIA_via1_7
* cell instance $19260 r0 *1 95.285,63.63
X$19260 1708 VIA_via1_4
* cell instance $19261 r0 *1 3.515,65.03
X$19261 1709 VIA_via2_5
* cell instance $19262 r0 *1 3.515,66.43
X$19262 1709 VIA_via1_4
* cell instance $19263 r0 *1 6.175,65.03
X$19263 1709 VIA_via1_4
* cell instance $19264 r0 *1 6.175,65.03
X$19264 1709 VIA_via2_5
* cell instance $19265 r0 *1 4.465,64.19
X$19265 1710 VIA_via1_7
* cell instance $19266 r0 *1 4.465,64.19
X$19266 1710 VIA_via2_5
* cell instance $19267 r0 *1 2.565,64.19
X$19267 1710 VIA_via2_5
* cell instance $19268 r0 *1 2.565,65.17
X$19268 1710 VIA_via1_4
* cell instance $19269 r0 *1 90.725,65.03
X$19269 1711 VIA_via2_5
* cell instance $19270 r0 *1 90.725,67.97
X$19270 1711 VIA_via1_4
* cell instance $19271 r0 *1 90.155,65.03
X$19271 1711 VIA_via1_4
* cell instance $19272 r0 *1 90.155,65.03
X$19272 1711 VIA_via2_5
* cell instance $19273 r0 *1 7.695,64.61
X$19273 1712 VIA_via1_7
* cell instance $19274 r0 *1 7.695,64.61
X$19274 1712 VIA_via2_5
* cell instance $19275 r0 *1 10.545,64.61
X$19275 1712 VIA_via2_5
* cell instance $19276 r0 *1 10.545,65.17
X$19276 1712 VIA_via1_4
* cell instance $19277 r0 *1 86.355,64.61
X$19277 1713 VIA_via1_7
* cell instance $19278 r0 *1 86.355,64.61
X$19278 1713 VIA_via2_5
* cell instance $19279 r0 *1 89.205,64.61
X$19279 1713 VIA_via2_5
* cell instance $19280 r0 *1 89.205,62.37
X$19280 1713 VIA_via1_4
* cell instance $19281 r0 *1 86.165,65.03
X$19281 1714 VIA_via2_5
* cell instance $19282 r0 *1 91.485,68.11
X$19282 1714 VIA_via2_5
* cell instance $19283 r0 *1 86.165,68.11
X$19283 1714 VIA_via2_5
* cell instance $19284 r0 *1 94.525,69.23
X$19284 1714 VIA_via2_5
* cell instance $19285 r0 *1 83.125,65.03
X$19285 1714 VIA_via2_5
* cell instance $19286 r0 *1 89.395,68.11
X$19286 1714 VIA_via1_4
* cell instance $19287 r0 *1 89.395,68.11
X$19287 1714 VIA_via2_5
* cell instance $19288 r0 *1 86.355,72.03
X$19288 1714 VIA_via1_4
* cell instance $19289 r0 *1 86.545,69.23
X$19289 1714 VIA_via1_4
* cell instance $19290 r0 *1 89.965,67.97
X$19290 1714 VIA_via1_4
* cell instance $19291 r0 *1 89.965,68.11
X$19291 1714 VIA_via2_5
* cell instance $19292 r0 *1 94.525,67.97
X$19292 1714 VIA_via1_4
* cell instance $19293 r0 *1 91.485,69.23
X$19293 1714 VIA_via1_4
* cell instance $19294 r0 *1 91.485,69.23
X$19294 1714 VIA_via2_5
* cell instance $19295 r0 *1 90.345,66.43
X$19295 1714 VIA_via1_4
* cell instance $19296 r0 *1 83.125,62.37
X$19296 1714 VIA_via1_4
* cell instance $19297 r0 *1 76.665,64.19
X$19297 1715 VIA_via1_7
* cell instance $19298 r0 *1 76.665,64.19
X$19298 1715 VIA_via2_5
* cell instance $19299 r0 *1 75.715,64.19
X$19299 1715 VIA_via2_5
* cell instance $19300 r0 *1 75.715,65.17
X$19300 1715 VIA_via1_4
* cell instance $19301 r0 *1 24.415,64.19
X$19301 1716 VIA_via1_7
* cell instance $19302 r0 *1 23.085,64.75
X$19302 1716 VIA_via2_5
* cell instance $19303 r0 *1 24.415,64.75
X$19303 1716 VIA_via2_5
* cell instance $19304 r0 *1 23.085,65.17
X$19304 1716 VIA_via1_4
* cell instance $19305 r0 *1 9.975,67.97
X$19305 1717 VIA_via2_5
* cell instance $19306 r0 *1 9.785,69.23
X$19306 1717 VIA_via1_4
* cell instance $19307 r0 *1 10.925,67.97
X$19307 1717 VIA_via1_4
* cell instance $19308 r0 *1 10.925,67.97
X$19308 1717 VIA_via2_5
* cell instance $19309 r0 *1 10.165,66.85
X$19309 1717 VIA_via1_4
* cell instance $19310 r0 *1 32.395,66.71
X$19310 1718 VIA_via1_7
* cell instance $19311 r0 *1 7.885,65.59
X$19311 1718 VIA_via2_5
* cell instance $19312 r0 *1 32.395,65.45
X$19312 1718 VIA_via2_5
* cell instance $19313 r0 *1 7.885,65.17
X$19313 1718 VIA_via1_4
* cell instance $19314 r0 *1 13.775,65.59
X$19314 1719 VIA_via1_7
* cell instance $19315 r0 *1 13.585,66.43
X$19315 1719 VIA_via1_4
* cell instance $19316 r0 *1 29.545,65.31
X$19316 1720 VIA_via2_5
* cell instance $19317 r0 *1 12.255,65.45
X$19317 1720 VIA_via1_4
* cell instance $19318 r0 *1 12.255,65.45
X$19318 1720 VIA_via2_5
* cell instance $19319 r0 *1 29.545,66.43
X$19319 1720 VIA_via1_4
* cell instance $19320 r0 *1 29.545,66.43
X$19320 1720 VIA_via2_5
* cell instance $19321 r0 *1 30.875,66.43
X$19321 1720 VIA_via1_4
* cell instance $19322 r0 *1 30.875,66.43
X$19322 1720 VIA_via2_5
* cell instance $19323 r0 *1 15.105,65.59
X$19323 1721 VIA_via1_7
* cell instance $19324 r0 *1 14.915,66.43
X$19324 1721 VIA_via1_4
* cell instance $19325 r0 *1 19.285,66.01
X$19325 1722 VIA_via1_7
* cell instance $19326 r0 *1 18.905,65.17
X$19326 1722 VIA_via1_4
* cell instance $19327 r0 *1 20.235,66.15
X$19327 1723 VIA_via2_5
* cell instance $19328 r0 *1 24.415,66.15
X$19328 1723 VIA_via1_4
* cell instance $19329 r0 *1 24.415,66.15
X$19329 1723 VIA_via2_5
* cell instance $19330 r0 *1 20.235,66.43
X$19330 1723 VIA_via1_4
* cell instance $19331 r0 *1 20.045,67.97
X$19331 1723 VIA_via1_4
* cell instance $19332 r0 *1 21.185,66.29
X$19332 1724 VIA_via2_5
* cell instance $19333 r0 *1 18.335,66.43
X$19333 1724 VIA_via1_4
* cell instance $19334 r0 *1 18.335,66.29
X$19334 1724 VIA_via2_5
* cell instance $19335 r0 *1 21.185,65.45
X$19335 1724 VIA_via1_4
* cell instance $19336 r0 *1 20.805,66.43
X$19336 1724 VIA_via1_4
* cell instance $19337 r0 *1 20.805,66.29
X$19337 1724 VIA_via2_5
* cell instance $19338 r0 *1 31.635,84.21
X$19338 1725 VIA_via1_7
* cell instance $19339 r0 *1 31.635,84.21
X$19339 1725 VIA_via2_5
* cell instance $19340 r0 *1 27.645,86.03
X$19340 1725 VIA_via2_5
* cell instance $19341 r0 *1 33.535,84.21
X$19341 1725 VIA_via2_5
* cell instance $19342 r0 *1 26.885,84.35
X$19342 1725 VIA_via2_5
* cell instance $19343 r0 *1 33.535,83.23
X$19343 1725 VIA_via2_5
* cell instance $19344 r0 *1 28.405,84.35
X$19344 1725 VIA_via2_5
* cell instance $19345 r0 *1 30.305,84.35
X$19345 1725 VIA_via2_5
* cell instance $19346 r0 *1 26.695,66.85
X$19346 1725 VIA_via2_5
* cell instance $19347 r0 *1 33.535,66.85
X$19347 1725 VIA_via2_5
* cell instance $19348 r0 *1 28.215,66.85
X$19348 1725 VIA_via2_5
* cell instance $19349 r0 *1 30.305,86.03
X$19349 1725 VIA_via1_4
* cell instance $19350 r0 *1 26.885,86.03
X$19350 1725 VIA_via1_4
* cell instance $19351 r0 *1 26.885,86.03
X$19351 1725 VIA_via2_5
* cell instance $19352 r0 *1 27.645,88.83
X$19352 1725 VIA_via1_4
* cell instance $19353 r0 *1 28.975,88.83
X$19353 1725 VIA_via1_4
* cell instance $19354 r0 *1 28.405,80.43
X$19354 1725 VIA_via1_4
* cell instance $19355 r0 *1 34.295,83.23
X$19355 1725 VIA_via1_4
* cell instance $19356 r0 *1 34.295,83.23
X$19356 1725 VIA_via2_5
* cell instance $19357 r0 *1 26.695,66.43
X$19357 1725 VIA_via1_4
* cell instance $19358 r0 *1 28.215,66.43
X$19358 1725 VIA_via1_4
* cell instance $19359 r0 *1 33.915,67.97
X$19359 1725 VIA_via1_4
* cell instance $19360 r0 *1 33.535,70.77
X$19360 1725 VIA_via1_4
* cell instance $19361 r0 *1 31.065,66.57
X$19361 1726 VIA_via1_7
* cell instance $19362 r0 *1 22.325,66.29
X$19362 1726 VIA_via2_5
* cell instance $19363 r0 *1 31.255,66.29
X$19363 1726 VIA_via2_5
* cell instance $19364 r0 *1 22.325,62.65
X$19364 1726 VIA_via1_4
* cell instance $19365 r0 *1 29.355,66.43
X$19365 1726 VIA_via1_4
* cell instance $19366 r0 *1 29.355,66.29
X$19366 1726 VIA_via2_5
* cell instance $19367 r0 *1 66.975,74.41
X$19367 1727 VIA_via1_7
* cell instance $19368 r0 *1 66.975,74.41
X$19368 1727 VIA_via2_5
* cell instance $19369 r0 *1 36.765,73.99
X$19369 1727 VIA_via2_5
* cell instance $19370 r0 *1 36.765,75.53
X$19370 1727 VIA_via2_5
* cell instance $19371 r0 *1 31.635,73.99
X$19371 1727 VIA_via2_5
* cell instance $19372 r0 *1 29.545,73.99
X$19372 1727 VIA_via2_5
* cell instance $19373 r0 *1 29.545,74.69
X$19373 1727 VIA_via2_5
* cell instance $19374 r0 *1 28.595,74.69
X$19374 1727 VIA_via2_5
* cell instance $19375 r0 *1 42.085,75.67
X$19375 1727 VIA_via2_5
* cell instance $19376 r0 *1 55.385,67.13
X$19376 1727 VIA_via2_5
* cell instance $19377 r0 *1 55.765,76.09
X$19377 1727 VIA_via2_5
* cell instance $19378 r0 *1 51.965,75.67
X$19378 1727 VIA_via2_5
* cell instance $19379 r0 *1 51.965,76.09
X$19379 1727 VIA_via2_5
* cell instance $19380 r0 *1 68.495,74.41
X$19380 1727 VIA_via2_5
* cell instance $19381 r0 *1 51.965,76.37
X$19381 1727 VIA_via1_4
* cell instance $19382 r0 *1 55.955,76.37
X$19382 1727 VIA_via1_4
* cell instance $19383 r0 *1 69.065,67.97
X$19383 1727 VIA_via1_4
* cell instance $19384 r0 *1 42.085,76.37
X$19384 1727 VIA_via1_4
* cell instance $19385 r0 *1 36.765,76.37
X$19385 1727 VIA_via1_4
* cell instance $19386 r0 *1 28.785,76.37
X$19386 1727 VIA_via1_4
* cell instance $19387 r0 *1 29.735,74.83
X$19387 1727 VIA_via1_4
* cell instance $19388 r0 *1 30.305,66.43
X$19388 1727 VIA_via1_4
* cell instance $19389 r0 *1 55.385,66.43
X$19389 1727 VIA_via1_4
* cell instance $19390 r0 *1 31.635,73.57
X$19390 1727 VIA_via1_4
* cell instance $19391 r0 *1 55.535,76.09
X$19391 1727 VIA_via3_2
* cell instance $19392 r0 *1 55.535,74.41
X$19392 1727 VIA_via3_2
* cell instance $19393 r0 *1 55.535,67.13
X$19393 1727 VIA_via3_2
* cell instance $19394 r0 *1 35.435,76.65
X$19394 1728 VIA_via2_5
* cell instance $19395 r0 *1 34.485,76.93
X$19395 1728 VIA_via2_5
* cell instance $19396 r0 *1 35.435,76.93
X$19396 1728 VIA_via2_5
* cell instance $19397 r0 *1 35.435,73.71
X$19397 1728 VIA_via2_5
* cell instance $19398 r0 *1 56.335,70.21
X$19398 1728 VIA_via2_5
* cell instance $19399 r0 *1 58.615,76.65
X$19399 1728 VIA_via2_5
* cell instance $19400 r0 *1 63.935,70.21
X$19400 1728 VIA_via2_5
* cell instance $19401 r0 *1 33.725,73.29
X$19401 1728 VIA_via2_5
* cell instance $19402 r0 *1 43.985,71.33
X$19402 1728 VIA_via2_5
* cell instance $19403 r0 *1 44.745,71.33
X$19403 1728 VIA_via2_5
* cell instance $19404 r0 *1 52.915,76.37
X$19404 1728 VIA_via1_4
* cell instance $19405 r0 *1 52.915,76.51
X$19405 1728 VIA_via2_5
* cell instance $19406 r0 *1 58.805,77.63
X$19406 1728 VIA_via1_4
* cell instance $19407 r0 *1 64.505,67.97
X$19407 1728 VIA_via1_4
* cell instance $19408 r0 *1 56.335,70.77
X$19408 1728 VIA_via1_4
* cell instance $19409 r0 *1 39.045,76.37
X$19409 1728 VIA_via1_4
* cell instance $19410 r0 *1 39.045,76.51
X$19410 1728 VIA_via2_5
* cell instance $19411 r0 *1 43.795,76.37
X$19411 1728 VIA_via1_4
* cell instance $19412 r0 *1 43.795,76.23
X$19412 1728 VIA_via2_5
* cell instance $19413 r0 *1 34.295,79.17
X$19413 1728 VIA_via1_4
* cell instance $19414 r0 *1 34.485,77.63
X$19414 1728 VIA_via1_4
* cell instance $19415 r0 *1 44.745,71.05
X$19415 1728 VIA_via1_4
* cell instance $19416 r0 *1 33.915,66.43
X$19416 1728 VIA_via1_4
* cell instance $19417 r0 *1 32.965,73.57
X$19417 1728 VIA_via1_4
* cell instance $19418 r0 *1 32.965,73.71
X$19418 1728 VIA_via2_5
* cell instance $19419 r0 *1 54.975,76.51
X$19419 1728 VIA_via3_2
* cell instance $19420 r0 *1 54.975,70.21
X$19420 1728 VIA_via3_2
* cell instance $19421 r0 *1 54.975,71.33
X$19421 1728 VIA_via3_2
* cell instance $19422 r0 *1 39.805,65.45
X$19422 1729 VIA_via2_5
* cell instance $19423 r0 *1 36.575,65.45
X$19423 1729 VIA_via2_5
* cell instance $19424 r0 *1 36.575,66.43
X$19424 1729 VIA_via1_4
* cell instance $19425 r0 *1 38.285,65.45
X$19425 1729 VIA_via1_4
* cell instance $19426 r0 *1 38.285,65.45
X$19426 1729 VIA_via2_5
* cell instance $19427 r0 *1 39.805,66.43
X$19427 1729 VIA_via1_4
* cell instance $19428 r0 *1 38.665,85.61
X$19428 1730 VIA_via1_7
* cell instance $19429 r0 *1 38.665,85.61
X$19429 1730 VIA_via2_5
* cell instance $19430 r0 *1 38.665,86.59
X$19430 1730 VIA_via1_7
* cell instance $19431 r0 *1 38.665,86.59
X$19431 1730 VIA_via2_5
* cell instance $19432 r0 *1 40.755,81.83
X$19432 1730 VIA_via2_5
* cell instance $19433 r0 *1 38.095,85.61
X$19433 1730 VIA_via2_5
* cell instance $19434 r0 *1 38.095,81.83
X$19434 1730 VIA_via2_5
* cell instance $19435 r0 *1 40.565,86.59
X$19435 1730 VIA_via2_5
* cell instance $19436 r0 *1 38.285,86.59
X$19436 1730 VIA_via2_5
* cell instance $19437 r0 *1 37.905,90.51
X$19437 1730 VIA_via2_5
* cell instance $19438 r0 *1 40.945,71.47
X$19438 1730 VIA_via2_5
* cell instance $19439 r0 *1 41.135,66.57
X$19439 1730 VIA_via2_5
* cell instance $19440 r0 *1 40.375,71.47
X$19440 1730 VIA_via2_5
* cell instance $19441 r0 *1 39.995,71.47
X$19441 1730 VIA_via2_5
* cell instance $19442 r0 *1 40.755,80.43
X$19442 1730 VIA_via1_4
* cell instance $19443 r0 *1 37.145,81.97
X$19443 1730 VIA_via1_4
* cell instance $19444 r0 *1 37.145,81.83
X$19444 1730 VIA_via2_5
* cell instance $19445 r0 *1 38.285,88.83
X$19445 1730 VIA_via1_4
* cell instance $19446 r0 *1 40.565,87.57
X$19446 1730 VIA_via1_4
* cell instance $19447 r0 *1 40.565,87.71
X$19447 1730 VIA_via2_5
* cell instance $19448 r0 *1 42.275,87.57
X$19448 1730 VIA_via1_4
* cell instance $19449 r0 *1 42.275,87.71
X$19449 1730 VIA_via2_5
* cell instance $19450 r0 *1 36.385,90.37
X$19450 1730 VIA_via1_4
* cell instance $19451 r0 *1 36.385,90.51
X$19451 1730 VIA_via2_5
* cell instance $19452 r0 *1 41.515,69.23
X$19452 1730 VIA_via1_4
* cell instance $19453 r0 *1 39.995,70.77
X$19453 1730 VIA_via1_4
* cell instance $19454 r0 *1 38.475,66.43
X$19454 1730 VIA_via1_4
* cell instance $19455 r0 *1 38.475,66.57
X$19455 1730 VIA_via2_5
* cell instance $19456 r0 *1 37.145,66.43
X$19456 1730 VIA_via1_4
* cell instance $19457 r0 *1 37.145,66.57
X$19457 1730 VIA_via2_5
* cell instance $19458 r0 *1 41.515,66.43
X$19458 1731 VIA_via2_5
* cell instance $19459 r0 *1 39.235,66.43
X$19459 1731 VIA_via1_4
* cell instance $19460 r0 *1 39.235,66.43
X$19460 1731 VIA_via2_5
* cell instance $19461 r0 *1 41.515,65.45
X$19461 1731 VIA_via1_4
* cell instance $19462 r0 *1 37.905,66.43
X$19462 1731 VIA_via1_4
* cell instance $19463 r0 *1 37.905,66.43
X$19463 1731 VIA_via2_5
* cell instance $19464 r0 *1 39.615,67.27
X$19464 1732 VIA_via2_5
* cell instance $19465 r0 *1 40.375,67.27
X$19465 1732 VIA_via2_5
* cell instance $19466 r0 *1 40.185,66.85
X$19466 1732 VIA_via1_4
* cell instance $19467 r0 *1 39.615,67.97
X$19467 1732 VIA_via1_4
* cell instance $19468 r0 *1 46.455,66.85
X$19468 1733 VIA_via2_5
* cell instance $19469 r0 *1 41.705,66.85
X$19469 1733 VIA_via2_5
* cell instance $19470 r0 *1 41.705,67.97
X$19470 1733 VIA_via1_4
* cell instance $19471 r0 *1 45.315,66.85
X$19471 1733 VIA_via1_4
* cell instance $19472 r0 *1 45.315,66.85
X$19472 1733 VIA_via2_5
* cell instance $19473 r0 *1 46.455,66.43
X$19473 1733 VIA_via1_4
* cell instance $19474 r0 *1 51.205,66.15
X$19474 1734 VIA_via2_5
* cell instance $19475 r0 *1 48.165,66.15
X$19475 1734 VIA_via2_5
* cell instance $19476 r0 *1 51.205,66.43
X$19476 1734 VIA_via1_4
* cell instance $19477 r0 *1 50.825,66.15
X$19477 1734 VIA_via1_4
* cell instance $19478 r0 *1 50.825,66.15
X$19478 1734 VIA_via2_5
* cell instance $19479 r0 *1 48.165,65.17
X$19479 1734 VIA_via1_4
* cell instance $19480 r0 *1 53.105,66.29
X$19480 1735 VIA_via1_7
* cell instance $19481 r0 *1 57.475,67.27
X$19481 1735 VIA_via2_5
* cell instance $19482 r0 *1 57.475,69.23
X$19482 1735 VIA_via2_5
* cell instance $19483 r0 *1 51.395,65.17
X$19483 1735 VIA_via2_5
* cell instance $19484 r0 *1 51.015,65.17
X$19484 1735 VIA_via2_5
* cell instance $19485 r0 *1 53.105,67.27
X$19485 1735 VIA_via2_5
* cell instance $19486 r0 *1 50.825,70.77
X$19486 1735 VIA_via2_5
* cell instance $19487 r0 *1 51.015,72.03
X$19487 1735 VIA_via1_4
* cell instance $19488 r0 *1 53.105,65.17
X$19488 1735 VIA_via1_4
* cell instance $19489 r0 *1 53.105,65.17
X$19489 1735 VIA_via2_5
* cell instance $19490 r0 *1 51.015,62.37
X$19490 1735 VIA_via1_4
* cell instance $19491 r0 *1 51.015,67.97
X$19491 1735 VIA_via1_4
* cell instance $19492 r0 *1 49.495,70.77
X$19492 1735 VIA_via1_4
* cell instance $19493 r0 *1 49.495,70.77
X$19493 1735 VIA_via2_5
* cell instance $19494 r0 *1 56.335,69.23
X$19494 1735 VIA_via1_4
* cell instance $19495 r0 *1 56.335,69.23
X$19495 1735 VIA_via2_5
* cell instance $19496 r0 *1 57.475,67.97
X$19496 1735 VIA_via1_4
* cell instance $19497 r0 *1 57.285,62.37
X$19497 1735 VIA_via1_4
* cell instance $19498 r0 *1 54.625,67.41
X$19498 1736 VIA_via2_5
* cell instance $19499 r0 *1 53.865,67.41
X$19499 1736 VIA_via2_5
* cell instance $19500 r0 *1 54.625,66.43
X$19500 1736 VIA_via1_4
* cell instance $19501 r0 *1 53.865,67.97
X$19501 1736 VIA_via1_4
* cell instance $19502 r0 *1 55.385,65.31
X$19502 1736 VIA_via1_4
* cell instance $19503 r0 *1 56.905,66.01
X$19503 1737 VIA_via2_5
* cell instance $19504 r0 *1 58.425,66.01
X$19504 1737 VIA_via2_5
* cell instance $19505 r0 *1 58.995,66.01
X$19505 1737 VIA_via2_5
* cell instance $19506 r0 *1 58.425,65.17
X$19506 1737 VIA_via1_4
* cell instance $19507 r0 *1 58.995,67.55
X$19507 1737 VIA_via1_4
* cell instance $19508 r0 *1 56.905,66.43
X$19508 1737 VIA_via1_4
* cell instance $19509 r0 *1 61.465,66.71
X$19509 1738 VIA_via2_5
* cell instance $19510 r0 *1 63.365,66.71
X$19510 1738 VIA_via2_5
* cell instance $19511 r0 *1 61.465,67.97
X$19511 1738 VIA_via1_4
* cell instance $19512 r0 *1 62.985,66.71
X$19512 1738 VIA_via1_4
* cell instance $19513 r0 *1 62.985,66.71
X$19513 1738 VIA_via2_5
* cell instance $19514 r0 *1 63.365,66.43
X$19514 1738 VIA_via1_4
* cell instance $19515 r0 *1 63.555,65.45
X$19515 1739 VIA_via2_5
* cell instance $19516 r0 *1 63.935,65.45
X$19516 1739 VIA_via2_5
* cell instance $19517 r0 *1 63.935,66.43
X$19517 1739 VIA_via1_4
* cell instance $19518 r0 *1 63.175,65.45
X$19518 1739 VIA_via1_4
* cell instance $19519 r0 *1 63.555,65.17
X$19519 1739 VIA_via1_4
* cell instance $19520 r0 *1 85.785,66.43
X$19520 1740 VIA_via1_4
* cell instance $19521 r0 *1 85.215,67.97
X$19521 1740 VIA_via1_4
* cell instance $19522 r0 *1 85.025,66.85
X$19522 1740 VIA_via1_4
* cell instance $19523 r0 *1 86.545,67.97
X$19523 1741 VIA_via1_4
* cell instance $19524 r0 *1 88.065,68.95
X$19524 1741 VIA_via1_4
* cell instance $19525 r0 *1 87.685,66.43
X$19525 1741 VIA_via1_4
* cell instance $19526 r0 *1 94.715,66.29
X$19526 1742 VIA_via2_5
* cell instance $19527 r0 *1 92.435,67.97
X$19527 1742 VIA_via2_5
* cell instance $19528 r0 *1 93.005,67.97
X$19528 1742 VIA_via2_5
* cell instance $19529 r0 *1 91.865,67.97
X$19529 1742 VIA_via1_4
* cell instance $19530 r0 *1 91.865,67.97
X$19530 1742 VIA_via2_5
* cell instance $19531 r0 *1 93.005,68.95
X$19531 1742 VIA_via1_4
* cell instance $19532 r0 *1 94.715,65.17
X$19532 1742 VIA_via1_4
* cell instance $19533 r0 *1 92.435,66.43
X$19533 1742 VIA_via1_4
* cell instance $19534 r0 *1 92.435,66.29
X$19534 1742 VIA_via2_5
* cell instance $19535 r0 *1 31.255,75.39
X$19535 1743 VIA_via2_5
* cell instance $19536 r0 *1 55.765,71.05
X$19536 1743 VIA_via2_5
* cell instance $19537 r0 *1 54.815,71.05
X$19537 1743 VIA_via2_5
* cell instance $19538 r0 *1 55.575,75.53
X$19538 1743 VIA_via2_5
* cell instance $19539 r0 *1 53.295,76.65
X$19539 1743 VIA_via2_5
* cell instance $19540 r0 *1 54.245,75.53
X$19540 1743 VIA_via2_5
* cell instance $19541 r0 *1 54.245,76.37
X$19541 1743 VIA_via2_5
* cell instance $19542 r0 *1 36.955,75.67
X$19542 1743 VIA_via2_5
* cell instance $19543 r0 *1 90.345,68.67
X$19543 1743 VIA_via2_5
* cell instance $19544 r0 *1 92.815,68.67
X$19544 1743 VIA_via2_5
* cell instance $19545 r0 *1 78.185,68.53
X$19545 1743 VIA_via2_5
* cell instance $19546 r0 *1 77.995,70.91
X$19546 1743 VIA_via2_5
* cell instance $19547 r0 *1 55.575,74.83
X$19547 1743 VIA_via1_4
* cell instance $19548 r0 *1 54.815,70.77
X$19548 1743 VIA_via1_4
* cell instance $19549 r0 *1 53.485,77.63
X$19549 1743 VIA_via1_4
* cell instance $19550 r0 *1 42.275,76.37
X$19550 1743 VIA_via1_4
* cell instance $19551 r0 *1 42.275,76.51
X$19551 1743 VIA_via2_5
* cell instance $19552 r0 *1 36.955,76.37
X$19552 1743 VIA_via1_4
* cell instance $19553 r0 *1 36.955,76.37
X$19553 1743 VIA_via2_5
* cell instance $19554 r0 *1 37.055,76.37
X$19554 1743 VIA_via3_2
* cell instance $19555 r0 *1 37.055,76.51
X$19555 1743 VIA_via4_0
* cell instance $19556 r0 *1 31.255,74.83
X$19556 1743 VIA_via1_4
* cell instance $19557 r0 *1 30.685,79.17
X$19557 1743 VIA_via1_4
* cell instance $19558 r0 *1 90.345,67.97
X$19558 1743 VIA_via1_4
* cell instance $19559 r0 *1 91.105,73.15
X$19559 1743 VIA_via1_4
* cell instance $19560 r0 *1 93.005,66.43
X$19560 1743 VIA_via1_4
* cell instance $19561 r0 *1 77.805,67.97
X$19561 1743 VIA_via1_4
* cell instance $19562 r0 *1 42.095,76.51
X$19562 1743 VIA_via3_2
* cell instance $19563 r0 *1 42.095,76.51
X$19563 1743 VIA_via4_0
* cell instance $19564 r0 *1 94.335,65.31
X$19564 1744 VIA_via1_4
* cell instance $19565 r0 *1 93.955,66.43
X$19565 1744 VIA_via1_4
* cell instance $19566 r0 *1 95.665,66.57
X$19566 1745 VIA_via2_5
* cell instance $19567 r0 *1 96.045,66.57
X$19567 1745 VIA_via2_5
* cell instance $19568 r0 *1 96.045,67.55
X$19568 1745 VIA_via1_4
* cell instance $19569 r0 *1 94.525,66.43
X$19569 1745 VIA_via1_4
* cell instance $19570 r0 *1 94.525,66.57
X$19570 1745 VIA_via2_5
* cell instance $19571 r0 *1 94.145,65.17
X$19571 1745 VIA_via1_4
* cell instance $19572 r0 *1 94.145,65.17
X$19572 1745 VIA_via2_5
* cell instance $19573 r0 *1 95.665,65.17
X$19573 1745 VIA_via1_4
* cell instance $19574 r0 *1 95.665,65.17
X$19574 1745 VIA_via2_5
* cell instance $19575 r0 *1 7.315,65.17
X$19575 1746 VIA_via1_4
* cell instance $19576 r0 *1 7.315,65.17
X$19576 1746 VIA_via2_5
* cell instance $19577 r0 *1 5.795,66.15
X$19577 1746 VIA_via1_4
* cell instance $19578 r0 *1 5.795,65.17
X$19578 1746 VIA_via1_4
* cell instance $19579 r0 *1 5.795,65.17
X$19579 1746 VIA_via2_5
* cell instance $19580 r0 *1 11.875,67.41
X$19580 1747 VIA_via1_7
* cell instance $19581 r0 *1 11.875,66.71
X$19581 1747 VIA_via2_5
* cell instance $19582 r0 *1 7.885,66.71
X$19582 1747 VIA_via2_5
* cell instance $19583 r0 *1 7.885,66.43
X$19583 1747 VIA_via1_4
* cell instance $19584 r0 *1 93.195,66.43
X$19584 1748 VIA_via1_4
* cell instance $19585 r0 *1 93.195,66.43
X$19585 1748 VIA_via2_5
* cell instance $19586 r0 *1 94.335,66.43
X$19586 1748 VIA_via1_4
* cell instance $19587 r0 *1 94.335,66.43
X$19587 1748 VIA_via2_5
* cell instance $19588 r0 *1 13.775,66.01
X$19588 1749 VIA_via1_7
* cell instance $19589 r0 *1 13.775,65.87
X$19589 1749 VIA_via2_5
* cell instance $19590 r0 *1 11.305,65.87
X$19590 1749 VIA_via2_5
* cell instance $19591 r0 *1 11.305,65.17
X$19591 1749 VIA_via1_4
* cell instance $19592 r0 *1 88.255,67.83
X$19592 1750 VIA_via2_5
* cell instance $19593 r0 *1 87.875,67.97
X$19593 1750 VIA_via1_4
* cell instance $19594 r0 *1 87.875,67.83
X$19594 1750 VIA_via2_5
* cell instance $19595 r0 *1 88.255,66.43
X$19595 1750 VIA_via1_4
* cell instance $19596 r0 *1 88.255,66.43
X$19596 1750 VIA_via2_5
* cell instance $19597 r0 *1 91.865,66.43
X$19597 1750 VIA_via1_4
* cell instance $19598 r0 *1 91.865,66.43
X$19598 1750 VIA_via2_5
* cell instance $19599 r0 *1 86.735,66.43
X$19599 1751 VIA_via1_4
* cell instance $19600 r0 *1 86.735,66.43
X$19600 1751 VIA_via2_5
* cell instance $19601 r0 *1 82.745,66.43
X$19601 1751 VIA_via1_4
* cell instance $19602 r0 *1 82.745,66.43
X$19602 1751 VIA_via2_5
* cell instance $19603 r0 *1 28.595,66.01
X$19603 1752 VIA_via1_7
* cell instance $19604 r0 *1 28.595,65.17
X$19604 1752 VIA_via2_5
* cell instance $19605 r0 *1 26.315,65.17
X$19605 1752 VIA_via1_4
* cell instance $19606 r0 *1 26.315,65.17
X$19606 1752 VIA_via2_5
* cell instance $19607 r0 *1 79.895,64.19
X$19607 1753 VIA_via1_7
* cell instance $19608 r0 *1 79.895,65.17
X$19608 1753 VIA_via2_5
* cell instance $19609 r0 *1 78.945,65.17
X$19609 1753 VIA_via1_4
* cell instance $19610 r0 *1 78.945,65.17
X$19610 1753 VIA_via2_5
* cell instance $19611 r0 *1 32.205,66.43
X$19611 1754 VIA_via1_4
* cell instance $19612 r0 *1 32.015,66.43
X$19612 1754 VIA_via1_4
* cell instance $19613 r0 *1 79.325,67.69
X$19613 1755 VIA_via2_5
* cell instance $19614 r0 *1 77.615,67.83
X$19614 1755 VIA_via2_5
* cell instance $19615 r0 *1 77.615,68.11
X$19615 1755 VIA_via2_5
* cell instance $19616 r0 *1 79.325,66.15
X$19616 1755 VIA_via2_5
* cell instance $19617 r0 *1 64.125,67.97
X$19617 1755 VIA_via1_4
* cell instance $19618 r0 *1 64.125,68.11
X$19618 1755 VIA_via2_5
* cell instance $19619 r0 *1 79.705,67.97
X$19619 1755 VIA_via1_4
* cell instance $19620 r0 *1 79.705,67.83
X$19620 1755 VIA_via2_5
* cell instance $19621 r0 *1 80.085,67.97
X$19621 1755 VIA_via1_4
* cell instance $19622 r0 *1 79.705,66.15
X$19622 1755 VIA_via1_4
* cell instance $19623 r0 *1 79.705,66.15
X$19623 1755 VIA_via2_5
* cell instance $19624 r0 *1 78.185,67.69
X$19624 1756 VIA_via1_7
* cell instance $19625 r0 *1 77.425,66.71
X$19625 1756 VIA_via2_5
* cell instance $19626 r0 *1 78.185,66.71
X$19626 1756 VIA_via2_5
* cell instance $19627 r0 *1 77.425,66.43
X$19627 1756 VIA_via1_4
* cell instance $19628 r0 *1 32.965,66.43
X$19628 1757 VIA_via1_4
* cell instance $19629 r0 *1 32.965,66.43
X$19629 1757 VIA_via2_5
* cell instance $19630 r0 *1 33.725,66.43
X$19630 1757 VIA_via1_4
* cell instance $19631 r0 *1 33.725,66.43
X$19631 1757 VIA_via2_5
* cell instance $19632 r0 *1 37.525,66.01
X$19632 1758 VIA_via1_7
* cell instance $19633 r0 *1 37.525,65.17
X$19633 1758 VIA_via2_5
* cell instance $19634 r0 *1 36.005,65.17
X$19634 1758 VIA_via1_4
* cell instance $19635 r0 *1 36.005,65.17
X$19635 1758 VIA_via2_5
* cell instance $19636 r0 *1 66.785,65.45
X$19636 1759 VIA_via2_5
* cell instance $19637 r0 *1 68.115,65.45
X$19637 1759 VIA_via2_5
* cell instance $19638 r0 *1 66.785,66.43
X$19638 1759 VIA_via1_4
* cell instance $19639 r0 *1 68.115,65.03
X$19639 1759 VIA_via1_4
* cell instance $19640 r0 *1 53.485,64.19
X$19640 1760 VIA_via1_7
* cell instance $19641 r0 *1 53.485,65.31
X$19641 1760 VIA_via2_5
* cell instance $19642 r0 *1 52.345,65.17
X$19642 1760 VIA_via1_4
* cell instance $19643 r0 *1 52.345,65.31
X$19643 1760 VIA_via2_5
* cell instance $19644 r0 *1 54.055,64.19
X$19644 1761 VIA_via1_7
* cell instance $19645 r0 *1 54.055,65.17
X$19645 1761 VIA_via2_5
* cell instance $19646 r0 *1 55.195,65.17
X$19646 1761 VIA_via1_4
* cell instance $19647 r0 *1 55.195,65.17
X$19647 1761 VIA_via2_5
* cell instance $19648 r0 *1 12.825,66.99
X$19648 1762 VIA_via2_5
* cell instance $19649 r0 *1 12.825,65.17
X$19649 1762 VIA_via1_4
* cell instance $19650 r0 *1 13.395,66.85
X$19650 1762 VIA_via1_4
* cell instance $19651 r0 *1 13.395,66.99
X$19651 1762 VIA_via2_5
* cell instance $19652 r0 *1 12.825,67.97
X$19652 1762 VIA_via1_4
* cell instance $19653 r0 *1 27.075,66.99
X$19653 1763 VIA_via1_7
* cell instance $19654 r0 *1 26.695,67.97
X$19654 1763 VIA_via1_4
* cell instance $19655 r0 *1 26.125,67.55
X$19655 1764 VIA_via2_5
* cell instance $19656 r0 *1 29.925,67.55
X$19656 1764 VIA_via2_5
* cell instance $19657 r0 *1 26.125,66.43
X$19657 1764 VIA_via1_4
* cell instance $19658 r0 *1 28.975,67.55
X$19658 1764 VIA_via1_4
* cell instance $19659 r0 *1 28.975,67.55
X$19659 1764 VIA_via2_5
* cell instance $19660 r0 *1 29.925,67.97
X$19660 1764 VIA_via1_4
* cell instance $19661 r0 *1 46.265,68.95
X$19661 1765 VIA_via1_7
* cell instance $19662 r0 *1 46.265,68.81
X$19662 1765 VIA_via2_5
* cell instance $19663 r0 *1 51.015,69.79
X$19663 1765 VIA_via1_7
* cell instance $19664 r0 *1 51.015,69.79
X$19664 1765 VIA_via2_5
* cell instance $19665 r0 *1 53.865,69.79
X$19665 1765 VIA_via2_5
* cell instance $19666 r0 *1 32.965,68.81
X$19666 1765 VIA_via2_5
* cell instance $19667 r0 *1 32.855,68.81
X$19667 1765 VIA_via3_2
* cell instance $19668 r0 *1 64.505,69.37
X$19668 1765 VIA_via1_4
* cell instance $19669 r0 *1 64.505,69.51
X$19669 1765 VIA_via2_5
* cell instance $19670 r0 *1 53.865,70.63
X$19670 1765 VIA_via1_4
* cell instance $19671 r0 *1 32.775,79.03
X$19671 1765 VIA_via1_4
* cell instance $19672 r0 *1 32.775,74.83
X$19672 1765 VIA_via1_4
* cell instance $19673 r0 *1 32.775,74.69
X$19673 1765 VIA_via2_5
* cell instance $19674 r0 *1 32.855,74.69
X$19674 1765 VIA_via3_2
* cell instance $19675 r0 *1 33.155,66.57
X$19675 1765 VIA_via1_4
* cell instance $19676 r0 *1 42.655,67.41
X$19676 1766 VIA_via1_7
* cell instance $19677 r0 *1 43.035,66.43
X$19677 1766 VIA_via1_4
* cell instance $19678 r0 *1 56.525,84.21
X$19678 1767 VIA_via1_7
* cell instance $19679 r0 *1 56.525,84.21
X$19679 1767 VIA_via2_5
* cell instance $19680 r0 *1 48.355,84.21
X$19680 1767 VIA_via2_5
* cell instance $19681 r0 *1 51.965,72.03
X$19681 1767 VIA_via2_5
* cell instance $19682 r0 *1 52.535,84.21
X$19682 1767 VIA_via2_5
* cell instance $19683 r0 *1 49.495,84.21
X$19683 1767 VIA_via2_5
* cell instance $19684 r0 *1 52.155,77.21
X$19684 1767 VIA_via2_5
* cell instance $19685 r0 *1 50.825,84.21
X$19685 1767 VIA_via2_5
* cell instance $19686 r0 *1 57.095,78.05
X$19686 1767 VIA_via2_5
* cell instance $19687 r0 *1 51.395,78.05
X$19687 1767 VIA_via2_5
* cell instance $19688 r0 *1 51.395,77.21
X$19688 1767 VIA_via2_5
* cell instance $19689 r0 *1 57.095,76.37
X$19689 1767 VIA_via1_4
* cell instance $19690 r0 *1 52.345,70.77
X$19690 1767 VIA_via1_4
* cell instance $19691 r0 *1 49.495,86.03
X$19691 1767 VIA_via1_4
* cell instance $19692 r0 *1 50.825,84.77
X$19692 1767 VIA_via1_4
* cell instance $19693 r0 *1 52.535,83.23
X$19693 1767 VIA_via1_4
* cell instance $19694 r0 *1 51.585,80.43
X$19694 1767 VIA_via1_4
* cell instance $19695 r0 *1 48.355,84.77
X$19695 1767 VIA_via1_4
* cell instance $19696 r0 *1 48.925,67.97
X$19696 1767 VIA_via1_4
* cell instance $19697 r0 *1 48.925,72.03
X$19697 1767 VIA_via1_4
* cell instance $19698 r0 *1 48.925,72.03
X$19698 1767 VIA_via2_5
* cell instance $19699 r0 *1 48.735,65.17
X$19699 1767 VIA_via1_4
* cell instance $19700 r0 *1 57.285,66.99
X$19700 1768 VIA_via1_7
* cell instance $19701 r0 *1 56.715,67.97
X$19701 1768 VIA_via1_4
* cell instance $19702 r0 *1 64.315,66.99
X$19702 1769 VIA_via1_7
* cell instance $19703 r0 *1 64.695,67.97
X$19703 1769 VIA_via1_4
* cell instance $19704 r0 *1 86.735,70.21
X$19704 1770 VIA_via1_7
* cell instance $19705 r0 *1 72.675,67.27
X$19705 1770 VIA_via2_5
* cell instance $19706 r0 *1 79.895,72.17
X$19706 1770 VIA_via2_5
* cell instance $19707 r0 *1 83.125,68.81
X$19707 1770 VIA_via2_5
* cell instance $19708 r0 *1 88.445,68.67
X$19708 1770 VIA_via2_5
* cell instance $19709 r0 *1 86.735,69.23
X$19709 1770 VIA_via2_5
* cell instance $19710 r0 *1 87.115,68.67
X$19710 1770 VIA_via2_5
* cell instance $19711 r0 *1 86.355,67.41
X$19711 1770 VIA_via2_5
* cell instance $19712 r0 *1 87.115,67.41
X$19712 1770 VIA_via2_5
* cell instance $19713 r0 *1 74.575,67.27
X$19713 1770 VIA_via2_5
* cell instance $19714 r0 *1 76.475,71.47
X$19714 1770 VIA_via2_5
* cell instance $19715 r0 *1 79.895,68.81
X$19715 1770 VIA_via2_5
* cell instance $19716 r0 *1 75.715,71.47
X$19716 1770 VIA_via2_5
* cell instance $19717 r0 *1 75.145,67.27
X$19717 1770 VIA_via2_5
* cell instance $19718 r0 *1 72.675,67.97
X$19718 1770 VIA_via1_4
* cell instance $19719 r0 *1 76.285,73.57
X$19719 1770 VIA_via1_4
* cell instance $19720 r0 *1 88.445,67.97
X$19720 1770 VIA_via1_4
* cell instance $19721 r0 *1 87.115,67.97
X$19721 1770 VIA_via1_4
* cell instance $19722 r0 *1 86.355,66.43
X$19722 1770 VIA_via1_4
* cell instance $19723 r0 *1 76.475,72.03
X$19723 1770 VIA_via1_4
* cell instance $19724 r0 *1 76.475,72.17
X$19724 1770 VIA_via2_5
* cell instance $19725 r0 *1 77.995,72.03
X$19725 1770 VIA_via1_4
* cell instance $19726 r0 *1 77.995,72.17
X$19726 1770 VIA_via2_5
* cell instance $19727 r0 *1 74.575,66.43
X$19727 1770 VIA_via1_4
* cell instance $19728 r0 *1 83.125,67.97
X$19728 1770 VIA_via1_4
* cell instance $19729 r0 *1 79.895,70.77
X$19729 1770 VIA_via1_4
* cell instance $19730 r0 *1 74.955,66.99
X$19730 1771 VIA_via1_7
* cell instance $19731 r0 *1 74.575,67.97
X$19731 1771 VIA_via1_4
* cell instance $19732 r0 *1 69.065,67.69
X$19732 1772 VIA_via1_4
* cell instance $19733 r0 *1 69.065,67.69
X$19733 1772 VIA_via2_5
* cell instance $19734 r0 *1 78.185,67.97
X$19734 1772 VIA_via1_4
* cell instance $19735 r0 *1 78.185,67.97
X$19735 1772 VIA_via2_5
* cell instance $19736 r0 *1 85.595,67.41
X$19736 1773 VIA_via1_7
* cell instance $19737 r0 *1 85.975,65.17
X$19737 1773 VIA_via1_4
* cell instance $19738 r0 *1 88.825,67.41
X$19738 1774 VIA_via1_7
* cell instance $19739 r0 *1 89.585,66.43
X$19739 1774 VIA_via1_4
* cell instance $19740 r0 *1 93.765,67.97
X$19740 1775 VIA_via1_4
* cell instance $19741 r0 *1 93.765,66.71
X$19741 1775 VIA_via1_4
* cell instance $19742 r0 *1 91.295,67.97
X$19742 1776 VIA_via1_4
* cell instance $19743 r0 *1 91.295,67.83
X$19743 1776 VIA_via2_5
* cell instance $19744 r0 *1 92.055,67.83
X$19744 1776 VIA_via1_4
* cell instance $19745 r0 *1 92.055,67.83
X$19745 1776 VIA_via2_5
* cell instance $19746 r0 *1 92.245,66.99
X$19746 1777 VIA_via1_7
* cell instance $19747 r0 *1 92.245,66.99
X$19747 1777 VIA_via2_5
* cell instance $19748 r0 *1 90.535,66.99
X$19748 1777 VIA_via2_5
* cell instance $19749 r0 *1 90.535,67.97
X$19749 1777 VIA_via1_4
* cell instance $19750 r0 *1 10.925,68.81
X$19750 1778 VIA_via1_7
* cell instance $19751 r0 *1 11.115,67.13
X$19751 1778 VIA_via2_5
* cell instance $19752 r0 *1 11.495,67.13
X$19752 1778 VIA_via2_5
* cell instance $19753 r0 *1 11.495,65.17
X$19753 1778 VIA_via1_4
* cell instance $19754 r0 *1 13.775,67.41
X$19754 1779 VIA_via1_7
* cell instance $19755 r0 *1 11.115,66.85
X$19755 1779 VIA_via2_5
* cell instance $19756 r0 *1 13.775,66.85
X$19756 1779 VIA_via2_5
* cell instance $19757 r0 *1 11.115,66.43
X$19757 1779 VIA_via1_4
* cell instance $19758 r0 *1 21.185,66.99
X$19758 1780 VIA_via1_7
* cell instance $19759 r0 *1 21.185,67.97
X$19759 1780 VIA_via1_4
* cell instance $19760 r0 *1 20.995,67.41
X$19760 1781 VIA_via1_7
* cell instance $19761 r0 *1 20.995,67.41
X$19761 1781 VIA_via2_5
* cell instance $19762 r0 *1 22.135,67.41
X$19762 1781 VIA_via2_5
* cell instance $19763 r0 *1 22.135,66.43
X$19763 1781 VIA_via1_4
* cell instance $19764 r0 *1 47.025,67.83
X$19764 1782 VIA_via2_5
* cell instance $19765 r0 *1 47.215,67.83
X$19765 1782 VIA_via1_4
* cell instance $19766 r0 *1 47.215,67.83
X$19766 1782 VIA_via2_5
* cell instance $19767 r0 *1 43.035,67.97
X$19767 1782 VIA_via1_4
* cell instance $19768 r0 *1 43.035,67.83
X$19768 1782 VIA_via2_5
* cell instance $19769 r0 *1 47.025,66.43
X$19769 1782 VIA_via1_4
* cell instance $19770 r0 *1 43.985,67.97
X$19770 1783 VIA_via1_4
* cell instance $19771 r0 *1 43.985,67.97
X$19771 1783 VIA_via2_5
* cell instance $19772 r0 *1 44.935,67.97
X$19772 1783 VIA_via1_4
* cell instance $19773 r0 *1 44.935,67.97
X$19773 1783 VIA_via2_5
* cell instance $19774 r0 *1 51.775,67.97
X$19774 1784 VIA_via2_5
* cell instance $19775 r0 *1 51.775,66.43
X$19775 1784 VIA_via1_4
* cell instance $19776 r0 *1 52.535,67.97
X$19776 1784 VIA_via1_4
* cell instance $19777 r0 *1 52.535,67.97
X$19777 1784 VIA_via2_5
* cell instance $19778 r0 *1 48.355,67.97
X$19778 1784 VIA_via1_4
* cell instance $19779 r0 *1 48.355,67.97
X$19779 1784 VIA_via2_5
* cell instance $19780 r0 *1 66.975,68.95
X$19780 1785 VIA_via1_4
* cell instance $19781 r0 *1 68.115,67.97
X$19781 1785 VIA_via1_4
* cell instance $19782 r0 *1 68.115,67.97
X$19782 1785 VIA_via2_5
* cell instance $19783 r0 *1 66.975,67.97
X$19783 1785 VIA_via1_4
* cell instance $19784 r0 *1 66.975,67.97
X$19784 1785 VIA_via2_5
* cell instance $19785 r0 *1 52.155,66.99
X$19785 1786 VIA_via1_7
* cell instance $19786 r0 *1 52.155,67.69
X$19786 1786 VIA_via2_5
* cell instance $19787 r0 *1 52.915,67.69
X$19787 1786 VIA_via2_5
* cell instance $19788 r0 *1 52.915,70.77
X$19788 1786 VIA_via1_4
* cell instance $19789 r0 *1 60.135,74.41
X$19789 1787 VIA_via1_7
* cell instance $19790 r0 *1 60.135,74.27
X$19790 1787 VIA_via2_5
* cell instance $19791 r0 *1 31.445,73.71
X$19791 1787 VIA_via2_5
* cell instance $19792 r0 *1 30.115,76.93
X$19792 1787 VIA_via2_5
* cell instance $19793 r0 *1 37.145,77.07
X$19793 1787 VIA_via2_5
* cell instance $19794 r0 *1 42.275,77.07
X$19794 1787 VIA_via2_5
* cell instance $19795 r0 *1 60.135,73.57
X$19795 1787 VIA_via2_5
* cell instance $19796 r0 *1 56.145,77.07
X$19796 1787 VIA_via2_5
* cell instance $19797 r0 *1 51.585,77.07
X$19797 1787 VIA_via2_5
* cell instance $19798 r0 *1 67.545,74.27
X$19798 1787 VIA_via2_5
* cell instance $19799 r0 *1 51.585,77.63
X$19799 1787 VIA_via1_4
* cell instance $19800 r0 *1 56.145,77.63
X$19800 1787 VIA_via1_4
* cell instance $19801 r0 *1 67.545,67.97
X$19801 1787 VIA_via1_4
* cell instance $19802 r0 *1 54.625,67.97
X$19802 1787 VIA_via1_4
* cell instance $19803 r0 *1 54.625,67.97
X$19803 1787 VIA_via2_5
* cell instance $19804 r0 *1 54.695,67.97
X$19804 1787 VIA_via3_2
* cell instance $19805 r0 *1 42.275,77.63
X$19805 1787 VIA_via1_4
* cell instance $19806 r0 *1 37.145,77.63
X$19806 1787 VIA_via1_4
* cell instance $19807 r0 *1 30.305,77.63
X$19807 1787 VIA_via1_4
* cell instance $19808 r0 *1 30.115,76.37
X$19808 1787 VIA_via1_4
* cell instance $19809 r0 *1 31.635,66.43
X$19809 1787 VIA_via1_4
* cell instance $19810 r0 *1 30.115,73.57
X$19810 1787 VIA_via1_4
* cell instance $19811 r0 *1 30.115,73.71
X$19811 1787 VIA_via2_5
* cell instance $19812 r0 *1 55.255,73.57
X$19812 1787 VIA_via3_2
* cell instance $19813 r0 *1 54.695,73.57
X$19813 1787 VIA_via3_2
* cell instance $19814 r0 *1 55.255,77.07
X$19814 1787 VIA_via3_2
* cell instance $19815 r0 *1 62.415,67.41
X$19815 1788 VIA_via1_7
* cell instance $19816 r0 *1 62.415,67.41
X$19816 1788 VIA_via2_5
* cell instance $19817 r0 *1 60.705,67.41
X$19817 1788 VIA_via2_5
* cell instance $19818 r0 *1 60.705,66.43
X$19818 1788 VIA_via1_4
* cell instance $19819 r0 *1 5.415,69.23
X$19819 1789 VIA_via1_4
* cell instance $19820 r0 *1 5.985,70.77
X$19820 1789 VIA_via1_4
* cell instance $19821 r0 *1 5.035,68.95
X$19821 1789 VIA_via1_4
* cell instance $19822 r0 *1 10.355,69.23
X$19822 1790 VIA_via2_5
* cell instance $19823 r0 *1 10.355,68.25
X$19823 1790 VIA_via1_4
* cell instance $19824 r0 *1 9.215,69.23
X$19824 1790 VIA_via1_4
* cell instance $19825 r0 *1 9.215,69.23
X$19825 1790 VIA_via2_5
* cell instance $19826 r0 *1 7.885,69.23
X$19826 1790 VIA_via1_4
* cell instance $19827 r0 *1 7.885,69.23
X$19827 1790 VIA_via2_5
* cell instance $19828 r0 *1 10.735,76.51
X$19828 1791 VIA_via2_5
* cell instance $19829 r0 *1 16.815,68.39
X$19829 1791 VIA_via2_5
* cell instance $19830 r0 *1 7.885,76.09
X$19830 1791 VIA_via2_5
* cell instance $19831 r0 *1 16.815,76.51
X$19831 1791 VIA_via2_5
* cell instance $19832 r0 *1 18.905,68.39
X$19832 1791 VIA_via2_5
* cell instance $19833 r0 *1 10.735,76.09
X$19833 1791 VIA_via2_5
* cell instance $19834 r0 *1 20.615,68.39
X$19834 1791 VIA_via2_5
* cell instance $19835 r0 *1 10.735,72.73
X$19835 1791 VIA_via2_5
* cell instance $19836 r0 *1 7.885,69.79
X$19836 1791 VIA_via2_5
* cell instance $19837 r0 *1 5.985,69.79
X$19837 1791 VIA_via2_5
* cell instance $19838 r0 *1 11.495,72.73
X$19838 1791 VIA_via2_5
* cell instance $19839 r0 *1 18.905,66.43
X$19839 1791 VIA_via1_4
* cell instance $19840 r0 *1 20.615,67.97
X$19840 1791 VIA_via1_4
* cell instance $19841 r0 *1 16.815,69.23
X$19841 1791 VIA_via1_4
* cell instance $19842 r0 *1 7.885,70.77
X$19842 1791 VIA_via1_4
* cell instance $19843 r0 *1 5.985,69.23
X$19843 1791 VIA_via1_4
* cell instance $19844 r0 *1 11.495,72.03
X$19844 1791 VIA_via1_4
* cell instance $19845 r0 *1 16.815,77.63
X$19845 1791 VIA_via1_4
* cell instance $19846 r0 *1 10.735,74.83
X$19846 1791 VIA_via1_4
* cell instance $19847 r0 *1 7.885,76.37
X$19847 1791 VIA_via1_4
* cell instance $19848 r0 *1 11.875,76.37
X$19848 1791 VIA_via1_4
* cell instance $19849 r0 *1 11.875,76.51
X$19849 1791 VIA_via2_5
* cell instance $19850 r0 *1 16.815,73.57
X$19850 1791 VIA_via1_4
* cell instance $19851 r0 *1 19.095,70.21
X$19851 1792 VIA_via1_7
* cell instance $19852 r0 *1 18.905,69.23
X$19852 1792 VIA_via1_4
* cell instance $19853 r0 *1 21.375,68.39
X$19853 1793 VIA_via1_7
* cell instance $19854 r0 *1 21.375,73.71
X$19854 1793 VIA_via2_5
* cell instance $19855 r0 *1 20.045,73.57
X$19855 1793 VIA_via1_4
* cell instance $19856 r0 *1 20.045,73.71
X$19856 1793 VIA_via2_5
* cell instance $19857 r0 *1 25.365,69.23
X$19857 1794 VIA_via2_5
* cell instance $19858 r0 *1 30.115,69.23
X$19858 1794 VIA_via1_4
* cell instance $19859 r0 *1 30.115,69.23
X$19859 1794 VIA_via2_5
* cell instance $19860 r0 *1 25.935,69.23
X$19860 1794 VIA_via1_4
* cell instance $19861 r0 *1 25.935,69.23
X$19861 1794 VIA_via2_5
* cell instance $19862 r0 *1 25.365,72.03
X$19862 1794 VIA_via1_4
* cell instance $19863 r0 *1 34.485,72.03
X$19863 1795 VIA_via2_5
* cell instance $19864 r0 *1 34.675,69.23
X$19864 1795 VIA_via2_5
* cell instance $19865 r0 *1 36.765,69.23
X$19865 1795 VIA_via2_5
* cell instance $19866 r0 *1 32.395,72.03
X$19866 1795 VIA_via2_5
* cell instance $19867 r0 *1 32.395,76.37
X$19867 1795 VIA_via1_4
* cell instance $19868 r0 *1 32.395,77.63
X$19868 1795 VIA_via1_4
* cell instance $19869 r0 *1 30.495,72.03
X$19869 1795 VIA_via1_4
* cell instance $19870 r0 *1 30.495,72.03
X$19870 1795 VIA_via2_5
* cell instance $19871 r0 *1 36.765,65.17
X$19871 1795 VIA_via1_4
* cell instance $19872 r0 *1 35.055,69.23
X$19872 1795 VIA_via1_4
* cell instance $19873 r0 *1 35.055,69.23
X$19873 1795 VIA_via2_5
* cell instance $19874 r0 *1 32.775,72.03
X$19874 1795 VIA_via1_4
* cell instance $19875 r0 *1 32.775,72.03
X$19875 1795 VIA_via2_5
* cell instance $19876 r0 *1 34.675,72.03
X$19876 1795 VIA_via1_4
* cell instance $19877 r0 *1 34.675,72.03
X$19877 1795 VIA_via2_5
* cell instance $19878 r0 *1 34.485,73.15
X$19878 1795 VIA_via1_4
* cell instance $19879 r0 *1 39.805,68.39
X$19879 1796 VIA_via1_7
* cell instance $19880 r0 *1 40.185,76.37
X$19880 1796 VIA_via1_4
* cell instance $19881 r0 *1 56.525,69.09
X$19881 1797 VIA_via2_5
* cell instance $19882 r0 *1 54.625,69.23
X$19882 1797 VIA_via1_4
* cell instance $19883 r0 *1 54.625,69.09
X$19883 1797 VIA_via2_5
* cell instance $19884 r0 *1 55.955,70.77
X$19884 1797 VIA_via1_4
* cell instance $19885 r0 *1 56.525,70.77
X$19885 1797 VIA_via1_4
* cell instance $19886 r0 *1 57.855,69.09
X$19886 1797 VIA_via1_4
* cell instance $19887 r0 *1 57.855,69.09
X$19887 1797 VIA_via2_5
* cell instance $19888 r0 *1 64.505,68.39
X$19888 1798 VIA_via1_7
* cell instance $19889 r0 *1 64.885,69.23
X$19889 1798 VIA_via1_4
* cell instance $19890 r0 *1 69.825,68.39
X$19890 1799 VIA_via1_7
* cell instance $19891 r0 *1 69.825,68.39
X$19891 1799 VIA_via2_5
* cell instance $19892 r0 *1 67.165,68.39
X$19892 1799 VIA_via2_5
* cell instance $19893 r0 *1 66.975,69.23
X$19893 1799 VIA_via1_4
* cell instance $19894 r0 *1 69.825,71.61
X$19894 1800 VIA_via1_7
* cell instance $19895 r0 *1 69.635,67.97
X$19895 1800 VIA_via1_4
* cell instance $19896 r0 *1 72.105,68.95
X$19896 1801 VIA_via2_5
* cell instance $19897 r0 *1 74.385,68.95
X$19897 1801 VIA_via2_5
* cell instance $19898 r0 *1 72.105,67.97
X$19898 1801 VIA_via1_4
* cell instance $19899 r0 *1 74.385,69.23
X$19899 1801 VIA_via1_4
* cell instance $19900 r0 *1 74.005,68.95
X$19900 1801 VIA_via1_4
* cell instance $19901 r0 *1 74.005,68.95
X$19901 1801 VIA_via2_5
* cell instance $19902 r0 *1 76.855,68.67
X$19902 1802 VIA_via2_5
* cell instance $19903 r0 *1 74.005,68.67
X$19903 1802 VIA_via2_5
* cell instance $19904 r0 *1 74.955,68.67
X$19904 1802 VIA_via2_5
* cell instance $19905 r0 *1 74.955,69.23
X$19905 1802 VIA_via1_4
* cell instance $19906 r0 *1 74.005,66.43
X$19906 1802 VIA_via1_4
* cell instance $19907 r0 *1 76.855,68.25
X$19907 1802 VIA_via1_4
* cell instance $19908 r0 *1 75.715,69.23
X$19908 1803 VIA_via1_4
* cell instance $19909 r0 *1 75.335,69.37
X$19909 1803 VIA_via1_4
* cell instance $19910 r0 *1 31.825,75.11
X$19910 1804 VIA_via2_5
* cell instance $19911 r0 *1 43.985,75.95
X$19911 1804 VIA_via2_5
* cell instance $19912 r0 *1 43.985,77.21
X$19912 1804 VIA_via2_5
* cell instance $19913 r0 *1 42.845,75.95
X$19913 1804 VIA_via2_5
* cell instance $19914 r0 *1 55.385,70.35
X$19914 1804 VIA_via2_5
* cell instance $19915 r0 *1 55.385,71.33
X$19915 1804 VIA_via2_5
* cell instance $19916 r0 *1 56.145,71.33
X$19916 1804 VIA_via2_5
* cell instance $19917 r0 *1 56.145,75.25
X$19917 1804 VIA_via2_5
* cell instance $19918 r0 *1 90.915,68.95
X$19918 1804 VIA_via2_5
* cell instance $19919 r0 *1 87.495,69.23
X$19919 1804 VIA_via2_5
* cell instance $19920 r0 *1 31.825,71.33
X$19920 1804 VIA_via2_5
* cell instance $19921 r0 *1 30.875,71.33
X$19921 1804 VIA_via2_5
* cell instance $19922 r0 *1 56.145,74.83
X$19922 1804 VIA_via1_4
* cell instance $19923 r0 *1 55.385,70.77
X$19923 1804 VIA_via1_4
* cell instance $19924 r0 *1 54.055,77.63
X$19924 1804 VIA_via1_4
* cell instance $19925 r0 *1 86.735,75.11
X$19925 1804 VIA_via1_4
* cell instance $19926 r0 *1 37.525,76.37
X$19926 1804 VIA_via1_4
* cell instance $19927 r0 *1 37.525,76.37
X$19927 1804 VIA_via2_5
* cell instance $19928 r0 *1 42.845,76.37
X$19928 1804 VIA_via1_4
* cell instance $19929 r0 *1 31.825,74.83
X$19929 1804 VIA_via1_4
* cell instance $19930 r0 *1 31.255,79.17
X$19930 1804 VIA_via1_4
* cell instance $19931 r0 *1 31.255,79.17
X$19931 1804 VIA_via2_5
* cell instance $19932 r0 *1 30.875,70.77
X$19932 1804 VIA_via1_4
* cell instance $19933 r0 *1 90.915,67.97
X$19933 1804 VIA_via1_4
* cell instance $19934 r0 *1 78.375,67.97
X$19934 1804 VIA_via1_4
* cell instance $19935 r0 *1 32.015,75.11
X$19935 1804 VIA_via4_0
* cell instance $19936 r0 *1 32.015,75.11
X$19936 1804 VIA_via3_2
* cell instance $19937 r0 *1 30.335,75.11
X$19937 1804 VIA_via4_0
* cell instance $19938 r0 *1 37.335,75.95
X$19938 1804 VIA_via4_0
* cell instance $19939 r0 *1 37.335,75.11
X$19939 1804 VIA_via4_0
* cell instance $19940 r0 *1 42.655,75.95
X$19940 1804 VIA_via4_0
* cell instance $19941 r0 *1 42.655,75.95
X$19941 1804 VIA_via3_2
* cell instance $19942 r0 *1 87.735,68.95
X$19942 1804 VIA_via4_0
* cell instance $19943 r0 *1 87.735,68.95
X$19943 1804 VIA_via3_2
* cell instance $19944 r0 *1 78.495,68.95
X$19944 1804 VIA_via4_0
* cell instance $19945 r0 *1 54.135,75.25
X$19945 1804 VIA_via3_2
* cell instance $19946 r0 *1 30.335,79.17
X$19946 1804 VIA_via3_2
* cell instance $19947 r0 *1 78.495,70.21
X$19947 1804 VIA_via3_2
* cell instance $19948 r0 *1 78.495,68.25
X$19948 1804 VIA_via3_2
* cell instance $19949 r0 *1 78.375,68.25
X$19949 1804 VIA_via2_5
* cell instance $19950 r0 *1 54.135,77.35
X$19950 1804 VIA_via3_2
* cell instance $19951 r0 *1 54.055,77.35
X$19951 1804 VIA_via2_5
* cell instance $19952 r0 *1 37.335,76.37
X$19952 1804 VIA_via3_2
* cell instance $19953 r0 *1 82.555,67.97
X$19953 1805 VIA_via1_4
* cell instance $19954 r0 *1 82.555,68.11
X$19954 1805 VIA_via2_5
* cell instance $19955 r0 *1 84.835,68.95
X$19955 1805 VIA_via1_4
* cell instance $19956 r0 *1 84.645,67.97
X$19956 1805 VIA_via1_4
* cell instance $19957 r0 *1 84.645,68.11
X$19957 1805 VIA_via2_5
* cell instance $19958 r0 *1 90.725,69.23
X$19958 1806 VIA_via1_4
* cell instance $19959 r0 *1 91.105,68.11
X$19959 1806 VIA_via1_4
* cell instance $19960 r0 *1 87.495,68.39
X$19960 1807 VIA_via1_7
* cell instance $19961 r0 *1 87.495,68.39
X$19961 1807 VIA_via2_5
* cell instance $19962 r0 *1 85.785,68.39
X$19962 1807 VIA_via2_5
* cell instance $19963 r0 *1 85.785,69.23
X$19963 1807 VIA_via1_4
* cell instance $19964 r0 *1 83.505,68.39
X$19964 1808 VIA_via1_7
* cell instance $19965 r0 *1 83.505,68.39
X$19965 1808 VIA_via2_5
* cell instance $19966 r0 *1 82.555,68.39
X$19966 1808 VIA_via2_5
* cell instance $19967 r0 *1 82.555,69.23
X$19967 1808 VIA_via1_4
* cell instance $19968 r0 *1 78.755,68.25
X$19968 1809 VIA_via2_5
* cell instance $19969 r0 *1 78.755,67.97
X$19969 1809 VIA_via1_4
* cell instance $19970 r0 *1 80.465,68.25
X$19970 1809 VIA_via1_4
* cell instance $19971 r0 *1 80.465,68.25
X$19971 1809 VIA_via2_5
* cell instance $19972 r0 *1 33.345,68.95
X$19972 1810 VIA_via2_5
* cell instance $19973 r0 *1 35.815,68.95
X$19973 1810 VIA_via2_5
* cell instance $19974 r0 *1 36.575,68.95
X$19974 1810 VIA_via1_4
* cell instance $19975 r0 *1 36.575,68.95
X$19975 1810 VIA_via2_5
* cell instance $19976 r0 *1 35.815,70.77
X$19976 1810 VIA_via1_4
* cell instance $19977 r0 *1 33.345,67.97
X$19977 1810 VIA_via1_4
* cell instance $19978 r0 *1 77.995,67.97
X$19978 1811 VIA_via1_4
* cell instance $19979 r0 *1 77.995,68.11
X$19979 1811 VIA_via2_5
* cell instance $19980 r0 *1 79.515,68.11
X$19980 1811 VIA_via1_4
* cell instance $19981 r0 *1 79.515,68.11
X$19981 1811 VIA_via2_5
* cell instance $19982 r0 *1 34.295,68.39
X$19982 1812 VIA_via1_7
* cell instance $19983 r0 *1 34.295,69.23
X$19983 1812 VIA_via1_4
* cell instance $19984 r0 *1 49.875,82.81
X$19984 1813 VIA_via1_7
* cell instance $19985 r0 *1 49.875,83.79
X$19985 1813 VIA_via1_7
* cell instance $19986 r0 *1 45.315,82.25
X$19986 1813 VIA_via2_5
* cell instance $19987 r0 *1 48.165,88.55
X$19987 1813 VIA_via2_5
* cell instance $19988 r0 *1 46.455,88.55
X$19988 1813 VIA_via2_5
* cell instance $19989 r0 *1 45.505,74.83
X$19989 1813 VIA_via2_5
* cell instance $19990 r0 *1 44.365,73.71
X$19990 1813 VIA_via2_5
* cell instance $19991 r0 *1 42.845,73.71
X$19991 1813 VIA_via2_5
* cell instance $19992 r0 *1 50.255,88.55
X$19992 1813 VIA_via2_5
* cell instance $19993 r0 *1 49.685,88.55
X$19993 1813 VIA_via2_5
* cell instance $19994 r0 *1 49.875,88.55
X$19994 1813 VIA_via2_5
* cell instance $19995 r0 *1 49.875,82.25
X$19995 1813 VIA_via2_5
* cell instance $19996 r0 *1 50.255,88.83
X$19996 1813 VIA_via1_4
* cell instance $19997 r0 *1 49.875,90.37
X$19997 1813 VIA_via1_4
* cell instance $19998 r0 *1 47.595,74.83
X$19998 1813 VIA_via1_4
* cell instance $19999 r0 *1 47.595,74.69
X$19999 1813 VIA_via2_5
* cell instance $20000 r0 *1 45.315,79.17
X$20000 1813 VIA_via1_4
* cell instance $20001 r0 *1 44.365,74.83
X$20001 1813 VIA_via1_4
* cell instance $20002 r0 *1 44.365,74.83
X$20002 1813 VIA_via2_5
* cell instance $20003 r0 *1 48.165,88.83
X$20003 1813 VIA_via1_4
* cell instance $20004 r0 *1 46.455,90.37
X$20004 1813 VIA_via1_4
* cell instance $20005 r0 *1 42.655,72.03
X$20005 1813 VIA_via1_4
* cell instance $20006 r0 *1 43.605,67.97
X$20006 1813 VIA_via1_4
* cell instance $20007 r0 *1 43.605,68.11
X$20007 1813 VIA_via2_5
* cell instance $20008 r0 *1 42.275,67.97
X$20008 1813 VIA_via1_4
* cell instance $20009 r0 *1 42.275,68.11
X$20009 1813 VIA_via2_5
* cell instance $20010 r0 *1 71.535,70.21
X$20010 1814 VIA_via1_7
* cell instance $20011 r0 *1 71.535,69.23
X$20011 1814 VIA_via2_5
* cell instance $20012 r0 *1 68.305,69.23
X$20012 1814 VIA_via1_4
* cell instance $20013 r0 *1 68.305,69.23
X$20013 1814 VIA_via2_5
* cell instance $20014 r0 *1 73.055,68.39
X$20014 1815 VIA_via1_7
* cell instance $20015 r0 *1 73.055,68.39
X$20015 1815 VIA_via2_5
* cell instance $20016 r0 *1 71.725,68.39
X$20016 1815 VIA_via2_5
* cell instance $20017 r0 *1 71.725,69.23
X$20017 1815 VIA_via1_4
* cell instance $20018 r0 *1 50.255,67.97
X$20018 1816 VIA_via1_4
* cell instance $20019 r0 *1 50.255,68.11
X$20019 1816 VIA_via2_5
* cell instance $20020 r0 *1 49.305,68.11
X$20020 1816 VIA_via1_4
* cell instance $20021 r0 *1 49.305,68.11
X$20021 1816 VIA_via2_5
* cell instance $20022 r0 *1 64.125,68.81
X$20022 1817 VIA_via2_5
* cell instance $20023 r0 *1 67.355,68.81
X$20023 1817 VIA_via2_5
* cell instance $20024 r0 *1 64.125,69.23
X$20024 1817 VIA_via1_4
* cell instance $20025 r0 *1 67.355,68.11
X$20025 1817 VIA_via1_4
* cell instance $20026 r0 *1 64.885,68.39
X$20026 1818 VIA_via1_7
* cell instance $20027 r0 *1 64.885,68.53
X$20027 1818 VIA_via2_5
* cell instance $20028 r0 *1 66.215,68.53
X$20028 1818 VIA_via2_5
* cell instance $20029 r0 *1 66.215,69.23
X$20029 1818 VIA_via1_4
* cell instance $20030 r0 *1 5.605,70.77
X$20030 1819 VIA_via1_4
* cell instance $20031 r0 *1 5.605,70.77
X$20031 1819 VIA_via2_5
* cell instance $20032 r0 *1 6.555,70.77
X$20032 1819 VIA_via1_4
* cell instance $20033 r0 *1 6.555,70.77
X$20033 1819 VIA_via2_5
* cell instance $20034 r0 *1 7.315,70.77
X$20034 1819 VIA_via1_4
* cell instance $20035 r0 *1 7.315,70.77
X$20035 1819 VIA_via2_5
* cell instance $20036 r0 *1 13.965,85.61
X$20036 1820 VIA_via1_7
* cell instance $20037 r0 *1 13.965,85.75
X$20037 1820 VIA_via2_5
* cell instance $20038 r0 *1 18.525,72.31
X$20038 1820 VIA_via2_5
* cell instance $20039 r0 *1 7.505,85.75
X$20039 1820 VIA_via2_5
* cell instance $20040 r0 *1 6.555,88.27
X$20040 1820 VIA_via2_5
* cell instance $20041 r0 *1 10.165,88.27
X$20041 1820 VIA_via2_5
* cell instance $20042 r0 *1 11.305,88.55
X$20042 1820 VIA_via2_5
* cell instance $20043 r0 *1 18.525,77.63
X$20043 1820 VIA_via2_5
* cell instance $20044 r0 *1 15.485,77.77
X$20044 1820 VIA_via2_5
* cell instance $20045 r0 *1 14.915,80.43
X$20045 1820 VIA_via2_5
* cell instance $20046 r0 *1 16.055,77.77
X$20046 1820 VIA_via2_5
* cell instance $20047 r0 *1 14.915,85.75
X$20047 1820 VIA_via2_5
* cell instance $20048 r0 *1 20.045,72.31
X$20048 1820 VIA_via2_5
* cell instance $20049 r0 *1 6.555,85.89
X$20049 1820 VIA_via2_5
* cell instance $20050 r0 *1 20.045,72.03
X$20050 1820 VIA_via1_4
* cell instance $20051 r0 *1 18.715,70.77
X$20051 1820 VIA_via1_4
* cell instance $20052 r0 *1 11.305,88.83
X$20052 1820 VIA_via1_4
* cell instance $20053 r0 *1 7.695,81.97
X$20053 1820 VIA_via1_4
* cell instance $20054 r0 *1 5.795,86.03
X$20054 1820 VIA_via1_4
* cell instance $20055 r0 *1 5.795,85.89
X$20055 1820 VIA_via2_5
* cell instance $20056 r0 *1 10.165,87.57
X$20056 1820 VIA_via1_4
* cell instance $20057 r0 *1 6.555,88.83
X$20057 1820 VIA_via1_4
* cell instance $20058 r0 *1 16.055,74.83
X$20058 1820 VIA_via1_4
* cell instance $20059 r0 *1 18.715,77.63
X$20059 1820 VIA_via1_4
* cell instance $20060 r0 *1 18.715,77.63
X$20060 1820 VIA_via2_5
* cell instance $20061 r0 *1 15.485,80.43
X$20061 1820 VIA_via1_4
* cell instance $20062 r0 *1 15.485,80.43
X$20062 1820 VIA_via2_5
* cell instance $20063 r0 *1 25.935,72.03
X$20063 1821 VIA_via1_4
* cell instance $20064 r0 *1 25.555,71.05
X$20064 1821 VIA_via1_4
* cell instance $20065 r0 *1 25.935,70.77
X$20065 1821 VIA_via1_4
* cell instance $20066 r0 *1 24.605,73.15
X$20066 1822 VIA_via2_5
* cell instance $20067 r0 *1 19.095,80.57
X$20067 1822 VIA_via2_5
* cell instance $20068 r0 *1 19.665,88.55
X$20068 1822 VIA_via2_5
* cell instance $20069 r0 *1 19.665,87.29
X$20069 1822 VIA_via2_5
* cell instance $20070 r0 *1 14.535,88.55
X$20070 1822 VIA_via2_5
* cell instance $20071 r0 *1 16.815,88.55
X$20071 1822 VIA_via2_5
* cell instance $20072 r0 *1 21.945,87.29
X$20072 1822 VIA_via2_5
* cell instance $20073 r0 *1 26.505,73.15
X$20073 1822 VIA_via2_5
* cell instance $20074 r0 *1 16.815,87.57
X$20074 1822 VIA_via1_4
* cell instance $20075 r0 *1 14.535,88.83
X$20075 1822 VIA_via1_4
* cell instance $20076 r0 *1 19.665,88.83
X$20076 1822 VIA_via1_4
* cell instance $20077 r0 *1 21.945,87.57
X$20077 1822 VIA_via1_4
* cell instance $20078 r0 *1 26.505,69.23
X$20078 1822 VIA_via1_4
* cell instance $20079 r0 *1 26.505,70.77
X$20079 1822 VIA_via1_4
* cell instance $20080 r0 *1 24.605,74.83
X$20080 1822 VIA_via1_4
* cell instance $20081 r0 *1 23.465,76.37
X$20081 1822 VIA_via1_4
* cell instance $20082 r0 *1 19.285,84.35
X$20082 1822 VIA_via1_4
* cell instance $20083 r0 *1 23.655,80.43
X$20083 1822 VIA_via1_4
* cell instance $20084 r0 *1 23.655,80.57
X$20084 1822 VIA_via2_5
* cell instance $20085 r0 *1 18.715,80.43
X$20085 1822 VIA_via1_4
* cell instance $20086 r0 *1 18.715,80.57
X$20086 1822 VIA_via2_5
* cell instance $20087 r0 *1 31.825,70.77
X$20087 1823 VIA_via1_4
* cell instance $20088 r0 *1 32.015,71.75
X$20088 1823 VIA_via1_4
* cell instance $20089 r0 *1 32.205,70.77
X$20089 1823 VIA_via1_4
* cell instance $20090 r0 *1 32.585,73.57
X$20090 1823 VIA_via1_4
* cell instance $20091 r0 *1 32.015,70.35
X$20091 1824 VIA_via2_5
* cell instance $20092 r0 *1 30.495,70.35
X$20092 1824 VIA_via2_5
* cell instance $20093 r0 *1 30.495,70.77
X$20093 1824 VIA_via1_4
* cell instance $20094 r0 *1 31.825,71.05
X$20094 1824 VIA_via1_4
* cell instance $20095 r0 *1 41.325,70.77
X$20095 1825 VIA_via1_4
* cell instance $20096 r0 *1 40.565,69.65
X$20096 1825 VIA_via1_4
* cell instance $20097 r0 *1 40.945,69.23
X$20097 1825 VIA_via1_4
* cell instance $20098 r0 *1 63.365,70.77
X$20098 1826 VIA_via1_4
* cell instance $20099 r0 *1 62.985,72.03
X$20099 1826 VIA_via1_4
* cell instance $20100 r0 *1 62.985,71.05
X$20100 1826 VIA_via1_4
* cell instance $20101 r0 *1 69.255,70.63
X$20101 1827 VIA_via1_4
* cell instance $20102 r0 *1 69.255,70.63
X$20102 1827 VIA_via2_5
* cell instance $20103 r0 *1 65.645,70.77
X$20103 1827 VIA_via1_4
* cell instance $20104 r0 *1 65.645,70.77
X$20104 1827 VIA_via2_5
* cell instance $20105 r0 *1 69.445,70.77
X$20105 1828 VIA_via2_5
* cell instance $20106 r0 *1 70.775,70.77
X$20106 1828 VIA_via2_5
* cell instance $20107 r0 *1 71.155,70.77
X$20107 1828 VIA_via1_4
* cell instance $20108 r0 *1 71.155,70.77
X$20108 1828 VIA_via2_5
* cell instance $20109 r0 *1 69.445,72.03
X$20109 1828 VIA_via1_4
* cell instance $20110 r0 *1 70.585,69.65
X$20110 1828 VIA_via1_4
* cell instance $20111 r0 *1 75.715,73.57
X$20111 1829 VIA_via1_4
* cell instance $20112 r0 *1 75.335,73.57
X$20112 1829 VIA_via1_4
* cell instance $20113 r0 *1 74.955,70.77
X$20113 1829 VIA_via1_4
* cell instance $20114 r0 *1 75.905,70.21
X$20114 1830 VIA_via1_7
* cell instance $20115 r0 *1 76.285,69.23
X$20115 1830 VIA_via1_4
* cell instance $20116 r0 *1 77.425,69.23
X$20116 1831 VIA_via1_4
* cell instance $20117 r0 *1 76.665,69.65
X$20117 1831 VIA_via1_4
* cell instance $20118 r0 *1 78.755,69.51
X$20118 1832 VIA_via1_4
* cell instance $20119 r0 *1 78.375,69.23
X$20119 1832 VIA_via1_4
* cell instance $20120 r0 *1 82.555,71.05
X$20120 1833 VIA_via2_5
* cell instance $20121 r0 *1 80.465,70.77
X$20121 1833 VIA_via1_4
* cell instance $20122 r0 *1 80.465,70.77
X$20122 1833 VIA_via2_5
* cell instance $20123 r0 *1 84.075,71.05
X$20123 1833 VIA_via1_4
* cell instance $20124 r0 *1 84.075,71.05
X$20124 1833 VIA_via2_5
* cell instance $20125 r0 *1 82.555,72.03
X$20125 1833 VIA_via1_4
* cell instance $20126 r0 *1 6.365,69.37
X$20126 1834 VIA_via1_4
* cell instance $20127 r0 *1 6.365,69.37
X$20127 1834 VIA_via2_5
* cell instance $20128 r0 *1 2.755,69.23
X$20128 1834 VIA_via1_4
* cell instance $20129 r0 *1 2.755,69.37
X$20129 1834 VIA_via2_5
* cell instance $20130 r0 *1 3.325,70.77
X$20130 1835 VIA_via1_4
* cell instance $20131 r0 *1 3.325,70.91
X$20131 1835 VIA_via2_5
* cell instance $20132 r0 *1 8.265,70.91
X$20132 1835 VIA_via1_4
* cell instance $20133 r0 *1 8.265,70.91
X$20133 1835 VIA_via2_5
* cell instance $20134 r0 *1 10.165,69.37
X$20134 1836 VIA_via1_4
* cell instance $20135 r0 *1 10.165,69.37
X$20135 1836 VIA_via2_5
* cell instance $20136 r0 *1 10.735,69.23
X$20136 1836 VIA_via1_4
* cell instance $20137 r0 *1 10.735,69.37
X$20137 1836 VIA_via2_5
* cell instance $20138 r0 *1 83.505,71.61
X$20138 1837 VIA_via1_7
* cell instance $20139 r0 *1 78.565,69.79
X$20139 1837 VIA_via2_5
* cell instance $20140 r0 *1 83.505,69.79
X$20140 1837 VIA_via2_5
* cell instance $20141 r0 *1 78.565,69.23
X$20141 1837 VIA_via1_4
* cell instance $20142 r0 *1 8.075,69.37
X$20142 1838 VIA_via2_5
* cell instance $20143 r0 *1 8.835,69.37
X$20143 1838 VIA_via1_4
* cell instance $20144 r0 *1 8.835,69.37
X$20144 1838 VIA_via2_5
* cell instance $20145 r0 *1 8.075,67.97
X$20145 1838 VIA_via1_4
* cell instance $20146 r0 *1 80.845,70.91
X$20146 1839 VIA_via1_4
* cell instance $20147 r0 *1 80.845,70.91
X$20147 1839 VIA_via2_5
* cell instance $20148 r0 *1 81.795,70.77
X$20148 1839 VIA_via1_4
* cell instance $20149 r0 *1 81.795,70.91
X$20149 1839 VIA_via2_5
* cell instance $20150 r0 *1 6.935,70.63
X$20150 1840 VIA_via1_4
* cell instance $20151 r0 *1 6.935,70.63
X$20151 1840 VIA_via2_5
* cell instance $20152 r0 *1 11.495,70.77
X$20152 1840 VIA_via1_4
* cell instance $20153 r0 *1 11.495,70.63
X$20153 1840 VIA_via2_5
* cell instance $20154 r0 *1 17.195,69.79
X$20154 1841 VIA_via1_7
* cell instance $20155 r0 *1 14.915,70.07
X$20155 1841 VIA_via2_5
* cell instance $20156 r0 *1 17.195,70.07
X$20156 1841 VIA_via2_5
* cell instance $20157 r0 *1 14.915,70.77
X$20157 1841 VIA_via1_4
* cell instance $20158 r0 *1 16.245,70.35
X$20158 1842 VIA_via2_5
* cell instance $20159 r0 *1 17.195,72.03
X$20159 1842 VIA_via1_4
* cell instance $20160 r0 *1 17.195,70.35
X$20160 1842 VIA_via1_4
* cell instance $20161 r0 *1 17.195,70.35
X$20161 1842 VIA_via2_5
* cell instance $20162 r0 *1 16.245,69.23
X$20162 1842 VIA_via1_4
* cell instance $20163 r0 *1 21.185,70.91
X$20163 1843 VIA_via2_5
* cell instance $20164 r0 *1 21.375,72.03
X$20164 1843 VIA_via1_4
* cell instance $20165 r0 *1 21.185,69.23
X$20165 1843 VIA_via1_4
* cell instance $20166 r0 *1 18.145,70.77
X$20166 1843 VIA_via1_4
* cell instance $20167 r0 *1 18.145,70.91
X$20167 1843 VIA_via2_5
* cell instance $20168 r0 *1 78.185,70.21
X$20168 1844 VIA_via1_7
* cell instance $20169 r0 *1 78.185,69.23
X$20169 1844 VIA_via1_4
* cell instance $20170 r0 *1 20.425,71.61
X$20170 1845 VIA_via1_7
* cell instance $20171 r0 *1 20.425,70.77
X$20171 1845 VIA_via2_5
* cell instance $20172 r0 *1 20.045,70.77
X$20172 1845 VIA_via1_4
* cell instance $20173 r0 *1 20.045,70.77
X$20173 1845 VIA_via2_5
* cell instance $20174 r0 *1 77.615,69.65
X$20174 1846 VIA_via2_5
* cell instance $20175 r0 *1 76.095,69.65
X$20175 1846 VIA_via1_4
* cell instance $20176 r0 *1 76.095,69.65
X$20176 1846 VIA_via2_5
* cell instance $20177 r0 *1 77.615,69.23
X$20177 1846 VIA_via1_4
* cell instance $20178 r0 *1 23.275,70.77
X$20178 1847 VIA_via1_4
* cell instance $20179 r0 *1 23.275,70.91
X$20179 1847 VIA_via2_5
* cell instance $20180 r0 *1 26.885,70.91
X$20180 1847 VIA_via1_4
* cell instance $20181 r0 *1 26.885,70.91
X$20181 1847 VIA_via2_5
* cell instance $20182 r0 *1 15.865,76.37
X$20182 1848 VIA_via2_5
* cell instance $20183 r0 *1 15.105,76.37
X$20183 1848 VIA_via2_5
* cell instance $20184 r0 *1 19.285,76.37
X$20184 1848 VIA_via2_5
* cell instance $20185 r0 *1 23.465,74.83
X$20185 1848 VIA_via2_5
* cell instance $20186 r0 *1 19.475,76.37
X$20186 1848 VIA_via2_5
* cell instance $20187 r0 *1 23.465,70.77
X$20187 1848 VIA_via2_5
* cell instance $20188 r0 *1 24.035,70.77
X$20188 1848 VIA_via1_4
* cell instance $20189 r0 *1 24.035,70.77
X$20189 1848 VIA_via2_5
* cell instance $20190 r0 *1 20.805,70.77
X$20190 1848 VIA_via1_4
* cell instance $20191 r0 *1 20.805,70.77
X$20191 1848 VIA_via2_5
* cell instance $20192 r0 *1 15.675,76.37
X$20192 1848 VIA_via1_4
* cell instance $20193 r0 *1 15.675,76.37
X$20193 1848 VIA_via2_5
* cell instance $20194 r0 *1 14.915,77.63
X$20194 1848 VIA_via1_4
* cell instance $20195 r0 *1 18.905,76.37
X$20195 1848 VIA_via1_4
* cell instance $20196 r0 *1 18.905,76.37
X$20196 1848 VIA_via2_5
* cell instance $20197 r0 *1 19.475,74.83
X$20197 1848 VIA_via1_4
* cell instance $20198 r0 *1 19.475,74.83
X$20198 1848 VIA_via2_5
* cell instance $20199 r0 *1 22.135,74.83
X$20199 1848 VIA_via1_4
* cell instance $20200 r0 *1 22.135,74.83
X$20200 1848 VIA_via2_5
* cell instance $20201 r0 *1 19.285,77.63
X$20201 1848 VIA_via1_4
* cell instance $20202 r0 *1 16.245,81.97
X$20202 1848 VIA_via1_4
* cell instance $20203 r0 *1 27.835,69.23
X$20203 1849 VIA_via1_4
* cell instance $20204 r0 *1 27.835,69.37
X$20204 1849 VIA_via2_5
* cell instance $20205 r0 *1 26.885,69.37
X$20205 1849 VIA_via1_4
* cell instance $20206 r0 *1 26.885,69.37
X$20206 1849 VIA_via2_5
* cell instance $20207 r0 *1 30.685,70.49
X$20207 1850 VIA_via1_7
* cell instance $20208 r0 *1 30.685,70.49
X$20208 1850 VIA_via2_5
* cell instance $20209 r0 *1 29.735,70.49
X$20209 1850 VIA_via2_5
* cell instance $20210 r0 *1 29.735,72.03
X$20210 1850 VIA_via1_4
* cell instance $20211 r0 *1 30.305,68.39
X$20211 1851 VIA_via1_7
* cell instance $20212 r0 *1 30.305,69.65
X$20212 1851 VIA_via2_5
* cell instance $20213 r0 *1 34.105,69.65
X$20213 1851 VIA_via2_5
* cell instance $20214 r0 *1 34.105,70.77
X$20214 1851 VIA_via1_4
* cell instance $20215 r0 *1 32.395,70.77
X$20215 1852 VIA_via1_4
* cell instance $20216 r0 *1 32.395,70.77
X$20216 1852 VIA_via2_5
* cell instance $20217 r0 *1 31.255,70.77
X$20217 1852 VIA_via1_4
* cell instance $20218 r0 *1 31.255,70.77
X$20218 1852 VIA_via2_5
* cell instance $20219 r0 *1 68.875,70.77
X$20219 1853 VIA_via1_4
* cell instance $20220 r0 *1 68.875,70.77
X$20220 1853 VIA_via2_5
* cell instance $20221 r0 *1 68.875,72.03
X$20221 1853 VIA_via1_4
* cell instance $20222 r0 *1 67.925,70.77
X$20222 1853 VIA_via1_4
* cell instance $20223 r0 *1 67.925,70.77
X$20223 1853 VIA_via2_5
* cell instance $20224 r0 *1 38.285,69.23
X$20224 1854 VIA_via1_4
* cell instance $20225 r0 *1 38.285,69.37
X$20225 1854 VIA_via2_5
* cell instance $20226 r0 *1 41.895,69.37
X$20226 1854 VIA_via1_4
* cell instance $20227 r0 *1 41.895,69.37
X$20227 1854 VIA_via2_5
* cell instance $20228 r0 *1 36.195,70.77
X$20228 1855 VIA_via2_5
* cell instance $20229 r0 *1 32.965,70.77
X$20229 1855 VIA_via1_4
* cell instance $20230 r0 *1 32.965,70.77
X$20230 1855 VIA_via2_5
* cell instance $20231 r0 *1 36.195,71.75
X$20231 1855 VIA_via1_4
* cell instance $20232 r0 *1 36.385,70.77
X$20232 1855 VIA_via1_4
* cell instance $20233 r0 *1 36.385,70.77
X$20233 1855 VIA_via2_5
* cell instance $20234 r0 *1 39.425,70.77
X$20234 1856 VIA_via1_4
* cell instance $20235 r0 *1 39.425,70.77
X$20235 1856 VIA_via2_5
* cell instance $20236 r0 *1 40.755,70.77
X$20236 1856 VIA_via1_4
* cell instance $20237 r0 *1 40.755,70.77
X$20237 1856 VIA_via2_5
* cell instance $20238 r0 *1 40.755,71.75
X$20238 1856 VIA_via1_4
* cell instance $20239 r0 *1 64.315,69.51
X$20239 1857 VIA_via1_7
* cell instance $20240 r0 *1 64.315,69.79
X$20240 1857 VIA_via2_5
* cell instance $20241 r0 *1 64.315,94.43
X$20241 1857 VIA_via1_4
* cell instance $20242 r0 *1 64.315,94.43
X$20242 1857 VIA_via2_5
* cell instance $20243 r0 *1 63.655,94.43
X$20243 1857 VIA_via3_2
* cell instance $20244 r0 *1 63.655,69.79
X$20244 1857 VIA_via3_2
* cell instance $20245 r0 *1 64.315,70.77
X$20245 1858 VIA_via1_4
* cell instance $20246 r0 *1 64.315,70.77
X$20246 1858 VIA_via2_5
* cell instance $20247 r0 *1 60.705,70.77
X$20247 1858 VIA_via1_4
* cell instance $20248 r0 *1 60.705,70.77
X$20248 1858 VIA_via2_5
* cell instance $20249 r0 *1 47.405,66.99
X$20249 1859 VIA_via1_7
* cell instance $20250 r0 *1 47.405,70.7
X$20250 1859 VIA_via1_4
* cell instance $20251 r0 *1 56.715,70.77
X$20251 1860 VIA_via1_4
* cell instance $20252 r0 *1 56.715,70.77
X$20252 1860 VIA_via2_5
* cell instance $20253 r0 *1 55.765,70.77
X$20253 1860 VIA_via1_4
* cell instance $20254 r0 *1 55.765,70.77
X$20254 1860 VIA_via2_5
* cell instance $20255 r0 *1 55.575,69.23
X$20255 1861 VIA_via1_4
* cell instance $20256 r0 *1 55.575,70.49
X$20256 1861 VIA_via1_4
* cell instance $20257 r0 *1 54.245,70.77
X$20257 1862 VIA_via1_4
* cell instance $20258 r0 *1 54.245,70.91
X$20258 1862 VIA_via2_5
* cell instance $20259 r0 *1 56.145,70.91
X$20259 1862 VIA_via1_4
* cell instance $20260 r0 *1 56.145,70.91
X$20260 1862 VIA_via2_5
* cell instance $20261 r0 *1 55.005,69.37
X$20261 1863 VIA_via2_5
* cell instance $20262 r0 *1 53.485,69.37
X$20262 1863 VIA_via2_5
* cell instance $20263 r0 *1 55.005,68.11
X$20263 1863 VIA_via1_4
* cell instance $20264 r0 *1 53.485,70.77
X$20264 1863 VIA_via1_4
* cell instance $20265 r0 *1 55.195,70.77
X$20265 1864 VIA_via1_4
* cell instance $20266 r0 *1 55.195,66.71
X$20266 1864 VIA_via1_4
* cell instance $20267 r0 *1 54.435,70.77
X$20267 1865 VIA_via2_5
* cell instance $20268 r0 *1 54.435,69.23
X$20268 1865 VIA_via1_4
* cell instance $20269 r0 *1 55.005,70.77
X$20269 1865 VIA_via1_4
* cell instance $20270 r0 *1 55.005,70.77
X$20270 1865 VIA_via2_5
* cell instance $20271 r0 *1 53.675,70.49
X$20271 1866 VIA_via1_7
* cell instance $20272 r0 *1 53.675,70.49
X$20272 1866 VIA_via2_5
* cell instance $20273 r0 *1 53.675,95.97
X$20273 1866 VIA_via1_4
* cell instance $20274 r0 *1 53.675,95.97
X$20274 1866 VIA_via2_5
* cell instance $20275 r0 *1 53.855,95.97
X$20275 1866 VIA_via3_2
* cell instance $20276 r0 *1 53.855,70.49
X$20276 1866 VIA_via3_2
* cell instance $20277 r0 *1 1.615,71.75
X$20277 1867 VIA_via2_5
* cell instance $20278 r0 *1 1.615,72.03
X$20278 1867 VIA_via1_4
* cell instance $20279 r0 *1 0.935,71.75
X$20279 1867 VIA_via3_2
* cell instance $20280 r0 *1 0.935,71.75
X$20280 1867 VIA_via4_0
* cell instance $20281 r0 *1 10.925,73.57
X$20281 1868 VIA_via2_5
* cell instance $20282 r0 *1 10.925,72.03
X$20282 1868 VIA_via1_4
* cell instance $20283 r0 *1 10.545,72.45
X$20283 1868 VIA_via1_4
* cell instance $20284 r0 *1 12.445,73.57
X$20284 1868 VIA_via1_4
* cell instance $20285 r0 *1 12.445,73.57
X$20285 1868 VIA_via2_5
* cell instance $20286 r0 *1 11.685,71.19
X$20286 1869 VIA_via1_7
* cell instance $20287 r0 *1 12.255,74.83
X$20287 1869 VIA_via1_4
* cell instance $20288 r0 *1 16.625,72.03
X$20288 1870 VIA_via1_4
* cell instance $20289 r0 *1 15.865,72.45
X$20289 1870 VIA_via1_4
* cell instance $20290 r0 *1 16.245,73.57
X$20290 1870 VIA_via1_4
* cell instance $20291 r0 *1 22.325,72.03
X$20291 1871 VIA_via2_5
* cell instance $20292 r0 *1 19.475,72.03
X$20292 1871 VIA_via1_4
* cell instance $20293 r0 *1 19.475,72.03
X$20293 1871 VIA_via2_5
* cell instance $20294 r0 *1 22.325,71.05
X$20294 1871 VIA_via1_4
* cell instance $20295 r0 *1 20.805,72.03
X$20295 1871 VIA_via1_4
* cell instance $20296 r0 *1 20.805,72.03
X$20296 1871 VIA_via2_5
* cell instance $20297 r0 *1 21.755,72.59
X$20297 1872 VIA_via1_7
* cell instance $20298 r0 *1 21.565,73.57
X$20298 1872 VIA_via1_4
* cell instance $20299 r0 *1 36.765,71.19
X$20299 1873 VIA_via1_7
* cell instance $20300 r0 *1 36.955,72.03
X$20300 1873 VIA_via1_4
* cell instance $20301 r0 *1 41.705,71.19
X$20301 1874 VIA_via1_7
* cell instance $20302 r0 *1 41.135,72.03
X$20302 1874 VIA_via1_4
* cell instance $20303 r0 *1 47.595,71.19
X$20303 1875 VIA_via1_7
* cell instance $20304 r0 *1 48.165,76.37
X$20304 1875 VIA_via1_4
* cell instance $20305 r0 *1 51.015,71.75
X$20305 1876 VIA_via2_5
* cell instance $20306 r0 *1 52.915,72.03
X$20306 1876 VIA_via1_4
* cell instance $20307 r0 *1 52.915,71.89
X$20307 1876 VIA_via2_5
* cell instance $20308 r0 *1 51.015,71.05
X$20308 1876 VIA_via1_4
* cell instance $20309 r0 *1 48.355,72.03
X$20309 1876 VIA_via1_4
* cell instance $20310 r0 *1 48.355,72.03
X$20310 1876 VIA_via2_5
* cell instance $20311 r0 *1 49.305,72.31
X$20311 1877 VIA_via1_4
* cell instance $20312 r0 *1 48.735,70.77
X$20312 1877 VIA_via1_4
* cell instance $20313 r0 *1 51.775,71.75
X$20313 1878 VIA_via2_5
* cell instance $20314 r0 *1 53.485,71.75
X$20314 1878 VIA_via2_5
* cell instance $20315 r0 *1 51.775,70.77
X$20315 1878 VIA_via1_4
* cell instance $20316 r0 *1 52.535,71.75
X$20316 1878 VIA_via1_4
* cell instance $20317 r0 *1 52.535,71.75
X$20317 1878 VIA_via2_5
* cell instance $20318 r0 *1 53.485,72.03
X$20318 1878 VIA_via1_4
* cell instance $20319 r0 *1 54.055,74.83
X$20319 1879 VIA_via1_4
* cell instance $20320 r0 *1 54.245,72.31
X$20320 1879 VIA_via1_4
* cell instance $20321 r0 *1 63.555,72.45
X$20321 1880 VIA_via2_5
* cell instance $20322 r0 *1 61.465,72.45
X$20322 1880 VIA_via2_5
* cell instance $20323 r0 *1 63.555,72.03
X$20323 1880 VIA_via1_4
* cell instance $20324 r0 *1 62.605,72.45
X$20324 1880 VIA_via1_4
* cell instance $20325 r0 *1 62.605,72.45
X$20325 1880 VIA_via2_5
* cell instance $20326 r0 *1 61.465,73.57
X$20326 1880 VIA_via1_4
* cell instance $20327 r0 *1 65.835,71.61
X$20327 1881 VIA_via1_7
* cell instance $20328 r0 *1 66.025,69.23
X$20328 1881 VIA_via1_4
* cell instance $20329 r0 *1 66.595,71.61
X$20329 1882 VIA_via1_7
* cell instance $20330 r0 *1 66.785,69.23
X$20330 1882 VIA_via1_4
* cell instance $20331 r0 *1 75.905,72.03
X$20331 1883 VIA_via1_4
* cell instance $20332 r0 *1 75.525,71.75
X$20332 1883 VIA_via1_4
* cell instance $20333 r0 *1 75.525,70.77
X$20333 1883 VIA_via1_4
* cell instance $20334 r0 *1 78.945,72.59
X$20334 1884 VIA_via1_7
* cell instance $20335 r0 *1 78.755,73.57
X$20335 1884 VIA_via1_4
* cell instance $20336 r0 *1 79.705,73.71
X$20336 1885 VIA_via2_5
* cell instance $20337 r0 *1 78.565,73.71
X$20337 1885 VIA_via2_5
* cell instance $20338 r0 *1 81.035,73.71
X$20338 1885 VIA_via1_4
* cell instance $20339 r0 *1 81.035,73.71
X$20339 1885 VIA_via2_5
* cell instance $20340 r0 *1 79.515,72.03
X$20340 1885 VIA_via1_4
* cell instance $20341 r0 *1 78.565,72.03
X$20341 1885 VIA_via1_4
* cell instance $20342 r0 *1 81.795,72.59
X$20342 1886 VIA_via1_7
* cell instance $20343 r0 *1 81.985,73.57
X$20343 1886 VIA_via1_4
* cell instance $20344 r0 *1 85.405,71.75
X$20344 1887 VIA_via2_5
* cell instance $20345 r0 *1 83.125,71.75
X$20345 1887 VIA_via2_5
* cell instance $20346 r0 *1 87.875,71.75
X$20346 1887 VIA_via1_4
* cell instance $20347 r0 *1 87.875,71.75
X$20347 1887 VIA_via2_5
* cell instance $20348 r0 *1 83.125,72.03
X$20348 1887 VIA_via1_4
* cell instance $20349 r0 *1 85.405,70.77
X$20349 1887 VIA_via1_4
* cell instance $20350 r0 *1 85.785,71.19
X$20350 1888 VIA_via1_7
* cell instance $20351 r0 *1 85.595,72.03
X$20351 1888 VIA_via1_4
* cell instance $20352 r0 *1 94.145,71.75
X$20352 1889 VIA_via2_5
* cell instance $20353 r0 *1 94.145,72.03
X$20353 1889 VIA_via1_4
* cell instance $20354 r0 *1 94.455,71.75
X$20354 1889 VIA_via4_0
* cell instance $20355 r0 *1 94.455,71.75
X$20355 1889 VIA_via3_2
* cell instance $20356 r0 *1 8.265,72.03
X$20356 1890 VIA_via1_4
* cell instance $20357 r0 *1 8.265,71.89
X$20357 1890 VIA_via2_5
* cell instance $20358 r0 *1 11.875,71.89
X$20358 1890 VIA_via1_4
* cell instance $20359 r0 *1 11.875,71.89
X$20359 1890 VIA_via2_5
* cell instance $20360 r0 *1 18.715,72.03
X$20360 1891 VIA_via1_4
* cell instance $20361 r0 *1 18.715,72.03
X$20361 1891 VIA_via2_5
* cell instance $20362 r0 *1 17.575,72.03
X$20362 1891 VIA_via1_4
* cell instance $20363 r0 *1 17.575,72.03
X$20363 1891 VIA_via2_5
* cell instance $20364 r0 *1 80.465,71.61
X$20364 1892 VIA_via1_7
* cell instance $20365 r0 *1 80.465,71.05
X$20365 1892 VIA_via2_5
* cell instance $20366 r0 *1 77.805,71.05
X$20366 1892 VIA_via2_5
* cell instance $20367 r0 *1 77.805,70.77
X$20367 1892 VIA_via1_4
* cell instance $20368 r0 *1 73.245,72.03
X$20368 1893 VIA_via1_4
* cell instance $20369 r0 *1 73.245,72.03
X$20369 1893 VIA_via2_5
* cell instance $20370 r0 *1 76.855,72.03
X$20370 1893 VIA_via1_4
* cell instance $20371 r0 *1 76.855,72.03
X$20371 1893 VIA_via2_5
* cell instance $20372 r0 *1 33.915,71.19
X$20372 1894 VIA_via1_7
* cell instance $20373 r0 *1 33.915,72.03
X$20373 1894 VIA_via1_4
* cell instance $20374 r0 *1 40.375,71.19
X$20374 1895 VIA_via1_7
* cell instance $20375 r0 *1 40.375,71.19
X$20375 1895 VIA_via2_5
* cell instance $20376 r0 *1 38.475,71.19
X$20376 1895 VIA_via2_5
* cell instance $20377 r0 *1 38.475,72.03
X$20377 1895 VIA_via1_4
* cell instance $20378 r0 *1 69.255,71.75
X$20378 1896 VIA_via2_5
* cell instance $20379 r0 *1 68.115,71.75
X$20379 1896 VIA_via1_4
* cell instance $20380 r0 *1 68.115,71.75
X$20380 1896 VIA_via2_5
* cell instance $20381 r0 *1 69.445,73.57
X$20381 1896 VIA_via1_4
* cell instance $20382 r0 *1 68.115,73.01
X$20382 1897 VIA_via1_7
* cell instance $20383 r0 *1 68.115,72.03
X$20383 1897 VIA_via2_5
* cell instance $20384 r0 *1 66.405,72.03
X$20384 1897 VIA_via1_4
* cell instance $20385 r0 *1 66.405,72.03
X$20385 1897 VIA_via2_5
* cell instance $20386 r0 *1 52.725,71.19
X$20386 1898 VIA_via1_7
* cell instance $20387 r0 *1 50.255,71.47
X$20387 1898 VIA_via2_5
* cell instance $20388 r0 *1 52.725,71.47
X$20388 1898 VIA_via2_5
* cell instance $20389 r0 *1 50.255,72.03
X$20389 1898 VIA_via1_4
* cell instance $20390 r0 *1 54.055,72.03
X$20390 1899 VIA_via1_4
* cell instance $20391 r0 *1 53.865,72.03
X$20391 1899 VIA_via1_4
* cell instance $20392 r0 *1 65.645,72.03
X$20392 1900 VIA_via1_4
* cell instance $20393 r0 *1 65.645,72.03
X$20393 1900 VIA_via2_5
* cell instance $20394 r0 *1 63.935,72.03
X$20394 1900 VIA_via1_4
* cell instance $20395 r0 *1 63.935,72.03
X$20395 1900 VIA_via2_5
* cell instance $20396 r0 *1 62.415,73.01
X$20396 1901 VIA_via1_7
* cell instance $20397 r0 *1 62.415,72.03
X$20397 1901 VIA_via2_5
* cell instance $20398 r0 *1 60.325,72.03
X$20398 1901 VIA_via1_4
* cell instance $20399 r0 *1 60.325,72.03
X$20399 1901 VIA_via2_5
* cell instance $20400 r0 *1 3.895,77.63
X$20400 1902 VIA_via2_5
* cell instance $20401 r0 *1 3.515,77.63
X$20401 1902 VIA_via2_5
* cell instance $20402 r0 *1 13.965,79.17
X$20402 1902 VIA_via2_5
* cell instance $20403 r0 *1 7.505,77.91
X$20403 1902 VIA_via2_5
* cell instance $20404 r0 *1 9.595,77.77
X$20404 1902 VIA_via2_5
* cell instance $20405 r0 *1 9.595,79.31
X$20405 1902 VIA_via2_5
* cell instance $20406 r0 *1 3.515,80.43
X$20406 1902 VIA_via1_4
* cell instance $20407 r0 *1 3.895,76.37
X$20407 1902 VIA_via1_4
* cell instance $20408 r0 *1 3.705,81.97
X$20408 1902 VIA_via1_4
* cell instance $20409 r0 *1 5.035,77.63
X$20409 1902 VIA_via1_4
* cell instance $20410 r0 *1 5.035,77.63
X$20410 1902 VIA_via2_5
* cell instance $20411 r0 *1 13.015,79.17
X$20411 1902 VIA_via1_4
* cell instance $20412 r0 *1 13.015,79.17
X$20412 1902 VIA_via2_5
* cell instance $20413 r0 *1 8.265,77.63
X$20413 1902 VIA_via1_4
* cell instance $20414 r0 *1 8.265,77.77
X$20414 1902 VIA_via2_5
* cell instance $20415 r0 *1 7.505,78.75
X$20415 1902 VIA_via1_4
* cell instance $20416 r0 *1 14.155,83.23
X$20416 1902 VIA_via1_4
* cell instance $20417 r0 *1 9.975,73.57
X$20417 1902 VIA_via1_4
* cell instance $20418 r0 *1 11.875,73.85
X$20418 1903 VIA_via2_5
* cell instance $20419 r0 *1 10.165,73.85
X$20419 1903 VIA_via2_5
* cell instance $20420 r0 *1 10.165,74.83
X$20420 1903 VIA_via1_4
* cell instance $20421 r0 *1 11.495,73.85
X$20421 1903 VIA_via1_4
* cell instance $20422 r0 *1 11.495,73.85
X$20422 1903 VIA_via2_5
* cell instance $20423 r0 *1 11.875,73.57
X$20423 1903 VIA_via1_4
* cell instance $20424 r0 *1 19.095,72.59
X$20424 1904 VIA_via1_7
* cell instance $20425 r0 *1 20.235,73.57
X$20425 1904 VIA_via1_4
* cell instance $20426 r0 *1 30.685,73.85
X$20426 1905 VIA_via2_5
* cell instance $20427 r0 *1 28.975,73.85
X$20427 1905 VIA_via2_5
* cell instance $20428 r0 *1 28.975,73.43
X$20428 1905 VIA_via1_4
* cell instance $20429 r0 *1 20.995,73.85
X$20429 1905 VIA_via1_4
* cell instance $20430 r0 *1 20.995,73.85
X$20430 1905 VIA_via2_5
* cell instance $20431 r0 *1 30.685,73.57
X$20431 1905 VIA_via1_4
* cell instance $20432 r0 *1 31.065,73.29
X$20432 1906 VIA_via1_7
* cell instance $20433 r0 *1 30.685,70.77
X$20433 1906 VIA_via1_4
* cell instance $20434 r0 *1 30.305,74.41
X$20434 1907 VIA_via1_7
* cell instance $20435 r0 *1 31.445,74.83
X$20435 1907 VIA_via1_4
* cell instance $20436 r0 *1 32.965,73.99
X$20436 1908 VIA_via1_7
* cell instance $20437 r0 *1 33.155,74.83
X$20437 1908 VIA_via1_4
* cell instance $20438 r0 *1 25.745,77.21
X$20438 1909 VIA_via1_7
* cell instance $20439 r0 *1 25.745,77.21
X$20439 1909 VIA_via2_5
* cell instance $20440 r0 *1 33.915,75.67
X$20440 1909 VIA_via2_5
* cell instance $20441 r0 *1 29.165,87.85
X$20441 1909 VIA_via2_5
* cell instance $20442 r0 *1 29.165,77.21
X$20442 1909 VIA_via2_5
* cell instance $20443 r0 *1 28.785,77.21
X$20443 1909 VIA_via2_5
* cell instance $20444 r0 *1 29.165,75.81
X$20444 1909 VIA_via2_5
* cell instance $20445 r0 *1 25.745,75.67
X$20445 1909 VIA_via2_5
* cell instance $20446 r0 *1 32.205,87.85
X$20446 1909 VIA_via2_5
* cell instance $20447 r0 *1 8.075,79.17
X$20447 1909 VIA_via2_5
* cell instance $20448 r0 *1 15.105,79.03
X$20448 1909 VIA_via2_5
* cell instance $20449 r0 *1 19.095,75.67
X$20449 1909 VIA_via2_5
* cell instance $20450 r0 *1 42.845,84.77
X$20450 1909 VIA_via2_5
* cell instance $20451 r0 *1 22.515,87.85
X$20451 1909 VIA_via2_5
* cell instance $20452 r0 *1 15.105,87.57
X$20452 1909 VIA_via2_5
* cell instance $20453 r0 *1 15.105,91.63
X$20453 1909 VIA_via2_5
* cell instance $20454 r0 *1 43.415,84.77
X$20454 1909 VIA_via1_4
* cell instance $20455 r0 *1 43.415,84.77
X$20455 1909 VIA_via2_5
* cell instance $20456 r0 *1 13.965,91.63
X$20456 1909 VIA_via1_4
* cell instance $20457 r0 *1 13.965,91.63
X$20457 1909 VIA_via2_5
* cell instance $20458 r0 *1 22.515,87.57
X$20458 1909 VIA_via1_4
* cell instance $20459 r0 *1 22.515,87.57
X$20459 1909 VIA_via2_5
* cell instance $20460 r0 *1 32.015,95.97
X$20460 1909 VIA_via1_4
* cell instance $20461 r0 *1 42.465,91.63
X$20461 1909 VIA_via1_4
* cell instance $20462 r0 *1 29.165,83.23
X$20462 1909 VIA_via1_4
* cell instance $20463 r0 *1 8.075,86.03
X$20463 1909 VIA_via1_4
* cell instance $20464 r0 *1 19.095,74.83
X$20464 1909 VIA_via1_4
* cell instance $20465 r0 *1 6.745,79.17
X$20465 1909 VIA_via1_4
* cell instance $20466 r0 *1 6.745,79.17
X$20466 1909 VIA_via2_5
* cell instance $20467 r0 *1 33.725,73.57
X$20467 1909 VIA_via1_4
* cell instance $20468 r0 *1 33.975,77.63
X$20468 1909 VIA_via4_0
* cell instance $20469 r0 *1 40.135,77.63
X$20469 1909 VIA_via4_0
* cell instance $20470 r0 *1 40.135,77.63
X$20470 1909 VIA_via3_2
* cell instance $20471 r0 *1 40.185,77.63
X$20471 1909 VIA_via2_5
* cell instance $20472 r0 *1 40.185,77.63
X$20472 1909 VIA_via1_4
* cell instance $20473 r0 *1 40.415,84.77
X$20473 1909 VIA_via3_2
* cell instance $20474 r0 *1 33.975,75.81
X$20474 1909 VIA_via3_2
* cell instance $20475 r0 *1 37.335,72.59
X$20475 1910 VIA_via1_7
* cell instance $20476 r0 *1 37.335,72.59
X$20476 1910 VIA_via2_5
* cell instance $20477 r0 *1 34.105,72.59
X$20477 1910 VIA_via2_5
* cell instance $20478 r0 *1 34.295,76.37
X$20478 1910 VIA_via1_4
* cell instance $20479 r0 *1 34.295,71.19
X$20479 1911 VIA_via1_7
* cell instance $20480 r0 *1 34.485,76.37
X$20480 1911 VIA_via1_4
* cell instance $20481 r0 *1 42.085,72.03
X$20481 1912 VIA_via1_4
* cell instance $20482 r0 *1 42.275,73.15
X$20482 1912 VIA_via1_4
* cell instance $20483 r0 *1 42.655,73.57
X$20483 1912 VIA_via1_4
* cell instance $20484 r0 *1 66.785,73.15
X$20484 1913 VIA_via2_5
* cell instance $20485 r0 *1 64.885,73.15
X$20485 1913 VIA_via2_5
* cell instance $20486 r0 *1 67.165,73.15
X$20486 1913 VIA_via2_5
* cell instance $20487 r0 *1 64.885,72.03
X$20487 1913 VIA_via1_4
* cell instance $20488 r0 *1 67.165,73.57
X$20488 1913 VIA_via1_4
* cell instance $20489 r0 *1 66.785,73.57
X$20489 1913 VIA_via1_4
* cell instance $20490 r0 *1 71.725,73.71
X$20490 1914 VIA_via1_4
* cell instance $20491 r0 *1 71.725,73.71
X$20491 1914 VIA_via2_5
* cell instance $20492 r0 *1 67.735,72.03
X$20492 1914 VIA_via1_4
* cell instance $20493 r0 *1 67.735,73.57
X$20493 1914 VIA_via1_4
* cell instance $20494 r0 *1 67.735,73.71
X$20494 1914 VIA_via2_5
* cell instance $20495 r0 *1 65.265,76.51
X$20495 1915 VIA_via1_7
* cell instance $20496 r0 *1 65.265,76.37
X$20496 1915 VIA_via2_5
* cell instance $20497 r0 *1 69.065,73.57
X$20497 1915 VIA_via2_5
* cell instance $20498 r0 *1 59.945,76.37
X$20498 1915 VIA_via2_5
* cell instance $20499 r0 *1 63.175,76.37
X$20499 1915 VIA_via2_5
* cell instance $20500 r0 *1 59.755,76.37
X$20500 1915 VIA_via1_4
* cell instance $20501 r0 *1 59.755,76.37
X$20501 1915 VIA_via2_5
* cell instance $20502 r0 *1 65.645,76.37
X$20502 1915 VIA_via1_4
* cell instance $20503 r0 *1 65.645,76.37
X$20503 1915 VIA_via2_5
* cell instance $20504 r0 *1 69.065,69.23
X$20504 1915 VIA_via1_4
* cell instance $20505 r0 *1 63.175,80.43
X$20505 1915 VIA_via1_4
* cell instance $20506 r0 *1 70.205,73.57
X$20506 1915 VIA_via1_4
* cell instance $20507 r0 *1 70.205,73.57
X$20507 1915 VIA_via2_5
* cell instance $20508 r0 *1 65.265,73.57
X$20508 1915 VIA_via1_4
* cell instance $20509 r0 *1 65.265,73.57
X$20509 1915 VIA_via2_5
* cell instance $20510 r0 *1 59.945,80.43
X$20510 1915 VIA_via1_4
* cell instance $20511 r0 *1 80.085,73.85
X$20511 1916 VIA_via2_5
* cell instance $20512 r0 *1 84.075,73.71
X$20512 1916 VIA_via2_5
* cell instance $20513 r0 *1 81.415,73.71
X$20513 1916 VIA_via2_5
* cell instance $20514 r0 *1 80.085,72.03
X$20514 1916 VIA_via1_4
* cell instance $20515 r0 *1 84.265,73.29
X$20515 1916 VIA_via1_4
* cell instance $20516 r0 *1 81.415,72.03
X$20516 1916 VIA_via1_4
* cell instance $20517 r0 *1 84.455,79.17
X$20517 1917 VIA_via2_5
* cell instance $20518 r0 *1 84.265,73.57
X$20518 1917 VIA_via2_5
* cell instance $20519 r0 *1 84.075,79.17
X$20519 1917 VIA_via2_5
* cell instance $20520 r0 *1 84.265,83.23
X$20520 1917 VIA_via1_4
* cell instance $20521 r0 *1 88.445,73.57
X$20521 1917 VIA_via1_4
* cell instance $20522 r0 *1 88.445,73.57
X$20522 1917 VIA_via2_5
* cell instance $20523 r0 *1 82.745,73.57
X$20523 1917 VIA_via1_4
* cell instance $20524 r0 *1 82.745,73.57
X$20524 1917 VIA_via2_5
* cell instance $20525 r0 *1 79.515,73.57
X$20525 1917 VIA_via1_4
* cell instance $20526 r0 *1 79.515,73.57
X$20526 1917 VIA_via2_5
* cell instance $20527 r0 *1 84.265,77.35
X$20527 1917 VIA_via1_4
* cell instance $20528 r0 *1 84.835,77.63
X$20528 1917 VIA_via1_4
* cell instance $20529 r0 *1 82.555,79.17
X$20529 1917 VIA_via1_4
* cell instance $20530 r0 *1 82.555,79.17
X$20530 1917 VIA_via2_5
* cell instance $20531 r0 *1 85.785,79.17
X$20531 1917 VIA_via1_4
* cell instance $20532 r0 *1 85.785,79.17
X$20532 1917 VIA_via2_5
* cell instance $20533 r0 *1 86.735,73.99
X$20533 1918 VIA_via1_7
* cell instance $20534 r0 *1 86.925,74.83
X$20534 1918 VIA_via1_4
* cell instance $20535 r0 *1 87.305,74.41
X$20535 1919 VIA_via1_7
* cell instance $20536 r0 *1 87.685,73.57
X$20536 1919 VIA_via1_4
* cell instance $20537 r0 *1 89.965,73.15
X$20537 1920 VIA_via1_4
* cell instance $20538 r0 *1 89.015,72.03
X$20538 1920 VIA_via1_4
* cell instance $20539 r0 *1 94.905,72.87
X$20539 1921 VIA_via2_5
* cell instance $20540 r0 *1 94.905,72.03
X$20540 1921 VIA_via1_4
* cell instance $20541 r0 *1 97.815,72.87
X$20541 1921 VIA_via3_2
* cell instance $20542 r0 *1 97.815,72.87
X$20542 1921 VIA_via4_0
* cell instance $20543 r0 *1 13.205,73.99
X$20543 1922 VIA_via1_7
* cell instance $20544 r0 *1 13.205,73.99
X$20544 1922 VIA_via2_5
* cell instance $20545 r0 *1 12.065,73.99
X$20545 1922 VIA_via2_5
* cell instance $20546 r0 *1 12.065,74.83
X$20546 1922 VIA_via1_4
* cell instance $20547 r0 *1 17.195,73.01
X$20547 1923 VIA_via1_7
* cell instance $20548 r0 *1 17.195,73.01
X$20548 1923 VIA_via2_5
* cell instance $20549 r0 *1 13.585,73.01
X$20549 1923 VIA_via2_5
* cell instance $20550 r0 *1 13.585,72.03
X$20550 1923 VIA_via1_4
* cell instance $20551 r0 *1 13.015,73.57
X$20551 1924 VIA_via1_4
* cell instance $20552 r0 *1 12.825,73.57
X$20552 1924 VIA_via1_4
* cell instance $20553 r0 *1 20.045,77.21
X$20553 1925 VIA_via1_7
* cell instance $20554 r0 *1 19.665,73.57
X$20554 1925 VIA_via2_5
* cell instance $20555 r0 *1 20.995,73.57
X$20555 1925 VIA_via1_4
* cell instance $20556 r0 *1 20.995,73.57
X$20556 1925 VIA_via2_5
* cell instance $20557 r0 *1 26.315,72.59
X$20557 1926 VIA_via1_7
* cell instance $20558 r0 *1 26.315,73.57
X$20558 1926 VIA_via1_4
* cell instance $20559 r0 *1 29.355,74.13
X$20559 1927 VIA_via2_5
* cell instance $20560 r0 *1 13.015,74.13
X$20560 1927 VIA_via2_5
* cell instance $20561 r0 *1 13.015,74.55
X$20561 1927 VIA_via1_4
* cell instance $20562 r0 *1 29.355,73.57
X$20562 1927 VIA_via1_4
* cell instance $20563 r0 *1 29.355,73.57
X$20563 1927 VIA_via2_5
* cell instance $20564 r0 *1 30.875,73.57
X$20564 1927 VIA_via1_4
* cell instance $20565 r0 *1 30.875,73.57
X$20565 1927 VIA_via2_5
* cell instance $20566 r0 *1 32.015,73.43
X$20566 1928 VIA_via2_5
* cell instance $20567 r0 *1 32.395,74.83
X$20567 1928 VIA_via1_4
* cell instance $20568 r0 *1 30.495,73.43
X$20568 1928 VIA_via1_4
* cell instance $20569 r0 *1 30.495,73.43
X$20569 1928 VIA_via2_5
* cell instance $20570 r0 *1 73.055,73.57
X$20570 1929 VIA_via1_4
* cell instance $20571 r0 *1 73.055,73.43
X$20571 1929 VIA_via2_5
* cell instance $20572 r0 *1 76.665,73.43
X$20572 1929 VIA_via1_4
* cell instance $20573 r0 *1 76.665,73.43
X$20573 1929 VIA_via2_5
* cell instance $20574 r0 *1 43.035,72.59
X$20574 1930 VIA_via1_7
* cell instance $20575 r0 *1 43.035,72.59
X$20575 1930 VIA_via2_5
* cell instance $20576 r0 *1 39.995,72.59
X$20576 1930 VIA_via2_5
* cell instance $20577 r0 *1 39.995,73.57
X$20577 1930 VIA_via1_4
* cell instance $20578 r0 *1 65.265,72.59
X$20578 1931 VIA_via1_7
* cell instance $20579 r0 *1 65.265,72.59
X$20579 1931 VIA_via2_5
* cell instance $20580 r0 *1 64.505,72.59
X$20580 1931 VIA_via2_5
* cell instance $20581 r0 *1 64.505,73.57
X$20581 1931 VIA_via1_4
* cell instance $20582 r0 *1 45.885,73.43
X$20582 1932 VIA_via2_5
* cell instance $20583 r0 *1 45.885,74.83
X$20583 1932 VIA_via1_4
* cell instance $20584 r0 *1 43.605,73.43
X$20584 1932 VIA_via1_4
* cell instance $20585 r0 *1 43.605,73.43
X$20585 1932 VIA_via2_5
* cell instance $20586 r0 *1 40.565,76.51
X$20586 1933 VIA_via2_5
* cell instance $20587 r0 *1 40.755,76.09
X$20587 1933 VIA_via2_5
* cell instance $20588 r0 *1 40.375,80.43
X$20588 1933 VIA_via2_5
* cell instance $20589 r0 *1 44.175,73.57
X$20589 1933 VIA_via2_5
* cell instance $20590 r0 *1 40.565,77.35
X$20590 1933 VIA_via1_4
* cell instance $20591 r0 *1 40.565,78.05
X$20591 1933 VIA_via1_4
* cell instance $20592 r0 *1 40.375,79.17
X$20592 1933 VIA_via1_4
* cell instance $20593 r0 *1 37.715,83.23
X$20593 1933 VIA_via1_4
* cell instance $20594 r0 *1 37.525,80.43
X$20594 1933 VIA_via1_4
* cell instance $20595 r0 *1 37.525,80.43
X$20595 1933 VIA_via2_5
* cell instance $20596 r0 *1 40.755,74.83
X$20596 1933 VIA_via1_4
* cell instance $20597 r0 *1 40.755,74.83
X$20597 1933 VIA_via2_5
* cell instance $20598 r0 *1 35.815,74.83
X$20598 1933 VIA_via1_4
* cell instance $20599 r0 *1 35.815,74.83
X$20599 1933 VIA_via2_5
* cell instance $20600 r0 *1 44.175,77.63
X$20600 1933 VIA_via1_4
* cell instance $20601 r0 *1 40.755,73.57
X$20601 1933 VIA_via1_4
* cell instance $20602 r0 *1 40.755,73.57
X$20602 1933 VIA_via2_5
* cell instance $20603 r0 *1 47.405,73.57
X$20603 1933 VIA_via1_4
* cell instance $20604 r0 *1 47.405,73.57
X$20604 1933 VIA_via2_5
* cell instance $20605 r0 *1 53.105,71.19
X$20605 1934 VIA_via1_7
* cell instance $20606 r0 *1 53.105,72.59
X$20606 1934 VIA_via2_5
* cell instance $20607 r0 *1 54.245,72.59
X$20607 1934 VIA_via2_5
* cell instance $20608 r0 *1 54.245,74.83
X$20608 1934 VIA_via1_4
* cell instance $20609 r0 *1 1.995,72.59
X$20609 1935 VIA_via1_7
* cell instance $20610 r0 *1 10.355,76.37
X$20610 1935 VIA_via2_5
* cell instance $20611 r0 *1 11.305,77.63
X$20611 1935 VIA_via2_5
* cell instance $20612 r0 *1 2.565,76.09
X$20612 1935 VIA_via2_5
* cell instance $20613 r0 *1 3.135,76.09
X$20613 1935 VIA_via2_5
* cell instance $20614 r0 *1 5.795,76.09
X$20614 1935 VIA_via2_5
* cell instance $20615 r0 *1 3.895,83.23
X$20615 1935 VIA_via1_4
* cell instance $20616 r0 *1 3.895,83.09
X$20616 1935 VIA_via2_5
* cell instance $20617 r0 *1 2.565,83.23
X$20617 1935 VIA_via1_4
* cell instance $20618 r0 *1 2.565,83.09
X$20618 1935 VIA_via2_5
* cell instance $20619 r0 *1 10.355,80.43
X$20619 1935 VIA_via1_4
* cell instance $20620 r0 *1 3.135,74.83
X$20620 1935 VIA_via1_4
* cell instance $20621 r0 *1 5.795,76.37
X$20621 1935 VIA_via1_4
* cell instance $20622 r0 *1 5.795,76.37
X$20622 1935 VIA_via2_5
* cell instance $20623 r0 *1 11.305,76.37
X$20623 1935 VIA_via1_4
* cell instance $20624 r0 *1 11.305,76.37
X$20624 1935 VIA_via2_5
* cell instance $20625 r0 *1 12.065,77.63
X$20625 1935 VIA_via1_4
* cell instance $20626 r0 *1 12.065,77.63
X$20626 1935 VIA_via2_5
* cell instance $20627 r0 *1 17.195,74.83
X$20627 1936 VIA_via2_5
* cell instance $20628 r0 *1 15.485,74.83
X$20628 1936 VIA_via1_4
* cell instance $20629 r0 *1 15.485,74.83
X$20629 1936 VIA_via2_5
* cell instance $20630 r0 *1 17.195,75.95
X$20630 1936 VIA_via1_4
* cell instance $20631 r0 *1 17.765,74.83
X$20631 1936 VIA_via1_4
* cell instance $20632 r0 *1 17.765,74.83
X$20632 1936 VIA_via2_5
* cell instance $20633 r0 *1 18.145,76.65
X$20633 1937 VIA_via2_5
* cell instance $20634 r0 *1 18.145,77.63
X$20634 1937 VIA_via1_4
* cell instance $20635 r0 *1 20.425,76.65
X$20635 1937 VIA_via1_4
* cell instance $20636 r0 *1 20.425,76.65
X$20636 1937 VIA_via2_5
* cell instance $20637 r0 *1 18.335,74.83
X$20637 1937 VIA_via1_4
* cell instance $20638 r0 *1 18.715,74.83
X$20638 1938 VIA_via1_4
* cell instance $20639 r0 *1 18.715,74.83
X$20639 1938 VIA_via2_5
* cell instance $20640 r0 *1 20.045,74.83
X$20640 1938 VIA_via1_4
* cell instance $20641 r0 *1 20.045,74.69
X$20641 1938 VIA_via2_5
* cell instance $20642 r0 *1 24.985,75.11
X$20642 1939 VIA_via2_5
* cell instance $20643 r0 *1 24.035,75.11
X$20643 1939 VIA_via2_5
* cell instance $20644 r0 *1 24.985,76.37
X$20644 1939 VIA_via1_4
* cell instance $20645 r0 *1 24.035,74.83
X$20645 1939 VIA_via1_4
* cell instance $20646 r0 *1 23.655,75.25
X$20646 1939 VIA_via1_4
* cell instance $20647 r0 *1 25.365,75.81
X$20647 1940 VIA_via1_7
* cell instance $20648 r0 *1 26.315,74.83
X$20648 1940 VIA_via1_4
* cell instance $20649 r0 *1 26.315,75.11
X$20649 1941 VIA_via2_5
* cell instance $20650 r0 *1 26.505,74.83
X$20650 1941 VIA_via2_5
* cell instance $20651 r0 *1 26.315,76.37
X$20651 1941 VIA_via1_4
* cell instance $20652 r0 *1 26.505,73.43
X$20652 1941 VIA_via1_4
* cell instance $20653 r0 *1 31.635,74.83
X$20653 1942 VIA_via1_4
* cell instance $20654 r0 *1 31.635,74.83
X$20654 1942 VIA_via2_5
* cell instance $20655 r0 *1 29.545,74.97
X$20655 1942 VIA_via1_4
* cell instance $20656 r0 *1 29.545,74.97
X$20656 1942 VIA_via2_5
* cell instance $20657 r0 *1 34.105,74.55
X$20657 1943 VIA_via1_4
* cell instance $20658 r0 *1 34.105,74.55
X$20658 1943 VIA_via2_5
* cell instance $20659 r0 *1 32.205,74.83
X$20659 1943 VIA_via1_4
* cell instance $20660 r0 *1 32.205,74.83
X$20660 1943 VIA_via2_5
* cell instance $20661 r0 *1 37.905,74.83
X$20661 1944 VIA_via1_4
* cell instance $20662 r0 *1 37.905,74.69
X$20662 1944 VIA_via2_5
* cell instance $20663 r0 *1 38.665,76.37
X$20663 1944 VIA_via1_4
* cell instance $20664 r0 *1 38.095,76.37
X$20664 1944 VIA_via1_4
* cell instance $20665 r0 *1 37.335,74.69
X$20665 1944 VIA_via1_4
* cell instance $20666 r0 *1 37.335,74.69
X$20666 1944 VIA_via2_5
* cell instance $20667 r0 *1 43.035,75.39
X$20667 1945 VIA_via2_5
* cell instance $20668 r0 *1 43.415,76.65
X$20668 1945 VIA_via2_5
* cell instance $20669 r0 *1 43.415,75.39
X$20669 1945 VIA_via2_5
* cell instance $20670 r0 *1 42.085,76.65
X$20670 1945 VIA_via2_5
* cell instance $20671 r0 *1 41.895,78.75
X$20671 1945 VIA_via1_4
* cell instance $20672 r0 *1 42.845,74.83
X$20672 1945 VIA_via1_4
* cell instance $20673 r0 *1 43.035,74.83
X$20673 1945 VIA_via1_4
* cell instance $20674 r0 *1 43.415,76.37
X$20674 1945 VIA_via1_4
* cell instance $20675 r0 *1 48.925,79.45
X$20675 1946 VIA_via2_5
* cell instance $20676 r0 *1 50.255,79.45
X$20676 1946 VIA_via2_5
* cell instance $20677 r0 *1 51.585,79.45
X$20677 1946 VIA_via1_4
* cell instance $20678 r0 *1 51.585,79.45
X$20678 1946 VIA_via2_5
* cell instance $20679 r0 *1 49.495,74.83
X$20679 1946 VIA_via1_4
* cell instance $20680 r0 *1 48.925,80.43
X$20680 1946 VIA_via1_4
* cell instance $20681 r0 *1 54.435,75.11
X$20681 1947 VIA_via1_4
* cell instance $20682 r0 *1 55.005,76.37
X$20682 1947 VIA_via1_4
* cell instance $20683 r0 *1 55.005,77.63
X$20683 1947 VIA_via1_4
* cell instance $20684 r0 *1 58.425,76.51
X$20684 1948 VIA_via2_5
* cell instance $20685 r0 *1 56.525,76.37
X$20685 1948 VIA_via1_4
* cell instance $20686 r0 *1 56.525,76.51
X$20686 1948 VIA_via2_5
* cell instance $20687 r0 *1 56.715,73.85
X$20687 1948 VIA_via1_4
* cell instance $20688 r0 *1 56.905,74.83
X$20688 1948 VIA_via1_4
* cell instance $20689 r0 *1 58.425,77.63
X$20689 1948 VIA_via1_4
* cell instance $20690 r0 *1 81.415,75.95
X$20690 1949 VIA_via2_5
* cell instance $20691 r0 *1 88.065,85.05
X$20691 1949 VIA_via2_5
* cell instance $20692 r0 *1 85.975,75.95
X$20692 1949 VIA_via2_5
* cell instance $20693 r0 *1 46.455,75.95
X$20693 1949 VIA_via2_5
* cell instance $20694 r0 *1 83.505,89.25
X$20694 1949 VIA_via2_5
* cell instance $20695 r0 *1 71.535,82.39
X$20695 1949 VIA_via2_5
* cell instance $20696 r0 *1 84.455,85.05
X$20696 1949 VIA_via2_5
* cell instance $20697 r0 *1 84.455,84.07
X$20697 1949 VIA_via2_5
* cell instance $20698 r0 *1 81.795,83.93
X$20698 1949 VIA_via2_5
* cell instance $20699 r0 *1 81.795,82.39
X$20699 1949 VIA_via2_5
* cell instance $20700 r0 *1 63.745,86.31
X$20700 1949 VIA_via2_5
* cell instance $20701 r0 *1 88.255,89.25
X$20701 1949 VIA_via2_5
* cell instance $20702 r0 *1 71.535,86.31
X$20702 1949 VIA_via2_5
* cell instance $20703 r0 *1 71.535,83.23
X$20703 1949 VIA_via1_4
* cell instance $20704 r0 *1 81.795,80.43
X$20704 1949 VIA_via1_4
* cell instance $20705 r0 *1 84.455,84.77
X$20705 1949 VIA_via1_4
* cell instance $20706 r0 *1 83.505,88.83
X$20706 1949 VIA_via1_4
* cell instance $20707 r0 *1 88.065,86.03
X$20707 1949 VIA_via1_4
* cell instance $20708 r0 *1 88.255,88.83
X$20708 1949 VIA_via1_4
* cell instance $20709 r0 *1 79.515,75.95
X$20709 1949 VIA_via1_4
* cell instance $20710 r0 *1 79.515,75.95
X$20710 1949 VIA_via2_5
* cell instance $20711 r0 *1 63.745,87.57
X$20711 1949 VIA_via1_4
* cell instance $20712 r0 *1 85.975,74.83
X$20712 1949 VIA_via1_4
* cell instance $20713 r0 *1 85.975,74.69
X$20713 1949 VIA_via2_5
* cell instance $20714 r0 *1 87.685,74.83
X$20714 1949 VIA_via1_4
* cell instance $20715 r0 *1 87.685,74.69
X$20715 1949 VIA_via2_5
* cell instance $20716 r0 *1 46.455,72.03
X$20716 1949 VIA_via1_4
* cell instance $20717 r0 *1 46.855,75.95
X$20717 1949 VIA_via3_2
* cell instance $20718 r0 *1 46.855,86.31
X$20718 1949 VIA_via3_2
* cell instance $20719 r0 *1 3.705,74.83
X$20719 1950 VIA_via1_4
* cell instance $20720 r0 *1 3.705,74.83
X$20720 1950 VIA_via2_5
* cell instance $20721 r0 *1 5.415,74.83
X$20721 1950 VIA_via1_4
* cell instance $20722 r0 *1 5.415,74.83
X$20722 1950 VIA_via2_5
* cell instance $20723 r0 *1 5.415,75.95
X$20723 1950 VIA_via1_4
* cell instance $20724 r0 *1 81.795,75.53
X$20724 1951 VIA_via2_5
* cell instance $20725 r0 *1 81.795,74.83
X$20725 1951 VIA_via2_5
* cell instance $20726 r0 *1 81.225,75.53
X$20726 1951 VIA_via2_5
* cell instance $20727 r0 *1 80.085,75.53
X$20727 1951 VIA_via2_5
* cell instance $20728 r0 *1 65.835,83.09
X$20728 1951 VIA_via2_5
* cell instance $20729 r0 *1 74.195,84.07
X$20729 1951 VIA_via2_5
* cell instance $20730 r0 *1 79.135,84.07
X$20730 1951 VIA_via2_5
* cell instance $20731 r0 *1 80.085,84.07
X$20731 1951 VIA_via2_5
* cell instance $20732 r0 *1 65.835,81.97
X$20732 1951 VIA_via2_5
* cell instance $20733 r0 *1 61.845,82.11
X$20733 1951 VIA_via2_5
* cell instance $20734 r0 *1 61.845,74.83
X$20734 1951 VIA_via1_4
* cell instance $20735 r0 *1 67.545,81.97
X$20735 1951 VIA_via1_4
* cell instance $20736 r0 *1 67.545,81.83
X$20736 1951 VIA_via2_5
* cell instance $20737 r0 *1 80.085,80.43
X$20737 1951 VIA_via1_4
* cell instance $20738 r0 *1 74.195,83.23
X$20738 1951 VIA_via1_4
* cell instance $20739 r0 *1 74.195,83.09
X$20739 1951 VIA_via2_5
* cell instance $20740 r0 *1 79.135,86.17
X$20740 1951 VIA_via1_4
* cell instance $20741 r0 *1 79.135,86.03
X$20741 1951 VIA_via2_5
* cell instance $20742 r0 *1 80.275,86.03
X$20742 1951 VIA_via1_4
* cell instance $20743 r0 *1 80.275,86.03
X$20743 1951 VIA_via2_5
* cell instance $20744 r0 *1 83.125,86.03
X$20744 1951 VIA_via1_4
* cell instance $20745 r0 *1 83.125,86.03
X$20745 1951 VIA_via2_5
* cell instance $20746 r0 *1 65.455,86.03
X$20746 1951 VIA_via1_4
* cell instance $20747 r0 *1 81.225,77.63
X$20747 1951 VIA_via1_4
* cell instance $20748 r0 *1 84.645,74.83
X$20748 1951 VIA_via1_4
* cell instance $20749 r0 *1 84.645,74.83
X$20749 1951 VIA_via2_5
* cell instance $20750 r0 *1 81.795,76.37
X$20750 1951 VIA_via1_4
* cell instance $20751 r0 *1 11.115,74.41
X$20751 1952 VIA_via1_7
* cell instance $20752 r0 *1 11.115,74.41
X$20752 1952 VIA_via2_5
* cell instance $20753 r0 *1 9.215,74.41
X$20753 1952 VIA_via2_5
* cell instance $20754 r0 *1 9.215,73.57
X$20754 1952 VIA_via1_4
* cell instance $20755 r0 *1 74.575,95.97
X$20755 1953 VIA_via1_4
* cell instance $20756 r0 *1 74.575,95.97
X$20756 1953 VIA_via3_2
* cell instance $20757 r0 *1 74.575,95.97
X$20757 1953 VIA_via2_5
* cell instance $20758 r0 *1 76.855,86.03
X$20758 1953 VIA_via1_4
* cell instance $20759 r0 *1 76.855,86.03
X$20759 1953 VIA_via2_5
* cell instance $20760 r0 *1 73.625,74.83
X$20760 1953 VIA_via1_4
* cell instance $20761 r0 *1 73.625,74.83
X$20761 1953 VIA_via2_5
* cell instance $20762 r0 *1 75.135,74.83
X$20762 1953 VIA_via3_2
* cell instance $20763 r0 *1 75.135,86.03
X$20763 1953 VIA_via3_2
* cell instance $20764 r0 *1 74.575,86.03
X$20764 1953 VIA_via3_2
* cell instance $20765 r0 *1 6.365,74.83
X$20765 1954 VIA_via1_4
* cell instance $20766 r0 *1 6.365,74.83
X$20766 1954 VIA_via2_5
* cell instance $20767 r0 *1 11.305,74.83
X$20767 1954 VIA_via1_4
* cell instance $20768 r0 *1 11.305,74.83
X$20768 1954 VIA_via2_5
* cell instance $20769 r0 *1 11.495,74.97
X$20769 1955 VIA_via1_4
* cell instance $20770 r0 *1 11.495,74.97
X$20770 1955 VIA_via2_5
* cell instance $20771 r0 *1 13.015,74.83
X$20771 1955 VIA_via1_4
* cell instance $20772 r0 *1 13.015,74.97
X$20772 1955 VIA_via2_5
* cell instance $20773 r0 *1 58.045,77.21
X$20773 1956 VIA_via1_7
* cell instance $20774 r0 *1 57.855,74.97
X$20774 1956 VIA_via2_5
* cell instance $20775 r0 *1 54.815,74.83
X$20775 1956 VIA_via1_4
* cell instance $20776 r0 *1 54.815,74.97
X$20776 1956 VIA_via2_5
* cell instance $20777 r0 *1 56.525,74.83
X$20777 1957 VIA_via1_4
* cell instance $20778 r0 *1 56.525,74.83
X$20778 1957 VIA_via2_5
* cell instance $20779 r0 *1 57.095,74.83
X$20779 1957 VIA_via1_4
* cell instance $20780 r0 *1 57.095,74.83
X$20780 1957 VIA_via2_5
* cell instance $20781 r0 *1 54.435,74.69
X$20781 1958 VIA_via2_5
* cell instance $20782 r0 *1 56.335,74.69
X$20782 1958 VIA_via1_4
* cell instance $20783 r0 *1 56.335,74.69
X$20783 1958 VIA_via2_5
* cell instance $20784 r0 *1 54.435,73.57
X$20784 1958 VIA_via1_4
* cell instance $20785 r0 *1 24.985,74.69
X$20785 1959 VIA_via1_4
* cell instance $20786 r0 *1 24.985,74.69
X$20786 1959 VIA_via2_5
* cell instance $20787 r0 *1 21.375,74.83
X$20787 1959 VIA_via1_4
* cell instance $20788 r0 *1 21.375,74.69
X$20788 1959 VIA_via2_5
* cell instance $20789 r0 *1 55.195,74.83
X$20789 1960 VIA_via2_5
* cell instance $20790 r0 *1 53.485,79.87
X$20790 1960 VIA_via2_5
* cell instance $20791 r0 *1 52.345,74.83
X$20791 1960 VIA_via2_5
* cell instance $20792 r0 *1 52.345,79.73
X$20792 1960 VIA_via2_5
* cell instance $20793 r0 *1 50.065,79.73
X$20793 1960 VIA_via2_5
* cell instance $20794 r0 *1 50.065,79.17
X$20794 1960 VIA_via1_4
* cell instance $20795 r0 *1 55.195,73.57
X$20795 1960 VIA_via1_4
* cell instance $20796 r0 *1 51.965,86.03
X$20796 1960 VIA_via1_4
* cell instance $20797 r0 *1 55.385,83.23
X$20797 1960 VIA_via1_4
* cell instance $20798 r0 *1 55.385,83.23
X$20798 1960 VIA_via2_5
* cell instance $20799 r0 *1 52.915,84.77
X$20799 1960 VIA_via1_4
* cell instance $20800 r0 *1 52.155,74.83
X$20800 1960 VIA_via1_4
* cell instance $20801 r0 *1 52.155,74.83
X$20801 1960 VIA_via2_5
* cell instance $20802 r0 *1 53.485,80.15
X$20802 1960 VIA_via1_4
* cell instance $20803 r0 *1 53.485,81.97
X$20803 1960 VIA_via1_4
* cell instance $20804 r0 *1 53.105,83.23
X$20804 1960 VIA_via1_4
* cell instance $20805 r0 *1 53.105,83.23
X$20805 1960 VIA_via2_5
* cell instance $20806 r0 *1 48.165,74.83
X$20806 1961 VIA_via1_4
* cell instance $20807 r0 *1 48.165,74.83
X$20807 1961 VIA_via2_5
* cell instance $20808 r0 *1 48.925,73.85
X$20808 1961 VIA_via1_4
* cell instance $20809 r0 *1 48.925,74.83
X$20809 1961 VIA_via1_4
* cell instance $20810 r0 *1 48.925,74.83
X$20810 1961 VIA_via2_5
* cell instance $20811 r0 *1 48.545,74.41
X$20811 1962 VIA_via1_7
* cell instance $20812 r0 *1 48.545,74.41
X$20812 1962 VIA_via2_5
* cell instance $20813 r0 *1 46.645,74.41
X$20813 1962 VIA_via2_5
* cell instance $20814 r0 *1 46.645,73.57
X$20814 1962 VIA_via1_4
* cell instance $20815 r0 *1 33.725,74.83
X$20815 1963 VIA_via1_4
* cell instance $20816 r0 *1 33.725,74.97
X$20816 1963 VIA_via2_5
* cell instance $20817 r0 *1 33.915,76.65
X$20817 1963 VIA_via1_4
* cell instance $20818 r0 *1 34.105,77.63
X$20818 1963 VIA_via1_4
* cell instance $20819 r0 *1 30.305,74.83
X$20819 1963 VIA_via1_4
* cell instance $20820 r0 *1 30.305,74.97
X$20820 1963 VIA_via2_5
* cell instance $20821 r0 *1 43.225,74.83
X$20821 1964 VIA_via2_5
* cell instance $20822 r0 *1 42.275,74.83
X$20822 1964 VIA_via1_4
* cell instance $20823 r0 *1 42.275,74.83
X$20823 1964 VIA_via2_5
* cell instance $20824 r0 *1 43.795,74.83
X$20824 1964 VIA_via1_4
* cell instance $20825 r0 *1 43.795,74.83
X$20825 1964 VIA_via2_5
* cell instance $20826 r0 *1 43.225,73.57
X$20826 1964 VIA_via1_4
* cell instance $20827 r0 *1 39.995,74.83
X$20827 1965 VIA_via1_4
* cell instance $20828 r0 *1 39.995,74.69
X$20828 1965 VIA_via2_5
* cell instance $20829 r0 *1 44.745,74.69
X$20829 1965 VIA_via1_4
* cell instance $20830 r0 *1 44.745,74.69
X$20830 1965 VIA_via2_5
* cell instance $20831 r0 *1 37.335,76.09
X$20831 1966 VIA_via1_7
* cell instance $20832 r0 *1 37.335,74.97
X$20832 1966 VIA_via2_5
* cell instance $20833 r0 *1 35.055,74.83
X$20833 1966 VIA_via1_4
* cell instance $20834 r0 *1 35.055,74.97
X$20834 1966 VIA_via2_5
* cell instance $20835 r0 *1 4.085,75.39
X$20835 1967 VIA_via1_7
* cell instance $20836 r0 *1 3.135,76.37
X$20836 1967 VIA_via1_4
* cell instance $20837 r0 *1 5.985,74.83
X$20837 1968 VIA_via1_4
* cell instance $20838 r0 *1 6.365,76.37
X$20838 1968 VIA_via1_4
* cell instance $20839 r0 *1 6.555,77.35
X$20839 1968 VIA_via1_4
* cell instance $20840 r0 *1 18.335,77.77
X$20840 1969 VIA_via2_5
* cell instance $20841 r0 *1 19.095,77.77
X$20841 1969 VIA_via1_4
* cell instance $20842 r0 *1 19.095,77.77
X$20842 1969 VIA_via2_5
* cell instance $20843 r0 *1 18.145,76.37
X$20843 1969 VIA_via1_4
* cell instance $20844 r0 *1 20.615,77.21
X$20844 1970 VIA_via1_7
* cell instance $20845 r0 *1 20.805,73.57
X$20845 1970 VIA_via1_4
* cell instance $20846 r0 *1 26.695,76.23
X$20846 1971 VIA_via1_4
* cell instance $20847 r0 *1 26.695,76.23
X$20847 1971 VIA_via2_5
* cell instance $20848 r0 *1 28.975,76.23
X$20848 1971 VIA_via1_4
* cell instance $20849 r0 *1 28.975,76.23
X$20849 1971 VIA_via2_5
* cell instance $20850 r0 *1 28.785,74.83
X$20850 1971 VIA_via1_4
* cell instance $20851 r0 *1 29.355,79.59
X$20851 1972 VIA_via2_5
* cell instance $20852 r0 *1 19.855,79.59
X$20852 1972 VIA_via2_5
* cell instance $20853 r0 *1 20.045,90.09
X$20853 1972 VIA_via1_4
* cell instance $20854 r0 *1 29.355,76.37
X$20854 1972 VIA_via1_4
* cell instance $20855 r0 *1 28.975,74.83
X$20855 1972 VIA_via1_4
* cell instance $20856 r0 *1 33.155,75.39
X$20856 1973 VIA_via1_7
* cell instance $20857 r0 *1 32.775,92.33
X$20857 1973 VIA_via2_5
* cell instance $20858 r0 *1 31.635,92.33
X$20858 1973 VIA_via2_5
* cell instance $20859 r0 *1 31.445,95.97
X$20859 1973 VIA_via1_4
* cell instance $20860 r0 *1 42.465,78.61
X$20860 1974 VIA_via1_7
* cell instance $20861 r0 *1 42.465,78.61
X$20861 1974 VIA_via2_5
* cell instance $20862 r0 *1 40.945,78.61
X$20862 1974 VIA_via2_5
* cell instance $20863 r0 *1 40.725,76.405
X$20863 1974 VIA_via1_4
* cell instance $20864 r0 *1 42.655,75.39
X$20864 1975 VIA_via1_7
* cell instance $20865 r0 *1 42.465,76.37
X$20865 1975 VIA_via1_4
* cell instance $20866 r0 *1 50.445,76.37
X$20866 1976 VIA_via2_5
* cell instance $20867 r0 *1 50.445,77.63
X$20867 1976 VIA_via1_4
* cell instance $20868 r0 *1 51.015,76.37
X$20868 1976 VIA_via1_4
* cell instance $20869 r0 *1 51.015,76.37
X$20869 1976 VIA_via2_5
* cell instance $20870 r0 *1 48.545,76.09
X$20870 1976 VIA_via1_4
* cell instance $20871 r0 *1 48.545,76.09
X$20871 1976 VIA_via2_5
* cell instance $20872 r0 *1 53.485,76.37
X$20872 1977 VIA_via1_4
* cell instance $20873 r0 *1 53.485,76.23
X$20873 1977 VIA_via2_5
* cell instance $20874 r0 *1 53.675,75.25
X$20874 1977 VIA_via1_4
* cell instance $20875 r0 *1 52.535,76.37
X$20875 1977 VIA_via1_4
* cell instance $20876 r0 *1 52.535,76.23
X$20876 1977 VIA_via2_5
* cell instance $20877 r0 *1 53.675,76.37
X$20877 1977 VIA_via1_4
* cell instance $20878 r0 *1 54.815,75.81
X$20878 1978 VIA_via1_7
* cell instance $20879 r0 *1 55.005,74.83
X$20879 1978 VIA_via1_4
* cell instance $20880 r0 *1 57.665,74.83
X$20880 1979 VIA_via1_4
* cell instance $20881 r0 *1 57.665,76.37
X$20881 1979 VIA_via1_4
* cell instance $20882 r0 *1 57.665,76.23
X$20882 1979 VIA_via2_5
* cell instance $20883 r0 *1 61.275,76.23
X$20883 1979 VIA_via1_4
* cell instance $20884 r0 *1 61.275,76.23
X$20884 1979 VIA_via2_5
* cell instance $20885 r0 *1 71.345,86.59
X$20885 1980 VIA_via1_7
* cell instance $20886 r0 *1 71.345,88.83
X$20886 1980 VIA_via2_5
* cell instance $20887 r0 *1 69.445,76.37
X$20887 1980 VIA_via1_4
* cell instance $20888 r0 *1 69.635,88.83
X$20888 1980 VIA_via1_4
* cell instance $20889 r0 *1 69.635,88.83
X$20889 1980 VIA_via2_5
* cell instance $20890 r0 *1 74.385,81.97
X$20890 1981 VIA_via2_5
* cell instance $20891 r0 *1 73.055,83.23
X$20891 1981 VIA_via2_5
* cell instance $20892 r0 *1 70.965,83.23
X$20892 1981 VIA_via2_5
* cell instance $20893 r0 *1 70.965,81.97
X$20893 1981 VIA_via2_5
* cell instance $20894 r0 *1 74.385,83.23
X$20894 1981 VIA_via2_5
* cell instance $20895 r0 *1 70.205,76.37
X$20895 1981 VIA_via1_4
* cell instance $20896 r0 *1 71.345,77.63
X$20896 1981 VIA_via1_4
* cell instance $20897 r0 *1 70.775,79.17
X$20897 1981 VIA_via1_4
* cell instance $20898 r0 *1 69.065,83.23
X$20898 1981 VIA_via1_4
* cell instance $20899 r0 *1 69.065,83.23
X$20899 1981 VIA_via2_5
* cell instance $20900 r0 *1 71.915,81.97
X$20900 1981 VIA_via1_4
* cell instance $20901 r0 *1 71.915,81.97
X$20901 1981 VIA_via2_5
* cell instance $20902 r0 *1 76.855,84.77
X$20902 1981 VIA_via1_4
* cell instance $20903 r0 *1 74.385,82.25
X$20903 1981 VIA_via1_4
* cell instance $20904 r0 *1 76.665,81.97
X$20904 1981 VIA_via1_4
* cell instance $20905 r0 *1 76.665,81.97
X$20905 1981 VIA_via2_5
* cell instance $20906 r0 *1 73.055,86.03
X$20906 1981 VIA_via1_4
* cell instance $20907 r0 *1 71.915,76.37
X$20907 1982 VIA_via1_4
* cell instance $20908 r0 *1 72.295,78.75
X$20908 1982 VIA_via1_4
* cell instance $20909 r0 *1 79.895,76.37
X$20909 1983 VIA_via2_5
* cell instance $20910 r0 *1 78.755,76.37
X$20910 1983 VIA_via1_4
* cell instance $20911 r0 *1 78.755,76.37
X$20911 1983 VIA_via2_5
* cell instance $20912 r0 *1 79.135,79.17
X$20912 1983 VIA_via1_4
* cell instance $20913 r0 *1 79.135,76.37
X$20913 1983 VIA_via1_4
* cell instance $20914 r0 *1 79.135,76.37
X$20914 1983 VIA_via2_5
* cell instance $20915 r0 *1 79.895,77.63
X$20915 1983 VIA_via1_4
* cell instance $20916 r0 *1 80.275,76.37
X$20916 1983 VIA_via1_4
* cell instance $20917 r0 *1 80.275,76.37
X$20917 1983 VIA_via2_5
* cell instance $20918 r0 *1 72.105,80.57
X$20918 1984 VIA_via1_7
* cell instance $20919 r0 *1 72.105,80.71
X$20919 1984 VIA_via2_5
* cell instance $20920 r0 *1 70.015,80.57
X$20920 1984 VIA_via1_7
* cell instance $20921 r0 *1 70.015,80.71
X$20921 1984 VIA_via2_5
* cell instance $20922 r0 *1 71.345,85.89
X$20922 1984 VIA_via2_5
* cell instance $20923 r0 *1 80.655,85.89
X$20923 1984 VIA_via2_5
* cell instance $20924 r0 *1 86.355,85.61
X$20924 1984 VIA_via2_5
* cell instance $20925 r0 *1 71.155,80.71
X$20925 1984 VIA_via2_5
* cell instance $20926 r0 *1 80.655,85.61
X$20926 1984 VIA_via2_5
* cell instance $20927 r0 *1 80.655,86.17
X$20927 1984 VIA_via1_4
* cell instance $20928 r0 *1 70.205,86.03
X$20928 1984 VIA_via1_4
* cell instance $20929 r0 *1 70.205,85.89
X$20929 1984 VIA_via2_5
* cell instance $20930 r0 *1 87.305,74.83
X$20930 1984 VIA_via1_4
* cell instance $20931 r0 *1 96.615,76.37
X$20931 1985 VIA_via1_4
* cell instance $20932 r0 *1 96.615,75.25
X$20932 1985 VIA_via1_4
* cell instance $20933 r0 *1 96.235,76.37
X$20933 1985 VIA_via1_4
* cell instance $20934 r0 *1 94.335,76.09
X$20934 1986 VIA_via1_4
* cell instance $20935 r0 *1 94.335,74.83
X$20935 1986 VIA_via1_4
* cell instance $20936 r0 *1 58.615,75.39
X$20936 1987 VIA_via1_7
* cell instance $20937 r0 *1 58.615,75.39
X$20937 1987 VIA_via2_5
* cell instance $20938 r0 *1 54.435,75.39
X$20938 1987 VIA_via2_5
* cell instance $20939 r0 *1 54.435,76.37
X$20939 1987 VIA_via1_4
* cell instance $20940 r0 *1 16.435,75.39
X$20940 1988 VIA_via1_7
* cell instance $20941 r0 *1 16.435,75.39
X$20941 1988 VIA_via2_5
* cell instance $20942 r0 *1 14.915,75.39
X$20942 1988 VIA_via2_5
* cell instance $20943 r0 *1 14.915,76.37
X$20943 1988 VIA_via1_4
* cell instance $20944 r0 *1 56.335,75.81
X$20944 1989 VIA_via1_7
* cell instance $20945 r0 *1 56.335,75.81
X$20945 1989 VIA_via2_5
* cell instance $20946 r0 *1 55.765,75.81
X$20946 1989 VIA_via2_5
* cell instance $20947 r0 *1 55.765,74.83
X$20947 1989 VIA_via1_4
* cell instance $20948 r0 *1 55.955,76.09
X$20948 1990 VIA_via1_4
* cell instance $20949 r0 *1 55.955,74.83
X$20949 1990 VIA_via1_4
* cell instance $20950 r0 *1 20.995,75.11
X$20950 1991 VIA_via2_5
* cell instance $20951 r0 *1 20.235,75.11
X$20951 1991 VIA_via1_4
* cell instance $20952 r0 *1 20.235,75.11
X$20952 1991 VIA_via2_5
* cell instance $20953 r0 *1 20.995,76.37
X$20953 1991 VIA_via1_4
* cell instance $20954 r0 *1 21.755,73.99
X$20954 1992 VIA_via1_7
* cell instance $20955 r0 *1 21.755,75.81
X$20955 1992 VIA_via2_5
* cell instance $20956 r0 *1 20.805,75.81
X$20956 1992 VIA_via2_5
* cell instance $20957 r0 *1 20.805,76.37
X$20957 1992 VIA_via1_4
* cell instance $20958 r0 *1 53.865,75.11
X$20958 1993 VIA_via2_5
* cell instance $20959 r0 *1 51.395,75.11
X$20959 1993 VIA_via2_5
* cell instance $20960 r0 *1 51.395,74.83
X$20960 1993 VIA_via1_4
* cell instance $20961 r0 *1 54.245,77.49
X$20961 1993 VIA_via1_4
* cell instance $20962 r0 *1 49.875,75.39
X$20962 1994 VIA_via1_7
* cell instance $20963 r0 *1 49.875,75.53
X$20963 1994 VIA_via2_5
* cell instance $20964 r0 *1 49.305,75.53
X$20964 1994 VIA_via2_5
* cell instance $20965 r0 *1 49.305,76.37
X$20965 1994 VIA_via1_4
* cell instance $20966 r0 *1 49.115,75.95
X$20966 1995 VIA_via2_5
* cell instance $20967 r0 *1 49.685,75.95
X$20967 1995 VIA_via1_4
* cell instance $20968 r0 *1 49.685,75.95
X$20968 1995 VIA_via2_5
* cell instance $20969 r0 *1 49.115,76.37
X$20969 1995 VIA_via1_4
* cell instance $20970 r0 *1 48.355,75.11
X$20970 1996 VIA_via2_5
* cell instance $20971 r0 *1 46.075,75.11
X$20971 1996 VIA_via1_4
* cell instance $20972 r0 *1 46.075,75.11
X$20972 1996 VIA_via2_5
* cell instance $20973 r0 *1 48.355,76.37
X$20973 1996 VIA_via1_4
* cell instance $20974 r0 *1 36.385,76.09
X$20974 1997 VIA_via1_7
* cell instance $20975 r0 *1 36.385,75.81
X$20975 1997 VIA_via2_5
* cell instance $20976 r0 *1 37.715,75.81
X$20976 1997 VIA_via2_5
* cell instance $20977 r0 *1 37.335,76.37
X$20977 1997 VIA_via1_4
* cell instance $20978 r0 *1 41.325,75.11
X$20978 1998 VIA_via2_5
* cell instance $20979 r0 *1 39.995,75.11
X$20979 1998 VIA_via2_5
* cell instance $20980 r0 *1 39.995,76.37
X$20980 1998 VIA_via1_4
* cell instance $20981 r0 *1 41.325,72.31
X$20981 1998 VIA_via1_4
* cell instance $20982 r0 *1 37.715,75.39
X$20982 1999 VIA_via1_7
* cell instance $20983 r0 *1 37.715,75.39
X$20983 1999 VIA_via2_5
* cell instance $20984 r0 *1 37.145,75.39
X$20984 1999 VIA_via2_5
* cell instance $20985 r0 *1 37.145,76.37
X$20985 1999 VIA_via1_4
* cell instance $20986 r0 *1 8.455,77.35
X$20986 2000 VIA_via2_5
* cell instance $20987 r0 *1 8.455,76.37
X$20987 2000 VIA_via1_4
* cell instance $20988 r0 *1 10.165,77.63
X$20988 2000 VIA_via1_4
* cell instance $20989 r0 *1 9.785,77.35
X$20989 2000 VIA_via1_4
* cell instance $20990 r0 *1 9.785,77.35
X$20990 2000 VIA_via2_5
* cell instance $20991 r0 *1 21.375,77.21
X$20991 2001 VIA_via1_7
* cell instance $20992 r0 *1 21.565,76.37
X$20992 2001 VIA_via1_4
* cell instance $20993 r0 *1 24.795,77.35
X$20993 2002 VIA_via1_4
* cell instance $20994 r0 *1 22.895,76.37
X$20994 2002 VIA_via1_4
* cell instance $20995 r0 *1 22.895,76.37
X$20995 2002 VIA_via2_5
* cell instance $20996 r0 *1 24.415,76.37
X$20996 2002 VIA_via1_4
* cell instance $20997 r0 *1 24.415,76.37
X$20997 2002 VIA_via2_5
* cell instance $20998 r0 *1 26.125,77.21
X$20998 2003 VIA_via1_7
* cell instance $20999 r0 *1 27.075,76.37
X$20999 2003 VIA_via1_4
* cell instance $21000 r0 *1 27.075,77.21
X$21000 2004 VIA_via1_7
* cell instance $21001 r0 *1 27.265,76.37
X$21001 2004 VIA_via1_4
* cell instance $21002 r0 *1 27.835,77.49
X$21002 2005 VIA_via2_5
* cell instance $21003 r0 *1 29.165,77.63
X$21003 2005 VIA_via1_4
* cell instance $21004 r0 *1 29.165,77.49
X$21004 2005 VIA_via2_5
* cell instance $21005 r0 *1 27.835,76.37
X$21005 2005 VIA_via1_4
* cell instance $21006 r0 *1 27.835,76.51
X$21006 2005 VIA_via2_5
* cell instance $21007 r0 *1 21.185,76.51
X$21007 2005 VIA_via1_4
* cell instance $21008 r0 *1 21.185,76.51
X$21008 2005 VIA_via2_5
* cell instance $21009 r0 *1 35.245,76.37
X$21009 2006 VIA_via1_4
* cell instance $21010 r0 *1 34.865,77.35
X$21010 2006 VIA_via1_4
* cell instance $21011 r0 *1 35.815,76.37
X$21011 2007 VIA_via1_4
* cell instance $21012 r0 *1 35.815,76.51
X$21012 2007 VIA_via2_5
* cell instance $21013 r0 *1 34.675,76.51
X$21013 2007 VIA_via1_4
* cell instance $21014 r0 *1 34.675,76.51
X$21014 2007 VIA_via2_5
* cell instance $21015 r0 *1 36.005,77.63
X$21015 2007 VIA_via1_4
* cell instance $21016 r0 *1 36.195,88.55
X$21016 2008 VIA_via2_5
* cell instance $21017 r0 *1 36.005,76.37
X$21017 2008 VIA_via1_4
* cell instance $21018 r0 *1 36.385,77.63
X$21018 2008 VIA_via1_4
* cell instance $21019 r0 *1 33.535,88.55
X$21019 2008 VIA_via1_4
* cell instance $21020 r0 *1 33.535,88.55
X$21020 2008 VIA_via2_5
* cell instance $21021 r0 *1 38.095,77.21
X$21021 2009 VIA_via1_7
* cell instance $21022 r0 *1 38.285,76.37
X$21022 2009 VIA_via2_5
* cell instance $21023 r0 *1 40.945,76.37
X$21023 2009 VIA_via1_4
* cell instance $21024 r0 *1 40.945,76.37
X$21024 2009 VIA_via2_5
* cell instance $21025 r0 *1 32.585,79.59
X$21025 2010 VIA_via2_5
* cell instance $21026 r0 *1 38.855,79.59
X$21026 2010 VIA_via2_5
* cell instance $21027 r0 *1 52.535,79.03
X$21027 2010 VIA_via2_5
* cell instance $21028 r0 *1 49.685,77.77
X$21028 2010 VIA_via2_5
* cell instance $21029 r0 *1 52.535,77.63
X$21029 2010 VIA_via1_4
* cell instance $21030 r0 *1 52.535,77.77
X$21030 2010 VIA_via2_5
* cell instance $21031 r0 *1 55.385,79.03
X$21031 2010 VIA_via1_4
* cell instance $21032 r0 *1 55.385,79.03
X$21032 2010 VIA_via2_5
* cell instance $21033 r0 *1 38.855,77.63
X$21033 2010 VIA_via1_4
* cell instance $21034 r0 *1 38.855,77.49
X$21034 2010 VIA_via2_5
* cell instance $21035 r0 *1 43.225,77.63
X$21035 2010 VIA_via1_4
* cell instance $21036 r0 *1 43.225,77.63
X$21036 2010 VIA_via2_5
* cell instance $21037 r0 *1 47.025,77.63
X$21037 2010 VIA_via1_4
* cell instance $21038 r0 *1 47.025,77.63
X$21038 2010 VIA_via2_5
* cell instance $21039 r0 *1 49.685,77.35
X$21039 2010 VIA_via1_4
* cell instance $21040 r0 *1 32.585,80.57
X$21040 2010 VIA_via1_4
* cell instance $21041 r0 *1 39.045,76.79
X$21041 2011 VIA_via1_7
* cell instance $21042 r0 *1 39.235,77.63
X$21042 2011 VIA_via1_4
* cell instance $21043 r0 *1 41.135,77.63
X$21043 2012 VIA_via1_4
* cell instance $21044 r0 *1 40.945,76.65
X$21044 2012 VIA_via1_4
* cell instance $21045 r0 *1 41.135,76.37
X$21045 2012 VIA_via1_4
* cell instance $21046 r0 *1 41.515,77.63
X$21046 2013 VIA_via1_4
* cell instance $21047 r0 *1 41.325,76.37
X$21047 2013 VIA_via1_4
* cell instance $21048 r0 *1 40.945,90.09
X$21048 2013 VIA_via1_4
* cell instance $21049 r0 *1 39.615,78.33
X$21049 2014 VIA_via2_5
* cell instance $21050 r0 *1 42.465,78.33
X$21050 2014 VIA_via2_5
* cell instance $21051 r0 *1 39.615,79.17
X$21051 2014 VIA_via1_4
* cell instance $21052 r0 *1 43.035,76.51
X$21052 2014 VIA_via1_4
* cell instance $21053 r0 *1 50.065,76.79
X$21053 2015 VIA_via1_7
* cell instance $21054 r0 *1 48.925,76.65
X$21054 2015 VIA_via2_5
* cell instance $21055 r0 *1 49.875,76.65
X$21055 2015 VIA_via2_5
* cell instance $21056 r0 *1 48.925,76.37
X$21056 2015 VIA_via1_4
* cell instance $21057 r0 *1 51.205,76.37
X$21057 2016 VIA_via1_4
* cell instance $21058 r0 *1 50.825,77.63
X$21058 2016 VIA_via1_4
* cell instance $21059 r0 *1 51.015,91.49
X$21059 2016 VIA_via1_4
* cell instance $21060 r0 *1 53.485,76.79
X$21060 2017 VIA_via1_7
* cell instance $21061 r0 *1 53.675,77.63
X$21061 2017 VIA_via1_4
* cell instance $21062 r0 *1 54.055,76.79
X$21062 2018 VIA_via1_7
* cell instance $21063 r0 *1 54.435,77.63
X$21063 2018 VIA_via1_4
* cell instance $21064 r0 *1 55.385,77.63
X$21064 2019 VIA_via1_4
* cell instance $21065 r0 *1 55.195,76.37
X$21065 2019 VIA_via1_4
* cell instance $21066 r0 *1 55.575,85.89
X$21066 2019 VIA_via1_4
* cell instance $21067 r0 *1 58.425,80.15
X$21067 2020 VIA_via2_5
* cell instance $21068 r0 *1 58.235,74.83
X$21068 2020 VIA_via1_4
* cell instance $21069 r0 *1 61.465,80.15
X$21069 2020 VIA_via1_4
* cell instance $21070 r0 *1 61.465,80.15
X$21070 2020 VIA_via2_5
* cell instance $21071 r0 *1 58.425,81.97
X$21071 2020 VIA_via1_4
* cell instance $21072 r0 *1 72.865,77.49
X$21072 2021 VIA_via1_4
* cell instance $21073 r0 *1 72.865,77.49
X$21073 2021 VIA_via2_5
* cell instance $21074 r0 *1 66.785,77.63
X$21074 2021 VIA_via1_4
* cell instance $21075 r0 *1 66.785,77.63
X$21075 2021 VIA_via2_5
* cell instance $21076 r0 *1 87.495,77.77
X$21076 2022 VIA_via2_5
* cell instance $21077 r0 *1 96.045,80.43
X$21077 2022 VIA_via1_4
* cell instance $21078 r0 *1 96.045,80.29
X$21078 2022 VIA_via2_5
* cell instance $21079 r0 *1 89.965,80.43
X$21079 2022 VIA_via1_4
* cell instance $21080 r0 *1 89.965,80.29
X$21080 2022 VIA_via2_5
* cell instance $21081 r0 *1 88.825,80.43
X$21081 2022 VIA_via1_4
* cell instance $21082 r0 *1 88.825,80.29
X$21082 2022 VIA_via2_5
* cell instance $21083 r0 *1 88.825,79.17
X$21083 2022 VIA_via1_4
* cell instance $21084 r0 *1 88.825,79.17
X$21084 2022 VIA_via2_5
* cell instance $21085 r0 *1 87.495,79.17
X$21085 2022 VIA_via1_4
* cell instance $21086 r0 *1 87.495,79.17
X$21086 2022 VIA_via2_5
* cell instance $21087 r0 *1 86.735,77.63
X$21087 2022 VIA_via1_4
* cell instance $21088 r0 *1 86.735,77.63
X$21088 2022 VIA_via2_5
* cell instance $21089 r0 *1 88.635,78.89
X$21089 2023 VIA_via1_7
* cell instance $21090 r0 *1 94.715,77.49
X$21090 2023 VIA_via2_5
* cell instance $21091 r0 *1 88.445,77.35
X$21091 2023 VIA_via2_5
* cell instance $21092 r0 *1 94.905,80.43
X$21092 2023 VIA_via1_4
* cell instance $21093 r0 *1 88.635,80.43
X$21093 2023 VIA_via1_4
* cell instance $21094 r0 *1 88.635,80.43
X$21094 2023 VIA_via2_5
* cell instance $21095 r0 *1 90.155,80.43
X$21095 2023 VIA_via1_4
* cell instance $21096 r0 *1 90.155,80.43
X$21096 2023 VIA_via2_5
* cell instance $21097 r0 *1 88.445,76.37
X$21097 2023 VIA_via1_4
* cell instance $21098 r0 *1 92.625,77.49
X$21098 2023 VIA_via1_4
* cell instance $21099 r0 *1 92.625,77.49
X$21099 2023 VIA_via2_5
* cell instance $21100 r0 *1 89.015,76.79
X$21100 2024 VIA_via1_7
* cell instance $21101 r0 *1 88.825,77.63
X$21101 2024 VIA_via1_4
* cell instance $21102 r0 *1 88.065,77.77
X$21102 2025 VIA_via1_7
* cell instance $21103 r0 *1 88.065,77.91
X$21103 2025 VIA_via2_5
* cell instance $21104 r0 *1 85.405,78.75
X$21104 2025 VIA_via2_5
* cell instance $21105 r0 *1 82.935,78.75
X$21105 2025 VIA_via2_5
* cell instance $21106 r0 *1 85.405,77.91
X$21106 2025 VIA_via2_5
* cell instance $21107 r0 *1 94.335,77.91
X$21107 2025 VIA_via2_5
* cell instance $21108 r0 *1 82.935,81.83
X$21108 2025 VIA_via1_4
* cell instance $21109 r0 *1 85.405,77.63
X$21109 2025 VIA_via1_4
* cell instance $21110 r0 *1 94.525,80.43
X$21110 2025 VIA_via1_4
* cell instance $21111 r0 *1 94.525,76.37
X$21111 2025 VIA_via1_4
* cell instance $21112 r0 *1 95.095,81.97
X$21112 2026 VIA_via2_5
* cell instance $21113 r0 *1 94.905,77.63
X$21113 2026 VIA_via2_5
* cell instance $21114 r0 *1 95.095,77.63
X$21114 2026 VIA_via2_5
* cell instance $21115 r0 *1 94.905,81.97
X$21115 2026 VIA_via2_5
* cell instance $21116 r0 *1 94.145,87.57
X$21116 2026 VIA_via2_5
* cell instance $21117 r0 *1 89.965,87.57
X$21117 2026 VIA_via1_4
* cell instance $21118 r0 *1 89.965,87.57
X$21118 2026 VIA_via2_5
* cell instance $21119 r0 *1 94.335,81.97
X$21119 2026 VIA_via1_4
* cell instance $21120 r0 *1 94.335,81.97
X$21120 2026 VIA_via2_5
* cell instance $21121 r0 *1 94.525,81.97
X$21121 2026 VIA_via1_4
* cell instance $21122 r0 *1 94.525,81.97
X$21122 2026 VIA_via2_5
* cell instance $21123 r0 *1 94.905,83.23
X$21123 2026 VIA_via1_4
* cell instance $21124 r0 *1 94.145,84.77
X$21124 2026 VIA_via1_4
* cell instance $21125 r0 *1 94.525,77.63
X$21125 2026 VIA_via1_4
* cell instance $21126 r0 *1 94.525,77.63
X$21126 2026 VIA_via2_5
* cell instance $21127 r0 *1 90.915,77.63
X$21127 2026 VIA_via1_4
* cell instance $21128 r0 *1 90.915,77.63
X$21128 2026 VIA_via2_5
* cell instance $21129 r0 *1 95.095,74.83
X$21129 2026 VIA_via1_4
* cell instance $21130 r0 *1 94.905,79.17
X$21130 2026 VIA_via1_4
* cell instance $21131 r0 *1 96.805,77.21
X$21131 2027 VIA_via1_7
* cell instance $21132 r0 *1 95.855,76.37
X$21132 2027 VIA_via1_4
* cell instance $21133 r0 *1 96.995,76.79
X$21133 2028 VIA_via1_7
* cell instance $21134 r0 *1 96.995,76.79
X$21134 2028 VIA_via2_5
* cell instance $21135 r0 *1 97.255,77.35
X$21135 2028 VIA_via4_0
* cell instance $21136 r0 *1 97.255,76.79
X$21136 2028 VIA_via3_2
* cell instance $21137 r0 *1 6.745,76.79
X$21137 2029 VIA_via1_7
* cell instance $21138 r0 *1 6.745,76.79
X$21138 2029 VIA_via2_5
* cell instance $21139 r0 *1 4.275,76.79
X$21139 2029 VIA_via2_5
* cell instance $21140 r0 *1 4.275,77.63
X$21140 2029 VIA_via1_4
* cell instance $21141 r0 *1 94.145,76.37
X$21141 2030 VIA_via1_4
* cell instance $21142 r0 *1 94.145,76.37
X$21142 2030 VIA_via2_5
* cell instance $21143 r0 *1 96.045,76.37
X$21143 2030 VIA_via1_4
* cell instance $21144 r0 *1 96.045,76.37
X$21144 2030 VIA_via2_5
* cell instance $21145 r0 *1 8.835,76.79
X$21145 2031 VIA_via1_7
* cell instance $21146 r0 *1 8.835,76.79
X$21146 2031 VIA_via2_5
* cell instance $21147 r0 *1 7.505,76.79
X$21147 2031 VIA_via2_5
* cell instance $21148 r0 *1 7.505,77.63
X$21148 2031 VIA_via1_4
* cell instance $21149 r0 *1 86.165,77.63
X$21149 2032 VIA_via1_4
* cell instance $21150 r0 *1 86.165,77.49
X$21150 2032 VIA_via2_5
* cell instance $21151 r0 *1 87.305,77.49
X$21151 2032 VIA_via1_4
* cell instance $21152 r0 *1 87.305,77.49
X$21152 2032 VIA_via2_5
* cell instance $21153 r0 *1 16.435,77.49
X$21153 2033 VIA_via2_5
* cell instance $21154 r0 *1 17.385,77.63
X$21154 2033 VIA_via1_4
* cell instance $21155 r0 *1 17.385,77.49
X$21155 2033 VIA_via2_5
* cell instance $21156 r0 *1 16.435,78.05
X$21156 2033 VIA_via1_4
* cell instance $21157 r0 *1 16.245,79.17
X$21157 2033 VIA_via1_4
* cell instance $21158 r0 *1 58.045,76.37
X$21158 2034 VIA_via1_4
* cell instance $21159 r0 *1 58.045,76.37
X$21159 2034 VIA_via2_5
* cell instance $21160 r0 *1 58.995,76.37
X$21160 2034 VIA_via1_4
* cell instance $21161 r0 *1 58.995,76.37
X$21161 2034 VIA_via2_5
* cell instance $21162 r0 *1 21.755,77.07
X$21162 2035 VIA_via2_5
* cell instance $21163 r0 *1 19.475,77.07
X$21163 2035 VIA_via2_5
* cell instance $21164 r0 *1 21.755,76.37
X$21164 2035 VIA_via1_4
* cell instance $21165 r0 *1 19.475,78.89
X$21165 2035 VIA_via1_4
* cell instance $21166 r0 *1 23.845,76.79
X$21166 2036 VIA_via1_7
* cell instance $21167 r0 *1 23.845,76.79
X$21167 2036 VIA_via2_5
* cell instance $21168 r0 *1 22.515,76.79
X$21168 2036 VIA_via2_5
* cell instance $21169 r0 *1 22.515,77.63
X$21169 2036 VIA_via1_4
* cell instance $21170 r0 *1 26.505,75.11
X$21170 2037 VIA_via1_4
* cell instance $21171 r0 *1 26.505,76.37
X$21171 2037 VIA_via1_4
* cell instance $21172 r0 *1 31.635,75.11
X$21172 2038 VIA_via1_7
* cell instance $21173 r0 *1 31.635,76.37
X$21173 2038 VIA_via1_4
* cell instance $21174 r0 *1 31.065,78.61
X$21174 2039 VIA_via2_5
* cell instance $21175 r0 *1 30.495,78.61
X$21175 2039 VIA_via2_5
* cell instance $21176 r0 *1 30.685,76.51
X$21176 2039 VIA_via2_5
* cell instance $21177 r0 *1 31.065,79.17
X$21177 2039 VIA_via1_4
* cell instance $21178 r0 *1 28.595,76.51
X$21178 2039 VIA_via1_4
* cell instance $21179 r0 *1 28.595,76.51
X$21179 2039 VIA_via2_5
* cell instance $21180 r0 *1 35.625,77.21
X$21180 2040 VIA_via1_7
* cell instance $21181 r0 *1 35.625,76.37
X$21181 2040 VIA_via2_5
* cell instance $21182 r0 *1 35.055,76.37
X$21182 2040 VIA_via1_4
* cell instance $21183 r0 *1 35.055,76.37
X$21183 2040 VIA_via2_5
* cell instance $21184 r0 *1 38.475,76.79
X$21184 2041 VIA_via1_7
* cell instance $21185 r0 *1 38.475,76.93
X$21185 2041 VIA_via2_5
* cell instance $21186 r0 *1 37.905,76.93
X$21186 2041 VIA_via2_5
* cell instance $21187 r0 *1 37.905,76.37
X$21187 2041 VIA_via1_4
* cell instance $21188 r0 *1 43.225,75.39
X$21188 2042 VIA_via1_7
* cell instance $21189 r0 *1 43.225,76.37
X$21189 2042 VIA_via1_4
* cell instance $21190 r0 *1 41.895,76.37
X$21190 2043 VIA_via1_4
* cell instance $21191 r0 *1 41.895,76.37
X$21191 2043 VIA_via2_5
* cell instance $21192 r0 *1 42.655,76.37
X$21192 2043 VIA_via1_4
* cell instance $21193 r0 *1 42.655,76.37
X$21193 2043 VIA_via2_5
* cell instance $21194 r0 *1 48.355,78.61
X$21194 2044 VIA_via1_7
* cell instance $21195 r0 *1 48.545,76.37
X$21195 2044 VIA_via2_5
* cell instance $21196 r0 *1 49.875,76.37
X$21196 2044 VIA_via1_4
* cell instance $21197 r0 *1 49.875,76.37
X$21197 2044 VIA_via2_5
* cell instance $21198 r0 *1 7.695,84.07
X$21198 2045 VIA_via2_5
* cell instance $21199 r0 *1 8.265,88.83
X$21199 2045 VIA_via2_5
* cell instance $21200 r0 *1 7.125,88.83
X$21200 2045 VIA_via2_5
* cell instance $21201 r0 *1 3.895,88.83
X$21201 2045 VIA_via2_5
* cell instance $21202 r0 *1 8.835,84.07
X$21202 2045 VIA_via2_5
* cell instance $21203 r0 *1 9.595,85.89
X$21203 2045 VIA_via2_5
* cell instance $21204 r0 *1 7.695,85.89
X$21204 2045 VIA_via2_5
* cell instance $21205 r0 *1 9.595,84.77
X$21205 2045 VIA_via1_4
* cell instance $21206 r0 *1 7.695,83.23
X$21206 2045 VIA_via1_4
* cell instance $21207 r0 *1 3.895,87.57
X$21207 2045 VIA_via1_4
* cell instance $21208 r0 *1 8.455,86.03
X$21208 2045 VIA_via1_4
* cell instance $21209 r0 *1 8.455,85.89
X$21209 2045 VIA_via2_5
* cell instance $21210 r0 *1 7.125,87.57
X$21210 2045 VIA_via1_4
* cell instance $21211 r0 *1 6.745,91.63
X$21211 2045 VIA_via1_4
* cell instance $21212 r0 *1 10.545,86.03
X$21212 2045 VIA_via1_4
* cell instance $21213 r0 *1 10.545,85.89
X$21213 2045 VIA_via2_5
* cell instance $21214 r0 *1 8.835,88.83
X$21214 2045 VIA_via1_4
* cell instance $21215 r0 *1 8.835,88.83
X$21215 2045 VIA_via2_5
* cell instance $21216 r0 *1 9.215,79.17
X$21216 2045 VIA_via1_4
* cell instance $21217 r0 *1 10.925,80.43
X$21217 2046 VIA_via1_4
* cell instance $21218 r0 *1 10.735,77.63
X$21218 2046 VIA_via1_4
* cell instance $21219 r0 *1 10.735,79.45
X$21219 2046 VIA_via1_4
* cell instance $21220 r0 *1 12.635,78.75
X$21220 2047 VIA_via2_5
* cell instance $21221 r0 *1 16.815,78.75
X$21221 2047 VIA_via2_5
* cell instance $21222 r0 *1 14.535,78.75
X$21222 2047 VIA_via1_4
* cell instance $21223 r0 *1 14.535,78.75
X$21223 2047 VIA_via2_5
* cell instance $21224 r0 *1 12.635,77.63
X$21224 2047 VIA_via1_4
* cell instance $21225 r0 *1 16.815,79.17
X$21225 2047 VIA_via1_4
* cell instance $21226 r0 *1 17.195,78.61
X$21226 2048 VIA_via1_7
* cell instance $21227 r0 *1 17.195,78.61
X$21227 2048 VIA_via2_5
* cell instance $21228 r0 *1 20.045,78.61
X$21228 2048 VIA_via2_5
* cell instance $21229 r0 *1 19.855,77.63
X$21229 2048 VIA_via1_4
* cell instance $21230 r0 *1 26.695,80.01
X$21230 2049 VIA_via1_7
* cell instance $21231 r0 *1 26.885,77.63
X$21231 2049 VIA_via1_4
* cell instance $21232 r0 *1 33.345,79.17
X$21232 2050 VIA_via1_4
* cell instance $21233 r0 *1 33.345,79.03
X$21233 2050 VIA_via2_5
* cell instance $21234 r0 *1 33.345,79.31
X$21234 2050 VIA_via2_5
* cell instance $21235 r0 *1 30.495,79.17
X$21235 2050 VIA_via1_4
* cell instance $21236 r0 *1 30.495,79.31
X$21236 2050 VIA_via2_5
* cell instance $21237 r0 *1 33.915,79.17
X$21237 2050 VIA_via1_4
* cell instance $21238 r0 *1 33.915,79.03
X$21238 2050 VIA_via2_5
* cell instance $21239 r0 *1 33.915,78.05
X$21239 2050 VIA_via1_4
* cell instance $21240 r0 *1 35.625,80.01
X$21240 2051 VIA_via1_7
* cell instance $21241 r0 *1 35.435,77.63
X$21241 2051 VIA_via1_4
* cell instance $21242 r0 *1 43.035,77.91
X$21242 2052 VIA_via1_7
* cell instance $21243 r0 *1 42.275,94.43
X$21243 2052 VIA_via1_4
* cell instance $21244 r0 *1 55.385,78.19
X$21244 2053 VIA_via1_7
* cell instance $21245 r0 *1 55.005,79.17
X$21245 2053 VIA_via1_4
* cell instance $21246 r0 *1 56.525,80.01
X$21246 2054 VIA_via1_7
* cell instance $21247 r0 *1 56.715,77.63
X$21247 2054 VIA_via2_5
* cell instance $21248 r0 *1 57.855,77.63
X$21248 2054 VIA_via1_4
* cell instance $21249 r0 *1 57.855,77.63
X$21249 2054 VIA_via2_5
* cell instance $21250 r0 *1 65.455,80.15
X$21250 2055 VIA_via1_7
* cell instance $21251 r0 *1 65.455,80.15
X$21251 2055 VIA_via2_5
* cell instance $21252 r0 *1 67.545,80.15
X$21252 2055 VIA_via2_5
* cell instance $21253 r0 *1 67.735,79.17
X$21253 2055 VIA_via1_4
* cell instance $21254 r0 *1 73.245,81.69
X$21254 2056 VIA_via1_7
* cell instance $21255 r0 *1 73.435,79.17
X$21255 2056 VIA_via1_4
* cell instance $21256 r0 *1 79.515,92.61
X$21256 2057 VIA_via1_7
* cell instance $21257 r0 *1 79.515,93.59
X$21257 2057 VIA_via1_7
* cell instance $21258 r0 *1 85.785,92.47
X$21258 2057 VIA_via2_5
* cell instance $21259 r0 *1 88.255,92.19
X$21259 2057 VIA_via2_5
* cell instance $21260 r0 *1 86.925,79.87
X$21260 2057 VIA_via2_5
* cell instance $21261 r0 *1 79.515,92.19
X$21261 2057 VIA_via2_5
* cell instance $21262 r0 *1 70.585,79.73
X$21262 2057 VIA_via2_5
* cell instance $21263 r0 *1 67.925,79.73
X$21263 2057 VIA_via2_5
* cell instance $21264 r0 *1 70.965,84.63
X$21264 2057 VIA_via2_5
* cell instance $21265 r0 *1 69.825,84.63
X$21265 2057 VIA_via2_5
* cell instance $21266 r0 *1 69.445,90.37
X$21266 2057 VIA_via2_5
* cell instance $21267 r0 *1 83.695,92.19
X$21267 2057 VIA_via2_5
* cell instance $21268 r0 *1 67.925,79.17
X$21268 2057 VIA_via1_4
* cell instance $21269 r0 *1 79.325,94.43
X$21269 2057 VIA_via1_4
* cell instance $21270 r0 *1 74.765,84.77
X$21270 2057 VIA_via1_4
* cell instance $21271 r0 *1 74.765,84.63
X$21271 2057 VIA_via2_5
* cell instance $21272 r0 *1 83.695,91.63
X$21272 2057 VIA_via1_4
* cell instance $21273 r0 *1 88.255,91.63
X$21273 2057 VIA_via1_4
* cell instance $21274 r0 *1 85.785,93.17
X$21274 2057 VIA_via1_4
* cell instance $21275 r0 *1 68.305,90.37
X$21275 2057 VIA_via1_4
* cell instance $21276 r0 *1 68.305,90.37
X$21276 2057 VIA_via2_5
* cell instance $21277 r0 *1 69.825,87.57
X$21277 2057 VIA_via1_4
* cell instance $21278 r0 *1 87.685,80.43
X$21278 2057 VIA_via1_4
* cell instance $21279 r0 *1 87.685,80.43
X$21279 2057 VIA_via2_5
* cell instance $21280 r0 *1 86.925,80.43
X$21280 2057 VIA_via1_4
* cell instance $21281 r0 *1 86.925,80.43
X$21281 2057 VIA_via2_5
* cell instance $21282 r0 *1 79.055,92.19
X$21282 2057 VIA_via4_0
* cell instance $21283 r0 *1 79.055,92.19
X$21283 2057 VIA_via3_2
* cell instance $21284 r0 *1 71.215,92.19
X$21284 2057 VIA_via4_0
* cell instance $21285 r0 *1 71.215,90.37
X$21285 2057 VIA_via3_2
* cell instance $21286 r0 *1 74.195,80.01
X$21286 2058 VIA_via1_7
* cell instance $21287 r0 *1 74.195,80.01
X$21287 2058 VIA_via2_5
* cell instance $21288 r0 *1 74.005,80.29
X$21288 2058 VIA_via1_7
* cell instance $21289 r0 *1 86.615,82.11
X$21289 2058 VIA_via5_0
* cell instance $21290 r0 *1 86.355,92.47
X$21290 2058 VIA_via2_5
* cell instance $21291 r0 *1 83.315,80.01
X$21291 2058 VIA_via2_5
* cell instance $21292 r0 *1 83.315,81.83
X$21292 2058 VIA_via2_5
* cell instance $21293 r0 *1 71.535,80.01
X$21293 2058 VIA_via2_5
* cell instance $21294 r0 *1 54.055,80.43
X$21294 2058 VIA_via2_5
* cell instance $21295 r0 *1 64.695,80.43
X$21295 2058 VIA_via2_5
* cell instance $21296 r0 *1 71.535,80.43
X$21296 2058 VIA_via1_4
* cell instance $21297 r0 *1 71.535,80.29
X$21297 2058 VIA_via2_5
* cell instance $21298 r0 *1 64.695,76.37
X$21298 2058 VIA_via1_4
* cell instance $21299 r0 *1 74.005,81.97
X$21299 2058 VIA_via1_4
* cell instance $21300 r0 *1 86.355,93.17
X$21300 2058 VIA_via1_4
* cell instance $21301 r0 *1 64.885,88.83
X$21301 2058 VIA_via1_4
* cell instance $21302 r0 *1 53.105,80.43
X$21302 2058 VIA_via1_4
* cell instance $21303 r0 *1 53.105,80.43
X$21303 2058 VIA_via2_5
* cell instance $21304 r0 *1 54.055,91.63
X$21304 2058 VIA_via1_4
* cell instance $21305 r0 *1 83.885,77.63
X$21305 2058 VIA_via1_4
* cell instance $21306 r0 *1 93.575,81.97
X$21306 2058 VIA_via1_4
* cell instance $21307 r0 *1 93.575,81.97
X$21307 2058 VIA_via2_5
* cell instance $21308 r0 *1 86.615,92.47
X$21308 2058 VIA_via4_0
* cell instance $21309 r0 *1 86.615,92.47
X$21309 2058 VIA_via5_0
* cell instance $21310 r0 *1 86.615,92.47
X$21310 2058 VIA_via3_2
* cell instance $21311 r0 *1 87.735,82.11
X$21311 2058 VIA_via4_0
* cell instance $21312 r0 *1 87.735,81.97
X$21312 2058 VIA_via3_2
* cell instance $21313 r0 *1 84.265,94.57
X$21313 2059 VIA_via2_5
* cell instance $21314 r0 *1 82.935,94.57
X$21314 2059 VIA_via2_5
* cell instance $21315 r0 *1 84.265,95.97
X$21315 2059 VIA_via1_4
* cell instance $21316 r0 *1 84.645,80.43
X$21316 2059 VIA_via1_4
* cell instance $21317 r0 *1 84.645,80.57
X$21317 2059 VIA_via2_5
* cell instance $21318 r0 *1 83.695,80.43
X$21318 2059 VIA_via1_4
* cell instance $21319 r0 *1 83.695,80.57
X$21319 2059 VIA_via2_5
* cell instance $21320 r0 *1 82.175,80.43
X$21320 2059 VIA_via1_4
* cell instance $21321 r0 *1 82.175,80.57
X$21321 2059 VIA_via2_5
* cell instance $21322 r0 *1 84.075,78.89
X$21322 2059 VIA_via1_4
* cell instance $21323 r0 *1 86.735,80.43
X$21323 2060 VIA_via1_4
* cell instance $21324 r0 *1 87.115,79.45
X$21324 2060 VIA_via1_4
* cell instance $21325 r0 *1 87.875,79.45
X$21325 2061 VIA_via1_7
* cell instance $21326 r0 *1 87.495,80.43
X$21326 2061 VIA_via1_4
* cell instance $21327 r0 *1 89.585,79.59
X$21327 2062 VIA_via1_7
* cell instance $21328 r0 *1 89.585,79.59
X$21328 2062 VIA_via2_5
* cell instance $21329 r0 *1 90.345,79.59
X$21329 2062 VIA_via2_5
* cell instance $21330 r0 *1 88.445,79.59
X$21330 2062 VIA_via2_5
* cell instance $21331 r0 *1 82.365,82.11
X$21331 2062 VIA_via1_4
* cell instance $21332 r0 *1 82.385,81.97
X$21332 2062 VIA_via2_5
* cell instance $21333 r0 *1 90.345,79.17
X$21333 2062 VIA_via1_4
* cell instance $21334 r0 *1 88.635,81.97
X$21334 2062 VIA_via1_4
* cell instance $21335 r0 *1 88.635,82.11
X$21335 2062 VIA_via2_5
* cell instance $21336 r0 *1 85.595,80.99
X$21336 2063 VIA_via1_7
* cell instance $21337 r0 *1 86.165,83.37
X$21337 2063 VIA_via2_5
* cell instance $21338 r0 *1 90.535,83.51
X$21338 2063 VIA_via2_5
* cell instance $21339 r0 *1 85.595,83.37
X$21339 2063 VIA_via2_5
* cell instance $21340 r0 *1 87.875,89.39
X$21340 2063 VIA_via2_5
* cell instance $21341 r0 *1 87.115,89.39
X$21341 2063 VIA_via2_5
* cell instance $21342 r0 *1 86.355,89.11
X$21342 2063 VIA_via2_5
* cell instance $21343 r0 *1 87.115,89.11
X$21343 2063 VIA_via2_5
* cell instance $21344 r0 *1 86.735,88.27
X$21344 2063 VIA_via2_5
* cell instance $21345 r0 *1 86.355,88.27
X$21345 2063 VIA_via2_5
* cell instance $21346 r0 *1 86.355,86.03
X$21346 2063 VIA_via2_5
* cell instance $21347 r0 *1 86.735,88.62
X$21347 2063 VIA_via1_4
* cell instance $21348 r0 *1 87.875,90.37
X$21348 2063 VIA_via1_4
* cell instance $21349 r0 *1 87.115,86.03
X$21349 2063 VIA_via1_4
* cell instance $21350 r0 *1 87.115,86.03
X$21350 2063 VIA_via2_5
* cell instance $21351 r0 *1 89.585,83.23
X$21351 2063 VIA_via1_4
* cell instance $21352 r0 *1 89.585,83.37
X$21352 2063 VIA_via2_5
* cell instance $21353 r0 *1 90.535,84.77
X$21353 2063 VIA_via1_4
* cell instance $21354 r0 *1 89.775,80.43
X$21354 2063 VIA_via1_4
* cell instance $21355 r0 *1 86.735,83.23
X$21355 2063 VIA_via1_4
* cell instance $21356 r0 *1 86.735,83.37
X$21356 2063 VIA_via2_5
* cell instance $21357 r0 *1 89.965,79.17
X$21357 2063 VIA_via1_4
* cell instance $21358 r0 *1 96.615,79.87
X$21358 2064 VIA_via2_5
* cell instance $21359 r0 *1 96.045,79.87
X$21359 2064 VIA_via2_5
* cell instance $21360 r0 *1 93.765,79.87
X$21360 2064 VIA_via2_5
* cell instance $21361 r0 *1 90.155,79.87
X$21361 2064 VIA_via2_5
* cell instance $21362 r0 *1 89.015,79.87
X$21362 2064 VIA_via2_5
* cell instance $21363 r0 *1 96.615,80.43
X$21363 2064 VIA_via1_4
* cell instance $21364 r0 *1 89.015,80.43
X$21364 2064 VIA_via1_4
* cell instance $21365 r0 *1 88.825,81.97
X$21365 2064 VIA_via1_4
* cell instance $21366 r0 *1 91.295,80.43
X$21366 2064 VIA_via1_4
* cell instance $21367 r0 *1 91.295,80.57
X$21367 2064 VIA_via2_5
* cell instance $21368 r0 *1 93.765,80.43
X$21368 2064 VIA_via1_4
* cell instance $21369 r0 *1 93.765,80.57
X$21369 2064 VIA_via2_5
* cell instance $21370 r0 *1 90.155,79.17
X$21370 2064 VIA_via1_4
* cell instance $21371 r0 *1 96.045,78.05
X$21371 2064 VIA_via1_4
* cell instance $21372 r0 *1 87.685,90.09
X$21372 2065 VIA_via2_5
* cell instance $21373 r0 *1 89.015,90.09
X$21373 2065 VIA_via2_5
* cell instance $21374 r0 *1 81.035,88.69
X$21374 2065 VIA_via2_5
* cell instance $21375 r0 *1 80.465,88.69
X$21375 2065 VIA_via2_5
* cell instance $21376 r0 *1 65.835,88.55
X$21376 2065 VIA_via2_5
* cell instance $21377 r0 *1 88.065,88.27
X$21377 2065 VIA_via2_5
* cell instance $21378 r0 *1 87.305,88.27
X$21378 2065 VIA_via2_5
* cell instance $21379 r0 *1 91.295,88.27
X$21379 2065 VIA_via2_5
* cell instance $21380 r0 *1 81.035,80.85
X$21380 2065 VIA_via1_4
* cell instance $21381 r0 *1 80.465,90.37
X$21381 2065 VIA_via1_4
* cell instance $21382 r0 *1 80.465,90.23
X$21382 2065 VIA_via2_5
* cell instance $21383 r0 *1 84.455,90.3
X$21383 2065 VIA_via1_4
* cell instance $21384 r0 *1 84.455,90.23
X$21384 2065 VIA_via2_5
* cell instance $21385 r0 *1 87.875,88.83
X$21385 2065 VIA_via1_4
* cell instance $21386 r0 *1 87.305,87.57
X$21386 2065 VIA_via1_4
* cell instance $21387 r0 *1 91.485,86.03
X$21387 2065 VIA_via1_4
* cell instance $21388 r0 *1 89.015,90.37
X$21388 2065 VIA_via1_4
* cell instance $21389 r0 *1 65.835,88.83
X$21389 2065 VIA_via1_4
* cell instance $21390 r0 *1 90.725,83.23
X$21390 2065 VIA_via1_4
* cell instance $21391 r0 *1 90.915,80.43
X$21391 2065 VIA_via1_4
* cell instance $21392 r0 *1 91.675,79.17
X$21392 2065 VIA_via1_4
* cell instance $21393 r0 *1 93.005,81.69
X$21393 2066 VIA_via1_4
* cell instance $21394 r0 *1 92.815,79.17
X$21394 2066 VIA_via1_4
* cell instance $21395 r0 *1 93.195,80.01
X$21395 2067 VIA_via1_7
* cell instance $21396 r0 *1 93.765,77.63
X$21396 2067 VIA_via1_4
* cell instance $21397 r0 *1 96.995,78.61
X$21397 2068 VIA_via1_7
* cell instance $21398 r0 *1 96.615,77.63
X$21398 2068 VIA_via1_4
* cell instance $21399 r0 *1 96.615,81.97
X$21399 2069 VIA_via1_4
* cell instance $21400 r0 *1 96.615,82.11
X$21400 2069 VIA_via2_5
* cell instance $21401 r0 *1 91.485,81.97
X$21401 2069 VIA_via1_4
* cell instance $21402 r0 *1 91.485,82.11
X$21402 2069 VIA_via2_5
* cell instance $21403 r0 *1 89.015,81.97
X$21403 2069 VIA_via1_4
* cell instance $21404 r0 *1 89.015,82.11
X$21404 2069 VIA_via2_5
* cell instance $21405 r0 *1 89.205,80.43
X$21405 2069 VIA_via1_4
* cell instance $21406 r0 *1 93.195,81.97
X$21406 2069 VIA_via1_4
* cell instance $21407 r0 *1 93.195,82.11
X$21407 2069 VIA_via2_5
* cell instance $21408 r0 *1 96.425,79.45
X$21408 2069 VIA_via1_4
* cell instance $21409 r0 *1 94.335,80.01
X$21409 2070 VIA_via1_7
* cell instance $21410 r0 *1 94.335,80.01
X$21410 2070 VIA_via2_5
* cell instance $21411 r0 *1 97.815,79.59
X$21411 2070 VIA_via4_0
* cell instance $21412 r0 *1 97.815,80.01
X$21412 2070 VIA_via3_2
* cell instance $21413 r0 *1 96.615,79.17
X$21413 2071 VIA_via1_4
* cell instance $21414 r0 *1 96.615,79.03
X$21414 2071 VIA_via2_5
* cell instance $21415 r0 *1 97.815,79.03
X$21415 2071 VIA_via4_0
* cell instance $21416 r0 *1 97.815,79.03
X$21416 2071 VIA_via3_2
* cell instance $21417 r0 *1 13.015,78.19
X$21417 2072 VIA_via1_7
* cell instance $21418 r0 *1 13.015,78.19
X$21418 2072 VIA_via2_5
* cell instance $21419 r0 *1 12.255,78.19
X$21419 2072 VIA_via2_5
* cell instance $21420 r0 *1 12.255,79.17
X$21420 2072 VIA_via1_4
* cell instance $21421 r0 *1 93.195,79.17
X$21421 2073 VIA_via1_4
* cell instance $21422 r0 *1 93.195,79.17
X$21422 2073 VIA_via2_5
* cell instance $21423 r0 *1 94.145,79.17
X$21423 2073 VIA_via1_4
* cell instance $21424 r0 *1 94.145,79.17
X$21424 2073 VIA_via2_5
* cell instance $21425 r0 *1 90.535,79.17
X$21425 2074 VIA_via1_4
* cell instance $21426 r0 *1 91.295,79.17
X$21426 2074 VIA_via1_4
* cell instance $21427 r0 *1 17.765,77.63
X$21427 2075 VIA_via1_4
* cell instance $21428 r0 *1 17.765,77.63
X$21428 2075 VIA_via2_5
* cell instance $21429 r0 *1 14.155,77.63
X$21429 2075 VIA_via1_4
* cell instance $21430 r0 *1 14.155,77.63
X$21430 2075 VIA_via2_5
* cell instance $21431 r0 *1 92.055,79.03
X$21431 2076 VIA_via1_7
* cell instance $21432 r0 *1 91.865,79.03
X$21432 2076 VIA_via1_4
* cell instance $21433 r0 *1 17.765,80.01
X$21433 2077 VIA_via1_7
* cell instance $21434 r0 *1 17.765,79.17
X$21434 2077 VIA_via2_5
* cell instance $21435 r0 *1 19.285,79.17
X$21435 2077 VIA_via1_4
* cell instance $21436 r0 *1 19.285,79.17
X$21436 2077 VIA_via2_5
* cell instance $21437 r0 *1 20.425,77.91
X$21437 2078 VIA_via2_5
* cell instance $21438 r0 *1 20.425,77.63
X$21438 2078 VIA_via1_4
* cell instance $21439 r0 *1 11.115,77.91
X$21439 2078 VIA_via1_4
* cell instance $21440 r0 *1 11.115,77.91
X$21440 2078 VIA_via2_5
* cell instance $21441 r0 *1 89.205,77.77
X$21441 2079 VIA_via1_4
* cell instance $21442 r0 *1 89.205,77.77
X$21442 2079 VIA_via2_5
* cell instance $21443 r0 *1 90.345,77.63
X$21443 2079 VIA_via1_4
* cell instance $21444 r0 *1 90.345,77.77
X$21444 2079 VIA_via2_5
* cell instance $21445 r0 *1 22.135,80.01
X$21445 2080 VIA_via1_7
* cell instance $21446 r0 *1 25.935,78.33
X$21446 2080 VIA_via2_5
* cell instance $21447 r0 *1 22.135,78.33
X$21447 2080 VIA_via2_5
* cell instance $21448 r0 *1 25.935,77.63
X$21448 2080 VIA_via1_4
* cell instance $21449 r0 *1 27.645,85.05
X$21449 2081 VIA_via2_5
* cell instance $21450 r0 *1 28.025,77.63
X$21450 2081 VIA_via2_5
* cell instance $21451 r0 *1 12.825,85.05
X$21451 2081 VIA_via2_5
* cell instance $21452 r0 *1 12.635,90.09
X$21452 2081 VIA_via1_4
* cell instance $21453 r0 *1 29.545,77.63
X$21453 2081 VIA_via1_4
* cell instance $21454 r0 *1 29.545,77.63
X$21454 2081 VIA_via2_5
* cell instance $21455 r0 *1 28.025,76.37
X$21455 2081 VIA_via1_4
* cell instance $21456 r0 *1 29.545,78.19
X$21456 2082 VIA_via1_7
* cell instance $21457 r0 *1 29.545,79.73
X$21457 2082 VIA_via2_5
* cell instance $21458 r0 *1 31.635,79.73
X$21458 2082 VIA_via2_5
* cell instance $21459 r0 *1 31.635,80.43
X$21459 2082 VIA_via1_4
* cell instance $21460 r0 *1 30.495,79.59
X$21460 2083 VIA_via1_7
* cell instance $21461 r0 *1 30.495,79.59
X$21461 2083 VIA_via2_5
* cell instance $21462 r0 *1 30.875,79.59
X$21462 2083 VIA_via2_5
* cell instance $21463 r0 *1 30.875,79.17
X$21463 2083 VIA_via1_4
* cell instance $21464 r0 *1 31.825,77.77
X$21464 2084 VIA_via2_5
* cell instance $21465 r0 *1 30.495,77.77
X$21465 2084 VIA_via2_5
* cell instance $21466 r0 *1 31.825,79.17
X$21466 2084 VIA_via1_4
* cell instance $21467 r0 *1 30.495,76.51
X$21467 2084 VIA_via1_4
* cell instance $21468 r0 *1 32.585,77.63
X$21468 2085 VIA_via2_5
* cell instance $21469 r0 *1 32.585,79.17
X$21469 2085 VIA_via1_4
* cell instance $21470 r0 *1 34.295,77.63
X$21470 2085 VIA_via1_4
* cell instance $21471 r0 *1 34.295,77.63
X$21471 2085 VIA_via2_5
* cell instance $21472 r0 *1 31.635,78.61
X$21472 2086 VIA_via1_7
* cell instance $21473 r0 *1 31.635,77.63
X$21473 2086 VIA_via1_4
* cell instance $21474 r0 *1 33.535,79.17
X$21474 2087 VIA_via1_4
* cell instance $21475 r0 *1 33.535,79.17
X$21475 2087 VIA_via2_5
* cell instance $21476 r0 *1 31.635,79.17
X$21476 2087 VIA_via1_4
* cell instance $21477 r0 *1 31.635,79.17
X$21477 2087 VIA_via2_5
* cell instance $21478 r0 *1 30.685,80.01
X$21478 2088 VIA_via1_7
* cell instance $21479 r0 *1 34.675,79.45
X$21479 2088 VIA_via2_5
* cell instance $21480 r0 *1 30.685,79.45
X$21480 2088 VIA_via2_5
* cell instance $21481 r0 *1 34.675,77.63
X$21481 2088 VIA_via1_4
* cell instance $21482 r0 *1 87.305,80.01
X$21482 2089 VIA_via1_7
* cell instance $21483 r0 *1 85.595,78.61
X$21483 2089 VIA_via2_5
* cell instance $21484 r0 *1 87.305,78.61
X$21484 2089 VIA_via2_5
* cell instance $21485 r0 *1 85.595,77.63
X$21485 2089 VIA_via1_4
* cell instance $21486 r0 *1 38.475,77.63
X$21486 2090 VIA_via1_4
* cell instance $21487 r0 *1 38.475,77.77
X$21487 2090 VIA_via2_5
* cell instance $21488 r0 *1 37.525,77.77
X$21488 2090 VIA_via1_4
* cell instance $21489 r0 *1 37.525,77.77
X$21489 2090 VIA_via2_5
* cell instance $21490 r0 *1 39.425,81.41
X$21490 2091 VIA_via1_7
* cell instance $21491 r0 *1 39.425,77.63
X$21491 2091 VIA_via2_5
* cell instance $21492 r0 *1 37.905,77.63
X$21492 2091 VIA_via1_4
* cell instance $21493 r0 *1 37.905,77.63
X$21493 2091 VIA_via2_5
* cell instance $21494 r0 *1 86.545,78.19
X$21494 2092 VIA_via1_7
* cell instance $21495 r0 *1 86.545,78.19
X$21495 2092 VIA_via2_5
* cell instance $21496 r0 *1 85.215,78.19
X$21496 2092 VIA_via2_5
* cell instance $21497 r0 *1 85.215,79.17
X$21497 2092 VIA_via1_4
* cell instance $21498 r0 *1 42.845,77.63
X$21498 2093 VIA_via1_4
* cell instance $21499 r0 *1 42.655,77.63
X$21499 2093 VIA_via1_4
* cell instance $21500 r0 *1 43.605,77.63
X$21500 2094 VIA_via1_4
* cell instance $21501 r0 *1 43.605,76.51
X$21501 2094 VIA_via1_4
* cell instance $21502 r0 *1 47.405,80.15
X$21502 2095 VIA_via1_4
* cell instance $21503 r0 *1 47.405,79.17
X$21503 2095 VIA_via1_4
* cell instance $21504 r0 *1 47.405,79.17
X$21504 2095 VIA_via2_5
* cell instance $21505 r0 *1 45.885,79.17
X$21505 2095 VIA_via1_4
* cell instance $21506 r0 *1 45.885,79.17
X$21506 2095 VIA_via2_5
* cell instance $21507 r0 *1 83.505,80.01
X$21507 2096 VIA_via1_7
* cell instance $21508 r0 *1 83.505,79.31
X$21508 2096 VIA_via2_5
* cell instance $21509 r0 *1 81.795,79.17
X$21509 2096 VIA_via1_4
* cell instance $21510 r0 *1 81.795,79.31
X$21510 2096 VIA_via2_5
* cell instance $21511 r0 *1 51.965,77.63
X$21511 2097 VIA_via1_4
* cell instance $21512 r0 *1 52.155,77.63
X$21512 2097 VIA_via1_4
* cell instance $21513 r0 *1 51.775,77.63
X$21513 2098 VIA_via2_5
* cell instance $21514 r0 *1 51.775,76.51
X$21514 2098 VIA_via1_4
* cell instance $21515 r0 *1 53.865,77.63
X$21515 2098 VIA_via1_4
* cell instance $21516 r0 *1 53.865,77.63
X$21516 2098 VIA_via2_5
* cell instance $21517 r0 *1 71.155,80.01
X$21517 2099 VIA_via1_7
* cell instance $21518 r0 *1 71.155,77.63
X$21518 2099 VIA_via2_5
* cell instance $21519 r0 *1 70.585,77.63
X$21519 2099 VIA_via1_4
* cell instance $21520 r0 *1 70.585,77.63
X$21520 2099 VIA_via2_5
* cell instance $21521 r0 *1 52.915,76.79
X$21521 2100 VIA_via1_7
* cell instance $21522 r0 *1 52.915,77.63
X$21522 2100 VIA_via1_4
* cell instance $21523 r0 *1 73.815,85.19
X$21523 2101 VIA_via1_7
* cell instance $21524 r0 *1 73.815,85.19
X$21524 2101 VIA_via2_5
* cell instance $21525 r0 *1 72.485,85.19
X$21525 2101 VIA_via2_5
* cell instance $21526 r0 *1 72.295,85.19
X$21526 2101 VIA_via2_5
* cell instance $21527 r0 *1 72.485,79.17
X$21527 2101 VIA_via2_5
* cell instance $21528 r0 *1 70.015,79.17
X$21528 2101 VIA_via1_4
* cell instance $21529 r0 *1 70.015,79.17
X$21529 2101 VIA_via2_5
* cell instance $21530 r0 *1 72.295,86.03
X$21530 2101 VIA_via1_4
* cell instance $21531 r0 *1 65.265,82.95
X$21531 2102 VIA_via2_5
* cell instance $21532 r0 *1 67.165,79.17
X$21532 2102 VIA_via2_5
* cell instance $21533 r0 *1 65.265,79.17
X$21533 2102 VIA_via2_5
* cell instance $21534 r0 *1 70.775,82.95
X$21534 2102 VIA_via1_4
* cell instance $21535 r0 *1 70.775,82.95
X$21535 2102 VIA_via2_5
* cell instance $21536 r0 *1 64.315,79.17
X$21536 2102 VIA_via1_4
* cell instance $21537 r0 *1 64.315,79.17
X$21537 2102 VIA_via2_5
* cell instance $21538 r0 *1 67.165,80.43
X$21538 2102 VIA_via1_4
* cell instance $21539 r0 *1 65.265,84.77
X$21539 2102 VIA_via1_4
* cell instance $21540 r0 *1 65.265,84.77
X$21540 2102 VIA_via2_5
* cell instance $21541 r0 *1 64.315,84.77
X$21541 2102 VIA_via1_4
* cell instance $21542 r0 *1 64.315,84.77
X$21542 2102 VIA_via2_5
* cell instance $21543 r0 *1 58.615,79.17
X$21543 2103 VIA_via2_5
* cell instance $21544 r0 *1 55.765,79.17
X$21544 2103 VIA_via1_4
* cell instance $21545 r0 *1 55.765,79.17
X$21545 2103 VIA_via2_5
* cell instance $21546 r0 *1 58.615,77.63
X$21546 2103 VIA_via1_4
* cell instance $21547 r0 *1 65.075,78.61
X$21547 2104 VIA_via1_7
* cell instance $21548 r0 *1 65.075,77.63
X$21548 2104 VIA_via1_4
* cell instance $21549 r0 *1 17.765,80.43
X$21549 2105 VIA_via2_5
* cell instance $21550 r0 *1 16.055,80.43
X$21550 2105 VIA_via1_4
* cell instance $21551 r0 *1 16.055,80.43
X$21551 2105 VIA_via2_5
* cell instance $21552 r0 *1 17.765,81.55
X$21552 2105 VIA_via1_4
* cell instance $21553 r0 *1 16.815,80.43
X$21553 2105 VIA_via1_4
* cell instance $21554 r0 *1 16.815,80.43
X$21554 2105 VIA_via2_5
* cell instance $21555 r0 *1 29.165,80.43
X$21555 2106 VIA_via2_5
* cell instance $21556 r0 *1 28.975,80.43
X$21556 2106 VIA_via1_4
* cell instance $21557 r0 *1 29.165,81.55
X$21557 2106 VIA_via1_4
* cell instance $21558 r0 *1 29.735,80.43
X$21558 2106 VIA_via1_4
* cell instance $21559 r0 *1 29.735,80.43
X$21559 2106 VIA_via2_5
* cell instance $21560 r0 *1 36.005,83.23
X$21560 2107 VIA_via2_5
* cell instance $21561 r0 *1 36.005,84.35
X$21561 2107 VIA_via1_4
* cell instance $21562 r0 *1 34.675,80.43
X$21562 2107 VIA_via1_4
* cell instance $21563 r0 *1 34.865,83.23
X$21563 2107 VIA_via1_4
* cell instance $21564 r0 *1 34.865,83.23
X$21564 2107 VIA_via2_5
* cell instance $21565 r0 *1 43.795,80.43
X$21565 2108 VIA_via2_5
* cell instance $21566 r0 *1 41.325,80.43
X$21566 2108 VIA_via1_4
* cell instance $21567 r0 *1 41.325,80.43
X$21567 2108 VIA_via2_5
* cell instance $21568 r0 *1 42.085,80.43
X$21568 2108 VIA_via1_4
* cell instance $21569 r0 *1 42.085,80.43
X$21569 2108 VIA_via2_5
* cell instance $21570 r0 *1 43.795,81.55
X$21570 2108 VIA_via1_4
* cell instance $21571 r0 *1 43.035,80.01
X$21571 2109 VIA_via1_7
* cell instance $21572 r0 *1 42.085,79.17
X$21572 2109 VIA_via1_4
* cell instance $21573 r0 *1 55.195,78.89
X$21573 2110 VIA_via1_7
* cell instance $21574 r0 *1 55.195,95.97
X$21574 2110 VIA_via1_4
* cell instance $21575 r0 *1 66.975,80.01
X$21575 2111 VIA_via1_7
* cell instance $21576 r0 *1 66.025,79.17
X$21576 2111 VIA_via1_4
* cell instance $21577 r0 *1 68.305,79.59
X$21577 2112 VIA_via1_7
* cell instance $21578 r0 *1 68.685,80.43
X$21578 2112 VIA_via1_4
* cell instance $21579 r0 *1 91.485,80.71
X$21579 2113 VIA_via2_5
* cell instance $21580 r0 *1 90.535,85.61
X$21580 2113 VIA_via2_5
* cell instance $21581 r0 *1 91.485,85.61
X$21581 2113 VIA_via2_5
* cell instance $21582 r0 *1 67.355,80.01
X$21582 2113 VIA_via2_5
* cell instance $21583 r0 *1 69.445,80.15
X$21583 2113 VIA_via2_5
* cell instance $21584 r0 *1 73.625,80.71
X$21584 2113 VIA_via2_5
* cell instance $21585 r0 *1 73.625,80.15
X$21585 2113 VIA_via2_5
* cell instance $21586 r0 *1 66.595,80.43
X$21586 2113 VIA_via2_5
* cell instance $21587 r0 *1 79.895,80.71
X$21587 2113 VIA_via2_5
* cell instance $21588 r0 *1 91.865,87.29
X$21588 2113 VIA_via2_5
* cell instance $21589 r0 *1 90.535,87.29
X$21589 2113 VIA_via2_5
* cell instance $21590 r0 *1 69.445,80.43
X$21590 2113 VIA_via1_4
* cell instance $21591 r0 *1 67.355,80.43
X$21591 2113 VIA_via1_4
* cell instance $21592 r0 *1 67.355,80.43
X$21592 2113 VIA_via2_5
* cell instance $21593 r0 *1 66.595,84.77
X$21593 2113 VIA_via1_4
* cell instance $21594 r0 *1 79.895,80.43
X$21594 2113 VIA_via1_4
* cell instance $21595 r0 *1 79.895,83.23
X$21595 2113 VIA_via1_4
* cell instance $21596 r0 *1 90.535,86.03
X$21596 2113 VIA_via1_4
* cell instance $21597 r0 *1 91.865,87.57
X$21597 2113 VIA_via1_4
* cell instance $21598 r0 *1 91.485,84.77
X$21598 2113 VIA_via1_4
* cell instance $21599 r0 *1 91.675,81.97
X$21599 2113 VIA_via1_4
* cell instance $21600 r0 *1 91.485,80.43
X$21600 2113 VIA_via1_4
* cell instance $21601 r0 *1 73.625,79.17
X$21601 2113 VIA_via1_4
* cell instance $21602 r0 *1 74.765,80.57
X$21602 2114 VIA_via1_7
* cell instance $21603 r0 *1 74.575,82.81
X$21603 2114 VIA_via1_7
* cell instance $21604 r0 *1 77.045,82.25
X$21604 2115 VIA_via2_5
* cell instance $21605 r0 *1 77.425,82.25
X$21605 2115 VIA_via2_5
* cell instance $21606 r0 *1 78.185,82.25
X$21606 2115 VIA_via1_4
* cell instance $21607 r0 *1 78.185,82.25
X$21607 2115 VIA_via2_5
* cell instance $21608 r0 *1 76.855,80.43
X$21608 2115 VIA_via1_4
* cell instance $21609 r0 *1 77.045,80.43
X$21609 2115 VIA_via1_4
* cell instance $21610 r0 *1 77.425,82.95
X$21610 2115 VIA_via1_4
* cell instance $21611 r0 *1 92.625,80.43
X$21611 2116 VIA_via2_5
* cell instance $21612 r0 *1 92.055,85.47
X$21612 2116 VIA_via2_5
* cell instance $21613 r0 *1 79.515,80.57
X$21613 2116 VIA_via2_5
* cell instance $21614 r0 *1 78.375,80.43
X$21614 2116 VIA_via2_5
* cell instance $21615 r0 *1 83.885,85.47
X$21615 2116 VIA_via2_5
* cell instance $21616 r0 *1 67.165,85.05
X$21616 2116 VIA_via2_5
* cell instance $21617 r0 *1 67.165,85.47
X$21617 2116 VIA_via2_5
* cell instance $21618 r0 *1 64.505,85.05
X$21618 2116 VIA_via2_5
* cell instance $21619 r0 *1 78.185,85.47
X$21619 2116 VIA_via2_5
* cell instance $21620 r0 *1 67.165,84.77
X$21620 2116 VIA_via1_4
* cell instance $21621 r0 *1 79.135,83.23
X$21621 2116 VIA_via1_4
* cell instance $21622 r0 *1 76.475,80.43
X$21622 2116 VIA_via1_4
* cell instance $21623 r0 *1 76.475,80.43
X$21623 2116 VIA_via2_5
* cell instance $21624 r0 *1 83.885,84.77
X$21624 2116 VIA_via1_4
* cell instance $21625 r0 *1 93.195,86.03
X$21625 2116 VIA_via1_4
* cell instance $21626 r0 *1 93.195,85.89
X$21626 2116 VIA_via2_5
* cell instance $21627 r0 *1 64.885,87.57
X$21627 2116 VIA_via1_4
* cell instance $21628 r0 *1 92.815,81.97
X$21628 2116 VIA_via1_4
* cell instance $21629 r0 *1 79.515,79.45
X$21629 2116 VIA_via1_4
* cell instance $21630 r0 *1 93.385,80.43
X$21630 2116 VIA_via1_4
* cell instance $21631 r0 *1 93.385,80.43
X$21631 2116 VIA_via2_5
* cell instance $21632 r0 *1 92.245,81.97
X$21632 2116 VIA_via1_4
* cell instance $21633 r0 *1 92.055,84.77
X$21633 2116 VIA_via1_4
* cell instance $21634 r0 *1 81.985,80.15
X$21634 2117 VIA_via1_4
* cell instance $21635 r0 *1 82.555,80.43
X$21635 2117 VIA_via1_4
* cell instance $21636 r0 *1 88.065,80.01
X$21636 2118 VIA_via1_7
* cell instance $21637 r0 *1 88.255,77.63
X$21637 2118 VIA_via1_4
* cell instance $21638 r0 *1 91.105,80.15
X$21638 2119 VIA_via1_4
* cell instance $21639 r0 *1 92.055,80.43
X$21639 2119 VIA_via1_4
* cell instance $21640 r0 *1 92.055,81.41
X$21640 2120 VIA_via1_7
* cell instance $21641 r0 *1 92.245,79.17
X$21641 2120 VIA_via1_4
* cell instance $21642 r0 *1 92.245,80.43
X$21642 2121 VIA_via1_4
* cell instance $21643 r0 *1 91.865,80.15
X$21643 2121 VIA_via1_4
* cell instance $21644 r0 *1 95.285,80.15
X$21644 2122 VIA_via1_4
* cell instance $21645 r0 *1 95.285,80.15
X$21645 2122 VIA_via2_5
* cell instance $21646 r0 *1 96.695,80.15
X$21646 2122 VIA_via4_0
* cell instance $21647 r0 *1 96.695,80.15
X$21647 2122 VIA_via3_2
* cell instance $21648 r0 *1 11.305,80.01
X$21648 2123 VIA_via1_7
* cell instance $21649 r0 *1 11.305,80.01
X$21649 2123 VIA_via2_5
* cell instance $21650 r0 *1 8.455,80.01
X$21650 2123 VIA_via2_5
* cell instance $21651 r0 *1 8.455,79.17
X$21651 2123 VIA_via1_4
* cell instance $21652 r0 *1 94.715,80.43
X$21652 2124 VIA_via1_4
* cell instance $21653 r0 *1 94.715,80.43
X$21653 2124 VIA_via2_5
* cell instance $21654 r0 *1 93.955,80.43
X$21654 2124 VIA_via1_4
* cell instance $21655 r0 *1 93.955,80.43
X$21655 2124 VIA_via2_5
* cell instance $21656 r0 *1 92.815,80.15
X$21656 2125 VIA_via2_5
* cell instance $21657 r0 *1 93.575,80.15
X$21657 2125 VIA_via1_4
* cell instance $21658 r0 *1 93.575,80.15
X$21658 2125 VIA_via2_5
* cell instance $21659 r0 *1 92.815,80.43
X$21659 2125 VIA_via1_4
* cell instance $21660 r0 *1 10.925,81.41
X$21660 2126 VIA_via1_7
* cell instance $21661 r0 *1 11.115,80.15
X$21661 2126 VIA_via2_5
* cell instance $21662 r0 *1 21.185,80.15
X$21662 2126 VIA_via2_5
* cell instance $21663 r0 *1 21.185,77.63
X$21663 2126 VIA_via1_4
* cell instance $21664 r0 *1 21.565,81.55
X$21664 2127 VIA_via1_4
* cell instance $21665 r0 *1 19.285,80.43
X$21665 2127 VIA_via1_4
* cell instance $21666 r0 *1 19.285,80.43
X$21666 2127 VIA_via2_5
* cell instance $21667 r0 *1 21.185,80.43
X$21667 2127 VIA_via1_4
* cell instance $21668 r0 *1 21.185,80.43
X$21668 2127 VIA_via2_5
* cell instance $21669 r0 *1 25.745,80.43
X$21669 2128 VIA_via1_4
* cell instance $21670 r0 *1 25.745,80.43
X$21670 2128 VIA_via2_5
* cell instance $21671 r0 *1 25.365,81.55
X$21671 2128 VIA_via1_4
* cell instance $21672 r0 *1 24.225,80.43
X$21672 2128 VIA_via1_4
* cell instance $21673 r0 *1 24.225,80.43
X$21673 2128 VIA_via2_5
* cell instance $21674 r0 *1 90.345,80.43
X$21674 2129 VIA_via1_4
* cell instance $21675 r0 *1 90.535,80.43
X$21675 2129 VIA_via1_4
* cell instance $21676 r0 *1 34.295,79.59
X$21676 2130 VIA_via1_7
* cell instance $21677 r0 *1 34.295,80.43
X$21677 2130 VIA_via2_5
* cell instance $21678 r0 *1 32.395,80.43
X$21678 2130 VIA_via1_4
* cell instance $21679 r0 *1 32.395,80.43
X$21679 2130 VIA_via2_5
* cell instance $21680 r0 *1 83.125,80.43
X$21680 2131 VIA_via1_4
* cell instance $21681 r0 *1 83.125,80.43
X$21681 2131 VIA_via2_5
* cell instance $21682 r0 *1 84.265,80.43
X$21682 2131 VIA_via1_4
* cell instance $21683 r0 *1 84.265,80.43
X$21683 2131 VIA_via2_5
* cell instance $21684 r0 *1 85.025,80.43
X$21684 2132 VIA_via1_4
* cell instance $21685 r0 *1 85.215,80.43
X$21685 2132 VIA_via1_4
* cell instance $21686 r0 *1 46.265,79.59
X$21686 2133 VIA_via1_7
* cell instance $21687 r0 *1 46.265,80.43
X$21687 2133 VIA_via2_5
* cell instance $21688 r0 *1 45.125,80.43
X$21688 2133 VIA_via1_4
* cell instance $21689 r0 *1 45.125,80.43
X$21689 2133 VIA_via2_5
* cell instance $21690 r0 *1 74.955,80.43
X$21690 2134 VIA_via1_4
* cell instance $21691 r0 *1 74.955,80.29
X$21691 2134 VIA_via2_5
* cell instance $21692 r0 *1 77.615,80.29
X$21692 2134 VIA_via1_4
* cell instance $21693 r0 *1 77.615,80.29
X$21693 2134 VIA_via2_5
* cell instance $21694 r0 *1 49.305,80.01
X$21694 2135 VIA_via1_7
* cell instance $21695 r0 *1 49.305,79.17
X$21695 2135 VIA_via1_4
* cell instance $21696 r0 *1 74.005,79.59
X$21696 2136 VIA_via1_7
* cell instance $21697 r0 *1 74.005,79.87
X$21697 2136 VIA_via2_5
* cell instance $21698 r0 *1 72.295,79.87
X$21698 2136 VIA_via2_5
* cell instance $21699 r0 *1 72.295,80.43
X$21699 2136 VIA_via1_4
* cell instance $21700 r0 *1 71.725,82.81
X$21700 2137 VIA_via1_7
* cell instance $21701 r0 *1 71.725,80.43
X$21701 2137 VIA_via2_5
* cell instance $21702 r0 *1 70.205,80.43
X$21702 2137 VIA_via1_4
* cell instance $21703 r0 *1 70.205,80.43
X$21703 2137 VIA_via2_5
* cell instance $21704 r0 *1 55.005,80.29
X$21704 2138 VIA_via2_5
* cell instance $21705 r0 *1 52.155,80.43
X$21705 2138 VIA_via1_4
* cell instance $21706 r0 *1 52.155,80.29
X$21706 2138 VIA_via2_5
* cell instance $21707 r0 *1 55.005,81.55
X$21707 2138 VIA_via1_4
* cell instance $21708 r0 *1 55.575,80.43
X$21708 2138 VIA_via1_4
* cell instance $21709 r0 *1 55.575,80.29
X$21709 2138 VIA_via2_5
* cell instance $21710 r0 *1 68.115,80.43
X$21710 2139 VIA_via1_4
* cell instance $21711 r0 *1 68.115,80.43
X$21711 2139 VIA_via2_5
* cell instance $21712 r0 *1 69.825,80.43
X$21712 2139 VIA_via1_4
* cell instance $21713 r0 *1 69.825,80.43
X$21713 2139 VIA_via2_5
* cell instance $21714 r0 *1 9.215,81.97
X$21714 2140 VIA_via2_5
* cell instance $21715 r0 *1 9.975,81.97
X$21715 2140 VIA_via1_4
* cell instance $21716 r0 *1 9.975,81.97
X$21716 2140 VIA_via2_5
* cell instance $21717 r0 *1 9.215,82.95
X$21717 2140 VIA_via1_4
* cell instance $21718 r0 *1 8.265,81.97
X$21718 2140 VIA_via1_4
* cell instance $21719 r0 *1 8.265,81.97
X$21719 2140 VIA_via2_5
* cell instance $21720 r0 *1 10.355,83.23
X$21720 2141 VIA_via2_5
* cell instance $21721 r0 *1 11.115,83.23
X$21721 2141 VIA_via2_5
* cell instance $21722 r0 *1 10.165,83.23
X$21722 2141 VIA_via1_4
* cell instance $21723 r0 *1 10.165,83.23
X$21723 2141 VIA_via2_5
* cell instance $21724 r0 *1 10.545,81.97
X$21724 2141 VIA_via1_4
* cell instance $21725 r0 *1 11.115,84.35
X$21725 2141 VIA_via1_4
* cell instance $21726 r0 *1 16.435,80.99
X$21726 2142 VIA_via1_7
* cell instance $21727 r0 *1 15.485,81.97
X$21727 2142 VIA_via1_4
* cell instance $21728 r0 *1 19.665,80.99
X$21728 2143 VIA_via1_7
* cell instance $21729 r0 *1 19.285,81.97
X$21729 2143 VIA_via1_4
* cell instance $21730 r0 *1 20.235,86.03
X$21730 2144 VIA_via2_5
* cell instance $21731 r0 *1 23.465,87.57
X$21731 2144 VIA_via2_5
* cell instance $21732 r0 *1 19.475,86.03
X$21732 2144 VIA_via2_5
* cell instance $21733 r0 *1 17.385,86.03
X$21733 2144 VIA_via1_4
* cell instance $21734 r0 *1 17.385,86.03
X$21734 2144 VIA_via2_5
* cell instance $21735 r0 *1 23.465,91.63
X$21735 2144 VIA_via1_4
* cell instance $21736 r0 *1 19.475,87.57
X$21736 2144 VIA_via1_4
* cell instance $21737 r0 *1 22.895,87.15
X$21737 2144 VIA_via1_4
* cell instance $21738 r0 *1 23.275,87.57
X$21738 2144 VIA_via1_4
* cell instance $21739 r0 *1 23.275,87.57
X$21739 2144 VIA_via2_5
* cell instance $21740 r0 *1 22.895,86.03
X$21740 2144 VIA_via1_4
* cell instance $21741 r0 *1 22.895,86.03
X$21741 2144 VIA_via2_5
* cell instance $21742 r0 *1 25.175,88.83
X$21742 2144 VIA_via1_4
* cell instance $21743 r0 *1 24.985,87.57
X$21743 2144 VIA_via1_4
* cell instance $21744 r0 *1 24.985,87.57
X$21744 2144 VIA_via2_5
* cell instance $21745 r0 *1 20.045,81.97
X$21745 2144 VIA_via1_4
* cell instance $21746 r0 *1 20.235,83.23
X$21746 2144 VIA_via1_4
* cell instance $21747 r0 *1 34.485,81.97
X$21747 2145 VIA_via2_5
* cell instance $21748 r0 *1 29.545,81.97
X$21748 2145 VIA_via2_5
* cell instance $21749 r0 *1 24.225,81.97
X$21749 2145 VIA_via2_5
* cell instance $21750 r0 *1 23.275,81.97
X$21750 2145 VIA_via2_5
* cell instance $21751 r0 *1 29.545,87.57
X$21751 2145 VIA_via1_4
* cell instance $21752 r0 *1 29.545,84.77
X$21752 2145 VIA_via1_4
* cell instance $21753 r0 *1 33.155,81.97
X$21753 2145 VIA_via1_4
* cell instance $21754 r0 *1 33.155,81.97
X$21754 2145 VIA_via2_5
* cell instance $21755 r0 *1 29.545,82.95
X$21755 2145 VIA_via1_4
* cell instance $21756 r0 *1 27.645,81.97
X$21756 2145 VIA_via1_4
* cell instance $21757 r0 *1 27.645,81.97
X$21757 2145 VIA_via2_5
* cell instance $21758 r0 *1 34.485,84.77
X$21758 2145 VIA_via1_4
* cell instance $21759 r0 *1 23.275,77.63
X$21759 2145 VIA_via1_4
* cell instance $21760 r0 *1 24.225,83.23
X$21760 2145 VIA_via1_4
* cell instance $21761 r0 *1 23.845,81.97
X$21761 2145 VIA_via1_4
* cell instance $21762 r0 *1 23.845,81.97
X$21762 2145 VIA_via2_5
* cell instance $21763 r0 *1 37.715,81.97
X$21763 2146 VIA_via1_4
* cell instance $21764 r0 *1 37.715,81.97
X$21764 2146 VIA_via2_5
* cell instance $21765 r0 *1 39.045,80.85
X$21765 2146 VIA_via1_4
* cell instance $21766 r0 *1 38.475,81.97
X$21766 2146 VIA_via1_4
* cell instance $21767 r0 *1 38.475,81.97
X$21767 2146 VIA_via2_5
* cell instance $21768 r0 *1 39.235,78.19
X$21768 2147 VIA_via1_7
* cell instance $21769 r0 *1 38.855,95.97
X$21769 2147 VIA_via1_4
* cell instance $21770 r0 *1 41.705,80.99
X$21770 2148 VIA_via1_7
* cell instance $21771 r0 *1 41.515,81.97
X$21771 2148 VIA_via1_4
* cell instance $21772 r0 *1 44.745,84.35
X$21772 2149 VIA_via2_5
* cell instance $21773 r0 *1 47.025,84.77
X$21773 2149 VIA_via2_5
* cell instance $21774 r0 *1 45.885,81.97
X$21774 2149 VIA_via2_5
* cell instance $21775 r0 *1 43.795,86.03
X$21775 2149 VIA_via2_5
* cell instance $21776 r0 *1 42.465,86.03
X$21776 2149 VIA_via2_5
* cell instance $21777 r0 *1 42.275,81.97
X$21777 2149 VIA_via1_4
* cell instance $21778 r0 *1 42.465,83.23
X$21778 2149 VIA_via1_4
* cell instance $21779 r0 *1 48.925,81.97
X$21779 2149 VIA_via1_4
* cell instance $21780 r0 *1 48.925,81.97
X$21780 2149 VIA_via2_5
* cell instance $21781 r0 *1 44.745,83.23
X$21781 2149 VIA_via1_4
* cell instance $21782 r0 *1 45.885,80.43
X$21782 2149 VIA_via1_4
* cell instance $21783 r0 *1 45.885,84.77
X$21783 2149 VIA_via1_4
* cell instance $21784 r0 *1 45.885,84.77
X$21784 2149 VIA_via2_5
* cell instance $21785 r0 *1 44.175,84.35
X$21785 2149 VIA_via1_4
* cell instance $21786 r0 *1 44.175,84.35
X$21786 2149 VIA_via2_5
* cell instance $21787 r0 *1 43.795,85.05
X$21787 2149 VIA_via1_4
* cell instance $21788 r0 *1 47.025,86.03
X$21788 2149 VIA_via1_4
* cell instance $21789 r0 *1 40.565,86.03
X$21789 2149 VIA_via1_4
* cell instance $21790 r0 *1 40.565,86.03
X$21790 2149 VIA_via2_5
* cell instance $21791 r0 *1 52.535,80.99
X$21791 2150 VIA_via1_7
* cell instance $21792 r0 *1 52.725,81.97
X$21792 2150 VIA_via1_4
* cell instance $21793 r0 *1 57.475,95.41
X$21793 2151 VIA_via1_7
* cell instance $21794 r0 *1 56.905,85.89
X$21794 2151 VIA_via2_5
* cell instance $21795 r0 *1 58.235,93.31
X$21795 2151 VIA_via2_5
* cell instance $21796 r0 *1 56.905,87.57
X$21796 2151 VIA_via2_5
* cell instance $21797 r0 *1 55.575,84.49
X$21797 2151 VIA_via2_5
* cell instance $21798 r0 *1 56.145,85.75
X$21798 2151 VIA_via2_5
* cell instance $21799 r0 *1 58.235,87.57
X$21799 2151 VIA_via2_5
* cell instance $21800 r0 *1 57.475,93.31
X$21800 2151 VIA_via2_5
* cell instance $21801 r0 *1 55.195,93.17
X$21801 2151 VIA_via1_4
* cell instance $21802 r0 *1 55.195,93.31
X$21802 2151 VIA_via2_5
* cell instance $21803 r0 *1 57.665,84.77
X$21803 2151 VIA_via1_4
* cell instance $21804 r0 *1 57.665,84.77
X$21804 2151 VIA_via2_5
* cell instance $21805 r0 *1 56.145,84.77
X$21805 2151 VIA_via1_4
* cell instance $21806 r0 *1 56.145,84.77
X$21806 2151 VIA_via2_5
* cell instance $21807 r0 *1 57.855,81.97
X$21807 2151 VIA_via1_4
* cell instance $21808 r0 *1 55.385,81.97
X$21808 2151 VIA_via1_4
* cell instance $21809 r0 *1 56.145,87.57
X$21809 2151 VIA_via1_4
* cell instance $21810 r0 *1 56.145,87.57
X$21810 2151 VIA_via2_5
* cell instance $21811 r0 *1 58.235,90.37
X$21811 2151 VIA_via1_4
* cell instance $21812 r0 *1 58.805,81.41
X$21812 2152 VIA_via1_7
* cell instance $21813 r0 *1 59.185,80.43
X$21813 2152 VIA_via1_4
* cell instance $21814 r0 *1 64.505,80.71
X$21814 2153 VIA_via1_7
* cell instance $21815 r0 *1 64.505,80.71
X$21815 2153 VIA_via2_5
* cell instance $21816 r0 *1 65.835,80.71
X$21816 2153 VIA_via1_7
* cell instance $21817 r0 *1 65.835,80.71
X$21817 2153 VIA_via2_5
* cell instance $21818 r0 *1 64.125,80.71
X$21818 2153 VIA_via2_5
* cell instance $21819 r0 *1 64.125,79.03
X$21819 2153 VIA_via1_4
* cell instance $21820 r0 *1 65.455,81.69
X$21820 2154 VIA_via1_7
* cell instance $21821 r0 *1 70.775,92.61
X$21821 2154 VIA_via2_5
* cell instance $21822 r0 *1 71.155,84.91
X$21822 2154 VIA_via2_5
* cell instance $21823 r0 *1 64.125,84.91
X$21823 2154 VIA_via2_5
* cell instance $21824 r0 *1 69.255,80.71
X$21824 2154 VIA_via2_5
* cell instance $21825 r0 *1 65.455,80.85
X$21825 2154 VIA_via2_5
* cell instance $21826 r0 *1 73.815,92.61
X$21826 2154 VIA_via2_5
* cell instance $21827 r0 *1 69.255,80.43
X$21827 2154 VIA_via1_4
* cell instance $21828 r0 *1 64.885,80.85
X$21828 2154 VIA_via1_4
* cell instance $21829 r0 *1 64.885,80.85
X$21829 2154 VIA_via2_5
* cell instance $21830 r0 *1 64.125,84.63
X$21830 2154 VIA_via1_4
* cell instance $21831 r0 *1 65.455,84.91
X$21831 2154 VIA_via1_4
* cell instance $21832 r0 *1 65.455,84.91
X$21832 2154 VIA_via2_5
* cell instance $21833 r0 *1 73.815,93.31
X$21833 2154 VIA_via1_4
* cell instance $21834 r0 *1 70.775,91.77
X$21834 2154 VIA_via1_4
* cell instance $21835 r0 *1 63.745,91.21
X$21835 2155 VIA_via1_7
* cell instance $21836 r0 *1 63.745,92.19
X$21836 2155 VIA_via1_7
* cell instance $21837 r0 *1 65.075,82.11
X$21837 2155 VIA_via2_5
* cell instance $21838 r0 *1 63.745,93.17
X$21838 2155 VIA_via2_5
* cell instance $21839 r0 *1 65.265,93.17
X$21839 2155 VIA_via2_5
* cell instance $21840 r0 *1 67.735,81.97
X$21840 2155 VIA_via1_4
* cell instance $21841 r0 *1 67.735,81.97
X$21841 2155 VIA_via2_5
* cell instance $21842 r0 *1 65.075,83.23
X$21842 2155 VIA_via1_4
* cell instance $21843 r0 *1 65.075,83.09
X$21843 2155 VIA_via2_5
* cell instance $21844 r0 *1 63.745,83.23
X$21844 2155 VIA_via1_4
* cell instance $21845 r0 *1 63.745,83.09
X$21845 2155 VIA_via2_5
* cell instance $21846 r0 *1 65.265,94.43
X$21846 2155 VIA_via1_4
* cell instance $21847 r0 *1 80.085,91.35
X$21847 2156 VIA_via2_5
* cell instance $21848 r0 *1 76.475,91.35
X$21848 2156 VIA_via2_5
* cell instance $21849 r0 *1 82.935,82.11
X$21849 2156 VIA_via2_5
* cell instance $21850 r0 *1 67.355,83.93
X$21850 2156 VIA_via2_5
* cell instance $21851 r0 *1 76.475,84.35
X$21851 2156 VIA_via2_5
* cell instance $21852 r0 *1 76.475,83.93
X$21852 2156 VIA_via2_5
* cell instance $21853 r0 *1 81.985,84.35
X$21853 2156 VIA_via2_5
* cell instance $21854 r0 *1 67.165,81.97
X$21854 2156 VIA_via1_4
* cell instance $21855 r0 *1 76.095,93.17
X$21855 2156 VIA_via1_4
* cell instance $21856 r0 *1 83.125,81.83
X$21856 2156 VIA_via1_4
* cell instance $21857 r0 *1 81.985,82.11
X$21857 2156 VIA_via1_4
* cell instance $21858 r0 *1 81.985,82.11
X$21858 2156 VIA_via2_5
* cell instance $21859 r0 *1 80.085,91.63
X$21859 2156 VIA_via1_4
* cell instance $21860 r0 *1 67.925,80.57
X$21860 2157 VIA_via1_7
* cell instance $21861 r0 *1 67.925,81.97
X$21861 2157 VIA_via1_4
* cell instance $21862 r0 *1 67.545,82.25
X$21862 2157 VIA_via1_4
* cell instance $21863 r0 *1 73.245,80.99
X$21863 2158 VIA_via1_7
* cell instance $21864 r0 *1 73.435,82.11
X$21864 2158 VIA_via2_5
* cell instance $21865 r0 *1 71.345,81.97
X$21865 2158 VIA_via1_4
* cell instance $21866 r0 *1 71.345,82.11
X$21866 2158 VIA_via2_5
* cell instance $21867 r0 *1 82.365,80.57
X$21867 2159 VIA_via1_7
* cell instance $21868 r0 *1 82.175,81.55
X$21868 2159 VIA_via1_4
* cell instance $21869 r0 *1 73.815,88.13
X$21869 2160 VIA_via2_5
* cell instance $21870 r0 *1 75.525,87.57
X$21870 2160 VIA_via2_5
* cell instance $21871 r0 *1 84.455,81.69
X$21871 2160 VIA_via2_5
* cell instance $21872 r0 *1 83.505,81.69
X$21872 2160 VIA_via2_5
* cell instance $21873 r0 *1 82.745,81.69
X$21873 2160 VIA_via2_5
* cell instance $21874 r0 *1 79.325,85.75
X$21874 2160 VIA_via2_5
* cell instance $21875 r0 *1 75.525,85.75
X$21875 2160 VIA_via2_5
* cell instance $21876 r0 *1 79.325,85.19
X$21876 2160 VIA_via2_5
* cell instance $21877 r0 *1 82.555,85.19
X$21877 2160 VIA_via2_5
* cell instance $21878 r0 *1 80.465,81.69
X$21878 2160 VIA_via2_5
* cell instance $21879 r0 *1 79.135,89.95
X$21879 2160 VIA_via1_4
* cell instance $21880 r0 *1 73.815,87.57
X$21880 2160 VIA_via1_4
* cell instance $21881 r0 *1 73.815,87.57
X$21881 2160 VIA_via2_5
* cell instance $21882 r0 *1 73.815,88.83
X$21882 2160 VIA_via1_4
* cell instance $21883 r0 *1 75.525,86.03
X$21883 2160 VIA_via1_4
* cell instance $21884 r0 *1 83.505,81.97
X$21884 2160 VIA_via1_4
* cell instance $21885 r0 *1 82.745,81.97
X$21885 2160 VIA_via1_4
* cell instance $21886 r0 *1 84.455,80.43
X$21886 2160 VIA_via1_4
* cell instance $21887 r0 *1 79.515,86.03
X$21887 2160 VIA_via1_4
* cell instance $21888 r0 *1 80.465,79.17
X$21888 2160 VIA_via1_4
* cell instance $21889 r0 *1 89.585,80.99
X$21889 2161 VIA_via1_7
* cell instance $21890 r0 *1 86.545,84.49
X$21890 2161 VIA_via2_5
* cell instance $21891 r0 *1 90.345,84.49
X$21891 2161 VIA_via2_5
* cell instance $21892 r0 *1 89.205,84.49
X$21892 2161 VIA_via2_5
* cell instance $21893 r0 *1 88.445,88.69
X$21893 2161 VIA_via2_5
* cell instance $21894 r0 *1 86.735,86.03
X$21894 2161 VIA_via1_4
* cell instance $21895 r0 *1 86.545,88.69
X$21895 2161 VIA_via1_4
* cell instance $21896 r0 *1 86.545,88.69
X$21896 2161 VIA_via2_5
* cell instance $21897 r0 *1 88.065,90.37
X$21897 2161 VIA_via1_4
* cell instance $21898 r0 *1 90.345,84.77
X$21898 2161 VIA_via1_4
* cell instance $21899 r0 *1 96.995,81.83
X$21899 2162 VIA_via1_4
* cell instance $21900 r0 *1 96.995,81.83
X$21900 2162 VIA_via2_5
* cell instance $21901 r0 *1 97.535,81.83
X$21901 2162 VIA_via3_2
* cell instance $21902 r0 *1 97.535,81.83
X$21902 2162 VIA_via4_0
* cell instance $21903 r0 *1 96.995,80.99
X$21903 2163 VIA_via1_7
* cell instance $21904 r0 *1 96.995,80.99
X$21904 2163 VIA_via2_5
* cell instance $21905 r0 *1 97.535,81.27
X$21905 2163 VIA_via4_0
* cell instance $21906 r0 *1 97.535,80.99
X$21906 2163 VIA_via3_2
* cell instance $21907 r0 *1 96.425,80.71
X$21907 2164 VIA_via1_4
* cell instance $21908 r0 *1 96.425,80.71
X$21908 2164 VIA_via2_5
* cell instance $21909 r0 *1 97.255,80.71
X$21909 2164 VIA_via4_0
* cell instance $21910 r0 *1 97.255,80.71
X$21910 2164 VIA_via3_2
* cell instance $21911 r0 *1 4.465,82.39
X$21911 2165 VIA_via2_5
* cell instance $21912 r0 *1 6.175,82.39
X$21912 2165 VIA_via2_5
* cell instance $21913 r0 *1 4.465,80.85
X$21913 2165 VIA_via2_5
* cell instance $21914 r0 *1 6.175,81.97
X$21914 2165 VIA_via1_4
* cell instance $21915 r0 *1 5.035,80.85
X$21915 2165 VIA_via1_4
* cell instance $21916 r0 *1 5.035,80.85
X$21916 2165 VIA_via2_5
* cell instance $21917 r0 *1 4.465,83.23
X$21917 2165 VIA_via1_4
* cell instance $21918 r0 *1 12.825,81.41
X$21918 2166 VIA_via1_7
* cell instance $21919 r0 *1 12.825,74.83
X$21919 2166 VIA_via1_4
* cell instance $21920 r0 *1 24.605,80.99
X$21920 2167 VIA_via1_7
* cell instance $21921 r0 *1 24.605,81.83
X$21921 2167 VIA_via2_5
* cell instance $21922 r0 *1 23.085,81.97
X$21922 2167 VIA_via1_4
* cell instance $21923 r0 *1 23.085,81.83
X$21923 2167 VIA_via2_5
* cell instance $21924 r0 *1 76.665,80.57
X$21924 2168 VIA_via1_4
* cell instance $21925 r0 *1 76.665,80.57
X$21925 2168 VIA_via2_5
* cell instance $21926 r0 *1 75.525,80.43
X$21926 2168 VIA_via1_4
* cell instance $21927 r0 *1 75.525,80.57
X$21927 2168 VIA_via2_5
* cell instance $21928 r0 *1 31.825,80.71
X$21928 2169 VIA_via1_7
* cell instance $21929 r0 *1 31.825,81.41
X$21929 2169 VIA_via2_5
* cell instance $21930 r0 *1 30.495,81.41
X$21930 2169 VIA_via2_5
* cell instance $21931 r0 *1 30.305,95.97
X$21931 2169 VIA_via1_4
* cell instance $21932 r0 *1 72.675,82.81
X$21932 2170 VIA_via1_7
* cell instance $21933 r0 *1 72.865,80.43
X$21933 2170 VIA_via1_4
* cell instance $21934 r0 *1 72.865,80.57
X$21934 2170 VIA_via2_5
* cell instance $21935 r0 *1 70.775,80.43
X$21935 2170 VIA_via1_4
* cell instance $21936 r0 *1 70.775,80.57
X$21936 2170 VIA_via2_5
* cell instance $21937 r0 *1 67.735,80.99
X$21937 2171 VIA_via1_7
* cell instance $21938 r0 *1 67.735,80.99
X$21938 2171 VIA_via2_5
* cell instance $21939 r0 *1 68.115,80.99
X$21939 2171 VIA_via2_5
* cell instance $21940 r0 *1 68.115,81.97
X$21940 2171 VIA_via1_4
* cell instance $21941 r0 *1 69.065,80.57
X$21941 2172 VIA_via1_4
* cell instance $21942 r0 *1 69.065,80.57
X$21942 2172 VIA_via2_5
* cell instance $21943 r0 *1 62.605,80.43
X$21943 2172 VIA_via1_4
* cell instance $21944 r0 *1 62.605,80.57
X$21944 2172 VIA_via2_5
* cell instance $21945 r0 *1 38.095,81.41
X$21945 2173 VIA_via1_7
* cell instance $21946 r0 *1 38.095,81.41
X$21946 2173 VIA_via2_5
* cell instance $21947 r0 *1 36.765,81.41
X$21947 2173 VIA_via2_5
* cell instance $21948 r0 *1 36.765,80.43
X$21948 2173 VIA_via1_4
* cell instance $21949 r0 *1 3.515,82.81
X$21949 2174 VIA_via1_7
* cell instance $21950 r0 *1 2.945,81.97
X$21950 2174 VIA_via1_4
* cell instance $21951 r0 *1 5.225,83.23
X$21951 2175 VIA_via2_5
* cell instance $21952 r0 *1 3.135,83.23
X$21952 2175 VIA_via1_4
* cell instance $21953 r0 *1 3.135,83.23
X$21953 2175 VIA_via2_5
* cell instance $21954 r0 *1 5.225,82.25
X$21954 2175 VIA_via1_4
* cell instance $21955 r0 *1 5.605,81.97
X$21955 2175 VIA_via1_4
* cell instance $21956 r0 *1 17.385,82.95
X$21956 2176 VIA_via2_5
* cell instance $21957 r0 *1 13.775,82.95
X$21957 2176 VIA_via2_5
* cell instance $21958 r0 *1 15.675,82.95
X$21958 2176 VIA_via1_4
* cell instance $21959 r0 *1 15.675,82.95
X$21959 2176 VIA_via2_5
* cell instance $21960 r0 *1 17.385,80.43
X$21960 2176 VIA_via1_4
* cell instance $21961 r0 *1 13.775,81.97
X$21961 2176 VIA_via1_4
* cell instance $21962 r0 *1 21.565,84.77
X$21962 2177 VIA_via1_4
* cell instance $21963 r0 *1 21.755,80.43
X$21963 2177 VIA_via1_4
* cell instance $21964 r0 *1 21.755,82.95
X$21964 2177 VIA_via1_4
* cell instance $21965 r0 *1 25.745,84.77
X$21965 2178 VIA_via2_5
* cell instance $21966 r0 *1 23.275,84.77
X$21966 2178 VIA_via2_5
* cell instance $21967 r0 *1 25.745,83.65
X$21967 2178 VIA_via1_4
* cell instance $21968 r0 *1 26.315,80.43
X$21968 2178 VIA_via1_4
* cell instance $21969 r0 *1 23.085,84.77
X$21969 2178 VIA_via1_4
* cell instance $21970 r0 *1 28.975,83.79
X$21970 2179 VIA_via1_7
* cell instance $21971 r0 *1 28.785,84.77
X$21971 2179 VIA_via1_4
* cell instance $21972 r0 *1 35.245,82.25
X$21972 2180 VIA_via2_5
* cell instance $21973 r0 *1 33.345,82.25
X$21973 2180 VIA_via2_5
* cell instance $21974 r0 *1 33.345,83.23
X$21974 2180 VIA_via1_4
* cell instance $21975 r0 *1 35.245,80.43
X$21975 2180 VIA_via1_4
* cell instance $21976 r0 *1 34.675,82.25
X$21976 2180 VIA_via1_4
* cell instance $21977 r0 *1 34.675,82.25
X$21977 2180 VIA_via2_5
* cell instance $21978 r0 *1 47.975,82.11
X$21978 2181 VIA_via2_5
* cell instance $21979 r0 *1 47.975,83.23
X$21979 2181 VIA_via2_5
* cell instance $21980 r0 *1 50.445,82.11
X$21980 2181 VIA_via1_4
* cell instance $21981 r0 *1 50.445,82.11
X$21981 2181 VIA_via2_5
* cell instance $21982 r0 *1 47.975,79.17
X$21982 2181 VIA_via1_4
* cell instance $21983 r0 *1 48.925,83.23
X$21983 2181 VIA_via1_4
* cell instance $21984 r0 *1 48.925,83.23
X$21984 2181 VIA_via2_5
* cell instance $21985 r0 *1 59.185,95.41
X$21985 2182 VIA_via1_7
* cell instance $21986 r0 *1 53.295,92.89
X$21986 2182 VIA_via2_5
* cell instance $21987 r0 *1 53.295,94.43
X$21987 2182 VIA_via2_5
* cell instance $21988 r0 *1 58.615,92.89
X$21988 2182 VIA_via2_5
* cell instance $21989 r0 *1 48.925,94.43
X$21989 2182 VIA_via2_5
* cell instance $21990 r0 *1 58.615,94.43
X$21990 2182 VIA_via1_4
* cell instance $21991 r0 *1 50.445,94.43
X$21991 2182 VIA_via1_4
* cell instance $21992 r0 *1 50.445,94.43
X$21992 2182 VIA_via2_5
* cell instance $21993 r0 *1 53.295,93.17
X$21993 2182 VIA_via1_4
* cell instance $21994 r0 *1 49.495,83.23
X$21994 2182 VIA_via1_4
* cell instance $21995 r0 *1 48.355,83.23
X$21995 2182 VIA_via1_4
* cell instance $21996 r0 *1 48.355,80.43
X$21996 2182 VIA_via1_4
* cell instance $21997 r0 *1 48.925,93.17
X$21997 2182 VIA_via1_4
* cell instance $21998 r0 *1 52.915,78.19
X$21998 2183 VIA_via1_7
* cell instance $21999 r0 *1 51.585,81.97
X$21999 2183 VIA_via2_5
* cell instance $22000 r0 *1 52.915,81.97
X$22000 2183 VIA_via2_5
* cell instance $22001 r0 *1 51.775,95.97
X$22001 2183 VIA_via1_4
* cell instance $22002 r0 *1 52.725,84.07
X$22002 2184 VIA_via2_5
* cell instance $22003 r0 *1 52.155,84.07
X$22003 2184 VIA_via2_5
* cell instance $22004 r0 *1 52.155,84.77
X$22004 2184 VIA_via1_4
* cell instance $22005 r0 *1 52.915,82.95
X$22005 2184 VIA_via1_4
* cell instance $22006 r0 *1 68.305,85.61
X$22006 2185 VIA_via1_7
* cell instance $22007 r0 *1 68.305,85.61
X$22007 2185 VIA_via2_5
* cell instance $22008 r0 *1 67.545,85.61
X$22008 2185 VIA_via2_5
* cell instance $22009 r0 *1 61.655,83.23
X$22009 2185 VIA_via2_5
* cell instance $22010 r0 *1 66.405,83.23
X$22010 2185 VIA_via2_5
* cell instance $22011 r0 *1 62.605,83.23
X$22011 2185 VIA_via2_5
* cell instance $22012 r0 *1 67.545,84.77
X$22012 2185 VIA_via1_4
* cell instance $22013 r0 *1 67.545,84.77
X$22013 2185 VIA_via2_5
* cell instance $22014 r0 *1 63.555,83.23
X$22014 2185 VIA_via1_4
* cell instance $22015 r0 *1 63.555,83.23
X$22015 2185 VIA_via2_5
* cell instance $22016 r0 *1 64.885,83.23
X$22016 2185 VIA_via1_4
* cell instance $22017 r0 *1 64.885,83.23
X$22017 2185 VIA_via2_5
* cell instance $22018 r0 *1 66.405,84.77
X$22018 2185 VIA_via1_4
* cell instance $22019 r0 *1 66.405,84.77
X$22019 2185 VIA_via2_5
* cell instance $22020 r0 *1 61.655,84.77
X$22020 2185 VIA_via1_4
* cell instance $22021 r0 *1 62.605,86.03
X$22021 2185 VIA_via1_4
* cell instance $22022 r0 *1 72.295,90.09
X$22022 2186 VIA_via1_7
* cell instance $22023 r0 *1 70.395,83.51
X$22023 2186 VIA_via1_7
* cell instance $22024 r0 *1 72.105,83.79
X$22024 2186 VIA_via2_5
* cell instance $22025 r0 *1 70.395,83.79
X$22025 2186 VIA_via2_5
* cell instance $22026 r0 *1 69.255,83.79
X$22026 2186 VIA_via2_5
* cell instance $22027 r0 *1 69.255,82.39
X$22027 2186 VIA_via2_5
* cell instance $22028 r0 *1 66.215,82.39
X$22028 2186 VIA_via2_5
* cell instance $22029 r0 *1 65.645,82.39
X$22029 2186 VIA_via2_5
* cell instance $22030 r0 *1 69.255,81.97
X$22030 2186 VIA_via1_4
* cell instance $22031 r0 *1 65.645,81.97
X$22031 2186 VIA_via1_4
* cell instance $22032 r0 *1 66.215,80.43
X$22032 2186 VIA_via1_4
* cell instance $22033 r0 *1 73.245,82.25
X$22033 2187 VIA_via2_5
* cell instance $22034 r0 *1 72.105,82.25
X$22034 2187 VIA_via2_5
* cell instance $22035 r0 *1 72.675,88.83
X$22035 2187 VIA_via2_5
* cell instance $22036 r0 *1 71.915,83.23
X$22036 2187 VIA_via1_4
* cell instance $22037 r0 *1 72.105,83.23
X$22037 2187 VIA_via1_4
* cell instance $22038 r0 *1 73.625,82.25
X$22038 2187 VIA_via1_4
* cell instance $22039 r0 *1 73.625,82.25
X$22039 2187 VIA_via2_5
* cell instance $22040 r0 *1 72.675,90.37
X$22040 2187 VIA_via1_4
* cell instance $22041 r0 *1 73.435,87.57
X$22041 2187 VIA_via1_4
* cell instance $22042 r0 *1 72.105,88.83
X$22042 2187 VIA_via1_4
* cell instance $22043 r0 *1 72.105,88.83
X$22043 2187 VIA_via2_5
* cell instance $22044 r0 *1 78.375,83.37
X$22044 2188 VIA_via1_4
* cell instance $22045 r0 *1 78.375,83.23
X$22045 2188 VIA_via2_5
* cell instance $22046 r0 *1 79.515,83.23
X$22046 2188 VIA_via1_4
* cell instance $22047 r0 *1 79.515,83.23
X$22047 2188 VIA_via2_5
* cell instance $22048 r0 *1 78.375,84.35
X$22048 2188 VIA_via1_4
* cell instance $22049 r0 *1 79.705,83.23
X$22049 2188 VIA_via1_4
* cell instance $22050 r0 *1 78.945,87.15
X$22050 2189 VIA_via2_5
* cell instance $22051 r0 *1 76.665,87.15
X$22051 2189 VIA_via2_5
* cell instance $22052 r0 *1 76.665,90.23
X$22052 2189 VIA_via1_4
* cell instance $22053 r0 *1 78.755,83.37
X$22053 2189 VIA_via1_4
* cell instance $22054 r0 *1 87.305,89.95
X$22054 2190 VIA_via2_5
* cell instance $22055 r0 *1 83.885,85.89
X$22055 2190 VIA_via2_5
* cell instance $22056 r0 *1 87.495,85.89
X$22056 2190 VIA_via2_5
* cell instance $22057 r0 *1 78.945,88.55
X$22057 2190 VIA_via2_5
* cell instance $22058 r0 *1 78.945,88.27
X$22058 2190 VIA_via2_5
* cell instance $22059 r0 *1 77.045,88.27
X$22059 2190 VIA_via2_5
* cell instance $22060 r0 *1 85.215,89.95
X$22060 2190 VIA_via2_5
* cell instance $22061 r0 *1 75.715,87.43
X$22061 2190 VIA_via2_5
* cell instance $22062 r0 *1 83.125,82.39
X$22062 2190 VIA_via2_5
* cell instance $22063 r0 *1 85.215,88.55
X$22063 2190 VIA_via2_5
* cell instance $22064 r0 *1 83.885,88.55
X$22064 2190 VIA_via2_5
* cell instance $22065 r0 *1 83.125,85.75
X$22065 2190 VIA_via2_5
* cell instance $22066 r0 *1 82.175,82.39
X$22066 2190 VIA_via2_5
* cell instance $22067 r0 *1 77.045,90.37
X$22067 2190 VIA_via1_4
* cell instance $22068 r0 *1 77.045,90.51
X$22068 2190 VIA_via2_5
* cell instance $22069 r0 *1 78.945,93.17
X$22069 2190 VIA_via1_4
* cell instance $22070 r0 *1 74.005,87.57
X$22070 2190 VIA_via1_4
* cell instance $22071 r0 *1 74.005,87.43
X$22071 2190 VIA_via2_5
* cell instance $22072 r0 *1 75.715,86.03
X$22072 2190 VIA_via1_4
* cell instance $22073 r0 *1 73.625,90.37
X$22073 2190 VIA_via1_4
* cell instance $22074 r0 *1 73.625,90.51
X$22074 2190 VIA_via2_5
* cell instance $22075 r0 *1 82.175,82.11
X$22075 2190 VIA_via1_4
* cell instance $22076 r0 *1 83.315,82.11
X$22076 2190 VIA_via1_4
* cell instance $22077 r0 *1 77.045,87.57
X$22077 2190 VIA_via1_4
* cell instance $22078 r0 *1 77.045,87.43
X$22078 2190 VIA_via2_5
* cell instance $22079 r0 *1 85.215,88.83
X$22079 2190 VIA_via1_4
* cell instance $22080 r0 *1 87.305,90.37
X$22080 2190 VIA_via1_4
* cell instance $22081 r0 *1 87.495,84.77
X$22081 2190 VIA_via1_4
* cell instance $22082 r0 *1 83.315,84.21
X$22082 2191 VIA_via1_7
* cell instance $22083 r0 *1 83.505,83.23
X$22083 2191 VIA_via1_4
* cell instance $22084 r0 *1 86.165,92.61
X$22084 2192 VIA_via2_5
* cell instance $22085 r0 *1 84.265,88.27
X$22085 2192 VIA_via2_5
* cell instance $22086 r0 *1 83.125,92.61
X$22086 2192 VIA_via2_5
* cell instance $22087 r0 *1 83.125,95.97
X$22087 2192 VIA_via1_4
* cell instance $22088 r0 *1 84.265,84.77
X$22088 2192 VIA_via1_4
* cell instance $22089 r0 *1 85.595,86.03
X$22089 2192 VIA_via1_4
* cell instance $22090 r0 *1 86.355,91.63
X$22090 2192 VIA_via1_4
* cell instance $22091 r0 *1 85.785,83.65
X$22091 2192 VIA_via1_4
* cell instance $22092 r0 *1 85.495,88.27
X$22092 2192 VIA_via3_2
* cell instance $22093 r0 *1 85.405,88.27
X$22093 2192 VIA_via2_5
* cell instance $22094 r0 *1 85.495,92.61
X$22094 2192 VIA_via3_2
* cell instance $22095 r0 *1 87.305,83.79
X$22095 2193 VIA_via1_7
* cell instance $22096 r0 *1 85.785,85.75
X$22096 2193 VIA_via2_5
* cell instance $22097 r0 *1 86.735,85.75
X$22097 2193 VIA_via2_5
* cell instance $22098 r0 *1 85.595,90.65
X$22098 2193 VIA_via2_5
* cell instance $22099 r0 *1 85.595,88.69
X$22099 2193 VIA_via2_5
* cell instance $22100 r0 *1 85.595,90.37
X$22100 2193 VIA_via1_4
* cell instance $22101 r0 *1 85.975,88.83
X$22101 2193 VIA_via1_4
* cell instance $22102 r0 *1 85.975,88.83
X$22102 2193 VIA_via2_5
* cell instance $22103 r0 *1 86.545,90.51
X$22103 2193 VIA_via1_4
* cell instance $22104 r0 *1 86.545,90.65
X$22104 2193 VIA_via2_5
* cell instance $22105 r0 *1 86.735,84.77
X$22105 2193 VIA_via1_4
* cell instance $22106 r0 *1 89.015,83.79
X$22106 2194 VIA_via1_7
* cell instance $22107 r0 *1 88.825,84.77
X$22107 2194 VIA_via1_4
* cell instance $22108 r0 *1 91.105,83.23
X$22108 2195 VIA_via1_4
* cell instance $22109 r0 *1 90.915,82.95
X$22109 2195 VIA_via1_4
* cell instance $22110 r0 *1 96.615,86.03
X$22110 2196 VIA_via1_4
* cell instance $22111 r0 *1 96.615,84.77
X$22111 2196 VIA_via1_4
* cell instance $22112 r0 *1 96.425,83.65
X$22112 2196 VIA_via1_4
* cell instance $22113 r0 *1 4.845,82.81
X$22113 2197 VIA_via1_7
* cell instance $22114 r0 *1 4.845,82.81
X$22114 2197 VIA_via2_5
* cell instance $22115 r0 *1 2.755,82.81
X$22115 2197 VIA_via2_5
* cell instance $22116 r0 *1 2.755,80.43
X$22116 2197 VIA_via1_4
* cell instance $22117 r0 *1 8.645,83.23
X$22117 2198 VIA_via2_5
* cell instance $22118 r0 *1 8.645,81.83
X$22118 2198 VIA_via1_4
* cell instance $22119 r0 *1 6.935,83.23
X$22119 2198 VIA_via1_4
* cell instance $22120 r0 *1 6.935,83.23
X$22120 2198 VIA_via2_5
* cell instance $22121 r0 *1 13.775,95.41
X$22121 2199 VIA_via1_7
* cell instance $22122 r0 *1 6.745,91.91
X$22122 2199 VIA_via2_5
* cell instance $22123 r0 *1 8.645,91.91
X$22123 2199 VIA_via2_5
* cell instance $22124 r0 *1 13.585,83.09
X$22124 2199 VIA_via2_5
* cell instance $22125 r0 *1 13.205,83.09
X$22125 2199 VIA_via2_5
* cell instance $22126 r0 *1 13.395,91.63
X$22126 2199 VIA_via2_5
* cell instance $22127 r0 *1 13.585,91.21
X$22127 2199 VIA_via2_5
* cell instance $22128 r0 *1 13.585,86.03
X$22128 2199 VIA_via1_4
* cell instance $22129 r0 *1 13.015,93.17
X$22129 2199 VIA_via1_4
* cell instance $22130 r0 *1 9.595,83.23
X$22130 2199 VIA_via1_4
* cell instance $22131 r0 *1 9.595,83.09
X$22131 2199 VIA_via2_5
* cell instance $22132 r0 *1 6.745,94.43
X$22132 2199 VIA_via1_4
* cell instance $22133 r0 *1 8.645,91.63
X$22133 2199 VIA_via1_4
* cell instance $22134 r0 *1 10.545,91.63
X$22134 2199 VIA_via1_4
* cell instance $22135 r0 *1 10.545,91.63
X$22135 2199 VIA_via2_5
* cell instance $22136 r0 *1 13.205,81.97
X$22136 2199 VIA_via1_4
* cell instance $22137 r0 *1 92.245,83.23
X$22137 2200 VIA_via1_4
* cell instance $22138 r0 *1 92.245,83.23
X$22138 2200 VIA_via2_5
* cell instance $22139 r0 *1 94.145,83.23
X$22139 2200 VIA_via1_4
* cell instance $22140 r0 *1 94.145,83.23
X$22140 2200 VIA_via2_5
* cell instance $22141 r0 *1 92.435,82.39
X$22141 2201 VIA_via2_5
* cell instance $22142 r0 *1 91.865,82.39
X$22142 2201 VIA_via2_5
* cell instance $22143 r0 *1 91.865,83.23
X$22143 2201 VIA_via1_4
* cell instance $22144 r0 *1 92.435,81.83
X$22144 2201 VIA_via1_4
* cell instance $22145 r0 *1 6.555,82.11
X$22145 2202 VIA_via1_4
* cell instance $22146 r0 *1 6.555,82.11
X$22146 2202 VIA_via2_5
* cell instance $22147 r0 *1 12.445,81.97
X$22147 2202 VIA_via1_4
* cell instance $22148 r0 *1 12.445,82.11
X$22148 2202 VIA_via2_5
* cell instance $22149 r0 *1 14.155,82.39
X$22149 2203 VIA_via1_7
* cell instance $22150 r0 *1 14.155,82.39
X$22150 2203 VIA_via2_5
* cell instance $22151 r0 *1 13.395,82.39
X$22151 2203 VIA_via2_5
* cell instance $22152 r0 *1 13.395,83.23
X$22152 2203 VIA_via1_4
* cell instance $22153 r0 *1 89.965,83.23
X$22153 2204 VIA_via1_4
* cell instance $22154 r0 *1 90.345,83.23
X$22154 2204 VIA_via1_4
* cell instance $22155 r0 *1 29.355,80.99
X$22155 2205 VIA_via1_7
* cell instance $22156 r0 *1 29.355,82.11
X$22156 2205 VIA_via2_5
* cell instance $22157 r0 *1 26.885,81.97
X$22157 2205 VIA_via1_4
* cell instance $22158 r0 *1 26.885,82.11
X$22158 2205 VIA_via2_5
* cell instance $22159 r0 *1 30.685,83.23
X$22159 2206 VIA_via2_5
* cell instance $22160 r0 *1 30.305,83.23
X$22160 2206 VIA_via2_5
* cell instance $22161 r0 *1 30.305,80.43
X$22161 2206 VIA_via1_4
* cell instance $22162 r0 *1 28.595,83.23
X$22162 2206 VIA_via1_4
* cell instance $22163 r0 *1 28.595,83.23
X$22163 2206 VIA_via2_5
* cell instance $22164 r0 *1 31.065,84.35
X$22164 2206 VIA_via1_4
* cell instance $22165 r0 *1 89.395,82.39
X$22165 2207 VIA_via1_7
* cell instance $22166 r0 *1 89.395,83.23
X$22166 2207 VIA_via1_4
* cell instance $22167 r0 *1 89.395,83.23
X$22167 2207 VIA_via2_5
* cell instance $22168 r0 *1 86.925,83.23
X$22168 2207 VIA_via1_4
* cell instance $22169 r0 *1 86.925,83.23
X$22169 2207 VIA_via2_5
* cell instance $22170 r0 *1 33.725,82.81
X$22170 2208 VIA_via1_7
* cell instance $22171 r0 *1 33.725,82.81
X$22171 2208 VIA_via2_5
* cell instance $22172 r0 *1 32.395,82.81
X$22172 2208 VIA_via2_5
* cell instance $22173 r0 *1 32.395,81.97
X$22173 2208 VIA_via1_4
* cell instance $22174 r0 *1 49.305,82.81
X$22174 2209 VIA_via1_7
* cell instance $22175 r0 *1 49.305,82.81
X$22175 2209 VIA_via2_5
* cell instance $22176 r0 *1 48.165,82.81
X$22176 2209 VIA_via2_5
* cell instance $22177 r0 *1 48.165,81.97
X$22177 2209 VIA_via1_4
* cell instance $22178 r0 *1 56.335,82.39
X$22178 2210 VIA_via1_7
* cell instance $22179 r0 *1 56.335,82.39
X$22179 2210 VIA_via2_5
* cell instance $22180 r0 *1 54.625,82.39
X$22180 2210 VIA_via2_5
* cell instance $22181 r0 *1 54.625,83.23
X$22181 2210 VIA_via1_4
* cell instance $22182 r0 *1 56.145,81.97
X$22182 2211 VIA_via2_5
* cell instance $22183 r0 *1 56.905,81.97
X$22183 2211 VIA_via2_5
* cell instance $22184 r0 *1 56.145,80.43
X$22184 2211 VIA_via1_4
* cell instance $22185 r0 *1 55.955,81.97
X$22185 2211 VIA_via1_4
* cell instance $22186 r0 *1 55.955,81.97
X$22186 2211 VIA_via2_5
* cell instance $22187 r0 *1 56.905,82.95
X$22187 2211 VIA_via1_4
* cell instance $22188 r0 *1 75.905,80.99
X$22188 2212 VIA_via1_7
* cell instance $22189 r0 *1 75.905,81.97
X$22189 2212 VIA_via1_4
* cell instance $22190 r0 *1 62.795,87.01
X$22190 2213 VIA_via1_7
* cell instance $22191 r0 *1 62.795,87.01
X$22191 2213 VIA_via2_5
* cell instance $22192 r0 *1 61.845,83.37
X$22192 2213 VIA_via2_5
* cell instance $22193 r0 *1 62.795,87.57
X$22193 2213 VIA_via2_5
* cell instance $22194 r0 *1 61.845,87.01
X$22194 2213 VIA_via2_5
* cell instance $22195 r0 *1 63.365,83.37
X$22195 2213 VIA_via1_4
* cell instance $22196 r0 *1 63.365,83.37
X$22196 2213 VIA_via2_5
* cell instance $22197 r0 *1 61.845,84.77
X$22197 2213 VIA_via1_4
* cell instance $22198 r0 *1 64.125,87.57
X$22198 2213 VIA_via1_4
* cell instance $22199 r0 *1 64.125,87.57
X$22199 2213 VIA_via2_5
* cell instance $22200 r0 *1 69.065,82.39
X$22200 2214 VIA_via1_7
* cell instance $22201 r0 *1 69.065,82.53
X$22201 2214 VIA_via2_5
* cell instance $22202 r0 *1 68.495,82.53
X$22202 2214 VIA_via2_5
* cell instance $22203 r0 *1 68.495,83.23
X$22203 2214 VIA_via1_4
* cell instance $22204 r0 *1 68.685,81.97
X$22204 2215 VIA_via1_4
* cell instance $22205 r0 *1 68.685,81.97
X$22205 2215 VIA_via2_5
* cell instance $22206 r0 *1 69.825,81.97
X$22206 2215 VIA_via1_4
* cell instance $22207 r0 *1 69.825,81.97
X$22207 2215 VIA_via2_5
* cell instance $22208 r0 *1 10.545,83.79
X$22208 2216 VIA_via1_7
* cell instance $22209 r0 *1 10.355,84.77
X$22209 2216 VIA_via2_5
* cell instance $22210 r0 *1 8.835,84.77
X$22210 2216 VIA_via1_4
* cell instance $22211 r0 *1 8.835,84.77
X$22211 2216 VIA_via2_5
* cell instance $22212 r0 *1 15.105,95.41
X$22212 2217 VIA_via1_7
* cell instance $22213 r0 *1 16.245,92.47
X$22213 2217 VIA_via2_5
* cell instance $22214 r0 *1 22.135,92.47
X$22214 2217 VIA_via2_5
* cell instance $22215 r0 *1 16.245,93.45
X$22215 2217 VIA_via2_5
* cell instance $22216 r0 *1 19.475,92.47
X$22216 2217 VIA_via2_5
* cell instance $22217 r0 *1 14.915,93.45
X$22217 2217 VIA_via2_5
* cell instance $22218 r0 *1 19.475,91.63
X$22218 2217 VIA_via1_4
* cell instance $22219 r0 *1 14.915,93.17
X$22219 2217 VIA_via1_4
* cell instance $22220 r0 *1 16.245,93.17
X$22220 2217 VIA_via1_4
* cell instance $22221 r0 *1 22.135,93.17
X$22221 2217 VIA_via1_4
* cell instance $22222 r0 *1 18.905,84.77
X$22222 2217 VIA_via1_4
* cell instance $22223 r0 *1 18.905,84.77
X$22223 2217 VIA_via2_5
* cell instance $22224 r0 *1 20.995,84.77
X$22224 2217 VIA_via1_4
* cell instance $22225 r0 *1 20.995,84.77
X$22225 2217 VIA_via2_5
* cell instance $22226 r0 *1 22.515,84.77
X$22226 2217 VIA_via1_4
* cell instance $22227 r0 *1 22.515,84.77
X$22227 2217 VIA_via2_5
* cell instance $22228 r0 *1 30.115,95.41
X$22228 2218 VIA_via1_7
* cell instance $22229 r0 *1 27.835,91.63
X$22229 2218 VIA_via2_5
* cell instance $22230 r0 *1 29.735,86.45
X$22230 2218 VIA_via2_5
* cell instance $22231 r0 *1 31.255,86.45
X$22231 2218 VIA_via2_5
* cell instance $22232 r0 *1 29.735,94.01
X$22232 2218 VIA_via2_5
* cell instance $22233 r0 *1 27.835,93.17
X$22233 2218 VIA_via2_5
* cell instance $22234 r0 *1 33.155,94.01
X$22234 2218 VIA_via2_5
* cell instance $22235 r0 *1 32.775,83.79
X$22235 2218 VIA_via2_5
* cell instance $22236 r0 *1 31.255,84.21
X$22236 2218 VIA_via2_5
* cell instance $22237 r0 *1 28.025,83.93
X$22237 2218 VIA_via2_5
* cell instance $22238 r0 *1 29.735,93.17
X$22238 2218 VIA_via1_4
* cell instance $22239 r0 *1 29.735,93.17
X$22239 2218 VIA_via2_5
* cell instance $22240 r0 *1 28.405,93.17
X$22240 2218 VIA_via1_4
* cell instance $22241 r0 *1 28.405,93.17
X$22241 2218 VIA_via2_5
* cell instance $22242 r0 *1 33.155,94.43
X$22242 2218 VIA_via1_4
* cell instance $22243 r0 *1 26.505,91.63
X$22243 2218 VIA_via1_4
* cell instance $22244 r0 *1 26.505,91.63
X$22244 2218 VIA_via2_5
* cell instance $22245 r0 *1 28.025,83.23
X$22245 2218 VIA_via1_4
* cell instance $22246 r0 *1 32.775,83.23
X$22246 2218 VIA_via1_4
* cell instance $22247 r0 *1 31.255,84.77
X$22247 2218 VIA_via1_4
* cell instance $22248 r0 *1 39.235,83.65
X$22248 2219 VIA_via1_4
* cell instance $22249 r0 *1 38.285,84.77
X$22249 2219 VIA_via1_4
* cell instance $22250 r0 *1 39.045,81.97
X$22250 2219 VIA_via1_4
* cell instance $22251 r0 *1 38.665,95.41
X$22251 2220 VIA_via1_7
* cell instance $22252 r0 *1 39.045,84.63
X$22252 2220 VIA_via2_5
* cell instance $22253 r0 *1 39.045,92.47
X$22253 2220 VIA_via2_5
* cell instance $22254 r0 *1 37.525,94.43
X$22254 2220 VIA_via2_5
* cell instance $22255 r0 *1 40.185,92.47
X$22255 2220 VIA_via2_5
* cell instance $22256 r0 *1 40.185,94.29
X$22256 2220 VIA_via2_5
* cell instance $22257 r0 *1 41.135,92.47
X$22257 2220 VIA_via2_5
* cell instance $22258 r0 *1 38.665,94.43
X$22258 2220 VIA_via2_5
* cell instance $22259 r0 *1 39.045,86.03
X$22259 2220 VIA_via2_5
* cell instance $22260 r0 *1 41.325,84.77
X$22260 2220 VIA_via1_4
* cell instance $22261 r0 *1 41.325,84.63
X$22261 2220 VIA_via2_5
* cell instance $22262 r0 *1 37.715,84.77
X$22262 2220 VIA_via1_4
* cell instance $22263 r0 *1 37.715,84.63
X$22263 2220 VIA_via2_5
* cell instance $22264 r0 *1 38.285,86.03
X$22264 2220 VIA_via1_4
* cell instance $22265 r0 *1 38.285,86.03
X$22265 2220 VIA_via2_5
* cell instance $22266 r0 *1 41.135,93.17
X$22266 2220 VIA_via1_4
* cell instance $22267 r0 *1 37.145,95.97
X$22267 2220 VIA_via1_4
* cell instance $22268 r0 *1 40.565,94.43
X$22268 2220 VIA_via1_4
* cell instance $22269 r0 *1 40.565,94.29
X$22269 2220 VIA_via2_5
* cell instance $22270 r0 *1 39.045,93.17
X$22270 2220 VIA_via1_4
* cell instance $22271 r0 *1 42.655,84.35
X$22271 2221 VIA_via2_5
* cell instance $22272 r0 *1 41.895,84.35
X$22272 2221 VIA_via2_5
* cell instance $22273 r0 *1 43.985,84.21
X$22273 2221 VIA_via2_5
* cell instance $22274 r0 *1 41.895,84.77
X$22274 2221 VIA_via1_4
* cell instance $22275 r0 *1 42.655,80.43
X$22275 2221 VIA_via1_4
* cell instance $22276 r0 *1 43.985,83.65
X$22276 2221 VIA_via1_4
* cell instance $22277 r0 *1 62.225,86.17
X$22277 2222 VIA_via2_5
* cell instance $22278 r0 *1 62.415,84.77
X$22278 2222 VIA_via1_4
* cell instance $22279 r0 *1 63.175,86.17
X$22279 2222 VIA_via1_4
* cell instance $22280 r0 *1 63.175,86.17
X$22280 2222 VIA_via2_5
* cell instance $22281 r0 *1 66.215,84.63
X$22281 2223 VIA_via2_5
* cell instance $22282 r0 *1 62.795,86.45
X$22282 2223 VIA_via2_5
* cell instance $22283 r0 *1 66.215,87.57
X$22283 2223 VIA_via2_5
* cell instance $22284 r0 *1 66.215,86.45
X$22284 2223 VIA_via2_5
* cell instance $22285 r0 *1 66.975,87.57
X$22285 2223 VIA_via2_5
* cell instance $22286 r0 *1 65.645,84.77
X$22286 2223 VIA_via1_4
* cell instance $22287 r0 *1 65.645,84.63
X$22287 2223 VIA_via2_5
* cell instance $22288 r0 *1 65.645,83.37
X$22288 2223 VIA_via1_4
* cell instance $22289 r0 *1 66.975,88.55
X$22289 2223 VIA_via1_4
* cell instance $22290 r0 *1 62.795,86.03
X$22290 2223 VIA_via1_4
* cell instance $22291 r0 *1 65.265,87.57
X$22291 2223 VIA_via1_4
* cell instance $22292 r0 *1 65.265,87.57
X$22292 2223 VIA_via2_5
* cell instance $22293 r0 *1 62.605,87.57
X$22293 2223 VIA_via1_4
* cell instance $22294 r0 *1 74.385,84.77
X$22294 2224 VIA_via1_4
* cell instance $22295 r0 *1 74.575,84.77
X$22295 2224 VIA_via1_4
* cell instance $22296 r0 *1 74.575,85.75
X$22296 2224 VIA_via1_4
* cell instance $22297 r0 *1 74.765,85.89
X$22297 2224 VIA_via1_4
* cell instance $22298 r0 *1 92.815,84.91
X$22298 2225 VIA_via2_5
* cell instance $22299 r0 *1 95.665,86.03
X$22299 2225 VIA_via2_5
* cell instance $22300 r0 *1 92.815,86.03
X$22300 2225 VIA_via2_5
* cell instance $22301 r0 *1 91.675,86.03
X$22301 2225 VIA_via2_5
* cell instance $22302 r0 *1 93.575,86.03
X$22302 2225 VIA_via1_4
* cell instance $22303 r0 *1 93.575,86.03
X$22303 2225 VIA_via2_5
* cell instance $22304 r0 *1 95.665,87.15
X$22304 2225 VIA_via1_4
* cell instance $22305 r0 *1 91.675,87.57
X$22305 2225 VIA_via1_4
* cell instance $22306 r0 *1 89.395,85.89
X$22306 2225 VIA_via1_4
* cell instance $22307 r0 *1 89.395,86.03
X$22307 2225 VIA_via2_5
* cell instance $22308 r0 *1 89.775,83.23
X$22308 2225 VIA_via1_4
* cell instance $22309 r0 *1 89.395,84.77
X$22309 2225 VIA_via1_4
* cell instance $22310 r0 *1 91.105,84.77
X$22310 2225 VIA_via1_4
* cell instance $22311 r0 *1 91.105,84.91
X$22311 2225 VIA_via2_5
* cell instance $22312 r0 *1 96.995,84.21
X$22312 2226 VIA_via1_7
* cell instance $22313 r0 *1 96.995,84.21
X$22313 2226 VIA_via2_5
* cell instance $22314 r0 *1 92.625,84.63
X$22314 2226 VIA_via2_5
* cell instance $22315 r0 *1 92.625,84.21
X$22315 2226 VIA_via2_5
* cell instance $22316 r0 *1 89.585,84.77
X$22316 2226 VIA_via1_4
* cell instance $22317 r0 *1 89.585,84.63
X$22317 2226 VIA_via2_5
* cell instance $22318 r0 *1 90.725,84.77
X$22318 2226 VIA_via1_4
* cell instance $22319 r0 *1 90.725,84.63
X$22319 2226 VIA_via2_5
* cell instance $22320 r0 *1 91.295,84.77
X$22320 2226 VIA_via1_4
* cell instance $22321 r0 *1 91.295,84.63
X$22321 2226 VIA_via2_5
* cell instance $22322 r0 *1 89.585,85.75
X$22322 2226 VIA_via1_4
* cell instance $22323 r0 *1 92.625,81.97
X$22323 2226 VIA_via1_4
* cell instance $22324 r0 *1 91.865,84.21
X$22324 2227 VIA_via1_7
* cell instance $22325 r0 *1 91.865,84.21
X$22325 2227 VIA_via2_5
* cell instance $22326 r0 *1 91.295,84.21
X$22326 2227 VIA_via2_5
* cell instance $22327 r0 *1 91.295,83.23
X$22327 2227 VIA_via1_4
* cell instance $22328 r0 *1 88.065,84.63
X$22328 2228 VIA_via1_7
* cell instance $22329 r0 *1 88.065,84.63
X$22329 2228 VIA_via2_5
* cell instance $22330 r0 *1 87.305,84.63
X$22330 2228 VIA_via1_4
* cell instance $22331 r0 *1 87.305,84.63
X$22331 2228 VIA_via2_5
* cell instance $22332 r0 *1 21.945,84.21
X$22332 2229 VIA_via1_7
* cell instance $22333 r0 *1 21.945,84.21
X$22333 2229 VIA_via2_5
* cell instance $22334 r0 *1 19.475,84.21
X$22334 2229 VIA_via2_5
* cell instance $22335 r0 *1 19.475,83.23
X$22335 2229 VIA_via1_4
* cell instance $22336 r0 *1 80.275,83.79
X$22336 2230 VIA_via1_7
* cell instance $22337 r0 *1 80.275,83.79
X$22337 2230 VIA_via2_5
* cell instance $22338 r0 *1 78.755,83.79
X$22338 2230 VIA_via2_5
* cell instance $22339 r0 *1 78.755,84.77
X$22339 2230 VIA_via1_4
* cell instance $22340 r0 *1 23.465,84.21
X$22340 2231 VIA_via1_7
* cell instance $22341 r0 *1 23.465,83.23
X$22341 2231 VIA_via1_4
* cell instance $22342 r0 *1 80.845,91.21
X$22342 2232 VIA_via1_7
* cell instance $22343 r0 *1 80.845,89.81
X$22343 2232 VIA_via2_5
* cell instance $22344 r0 *1 74.575,89.39
X$22344 2232 VIA_via2_5
* cell instance $22345 r0 *1 74.005,89.81
X$22345 2232 VIA_via2_5
* cell instance $22346 r0 *1 74.385,86.45
X$22346 2232 VIA_via2_5
* cell instance $22347 r0 *1 74.575,89.81
X$22347 2232 VIA_via2_5
* cell instance $22348 r0 *1 76.095,86.45
X$22348 2232 VIA_via2_5
* cell instance $22349 r0 *1 74.575,84.49
X$22349 2232 VIA_via2_5
* cell instance $22350 r0 *1 75.905,84.49
X$22350 2232 VIA_via2_5
* cell instance $22351 r0 *1 84.835,88.41
X$22351 2232 VIA_via2_5
* cell instance $22352 r0 *1 80.845,88.41
X$22352 2232 VIA_via2_5
* cell instance $22353 r0 *1 66.215,89.39
X$22353 2232 VIA_via2_5
* cell instance $22354 r0 *1 87.875,88.55
X$22354 2232 VIA_via2_5
* cell instance $22355 r0 *1 87.735,88.55
X$22355 2232 VIA_via3_2
* cell instance $22356 r0 *1 76.095,86.03
X$22356 2232 VIA_via1_4
* cell instance $22357 r0 *1 74.385,87.57
X$22357 2232 VIA_via1_4
* cell instance $22358 r0 *1 74.005,90.37
X$22358 2232 VIA_via1_4
* cell instance $22359 r0 *1 74.575,83.23
X$22359 2232 VIA_via1_4
* cell instance $22360 r0 *1 84.835,88.69
X$22360 2232 VIA_via1_4
* cell instance $22361 r0 *1 86.925,90.37
X$22361 2232 VIA_via1_4
* cell instance $22362 r0 *1 86.925,90.37
X$22362 2232 VIA_via2_5
* cell instance $22363 r0 *1 66.215,88.83
X$22363 2232 VIA_via1_4
* cell instance $22364 r0 *1 65.835,86.03
X$22364 2232 VIA_via1_4
* cell instance $22365 r0 *1 87.115,84.91
X$22365 2232 VIA_via1_4
* cell instance $22366 r0 *1 65.455,93.17
X$22366 2232 VIA_via1_4
* cell instance $22367 r0 *1 87.735,90.37
X$22367 2232 VIA_via3_2
* cell instance $22368 r0 *1 35.245,83.79
X$22368 2233 VIA_via1_7
* cell instance $22369 r0 *1 35.245,83.79
X$22369 2233 VIA_via2_5
* cell instance $22370 r0 *1 33.725,83.79
X$22370 2233 VIA_via2_5
* cell instance $22371 r0 *1 33.725,84.77
X$22371 2233 VIA_via1_4
* cell instance $22372 r0 *1 38.665,84.21
X$22372 2234 VIA_via1_7
* cell instance $22373 r0 *1 38.665,84.21
X$22373 2234 VIA_via2_5
* cell instance $22374 r0 *1 36.955,84.21
X$22374 2234 VIA_via2_5
* cell instance $22375 r0 *1 36.955,83.23
X$22375 2234 VIA_via1_4
* cell instance $22376 r0 *1 42.275,84.21
X$22376 2235 VIA_via1_7
* cell instance $22377 r0 *1 42.275,84.21
X$22377 2235 VIA_via2_5
* cell instance $22378 r0 *1 41.705,84.21
X$22378 2235 VIA_via2_5
* cell instance $22379 r0 *1 41.705,83.23
X$22379 2235 VIA_via1_4
* cell instance $22380 r0 *1 64.315,95.41
X$22380 2236 VIA_via1_7
* cell instance $22381 r0 *1 63.555,84.49
X$22381 2236 VIA_via2_5
* cell instance $22382 r0 *1 66.025,84.49
X$22382 2236 VIA_via2_5
* cell instance $22383 r0 *1 63.555,86.03
X$22383 2236 VIA_via2_5
* cell instance $22384 r0 *1 63.935,88.27
X$22384 2236 VIA_via2_5
* cell instance $22385 r0 *1 61.465,86.03
X$22385 2236 VIA_via2_5
* cell instance $22386 r0 *1 63.555,88.27
X$22386 2236 VIA_via2_5
* cell instance $22387 r0 *1 66.025,84.77
X$22387 2236 VIA_via1_4
* cell instance $22388 r0 *1 61.465,84.77
X$22388 2236 VIA_via1_4
* cell instance $22389 r0 *1 62.415,86.03
X$22389 2236 VIA_via1_4
* cell instance $22390 r0 *1 62.415,86.03
X$22390 2236 VIA_via2_5
* cell instance $22391 r0 *1 64.695,87.57
X$22391 2236 VIA_via1_4
* cell instance $22392 r0 *1 63.555,91.63
X$22392 2236 VIA_via1_4
* cell instance $22393 r0 *1 62.225,84.21
X$22393 2237 VIA_via1_7
* cell instance $22394 r0 *1 62.225,83.23
X$22394 2237 VIA_via1_4
* cell instance $22395 r0 *1 51.965,84.35
X$22395 2238 VIA_via2_5
* cell instance $22396 r0 *1 54.435,86.03
X$22396 2238 VIA_via1_4
* cell instance $22397 r0 *1 51.965,83.23
X$22397 2238 VIA_via1_4
* cell instance $22398 r0 *1 54.435,84.35
X$22398 2238 VIA_via1_4
* cell instance $22399 r0 *1 54.435,84.35
X$22399 2238 VIA_via2_5
* cell instance $22400 r0 *1 22.325,87.01
X$22400 2239 VIA_via1_7
* cell instance $22401 r0 *1 22.135,86.03
X$22401 2239 VIA_via1_4
* cell instance $22402 r0 *1 29.83,85.96
X$22402 2240 VIA_via1_7
* cell instance $22403 r0 *1 30.115,86.87
X$22403 2240 VIA_via2_5
* cell instance $22404 r0 *1 30.685,86.87
X$22404 2240 VIA_via2_5
* cell instance $22405 r0 *1 30.495,88.83
X$22405 2240 VIA_via1_4
* cell instance $22406 r0 *1 31.065,87.15
X$22406 2240 VIA_via1_4
* cell instance $22407 r0 *1 47.785,87.57
X$22407 2241 VIA_via2_5
* cell instance $22408 r0 *1 47.405,85.05
X$22408 2241 VIA_via1_4
* cell instance $22409 r0 *1 47.785,84.77
X$22409 2241 VIA_via1_4
* cell instance $22410 r0 *1 48.355,87.57
X$22410 2241 VIA_via1_4
* cell instance $22411 r0 *1 48.355,87.57
X$22411 2241 VIA_via2_5
* cell instance $22412 r0 *1 53.485,84.77
X$22412 2242 VIA_via2_5
* cell instance $22413 r0 *1 53.865,86.03
X$22413 2242 VIA_via1_4
* cell instance $22414 r0 *1 50.255,84.77
X$22414 2242 VIA_via1_4
* cell instance $22415 r0 *1 50.255,84.77
X$22415 2242 VIA_via2_5
* cell instance $22416 r0 *1 53.485,85.75
X$22416 2242 VIA_via1_4
* cell instance $22417 r0 *1 54.815,85.61
X$22417 2243 VIA_via1_7
* cell instance $22418 r0 *1 55.195,84.77
X$22418 2243 VIA_via1_4
* cell instance $22419 r0 *1 56.145,88.41
X$22419 2244 VIA_via1_7
* cell instance $22420 r0 *1 56.145,86.03
X$22420 2244 VIA_via1_4
* cell instance $22421 r0 *1 57.665,85.61
X$22421 2245 VIA_via1_7
* cell instance $22422 r0 *1 56.905,84.77
X$22422 2245 VIA_via1_4
* cell instance $22423 r0 *1 65.645,88.41
X$22423 2246 VIA_via1_7
* cell instance $22424 r0 *1 65.645,88.41
X$22424 2246 VIA_via2_5
* cell instance $22425 r0 *1 65.645,89.25
X$22425 2246 VIA_via1_4
* cell instance $22426 r0 *1 67.355,88.41
X$22426 2246 VIA_via2_5
* cell instance $22427 r0 *1 59.565,90.37
X$22427 2246 VIA_via2_5
* cell instance $22428 r0 *1 64.125,90.37
X$22428 2246 VIA_via2_5
* cell instance $22429 r0 *1 61.465,90.37
X$22429 2246 VIA_via2_5
* cell instance $22430 r0 *1 65.645,90.37
X$22430 2246 VIA_via2_5
* cell instance $22431 r0 *1 70.395,88.41
X$22431 2246 VIA_via2_5
* cell instance $22432 r0 *1 67.355,87.57
X$22432 2246 VIA_via1_4
* cell instance $22433 r0 *1 70.395,88.83
X$22433 2246 VIA_via1_4
* cell instance $22434 r0 *1 59.375,86.03
X$22434 2246 VIA_via1_4
* cell instance $22435 r0 *1 66.025,90.37
X$22435 2246 VIA_via1_4
* cell instance $22436 r0 *1 66.025,90.37
X$22436 2246 VIA_via2_5
* cell instance $22437 r0 *1 66.215,91.63
X$22437 2246 VIA_via1_4
* cell instance $22438 r0 *1 62.795,90.37
X$22438 2246 VIA_via1_4
* cell instance $22439 r0 *1 62.795,90.37
X$22439 2246 VIA_via2_5
* cell instance $22440 r0 *1 64.125,91.63
X$22440 2246 VIA_via1_4
* cell instance $22441 r0 *1 61.465,95.97
X$22441 2246 VIA_via1_4
* cell instance $22442 r0 *1 66.975,85.19
X$22442 2247 VIA_via1_7
* cell instance $22443 r0 *1 66.785,86.03
X$22443 2247 VIA_via1_4
* cell instance $22444 r0 *1 74.575,87.29
X$22444 2248 VIA_via2_5
* cell instance $22445 r0 *1 74.955,87.29
X$22445 2248 VIA_via2_5
* cell instance $22446 r0 *1 74.195,86.03
X$22446 2248 VIA_via1_4
* cell instance $22447 r0 *1 74.955,88.83
X$22447 2248 VIA_via1_4
* cell instance $22448 r0 *1 77.235,87.01
X$22448 2249 VIA_via1_7
* cell instance $22449 r0 *1 77.045,86.03
X$22449 2249 VIA_via1_7
* cell instance $22450 r0 *1 77.235,86.17
X$22450 2249 VIA_via2_5
* cell instance $22451 r0 *1 78.185,86.03
X$22451 2249 VIA_via1_4
* cell instance $22452 r0 *1 78.185,86.17
X$22452 2249 VIA_via2_5
* cell instance $22453 r0 *1 82.555,85.75
X$22453 2250 VIA_via1_7
* cell instance $22454 r0 *1 82.175,84.77
X$22454 2250 VIA_via1_4
* cell instance $22455 r0 *1 94.905,87.15
X$22455 2251 VIA_via2_5
* cell instance $22456 r0 *1 88.825,87.15
X$22456 2251 VIA_via2_5
* cell instance $22457 r0 *1 88.445,86.03
X$22457 2251 VIA_via1_4
* cell instance $22458 r0 *1 88.445,86.17
X$22458 2251 VIA_via2_5
* cell instance $22459 r0 *1 94.905,86.03
X$22459 2251 VIA_via1_4
* cell instance $22460 r0 *1 91.485,87.15
X$22460 2251 VIA_via1_4
* cell instance $22461 r0 *1 91.485,87.15
X$22461 2251 VIA_via2_5
* cell instance $22462 r0 *1 88.825,86.17
X$22462 2251 VIA_via1_4
* cell instance $22463 r0 *1 88.825,86.17
X$22463 2251 VIA_via2_5
* cell instance $22464 r0 *1 88.445,83.23
X$22464 2251 VIA_via1_4
* cell instance $22465 r0 *1 92.435,85.75
X$22465 2252 VIA_via2_5
* cell instance $22466 r0 *1 90.345,85.75
X$22466 2252 VIA_via2_5
* cell instance $22467 r0 *1 89.015,85.75
X$22467 2252 VIA_via2_5
* cell instance $22468 r0 *1 89.775,85.75
X$22468 2252 VIA_via2_5
* cell instance $22469 r0 *1 95.855,84.77
X$22469 2252 VIA_via2_5
* cell instance $22470 r0 *1 96.045,86.03
X$22470 2252 VIA_via1_4
* cell instance $22471 r0 *1 89.015,86.03
X$22471 2252 VIA_via1_4
* cell instance $22472 r0 *1 90.345,86.03
X$22472 2252 VIA_via1_4
* cell instance $22473 r0 *1 89.775,84.77
X$22473 2252 VIA_via1_4
* cell instance $22474 r0 *1 92.435,84.77
X$22474 2252 VIA_via1_4
* cell instance $22475 r0 *1 92.435,84.77
X$22475 2252 VIA_via2_5
* cell instance $22476 r0 *1 95.855,85.05
X$22476 2252 VIA_via1_4
* cell instance $22477 r0 *1 91.865,86.03
X$22477 2253 VIA_via1_4
* cell instance $22478 r0 *1 91.675,85.75
X$22478 2253 VIA_via1_4
* cell instance $22479 r0 *1 92.245,85.19
X$22479 2254 VIA_via1_7
* cell instance $22480 r0 *1 92.625,86.03
X$22480 2254 VIA_via1_4
* cell instance $22481 r0 *1 93.005,85.61
X$22481 2255 VIA_via1_7
* cell instance $22482 r0 *1 93.575,84.77
X$22482 2255 VIA_via1_4
* cell instance $22483 r0 *1 96.995,86.17
X$22483 2256 VIA_via1_4
* cell instance $22484 r0 *1 96.995,86.17
X$22484 2256 VIA_via2_5
* cell instance $22485 r0 *1 97.535,85.75
X$22485 2256 VIA_via4_0
* cell instance $22486 r0 *1 97.535,86.17
X$22486 2256 VIA_via3_2
* cell instance $22487 r0 *1 90.155,84.77
X$22487 2257 VIA_via1_4
* cell instance $22488 r0 *1 90.155,84.77
X$22488 2257 VIA_via2_5
* cell instance $22489 r0 *1 86.925,84.77
X$22489 2257 VIA_via1_4
* cell instance $22490 r0 *1 86.925,84.77
X$22490 2257 VIA_via2_5
* cell instance $22491 r0 *1 88.255,85.61
X$22491 2258 VIA_via1_7
* cell instance $22492 r0 *1 88.255,84.77
X$22492 2258 VIA_via1_4
* cell instance $22493 r0 *1 82.365,84.77
X$22493 2259 VIA_via1_4
* cell instance $22494 r0 *1 82.365,84.91
X$22494 2259 VIA_via2_5
* cell instance $22495 r0 *1 84.645,84.91
X$22495 2259 VIA_via1_4
* cell instance $22496 r0 *1 84.645,84.91
X$22496 2259 VIA_via2_5
* cell instance $22497 r0 *1 84.075,84.77
X$22497 2260 VIA_via1_4
* cell instance $22498 r0 *1 84.075,84.77
X$22498 2260 VIA_via2_5
* cell instance $22499 r0 *1 82.935,84.77
X$22499 2260 VIA_via1_4
* cell instance $22500 r0 *1 82.935,84.77
X$22500 2260 VIA_via2_5
* cell instance $22501 r0 *1 79.705,84.77
X$22501 2261 VIA_via1_4
* cell instance $22502 r0 *1 79.705,84.77
X$22502 2261 VIA_via2_5
* cell instance $22503 r0 *1 76.095,84.77
X$22503 2261 VIA_via1_4
* cell instance $22504 r0 *1 76.095,84.77
X$22504 2261 VIA_via2_5
* cell instance $22505 r0 *1 79.325,84.77
X$22505 2262 VIA_via1_4
* cell instance $22506 r0 *1 79.325,83.51
X$22506 2262 VIA_via1_4
* cell instance $22507 r0 *1 45.125,84.77
X$22507 2263 VIA_via1_4
* cell instance $22508 r0 *1 45.125,84.91
X$22508 2263 VIA_via2_5
* cell instance $22509 r0 *1 48.735,84.91
X$22509 2263 VIA_via1_4
* cell instance $22510 r0 *1 48.735,84.91
X$22510 2263 VIA_via2_5
* cell instance $22511 r0 *1 76.095,85.61
X$22511 2264 VIA_via1_7
* cell instance $22512 r0 *1 76.095,85.61
X$22512 2264 VIA_via2_5
* cell instance $22513 r0 *1 78.565,85.61
X$22513 2264 VIA_via2_5
* cell instance $22514 r0 *1 78.565,84.77
X$22514 2264 VIA_via1_4
* cell instance $22515 r0 *1 72.865,84.77
X$22515 2265 VIA_via1_4
* cell instance $22516 r0 *1 72.865,84.91
X$22516 2265 VIA_via2_5
* cell instance $22517 r0 *1 75.145,84.91
X$22517 2265 VIA_via1_4
* cell instance $22518 r0 *1 75.145,84.91
X$22518 2265 VIA_via2_5
* cell instance $22519 r0 *1 73.435,84.77
X$22519 2266 VIA_via1_4
* cell instance $22520 r0 *1 73.435,84.77
X$22520 2266 VIA_via2_5
* cell instance $22521 r0 *1 74.195,84.77
X$22521 2266 VIA_via1_4
* cell instance $22522 r0 *1 74.195,84.77
X$22522 2266 VIA_via2_5
* cell instance $22523 r0 *1 66.595,85.75
X$22523 2267 VIA_via2_5
* cell instance $22524 r0 *1 65.835,85.75
X$22524 2267 VIA_via1_4
* cell instance $22525 r0 *1 65.835,85.75
X$22525 2267 VIA_via2_5
* cell instance $22526 r0 *1 66.595,86.03
X$22526 2267 VIA_via1_4
* cell instance $22527 r0 *1 65.075,85.19
X$22527 2268 VIA_via1_7
* cell instance $22528 r0 *1 65.075,85.19
X$22528 2268 VIA_via2_5
* cell instance $22529 r0 *1 64.695,85.19
X$22529 2268 VIA_via2_5
* cell instance $22530 r0 *1 64.695,86.03
X$22530 2268 VIA_via1_4
* cell instance $22531 r0 *1 57.095,85.19
X$22531 2269 VIA_via1_7
* cell instance $22532 r0 *1 57.095,85.19
X$22532 2269 VIA_via2_5
* cell instance $22533 r0 *1 55.955,85.19
X$22533 2269 VIA_via2_5
* cell instance $22534 r0 *1 55.955,86.03
X$22534 2269 VIA_via1_4
* cell instance $22535 r0 *1 60.895,84.77
X$22535 2270 VIA_via2_5
* cell instance $22536 r0 *1 58.235,86.03
X$22536 2270 VIA_via2_5
* cell instance $22537 r0 *1 60.895,85.75
X$22537 2270 VIA_via1_4
* cell instance $22538 r0 *1 58.235,84.77
X$22538 2270 VIA_via1_4
* cell instance $22539 r0 *1 58.235,84.77
X$22539 2270 VIA_via2_5
* cell instance $22540 r0 *1 57.285,86.03
X$22540 2270 VIA_via1_4
* cell instance $22541 r0 *1 57.285,86.03
X$22541 2270 VIA_via2_5
* cell instance $22542 r0 *1 6.935,88.41
X$22542 2271 VIA_via1_7
* cell instance $22543 r0 *1 6.935,88.41
X$22543 2271 VIA_via2_5
* cell instance $22544 r0 *1 3.515,88.41
X$22544 2271 VIA_via2_5
* cell instance $22545 r0 *1 3.135,87.57
X$22545 2271 VIA_via1_4
* cell instance $22546 r0 *1 4.655,88.83
X$22546 2272 VIA_via1_4
* cell instance $22547 r0 *1 5.415,87.85
X$22547 2272 VIA_via1_4
* cell instance $22548 r0 *1 5.985,88.83
X$22548 2272 VIA_via1_4
* cell instance $22549 r0 *1 6.175,86.59
X$22549 2273 VIA_via1_7
* cell instance $22550 r0 *1 6.365,87.57
X$22550 2273 VIA_via1_4
* cell instance $22551 r0 *1 18.905,86.45
X$22551 2274 VIA_via2_5
* cell instance $22552 r0 *1 16.245,86.45
X$22552 2274 VIA_via2_5
* cell instance $22553 r0 *1 16.245,87.57
X$22553 2274 VIA_via1_4
* cell instance $22554 r0 *1 16.245,88.83
X$22554 2274 VIA_via1_4
* cell instance $22555 r0 *1 18.905,86.03
X$22555 2274 VIA_via1_4
* cell instance $22556 r0 *1 21.375,86.45
X$22556 2275 VIA_via2_5
* cell instance $22557 r0 *1 21.565,88.83
X$22557 2275 VIA_via1_4
* cell instance $22558 r0 *1 21.375,87.57
X$22558 2275 VIA_via1_4
* cell instance $22559 r0 *1 24.415,86.45
X$22559 2275 VIA_via1_4
* cell instance $22560 r0 *1 24.415,86.45
X$22560 2275 VIA_via2_5
* cell instance $22561 r0 *1 26.505,87.15
X$22561 2276 VIA_via1_4
* cell instance $22562 r0 *1 26.315,86.03
X$22562 2276 VIA_via1_4
* cell instance $22563 r0 *1 26.885,87.57
X$22563 2276 VIA_via1_4
* cell instance $22564 r0 *1 27.075,88.83
X$22564 2277 VIA_via1_4
* cell instance $22565 r0 *1 27.455,87.57
X$22565 2277 VIA_via1_4
* cell instance $22566 r0 *1 26.695,88.55
X$22566 2277 VIA_via1_4
* cell instance $22567 r0 *1 32.775,88.83
X$22567 2278 VIA_via1_4
* cell instance $22568 r0 *1 32.205,87.15
X$22568 2278 VIA_via1_4
* cell instance $22569 r0 *1 48.925,87.57
X$22569 2279 VIA_via1_4
* cell instance $22570 r0 *1 48.925,86.03
X$22570 2279 VIA_via1_4
* cell instance $22571 r0 *1 48.545,86.45
X$22571 2279 VIA_via1_4
* cell instance $22572 r0 *1 56.715,86.03
X$22572 2280 VIA_via1_4
* cell instance $22573 r0 *1 56.715,87.57
X$22573 2280 VIA_via1_4
* cell instance $22574 r0 *1 56.715,87.43
X$22574 2280 VIA_via2_5
* cell instance $22575 r0 *1 60.325,87.43
X$22575 2280 VIA_via1_4
* cell instance $22576 r0 *1 60.325,87.43
X$22576 2280 VIA_via2_5
* cell instance $22577 r0 *1 65.455,88.83
X$22577 2281 VIA_via2_5
* cell instance $22578 r0 *1 65.265,87.15
X$22578 2281 VIA_via1_4
* cell instance $22579 r0 *1 64.315,88.83
X$22579 2281 VIA_via1_4
* cell instance $22580 r0 *1 64.315,88.83
X$22580 2281 VIA_via2_5
* cell instance $22581 r0 *1 70.205,87.01
X$22581 2282 VIA_via1_7
* cell instance $22582 r0 *1 70.395,86.03
X$22582 2282 VIA_via1_4
* cell instance $22583 r0 *1 71.725,87.29
X$22583 2283 VIA_via1_7
* cell instance $22584 r0 *1 71.725,87.29
X$22584 2283 VIA_via2_5
* cell instance $22585 r0 *1 73.055,87.29
X$22585 2283 VIA_via2_5
* cell instance $22586 r0 *1 70.395,87.29
X$22586 2283 VIA_via2_5
* cell instance $22587 r0 *1 71.915,88.55
X$22587 2283 VIA_via1_4
* cell instance $22588 r0 *1 73.055,87.57
X$22588 2283 VIA_via1_4
* cell instance $22589 r0 *1 70.395,87.57
X$22589 2283 VIA_via1_4
* cell instance $22590 r0 *1 73.815,87.29
X$22590 2284 VIA_via2_5
* cell instance $22591 r0 *1 73.815,86.87
X$22591 2284 VIA_via2_5
* cell instance $22592 r0 *1 74.955,86.87
X$22592 2284 VIA_via2_5
* cell instance $22593 r0 *1 70.775,87.43
X$22593 2284 VIA_via2_5
* cell instance $22594 r0 *1 74.955,86.03
X$22594 2284 VIA_via1_4
* cell instance $22595 r0 *1 70.585,90.37
X$22595 2284 VIA_via1_4
* cell instance $22596 r0 *1 70.585,90.51
X$22596 2284 VIA_via2_5
* cell instance $22597 r0 *1 67.735,91.35
X$22597 2284 VIA_via1_4
* cell instance $22598 r0 *1 73.245,87.57
X$22598 2284 VIA_via1_4
* cell instance $22599 r0 *1 73.245,87.57
X$22599 2284 VIA_via2_5
* cell instance $22600 r0 *1 68.115,90.37
X$22600 2284 VIA_via1_4
* cell instance $22601 r0 *1 68.115,90.51
X$22601 2284 VIA_via2_5
* cell instance $22602 r0 *1 72.865,87.01
X$22602 2285 VIA_via1_7
* cell instance $22603 r0 *1 72.865,87.01
X$22603 2285 VIA_via2_5
* cell instance $22604 r0 *1 75.145,87.01
X$22604 2285 VIA_via2_5
* cell instance $22605 r0 *1 73.625,87.01
X$22605 2285 VIA_via2_5
* cell instance $22606 r0 *1 75.145,86.03
X$22606 2285 VIA_via1_4
* cell instance $22607 r0 *1 73.435,88.83
X$22607 2285 VIA_via1_4
* cell instance $22608 r0 *1 74.195,87.71
X$22608 2286 VIA_via2_5
* cell instance $22609 r0 *1 74.575,87.57
X$22609 2286 VIA_via1_4
* cell instance $22610 r0 *1 74.575,87.71
X$22610 2286 VIA_via2_5
* cell instance $22611 r0 *1 73.815,87.85
X$22611 2286 VIA_via1_4
* cell instance $22612 r0 *1 77.805,87.57
X$22612 2287 VIA_via2_5
* cell instance $22613 r0 *1 77.805,93.17
X$22613 2287 VIA_via1_4
* cell instance $22614 r0 *1 77.425,87.57
X$22614 2287 VIA_via1_4
* cell instance $22615 r0 *1 77.425,86.31
X$22615 2287 VIA_via1_4
* cell instance $22616 r0 *1 79.895,86.17
X$22616 2287 VIA_via1_4
* cell instance $22617 r0 *1 79.895,87.57
X$22617 2287 VIA_via1_4
* cell instance $22618 r0 *1 79.895,87.57
X$22618 2287 VIA_via2_5
* cell instance $22619 r0 *1 86.925,86.59
X$22619 2288 VIA_via1_7
* cell instance $22620 r0 *1 82.365,87.57
X$22620 2288 VIA_via2_5
* cell instance $22621 r0 *1 86.735,87.57
X$22621 2288 VIA_via2_5
* cell instance $22622 r0 *1 82.365,86.03
X$22622 2288 VIA_via1_4
* cell instance $22623 r0 *1 84.455,87.57
X$22623 2288 VIA_via1_4
* cell instance $22624 r0 *1 84.455,87.57
X$22624 2288 VIA_via2_5
* cell instance $22625 r0 *1 86.925,87.57
X$22625 2288 VIA_via1_4
* cell instance $22626 r0 *1 86.925,87.57
X$22626 2288 VIA_via2_5
* cell instance $22627 r0 *1 89.585,86.59
X$22627 2289 VIA_via1_7
* cell instance $22628 r0 *1 82.555,87.43
X$22628 2289 VIA_via2_5
* cell instance $22629 r0 *1 89.585,87.29
X$22629 2289 VIA_via2_5
* cell instance $22630 r0 *1 82.555,86.03
X$22630 2289 VIA_via1_4
* cell instance $22631 r0 *1 85.785,87.57
X$22631 2289 VIA_via1_4
* cell instance $22632 r0 *1 85.785,87.43
X$22632 2289 VIA_via2_5
* cell instance $22633 r0 *1 86.925,91.63
X$22633 2289 VIA_via1_4
* cell instance $22634 r0 *1 86.925,91.63
X$22634 2289 VIA_via2_5
* cell instance $22635 r0 *1 86.335,87.29
X$22635 2289 VIA_via3_2
* cell instance $22636 r0 *1 86.335,91.63
X$22636 2289 VIA_via3_2
* cell instance $22637 r0 *1 85.785,86.59
X$22637 2290 VIA_via1_7
* cell instance $22638 r0 *1 85.785,86.59
X$22638 2290 VIA_via2_5
* cell instance $22639 r0 *1 84.835,86.59
X$22639 2290 VIA_via2_5
* cell instance $22640 r0 *1 84.835,84.77
X$22640 2290 VIA_via1_4
* cell instance $22641 r0 *1 86.165,87.57
X$22641 2290 VIA_via1_4
* cell instance $22642 r0 *1 92.245,87.71
X$22642 2291 VIA_via1_4
* cell instance $22643 r0 *1 92.625,87.57
X$22643 2291 VIA_via1_4
* cell instance $22644 r0 *1 93.385,86.31
X$22644 2292 VIA_via1_4
* cell instance $22645 r0 *1 93.195,87.57
X$22645 2292 VIA_via1_4
* cell instance $22646 r0 *1 95.285,87.57
X$22646 2293 VIA_via1_4
* cell instance $22647 r0 *1 95.475,89.25
X$22647 2293 VIA_via1_4
* cell instance $22648 r0 *1 95.475,90.37
X$22648 2293 VIA_via1_4
* cell instance $22649 r0 *1 95.285,86.59
X$22649 2294 VIA_via1_7
* cell instance $22650 r0 *1 95.285,86.59
X$22650 2294 VIA_via2_5
* cell instance $22651 r0 *1 95.295,86.59
X$22651 2294 VIA_via3_2
* cell instance $22652 r0 *1 95.295,86.87
X$22652 2294 VIA_via4_0
* cell instance $22653 r0 *1 96.425,86.31
X$22653 2295 VIA_via1_4
* cell instance $22654 r0 *1 96.425,86.31
X$22654 2295 VIA_via2_5
* cell instance $22655 r0 *1 97.255,86.31
X$22655 2295 VIA_via4_0
* cell instance $22656 r0 *1 97.255,86.31
X$22656 2295 VIA_via3_2
* cell instance $22657 r0 *1 10.545,87.01
X$22657 2296 VIA_via1_7
* cell instance $22658 r0 *1 10.545,87.01
X$22658 2296 VIA_via2_5
* cell instance $22659 r0 *1 9.785,87.01
X$22659 2296 VIA_via2_5
* cell instance $22660 r0 *1 9.785,86.03
X$22660 2296 VIA_via1_4
* cell instance $22661 r0 *1 11.495,86.45
X$22661 2297 VIA_via2_5
* cell instance $22662 r0 *1 11.495,87.57
X$22662 2297 VIA_via1_4
* cell instance $22663 r0 *1 11.495,87.57
X$22663 2297 VIA_via2_5
* cell instance $22664 r0 *1 12.065,86.45
X$22664 2297 VIA_via1_4
* cell instance $22665 r0 *1 12.065,86.45
X$22665 2297 VIA_via2_5
* cell instance $22666 r0 *1 9.595,87.57
X$22666 2297 VIA_via1_4
* cell instance $22667 r0 *1 9.595,87.57
X$22667 2297 VIA_via2_5
* cell instance $22668 r0 *1 92.055,86.03
X$22668 2298 VIA_via1_4
* cell instance $22669 r0 *1 92.055,86.17
X$22669 2298 VIA_via2_5
* cell instance $22670 r0 *1 90.915,86.17
X$22670 2298 VIA_via1_4
* cell instance $22671 r0 *1 90.915,86.17
X$22671 2298 VIA_via2_5
* cell instance $22672 r0 *1 17.195,87.01
X$22672 2299 VIA_via1_7
* cell instance $22673 r0 *1 17.195,87.01
X$22673 2299 VIA_via2_5
* cell instance $22674 r0 *1 16.625,87.01
X$22674 2299 VIA_via2_5
* cell instance $22675 r0 *1 16.625,86.03
X$22675 2299 VIA_via1_4
* cell instance $22676 r0 *1 92.435,87.43
X$22676 2300 VIA_via1_7
* cell instance $22677 r0 *1 92.435,87.43
X$22677 2300 VIA_via2_5
* cell instance $22678 r0 *1 87.495,87.43
X$22678 2300 VIA_via1_4
* cell instance $22679 r0 *1 87.495,87.43
X$22679 2300 VIA_via2_5
* cell instance $22680 r0 *1 91.105,85.19
X$22680 2301 VIA_via1_7
* cell instance $22681 r0 *1 91.105,86.03
X$22681 2301 VIA_via1_4
* cell instance $22682 r0 *1 27.265,86.59
X$22682 2302 VIA_via1_7
* cell instance $22683 r0 *1 27.265,86.59
X$22683 2302 VIA_via2_5
* cell instance $22684 r0 *1 24.225,86.59
X$22684 2302 VIA_via2_5
* cell instance $22685 r0 *1 24.225,87.57
X$22685 2302 VIA_via1_4
* cell instance $22686 r0 *1 30.685,86.59
X$22686 2303 VIA_via1_7
* cell instance $22687 r0 *1 30.685,86.59
X$22687 2303 VIA_via2_5
* cell instance $22688 r0 *1 28.785,86.59
X$22688 2303 VIA_via2_5
* cell instance $22689 r0 *1 28.785,87.57
X$22689 2303 VIA_via1_4
* cell instance $22690 r0 *1 32.015,78.89
X$22690 2304 VIA_via1_7
* cell instance $22691 r0 *1 30.685,87.29
X$22691 2304 VIA_via2_5
* cell instance $22692 r0 *1 32.015,87.29
X$22692 2304 VIA_via2_5
* cell instance $22693 r0 *1 30.875,95.97
X$22693 2304 VIA_via1_4
* cell instance $22694 r0 *1 27.835,87.57
X$22694 2305 VIA_via1_4
* cell instance $22695 r0 *1 27.835,87.57
X$22695 2305 VIA_via2_5
* cell instance $22696 r0 *1 31.825,87.57
X$22696 2305 VIA_via1_4
* cell instance $22697 r0 *1 31.825,87.57
X$22697 2305 VIA_via2_5
* cell instance $22698 r0 *1 89.205,85.19
X$22698 2306 VIA_via1_7
* cell instance $22699 r0 *1 89.205,87.57
X$22699 2306 VIA_via1_4
* cell instance $22700 r0 *1 40.945,87.01
X$22700 2307 VIA_via1_7
* cell instance $22701 r0 *1 40.945,87.01
X$22701 2307 VIA_via2_5
* cell instance $22702 r0 *1 39.805,87.01
X$22702 2307 VIA_via2_5
* cell instance $22703 r0 *1 39.805,86.03
X$22703 2307 VIA_via1_4
* cell instance $22704 r0 *1 42.085,88.83
X$22704 2308 VIA_via2_5
* cell instance $22705 r0 *1 42.085,87.57
X$22705 2308 VIA_via2_5
* cell instance $22706 r0 *1 39.995,87.57
X$22706 2308 VIA_via1_4
* cell instance $22707 r0 *1 39.995,87.57
X$22707 2308 VIA_via2_5
* cell instance $22708 r0 *1 42.655,88.83
X$22708 2308 VIA_via1_4
* cell instance $22709 r0 *1 42.655,88.83
X$22709 2308 VIA_via2_5
* cell instance $22710 r0 *1 42.085,86.03
X$22710 2308 VIA_via1_4
* cell instance $22711 r0 *1 49.875,86.17
X$22711 2309 VIA_via1_4
* cell instance $22712 r0 *1 49.875,86.17
X$22712 2309 VIA_via2_5
* cell instance $22713 r0 *1 46.265,86.03
X$22713 2309 VIA_via1_4
* cell instance $22714 r0 *1 46.265,86.17
X$22714 2309 VIA_via2_5
* cell instance $22715 r0 *1 50.255,86.03
X$22715 2310 VIA_via2_5
* cell instance $22716 r0 *1 55.195,86.03
X$22716 2310 VIA_via1_4
* cell instance $22717 r0 *1 55.195,86.03
X$22717 2310 VIA_via2_5
* cell instance $22718 r0 *1 50.255,87.29
X$22718 2310 VIA_via1_4
* cell instance $22719 r0 *1 51.205,85.19
X$22719 2311 VIA_via1_7
* cell instance $22720 r0 *1 51.205,86.03
X$22720 2311 VIA_via1_4
* cell instance $22721 r0 *1 55.385,85.19
X$22721 2312 VIA_via1_7
* cell instance $22722 r0 *1 55.385,86.03
X$22722 2312 VIA_via1_4
* cell instance $22723 r0 *1 58.615,85.19
X$22723 2313 VIA_via1_7
* cell instance $22724 r0 *1 58.615,86.03
X$22724 2313 VIA_via1_4
* cell instance $22725 r0 *1 57.095,87.57
X$22725 2314 VIA_via1_4
* cell instance $22726 r0 *1 58.045,87.57
X$22726 2314 VIA_via1_4
* cell instance $22727 r0 *1 75.335,86.17
X$22727 2315 VIA_via1_4
* cell instance $22728 r0 *1 75.335,86.17
X$22728 2315 VIA_via2_5
* cell instance $22729 r0 *1 76.285,86.03
X$22729 2315 VIA_via1_4
* cell instance $22730 r0 *1 76.285,86.17
X$22730 2315 VIA_via2_5
* cell instance $22731 r0 *1 52.345,91.63
X$22731 2316 VIA_via2_5
* cell instance $22732 r0 *1 50.065,91.63
X$22732 2316 VIA_via2_5
* cell instance $22733 r0 *1 55.575,91.63
X$22733 2316 VIA_via2_5
* cell instance $22734 r0 *1 59.755,87.57
X$22734 2316 VIA_via2_5
* cell instance $22735 r0 *1 50.065,95.97
X$22735 2316 VIA_via1_4
* cell instance $22736 r0 *1 54.435,94.43
X$22736 2316 VIA_via1_4
* cell instance $22737 r0 *1 51.965,90.37
X$22737 2316 VIA_via1_4
* cell instance $22738 r0 *1 52.345,88.83
X$22738 2316 VIA_via1_4
* cell instance $22739 r0 *1 54.815,91.63
X$22739 2316 VIA_via1_4
* cell instance $22740 r0 *1 54.815,91.63
X$22740 2316 VIA_via2_5
* cell instance $22741 r0 *1 54.435,92.05
X$22741 2316 VIA_via1_4
* cell instance $22742 r0 *1 56.525,91.63
X$22742 2316 VIA_via1_4
* cell instance $22743 r0 *1 56.525,91.63
X$22743 2316 VIA_via2_5
* cell instance $22744 r0 *1 58.805,87.57
X$22744 2316 VIA_via1_4
* cell instance $22745 r0 *1 58.805,87.57
X$22745 2316 VIA_via2_5
* cell instance $22746 r0 *1 59.755,91.63
X$22746 2316 VIA_via1_4
* cell instance $22747 r0 *1 59.755,91.63
X$22747 2316 VIA_via2_5
* cell instance $22748 r0 *1 55.575,90.37
X$22748 2316 VIA_via1_4
* cell instance $22749 r0 *1 66.025,85.19
X$22749 2317 VIA_via1_7
* cell instance $22750 r0 *1 66.025,86.03
X$22750 2317 VIA_via1_4
* cell instance $22751 r0 *1 67.355,85.19
X$22751 2318 VIA_via1_7
* cell instance $22752 r0 *1 67.355,86.03
X$22752 2318 VIA_via1_4
* cell instance $22753 r0 *1 67.735,86.59
X$22753 2319 VIA_via1_7
* cell instance $22754 r0 *1 67.735,86.59
X$22754 2319 VIA_via2_5
* cell instance $22755 r0 *1 66.595,86.59
X$22755 2319 VIA_via2_5
* cell instance $22756 r0 *1 66.595,87.57
X$22756 2319 VIA_via1_4
* cell instance $22757 r0 *1 74.765,86.17
X$22757 2320 VIA_via2_5
* cell instance $22758 r0 *1 67.925,87.15
X$22758 2320 VIA_via2_5
* cell instance $22759 r0 *1 74.765,88.97
X$22759 2320 VIA_via1_4
* cell instance $22760 r0 *1 67.925,86.03
X$22760 2320 VIA_via1_4
* cell instance $22761 r0 *1 67.925,86.17
X$22761 2320 VIA_via2_5
* cell instance $22762 r0 *1 68.875,87.15
X$22762 2320 VIA_via1_4
* cell instance $22763 r0 *1 68.875,87.15
X$22763 2320 VIA_via2_5
* cell instance $22764 r0 *1 70.965,87.01
X$22764 2321 VIA_via1_7
* cell instance $22765 r0 *1 70.965,86.03
X$22765 2321 VIA_via1_4
* cell instance $22766 r0 *1 71.155,87.57
X$22766 2322 VIA_via1_4
* cell instance $22767 r0 *1 71.155,87.57
X$22767 2322 VIA_via2_5
* cell instance $22768 r0 *1 69.635,87.57
X$22768 2322 VIA_via1_4
* cell instance $22769 r0 *1 69.635,87.57
X$22769 2322 VIA_via2_5
* cell instance $22770 r0 *1 74.195,86.31
X$22770 2323 VIA_via2_5
* cell instance $22771 r0 *1 72.675,86.31
X$22771 2323 VIA_via2_5
* cell instance $22772 r0 *1 72.675,84.77
X$22772 2323 VIA_via1_4
* cell instance $22773 r0 *1 74.195,87.29
X$22773 2323 VIA_via1_4
* cell instance $22774 r0 *1 72.485,88.41
X$22774 2324 VIA_via1_7
* cell instance $22775 r0 *1 72.485,87.57
X$22775 2324 VIA_via2_5
* cell instance $22776 r0 *1 72.105,87.57
X$22776 2324 VIA_via1_4
* cell instance $22777 r0 *1 72.105,87.57
X$22777 2324 VIA_via2_5
* cell instance $22778 r0 *1 5.225,88.13
X$22778 2325 VIA_via2_5
* cell instance $22779 r0 *1 8.645,88.13
X$22779 2325 VIA_via2_5
* cell instance $22780 r0 *1 5.225,86.03
X$22780 2325 VIA_via1_4
* cell instance $22781 r0 *1 5.225,88.83
X$22781 2325 VIA_via1_4
* cell instance $22782 r0 *1 8.645,87.85
X$22782 2325 VIA_via1_4
* cell instance $22783 r0 *1 11.685,88.83
X$22783 2326 VIA_via1_4
* cell instance $22784 r0 *1 11.685,88.83
X$22784 2326 VIA_via2_5
* cell instance $22785 r0 *1 8.075,88.83
X$22785 2326 VIA_via1_4
* cell instance $22786 r0 *1 8.075,88.69
X$22786 2326 VIA_via2_5
* cell instance $22787 r0 *1 12.065,88.69
X$22787 2327 VIA_via2_5
* cell instance $22788 r0 *1 10.355,88.69
X$22788 2327 VIA_via1_4
* cell instance $22789 r0 *1 10.355,88.69
X$22789 2327 VIA_via2_5
* cell instance $22790 r0 *1 10.735,88.83
X$22790 2327 VIA_via1_4
* cell instance $22791 r0 *1 10.735,88.69
X$22791 2327 VIA_via2_5
* cell instance $22792 r0 *1 12.065,87.57
X$22792 2327 VIA_via1_4
* cell instance $22793 r0 *1 12.445,87.99
X$22793 2328 VIA_via1_7
* cell instance $22794 r0 *1 12.635,88.83
X$22794 2328 VIA_via1_4
* cell instance $22795 r0 *1 15.675,88.83
X$22795 2329 VIA_via1_4
* cell instance $22796 r0 *1 15.675,88.83
X$22796 2329 VIA_via2_5
* cell instance $22797 r0 *1 15.865,87.85
X$22797 2329 VIA_via1_4
* cell instance $22798 r0 *1 13.965,88.83
X$22798 2329 VIA_via1_4
* cell instance $22799 r0 *1 13.965,88.83
X$22799 2329 VIA_via2_5
* cell instance $22800 r0 *1 19.095,88.83
X$22800 2330 VIA_via1_4
* cell instance $22801 r0 *1 19.095,88.69
X$22801 2330 VIA_via2_5
* cell instance $22802 r0 *1 20.995,88.83
X$22802 2330 VIA_via1_4
* cell instance $22803 r0 *1 20.995,88.69
X$22803 2330 VIA_via2_5
* cell instance $22804 r0 *1 20.995,87.85
X$22804 2330 VIA_via1_4
* cell instance $22805 r0 *1 37.715,90.37
X$22805 2331 VIA_via1_4
* cell instance $22806 r0 *1 37.715,88.83
X$22806 2331 VIA_via1_4
* cell instance $22807 r0 *1 38.095,87.85
X$22807 2331 VIA_via1_4
* cell instance $22808 r0 *1 42.275,88.13
X$22808 2332 VIA_via2_5
* cell instance $22809 r0 *1 41.705,88.13
X$22809 2332 VIA_via2_5
* cell instance $22810 r0 *1 43.225,88.13
X$22810 2332 VIA_via2_5
* cell instance $22811 r0 *1 43.225,88.83
X$22811 2332 VIA_via1_4
* cell instance $22812 r0 *1 41.705,87.57
X$22812 2332 VIA_via1_4
* cell instance $22813 r0 *1 42.275,88.55
X$22813 2332 VIA_via1_4
* cell instance $22814 r0 *1 36.575,88.83
X$22814 2333 VIA_via2_5
* cell instance $22815 r0 *1 45.505,91.63
X$22815 2333 VIA_via2_5
* cell instance $22816 r0 *1 40.185,88.83
X$22816 2333 VIA_via2_5
* cell instance $22817 r0 *1 47.025,91.63
X$22817 2333 VIA_via2_5
* cell instance $22818 r0 *1 40.185,91.63
X$22818 2333 VIA_via2_5
* cell instance $22819 r0 *1 41.325,91.63
X$22819 2333 VIA_via2_5
* cell instance $22820 r0 *1 40.755,91.63
X$22820 2333 VIA_via1_4
* cell instance $22821 r0 *1 40.755,91.63
X$22821 2333 VIA_via2_5
* cell instance $22822 r0 *1 42.845,91.63
X$22822 2333 VIA_via1_4
* cell instance $22823 r0 *1 42.845,91.63
X$22823 2333 VIA_via2_5
* cell instance $22824 r0 *1 47.215,91.63
X$22824 2333 VIA_via1_4
* cell instance $22825 r0 *1 47.215,91.63
X$22825 2333 VIA_via2_5
* cell instance $22826 r0 *1 45.695,88.83
X$22826 2333 VIA_via1_4
* cell instance $22827 r0 *1 40.755,88.83
X$22827 2333 VIA_via1_4
* cell instance $22828 r0 *1 40.755,88.83
X$22828 2333 VIA_via2_5
* cell instance $22829 r0 *1 36.575,87.57
X$22829 2333 VIA_via1_4
* cell instance $22830 r0 *1 35.815,88.83
X$22830 2333 VIA_via1_4
* cell instance $22831 r0 *1 35.815,88.83
X$22831 2333 VIA_via2_5
* cell instance $22832 r0 *1 41.515,95.97
X$22832 2333 VIA_via1_4
* cell instance $22833 r0 *1 47.025,93.17
X$22833 2333 VIA_via1_4
* cell instance $22834 r0 *1 47.215,89.11
X$22834 2334 VIA_via1_4
* cell instance $22835 r0 *1 47.785,90.37
X$22835 2334 VIA_via1_4
* cell instance $22836 r0 *1 47.595,88.83
X$22836 2334 VIA_via1_4
* cell instance $22837 r0 *1 63.935,87.99
X$22837 2335 VIA_via1_7
* cell instance $22838 r0 *1 63.745,88.83
X$22838 2335 VIA_via1_4
* cell instance $22839 r0 *1 74.195,88.55
X$22839 2336 VIA_via1_7
* cell instance $22840 r0 *1 74.385,90.37
X$22840 2336 VIA_via2_5
* cell instance $22841 r0 *1 75.905,90.37
X$22841 2336 VIA_via2_5
* cell instance $22842 r0 *1 76.855,94.01
X$22842 2336 VIA_via2_5
* cell instance $22843 r0 *1 75.145,94.01
X$22843 2336 VIA_via2_5
* cell instance $22844 r0 *1 75.905,94.01
X$22844 2336 VIA_via2_5
* cell instance $22845 r0 *1 76.855,94.29
X$22845 2336 VIA_via1_4
* cell instance $22846 r0 *1 75.335,94.43
X$22846 2336 VIA_via1_4
* cell instance $22847 r0 *1 75.905,91.63
X$22847 2336 VIA_via1_4
* cell instance $22848 r0 *1 75.145,94.43
X$22848 2336 VIA_via1_4
* cell instance $22849 r0 *1 85.975,87.99
X$22849 2337 VIA_via1_7
* cell instance $22850 r0 *1 85.975,88.55
X$22850 2337 VIA_via2_5
* cell instance $22851 r0 *1 86.925,88.69
X$22851 2337 VIA_via1_4
* cell instance $22852 r0 *1 86.925,88.55
X$22852 2337 VIA_via2_5
* cell instance $22853 r0 *1 86.735,90.37
X$22853 2337 VIA_via1_4
* cell instance $22854 r0 *1 86.735,90.23
X$22854 2337 VIA_via2_5
* cell instance $22855 r0 *1 85.785,90.37
X$22855 2337 VIA_via1_4
* cell instance $22856 r0 *1 85.785,90.23
X$22856 2337 VIA_via2_5
* cell instance $22857 r0 *1 94.715,89.81
X$22857 2338 VIA_via1_7
* cell instance $22858 r0 *1 94.715,89.81
X$22858 2338 VIA_via2_5
* cell instance $22859 r0 *1 89.205,89.81
X$22859 2338 VIA_via2_5
* cell instance $22860 r0 *1 86.545,88.97
X$22860 2338 VIA_via2_5
* cell instance $22861 r0 *1 87.305,88.83
X$22861 2338 VIA_via1_4
* cell instance $22862 r0 *1 87.305,88.83
X$22862 2338 VIA_via2_5
* cell instance $22863 r0 *1 85.975,91.49
X$22863 2338 VIA_via1_4
* cell instance $22864 r0 *1 88.635,88.83
X$22864 2338 VIA_via1_4
* cell instance $22865 r0 *1 88.635,88.83
X$22865 2338 VIA_via2_5
* cell instance $22866 r0 *1 89.205,88.83
X$22866 2338 VIA_via1_4
* cell instance $22867 r0 *1 89.205,88.83
X$22867 2338 VIA_via2_5
* cell instance $22868 r0 *1 86.355,90.37
X$22868 2338 VIA_via1_4
* cell instance $22869 r0 *1 87.495,88.83
X$22869 2339 VIA_via1_4
* cell instance $22870 r0 *1 87.305,88.55
X$22870 2339 VIA_via1_4
* cell instance $22871 r0 *1 93.575,87.99
X$22871 2340 VIA_via1_7
* cell instance $22872 r0 *1 93.195,88.83
X$22872 2340 VIA_via1_4
* cell instance $22873 r0 *1 14.915,88.41
X$22873 2341 VIA_via1_7
* cell instance $22874 r0 *1 14.915,88.41
X$22874 2341 VIA_via2_5
* cell instance $22875 r0 *1 13.585,88.41
X$22875 2341 VIA_via2_5
* cell instance $22876 r0 *1 13.585,87.57
X$22876 2341 VIA_via1_4
* cell instance $22877 r0 *1 84.645,87.99
X$22877 2342 VIA_via1_7
* cell instance $22878 r0 *1 84.645,88.69
X$22878 2342 VIA_via1_4
* cell instance $22879 r0 *1 82.175,88.83
X$22879 2343 VIA_via1_4
* cell instance $22880 r0 *1 82.175,88.69
X$22880 2343 VIA_via2_5
* cell instance $22881 r0 *1 85.025,88.69
X$22881 2343 VIA_via1_4
* cell instance $22882 r0 *1 85.025,88.69
X$22882 2343 VIA_via2_5
* cell instance $22883 r0 *1 20.045,88.41
X$22883 2344 VIA_via1_7
* cell instance $22884 r0 *1 20.045,88.41
X$22884 2344 VIA_via2_5
* cell instance $22885 r0 *1 18.715,88.41
X$22885 2344 VIA_via2_5
* cell instance $22886 r0 *1 18.715,87.57
X$22886 2344 VIA_via1_4
* cell instance $22887 r0 *1 64.695,87.99
X$22887 2345 VIA_via1_7
* cell instance $22888 r0 *1 64.695,87.99
X$22888 2345 VIA_via2_5
* cell instance $22889 r0 *1 66.405,87.99
X$22889 2345 VIA_via2_5
* cell instance $22890 r0 *1 66.405,88.83
X$22890 2345 VIA_via1_4
* cell instance $22891 r0 *1 49.305,87.99
X$22891 2346 VIA_via1_7
* cell instance $22892 r0 *1 49.305,87.99
X$22892 2346 VIA_via2_5
* cell instance $22893 r0 *1 50.065,87.99
X$22893 2346 VIA_via2_5
* cell instance $22894 r0 *1 50.065,87.57
X$22894 2346 VIA_via1_4
* cell instance $22895 r0 *1 38.665,88.41
X$22895 2347 VIA_via1_7
* cell instance $22896 r0 *1 38.665,88.41
X$22896 2347 VIA_via2_5
* cell instance $22897 r0 *1 35.815,88.41
X$22897 2347 VIA_via2_5
* cell instance $22898 r0 *1 35.815,87.57
X$22898 2347 VIA_via1_4
* cell instance $22899 r0 *1 42.655,87.99
X$22899 2348 VIA_via1_7
* cell instance $22900 r0 *1 39.995,88.41
X$22900 2348 VIA_via2_5
* cell instance $22901 r0 *1 42.655,88.41
X$22901 2348 VIA_via2_5
* cell instance $22902 r0 *1 39.995,88.83
X$22902 2348 VIA_via1_4
* cell instance $22903 r0 *1 12.255,89.39
X$22903 2349 VIA_via1_7
* cell instance $22904 r0 *1 12.445,90.37
X$22904 2349 VIA_via1_4
* cell instance $22905 r0 *1 13.015,89.39
X$22905 2350 VIA_via1_7
* cell instance $22906 r0 *1 13.015,90.09
X$22906 2350 VIA_via2_5
* cell instance $22907 r0 *1 12.255,90.37
X$22907 2350 VIA_via1_4
* cell instance $22908 r0 *1 12.255,90.37
X$22908 2350 VIA_via2_5
* cell instance $22909 r0 *1 13.395,91.21
X$22909 2351 VIA_via1_7
* cell instance $22910 r0 *1 13.205,90.37
X$22910 2351 VIA_via1_4
* cell instance $22911 r0 *1 20.615,90.37
X$22911 2352 VIA_via1_4
* cell instance $22912 r0 *1 21.185,90.09
X$22912 2352 VIA_via1_4
* cell instance $22913 r0 *1 21.755,91.21
X$22913 2353 VIA_via1_7
* cell instance $22914 r0 *1 20.995,90.37
X$22914 2353 VIA_via1_4
* cell instance $22915 r0 *1 29.355,89.39
X$22915 2354 VIA_via1_7
* cell instance $22916 r0 *1 28.975,90.37
X$22916 2354 VIA_via1_4
* cell instance $22917 r0 *1 29.925,94.43
X$22917 2355 VIA_via2_5
* cell instance $22918 r0 *1 32.395,94.43
X$22918 2355 VIA_via2_5
* cell instance $22919 r0 *1 34.675,94.43
X$22919 2355 VIA_via2_5
* cell instance $22920 r0 *1 37.145,94.43
X$22920 2355 VIA_via2_5
* cell instance $22921 r0 *1 32.395,95.55
X$22921 2355 VIA_via1_4
* cell instance $22922 r0 *1 26.505,93.17
X$22922 2355 VIA_via1_4
* cell instance $22923 r0 *1 26.695,94.43
X$22923 2355 VIA_via1_4
* cell instance $22924 r0 *1 26.695,94.43
X$22924 2355 VIA_via2_5
* cell instance $22925 r0 *1 34.675,95.97
X$22925 2355 VIA_via1_4
* cell instance $22926 r0 *1 34.295,94.43
X$22926 2355 VIA_via1_4
* cell instance $22927 r0 *1 34.295,94.43
X$22927 2355 VIA_via2_5
* cell instance $22928 r0 *1 30.875,94.43
X$22928 2355 VIA_via1_4
* cell instance $22929 r0 *1 30.875,94.43
X$22929 2355 VIA_via2_5
* cell instance $22930 r0 *1 29.735,90.37
X$22930 2355 VIA_via1_4
* cell instance $22931 r0 *1 37.335,94.43
X$22931 2355 VIA_via1_4
* cell instance $22932 r0 *1 37.145,93.17
X$22932 2355 VIA_via1_4
* cell instance $22933 r0 *1 31.065,89.25
X$22933 2356 VIA_via2_5
* cell instance $22934 r0 *1 31.635,89.25
X$22934 2356 VIA_via2_5
* cell instance $22935 r0 *1 31.255,89.95
X$22935 2356 VIA_via1_4
* cell instance $22936 r0 *1 31.065,88.83
X$22936 2356 VIA_via1_4
* cell instance $22937 r0 *1 31.065,88.83
X$22937 2356 VIA_via2_5
* cell instance $22938 r0 *1 28.405,88.83
X$22938 2356 VIA_via1_4
* cell instance $22939 r0 *1 28.405,88.83
X$22939 2356 VIA_via2_5
* cell instance $22940 r0 *1 33.155,91.21
X$22940 2357 VIA_via1_7
* cell instance $22941 r0 *1 33.345,88.83
X$22941 2357 VIA_via1_4
* cell instance $22942 r0 *1 37.145,90.37
X$22942 2358 VIA_via1_4
* cell instance $22943 r0 *1 37.145,90.37
X$22943 2358 VIA_via2_5
* cell instance $22944 r0 *1 37.335,89.25
X$22944 2358 VIA_via1_4
* cell instance $22945 r0 *1 35.815,90.37
X$22945 2358 VIA_via1_4
* cell instance $22946 r0 *1 35.815,90.37
X$22946 2358 VIA_via2_5
* cell instance $22947 r0 *1 39.615,90.37
X$22947 2359 VIA_via1_4
* cell instance $22948 r0 *1 40.185,94.57
X$22948 2359 VIA_via1_4
* cell instance $22949 r0 *1 39.995,89.95
X$22949 2360 VIA_via1_4
* cell instance $22950 r0 *1 39.995,90.09
X$22950 2360 VIA_via2_5
* cell instance $22951 r0 *1 41.325,90.37
X$22951 2360 VIA_via1_4
* cell instance $22952 r0 *1 41.325,90.37
X$22952 2360 VIA_via2_5
* cell instance $22953 r0 *1 43.605,89.39
X$22953 2361 VIA_via1_7
* cell instance $22954 r0 *1 43.415,90.37
X$22954 2361 VIA_via1_4
* cell instance $22955 r0 *1 53.485,90.37
X$22955 2362 VIA_via1_4
* cell instance $22956 r0 *1 53.485,90.37
X$22956 2362 VIA_via2_5
* cell instance $22957 r0 *1 54.435,90.37
X$22957 2362 VIA_via1_4
* cell instance $22958 r0 *1 54.435,90.37
X$22958 2362 VIA_via2_5
* cell instance $22959 r0 *1 49.305,90.37
X$22959 2362 VIA_via1_4
* cell instance $22960 r0 *1 49.305,90.37
X$22960 2362 VIA_via2_5
* cell instance $22961 r0 *1 56.715,92.05
X$22961 2363 VIA_via2_5
* cell instance $22962 r0 *1 55.575,92.05
X$22962 2363 VIA_via2_5
* cell instance $22963 r0 *1 58.045,92.05
X$22963 2363 VIA_via1_4
* cell instance $22964 r0 *1 58.045,92.05
X$22964 2363 VIA_via2_5
* cell instance $22965 r0 *1 55.765,93.17
X$22965 2363 VIA_via1_4
* cell instance $22966 r0 *1 56.525,90.37
X$22966 2363 VIA_via1_4
* cell instance $22967 r0 *1 68.685,91.91
X$22967 2364 VIA_via1_7
* cell instance $22968 r0 *1 66.595,90.23
X$22968 2364 VIA_via2_5
* cell instance $22969 r0 *1 68.495,90.23
X$22969 2364 VIA_via2_5
* cell instance $22970 r0 *1 66.595,88.83
X$22970 2364 VIA_via1_4
* cell instance $22971 r0 *1 67.545,90.37
X$22971 2364 VIA_via1_4
* cell instance $22972 r0 *1 67.545,90.23
X$22972 2364 VIA_via2_5
* cell instance $22973 r0 *1 69.635,90.37
X$22973 2365 VIA_via1_4
* cell instance $22974 r0 *1 70.395,90.09
X$22974 2365 VIA_via1_4
* cell instance $22975 r0 *1 73.625,89.39
X$22975 2366 VIA_via1_7
* cell instance $22976 r0 *1 74.195,90.37
X$22976 2366 VIA_via1_4
* cell instance $22977 r0 *1 75.715,89.39
X$22977 2367 VIA_via1_7
* cell instance $22978 r0 *1 75.335,90.37
X$22978 2367 VIA_via1_4
* cell instance $22979 r0 *1 81.985,89.11
X$22979 2368 VIA_via1_4
* cell instance $22980 r0 *1 82.935,88.83
X$22980 2368 VIA_via1_4
* cell instance $22981 r0 *1 85.405,91.91
X$22981 2369 VIA_via2_5
* cell instance $22982 r0 *1 85.215,90.65
X$22982 2369 VIA_via2_5
* cell instance $22983 r0 *1 85.215,91.35
X$22983 2369 VIA_via2_5
* cell instance $22984 r0 *1 84.835,95.97
X$22984 2369 VIA_via1_4
* cell instance $22985 r0 *1 85.215,90.37
X$22985 2369 VIA_via1_4
* cell instance $22986 r0 *1 83.885,90.65
X$22986 2369 VIA_via1_4
* cell instance $22987 r0 *1 83.885,90.65
X$22987 2369 VIA_via2_5
* cell instance $22988 r0 *1 81.415,88.83
X$22988 2369 VIA_via1_4
* cell instance $22989 r0 *1 81.415,88.97
X$22989 2369 VIA_via2_5
* cell instance $22990 r0 *1 83.885,88.83
X$22990 2369 VIA_via1_4
* cell instance $22991 r0 *1 83.885,88.97
X$22991 2369 VIA_via2_5
* cell instance $22992 r0 *1 86.165,88.83
X$22992 2369 VIA_via1_4
* cell instance $22993 r0 *1 86.165,88.97
X$22993 2369 VIA_via2_5
* cell instance $22994 r0 *1 86.735,91.21
X$22994 2370 VIA_via1_7
* cell instance $22995 r0 *1 86.735,91.21
X$22995 2370 VIA_via2_5
* cell instance $22996 r0 *1 85.025,91.21
X$22996 2370 VIA_via2_5
* cell instance $22997 r0 *1 85.405,91.21
X$22997 2370 VIA_via2_5
* cell instance $22998 r0 *1 85.405,88.83
X$22998 2370 VIA_via2_5
* cell instance $22999 r0 *1 85.025,90.37
X$22999 2370 VIA_via1_4
* cell instance $23000 r0 *1 84.455,88.83
X$23000 2370 VIA_via1_4
* cell instance $23001 r0 *1 84.455,88.83
X$23001 2370 VIA_via2_5
* cell instance $23002 r0 *1 85.785,88.83
X$23002 2370 VIA_via1_4
* cell instance $23003 r0 *1 89.775,89.39
X$23003 2371 VIA_via1_7
* cell instance $23004 r0 *1 90.155,90.37
X$23004 2371 VIA_via1_4
* cell instance $23005 r0 *1 91.485,90.37
X$23005 2372 VIA_via1_4
* cell instance $23006 r0 *1 90.535,90.09
X$23006 2372 VIA_via1_4
* cell instance $23007 r0 *1 87.115,93.59
X$23007 2373 VIA_via1_7
* cell instance $23008 r0 *1 90.915,90.37
X$23008 2373 VIA_via2_5
* cell instance $23009 r0 *1 88.065,94.43
X$23009 2373 VIA_via2_5
* cell instance $23010 r0 *1 87.115,94.43
X$23010 2373 VIA_via2_5
* cell instance $23011 r0 *1 90.915,94.43
X$23011 2373 VIA_via2_5
* cell instance $23012 r0 *1 93.955,90.37
X$23012 2373 VIA_via2_5
* cell instance $23013 r0 *1 82.365,94.43
X$23013 2373 VIA_via2_5
* cell instance $23014 r0 *1 85.405,94.43
X$23014 2373 VIA_via1_4
* cell instance $23015 r0 *1 85.405,94.43
X$23015 2373 VIA_via2_5
* cell instance $23016 r0 *1 81.795,94.43
X$23016 2373 VIA_via1_4
* cell instance $23017 r0 *1 81.795,94.43
X$23017 2373 VIA_via2_5
* cell instance $23018 r0 *1 82.365,90.37
X$23018 2373 VIA_via1_4
* cell instance $23019 r0 *1 93.955,88.83
X$23019 2373 VIA_via1_4
* cell instance $23020 r0 *1 92.245,90.37
X$23020 2373 VIA_via1_4
* cell instance $23021 r0 *1 92.245,90.37
X$23021 2373 VIA_via2_5
* cell instance $23022 r0 *1 89.015,94.43
X$23022 2373 VIA_via1_4
* cell instance $23023 r0 *1 89.015,94.43
X$23023 2373 VIA_via2_5
* cell instance $23024 r0 *1 88.065,95.97
X$23024 2373 VIA_via1_4
* cell instance $23025 r0 *1 90.915,93.17
X$23025 2373 VIA_via1_4
* cell instance $23026 r0 *1 95.285,90.23
X$23026 2374 VIA_via1_4
* cell instance $23027 r0 *1 95.295,90.23
X$23027 2374 VIA_via3_2
* cell instance $23028 r0 *1 95.285,90.23
X$23028 2374 VIA_via2_5
* cell instance $23029 r0 *1 95.295,91.35
X$23029 2374 VIA_via4_0
* cell instance $23030 r0 *1 5.605,88.97
X$23030 2375 VIA_via1_4
* cell instance $23031 r0 *1 5.605,88.97
X$23031 2375 VIA_via2_5
* cell instance $23032 r0 *1 11.875,88.83
X$23032 2375 VIA_via1_4
* cell instance $23033 r0 *1 11.875,88.97
X$23033 2375 VIA_via2_5
* cell instance $23034 r0 *1 89.395,90.23
X$23034 2376 VIA_via1_7
* cell instance $23035 r0 *1 89.395,90.23
X$23035 2376 VIA_via2_5
* cell instance $23036 r0 *1 87.115,90.23
X$23036 2376 VIA_via1_4
* cell instance $23037 r0 *1 87.115,90.23
X$23037 2376 VIA_via2_5
* cell instance $23038 r0 *1 88.635,89.39
X$23038 2377 VIA_via1_7
* cell instance $23039 r0 *1 88.635,89.39
X$23039 2377 VIA_via2_5
* cell instance $23040 r0 *1 89.585,89.39
X$23040 2377 VIA_via2_5
* cell instance $23041 r0 *1 89.585,90.37
X$23041 2377 VIA_via1_4
* cell instance $23042 r0 *1 86.355,89.39
X$23042 2378 VIA_via1_7
* cell instance $23043 r0 *1 86.355,89.81
X$23043 2378 VIA_via2_5
* cell instance $23044 r0 *1 88.635,89.81
X$23044 2378 VIA_via2_5
* cell instance $23045 r0 *1 88.635,90.37
X$23045 2378 VIA_via1_4
* cell instance $23046 r0 *1 87.305,93.03
X$23046 2379 VIA_via1_7
* cell instance $23047 r0 *1 87.495,89.11
X$23047 2379 VIA_via2_5
* cell instance $23048 r0 *1 88.065,89.11
X$23048 2379 VIA_via1_4
* cell instance $23049 r0 *1 88.065,89.11
X$23049 2379 VIA_via2_5
* cell instance $23050 r0 *1 16.815,88.83
X$23050 2380 VIA_via1_4
* cell instance $23051 r0 *1 16.625,88.83
X$23051 2380 VIA_via1_4
* cell instance $23052 r0 *1 19.665,89.25
X$23052 2381 VIA_via2_5
* cell instance $23053 r0 *1 19.665,90.37
X$23053 2381 VIA_via1_4
* cell instance $23054 r0 *1 20.425,89.11
X$23054 2381 VIA_via1_4
* cell instance $23055 r0 *1 20.425,89.25
X$23055 2381 VIA_via2_5
* cell instance $23056 r0 *1 20.235,88.83
X$23056 2382 VIA_via1_4
* cell instance $23057 r0 *1 20.235,88.83
X$23057 2382 VIA_via2_5
* cell instance $23058 r0 *1 21.945,88.83
X$23058 2382 VIA_via1_4
* cell instance $23059 r0 *1 21.945,88.83
X$23059 2382 VIA_via2_5
* cell instance $23060 r0 *1 24.415,88.83
X$23060 2383 VIA_via1_4
* cell instance $23061 r0 *1 24.415,88.83
X$23061 2383 VIA_via2_5
* cell instance $23062 r0 *1 28.025,88.83
X$23062 2383 VIA_via1_4
* cell instance $23063 r0 *1 28.025,88.83
X$23063 2383 VIA_via2_5
* cell instance $23064 r0 *1 31.635,88.83
X$23064 2384 VIA_via1_4
* cell instance $23065 r0 *1 31.445,88.83
X$23065 2384 VIA_via1_4
* cell instance $23066 r0 *1 32.585,88.83
X$23066 2385 VIA_via1_4
* cell instance $23067 r0 *1 32.585,88.83
X$23067 2385 VIA_via2_5
* cell instance $23068 r0 *1 31.825,88.83
X$23068 2385 VIA_via1_4
* cell instance $23069 r0 *1 31.825,88.83
X$23069 2385 VIA_via2_5
* cell instance $23070 r0 *1 36.765,89.81
X$23070 2386 VIA_via1_7
* cell instance $23071 r0 *1 36.765,89.81
X$23071 2386 VIA_via2_5
* cell instance $23072 r0 *1 35.055,89.81
X$23072 2386 VIA_via2_5
* cell instance $23073 r0 *1 35.055,88.83
X$23073 2386 VIA_via1_4
* cell instance $23074 r0 *1 80.085,90.09
X$23074 2387 VIA_via2_5
* cell instance $23075 r0 *1 80.085,90.37
X$23075 2387 VIA_via1_4
* cell instance $23076 r0 *1 85.025,90.09
X$23076 2387 VIA_via1_4
* cell instance $23077 r0 *1 85.025,90.09
X$23077 2387 VIA_via2_5
* cell instance $23078 r0 *1 82.365,88.83
X$23078 2388 VIA_via1_4
* cell instance $23079 r0 *1 82.365,88.83
X$23079 2388 VIA_via2_5
* cell instance $23080 r0 *1 83.695,88.83
X$23080 2388 VIA_via1_4
* cell instance $23081 r0 *1 83.695,88.83
X$23081 2388 VIA_via2_5
* cell instance $23082 r0 *1 83.315,89.39
X$23082 2389 VIA_via1_7
* cell instance $23083 r0 *1 83.315,89.39
X$23083 2389 VIA_via2_5
* cell instance $23084 r0 *1 81.605,89.39
X$23084 2389 VIA_via2_5
* cell instance $23085 r0 *1 81.605,90.37
X$23085 2389 VIA_via1_4
* cell instance $23086 r0 *1 38.475,90.23
X$23086 2390 VIA_via1_4
* cell instance $23087 r0 *1 38.475,90.23
X$23087 2390 VIA_via2_5
* cell instance $23088 r0 *1 40.565,90.37
X$23088 2390 VIA_via1_4
* cell instance $23089 r0 *1 40.565,90.23
X$23089 2390 VIA_via2_5
* cell instance $23090 r0 *1 68.875,90.23
X$23090 2391 VIA_via1_7
* cell instance $23091 r0 *1 68.875,90.23
X$23091 2391 VIA_via2_5
* cell instance $23092 r0 *1 73.815,90.09
X$23092 2391 VIA_via1_4
* cell instance $23093 r0 *1 73.815,90.23
X$23093 2391 VIA_via2_5
* cell instance $23094 r0 *1 44.935,88.83
X$23094 2392 VIA_via1_4
* cell instance $23095 r0 *1 44.935,88.83
X$23095 2392 VIA_via2_5
* cell instance $23096 r0 *1 48.545,88.83
X$23096 2392 VIA_via1_4
* cell instance $23097 r0 *1 48.545,88.83
X$23097 2392 VIA_via2_5
* cell instance $23098 r0 *1 51.205,90.37
X$23098 2393 VIA_via1_4
* cell instance $23099 r0 *1 51.205,90.23
X$23099 2393 VIA_via2_5
* cell instance $23100 r0 *1 50.255,90.23
X$23100 2393 VIA_via1_4
* cell instance $23101 r0 *1 50.255,90.23
X$23101 2393 VIA_via2_5
* cell instance $23102 r0 *1 63.555,88.97
X$23102 2394 VIA_via1_7
* cell instance $23103 r0 *1 63.555,88.97
X$23103 2394 VIA_via2_5
* cell instance $23104 r0 *1 66.025,89.11
X$23104 2394 VIA_via1_4
* cell instance $23105 r0 *1 66.025,88.97
X$23105 2394 VIA_via2_5
* cell instance $23106 r0 *1 51.585,88.83
X$23106 2395 VIA_via1_4
* cell instance $23107 r0 *1 50.635,88.83
X$23107 2395 VIA_via1_4
* cell instance $23108 r0 *1 64.695,89.39
X$23108 2396 VIA_via1_7
* cell instance $23109 r0 *1 64.695,89.39
X$23109 2396 VIA_via2_5
* cell instance $23110 r0 *1 65.265,89.39
X$23110 2396 VIA_via2_5
* cell instance $23111 r0 *1 65.265,90.37
X$23111 2396 VIA_via1_4
* cell instance $23112 r0 *1 49.685,88.83
X$23112 2397 VIA_via1_4
* cell instance $23113 r0 *1 49.685,88.83
X$23113 2397 VIA_via2_5
* cell instance $23114 r0 *1 53.865,88.83
X$23114 2397 VIA_via1_4
* cell instance $23115 r0 *1 53.865,88.83
X$23115 2397 VIA_via2_5
* cell instance $23116 r0 *1 53.865,90.37
X$23116 2397 VIA_via1_4
* cell instance $23117 r0 *1 57.475,89.81
X$23117 2398 VIA_via1_7
* cell instance $23118 r0 *1 57.475,88.83
X$23118 2398 VIA_via2_5
* cell instance $23119 r0 *1 55.955,88.83
X$23119 2398 VIA_via1_4
* cell instance $23120 r0 *1 55.955,88.83
X$23120 2398 VIA_via2_5
* cell instance $23121 r0 *1 41.895,90.65
X$23121 2399 VIA_via1_4
* cell instance $23122 r0 *1 41.515,90.37
X$23122 2399 VIA_via1_4
* cell instance $23123 r0 *1 46.835,90.79
X$23123 2400 VIA_via1_7
* cell instance $23124 r0 *1 46.455,91.63
X$23124 2400 VIA_via1_4
* cell instance $23125 r0 *1 48.735,91.35
X$23125 2401 VIA_via1_4
* cell instance $23126 r0 *1 48.355,90.37
X$23126 2401 VIA_via1_4
* cell instance $23127 r0 *1 48.355,90.37
X$23127 2401 VIA_via2_5
* cell instance $23128 r0 *1 45.885,90.37
X$23128 2401 VIA_via1_4
* cell instance $23129 r0 *1 45.885,90.37
X$23129 2401 VIA_via2_5
* cell instance $23130 r0 *1 61.275,90.51
X$23130 2402 VIA_via2_5
* cell instance $23131 r0 *1 58.805,90.37
X$23131 2402 VIA_via1_4
* cell instance $23132 r0 *1 58.805,90.51
X$23132 2402 VIA_via2_5
* cell instance $23133 r0 *1 57.095,90.37
X$23133 2402 VIA_via1_4
* cell instance $23134 r0 *1 57.095,90.51
X$23134 2402 VIA_via2_5
* cell instance $23135 r0 *1 61.275,91.35
X$23135 2402 VIA_via1_4
* cell instance $23136 r0 *1 59.185,90.79
X$23136 2403 VIA_via1_7
* cell instance $23137 r0 *1 59.565,91.21
X$23137 2403 VIA_via2_5
* cell instance $23138 r0 *1 58.995,91.21
X$23138 2403 VIA_via2_5
* cell instance $23139 r0 *1 58.995,91.63
X$23139 2403 VIA_via1_4
* cell instance $23140 r0 *1 70.015,90.79
X$23140 2404 VIA_via1_7
* cell instance $23141 r0 *1 70.015,90.79
X$23141 2404 VIA_via2_5
* cell instance $23142 r0 *1 62.035,90.79
X$23142 2404 VIA_via2_5
* cell instance $23143 r0 *1 65.455,90.79
X$23143 2404 VIA_via2_5
* cell instance $23144 r0 *1 65.455,91.63
X$23144 2404 VIA_via1_4
* cell instance $23145 r0 *1 62.035,90.37
X$23145 2404 VIA_via1_4
* cell instance $23146 r0 *1 68.685,90.51
X$23146 2405 VIA_via1_4
* cell instance $23147 r0 *1 69.065,90.37
X$23147 2405 VIA_via1_4
* cell instance $23148 r0 *1 73.435,90.79
X$23148 2406 VIA_via1_7
* cell instance $23149 r0 *1 73.435,91.63
X$23149 2406 VIA_via1_4
* cell instance $23150 r0 *1 72.865,91.63
X$23150 2406 VIA_via1_4
* cell instance $23151 r0 *1 75.525,90.79
X$23151 2407 VIA_via1_7
* cell instance $23152 r0 *1 74.765,91.63
X$23152 2407 VIA_via1_4
* cell instance $23153 r0 *1 77.045,91.63
X$23153 2408 VIA_via1_4
* cell instance $23154 r0 *1 77.045,91.63
X$23154 2408 VIA_via2_5
* cell instance $23155 r0 *1 74.195,91.63
X$23155 2408 VIA_via1_4
* cell instance $23156 r0 *1 74.195,91.63
X$23156 2408 VIA_via2_5
* cell instance $23157 r0 *1 76.095,91.63
X$23157 2408 VIA_via1_4
* cell instance $23158 r0 *1 76.095,91.63
X$23158 2408 VIA_via2_5
* cell instance $23159 r0 *1 75.715,91.63
X$23159 2408 VIA_via1_4
* cell instance $23160 r0 *1 75.715,91.63
X$23160 2408 VIA_via2_5
* cell instance $23161 r0 *1 78.185,91.91
X$23161 2409 VIA_via1_7
* cell instance $23162 r0 *1 78.185,91.63
X$23162 2409 VIA_via2_5
* cell instance $23163 r0 *1 77.615,91.63
X$23163 2409 VIA_via2_5
* cell instance $23164 r0 *1 75.715,95.69
X$23164 2409 VIA_via2_5
* cell instance $23165 r0 *1 77.995,95.69
X$23165 2409 VIA_via2_5
* cell instance $23166 r0 *1 77.615,95.69
X$23166 2409 VIA_via2_5
* cell instance $23167 r0 *1 76.855,91.63
X$23167 2409 VIA_via1_4
* cell instance $23168 r0 *1 76.855,91.49
X$23168 2409 VIA_via2_5
* cell instance $23169 r0 *1 74.195,94.15
X$23169 2409 VIA_via1_4
* cell instance $23170 r0 *1 74.575,94.43
X$23170 2409 VIA_via1_4
* cell instance $23171 r0 *1 74.575,94.29
X$23171 2409 VIA_via2_5
* cell instance $23172 r0 *1 75.145,91.63
X$23172 2409 VIA_via1_4
* cell instance $23173 r0 *1 75.145,91.49
X$23173 2409 VIA_via2_5
* cell instance $23174 r0 *1 75.715,94.43
X$23174 2409 VIA_via1_4
* cell instance $23175 r0 *1 75.715,94.57
X$23175 2409 VIA_via2_5
* cell instance $23176 r0 *1 77.995,95.97
X$23176 2409 VIA_via1_4
* cell instance $23177 r0 *1 79.895,93.03
X$23177 2410 VIA_via1_7
* cell instance $23178 r0 *1 80.275,90.65
X$23178 2410 VIA_via1_7
* cell instance $23179 r0 *1 83.695,94.29
X$23179 2411 VIA_via2_5
* cell instance $23180 r0 *1 83.885,94.29
X$23180 2411 VIA_via2_5
* cell instance $23181 r0 *1 83.695,95.97
X$23181 2411 VIA_via1_4
* cell instance $23182 r0 *1 85.215,91.63
X$23182 2411 VIA_via1_4
* cell instance $23183 r0 *1 85.215,91.63
X$23183 2411 VIA_via2_5
* cell instance $23184 r0 *1 83.505,91.63
X$23184 2411 VIA_via1_4
* cell instance $23185 r0 *1 83.505,91.63
X$23185 2411 VIA_via2_5
* cell instance $23186 r0 *1 85.595,91.49
X$23186 2411 VIA_via1_4
* cell instance $23187 r0 *1 86.925,94.29
X$23187 2411 VIA_via1_4
* cell instance $23188 r0 *1 86.925,94.29
X$23188 2411 VIA_via2_5
* cell instance $23189 r0 *1 88.635,94.15
X$23189 2412 VIA_via2_5
* cell instance $23190 r0 *1 89.015,94.15
X$23190 2412 VIA_via2_5
* cell instance $23191 r0 *1 85.595,94.15
X$23191 2412 VIA_via2_5
* cell instance $23192 r0 *1 85.595,93.17
X$23192 2412 VIA_via1_4
* cell instance $23193 r0 *1 85.785,91.63
X$23193 2412 VIA_via1_4
* cell instance $23194 r0 *1 89.015,93.17
X$23194 2412 VIA_via1_4
* cell instance $23195 r0 *1 90.535,94.15
X$23195 2412 VIA_via1_4
* cell instance $23196 r0 *1 90.535,94.15
X$23196 2412 VIA_via2_5
* cell instance $23197 r0 *1 88.635,95.97
X$23197 2412 VIA_via1_4
* cell instance $23198 r0 *1 85.975,90.51
X$23198 2412 VIA_via1_4
* cell instance $23199 r0 *1 86.355,91.35
X$23199 2413 VIA_via1_4
* cell instance $23200 r0 *1 86.545,91.63
X$23200 2413 VIA_via1_4
* cell instance $23201 r0 *1 91.485,93.45
X$23201 2414 VIA_via2_5
* cell instance $23202 r0 *1 87.875,93.45
X$23202 2414 VIA_via2_5
* cell instance $23203 r0 *1 87.875,91.63
X$23203 2414 VIA_via1_4
* cell instance $23204 r0 *1 87.685,90.37
X$23204 2414 VIA_via1_4
* cell instance $23205 r0 *1 88.065,91.63
X$23205 2414 VIA_via1_4
* cell instance $23206 r0 *1 92.435,93.45
X$23206 2414 VIA_via1_4
* cell instance $23207 r0 *1 92.435,93.45
X$23207 2414 VIA_via2_5
* cell instance $23208 r0 *1 91.485,95.97
X$23208 2414 VIA_via1_4
* cell instance $23209 r0 *1 88.635,91.35
X$23209 2415 VIA_via1_4
* cell instance $23210 r0 *1 89.015,91.63
X$23210 2415 VIA_via1_4
* cell instance $23211 r0 *1 94.335,90.37
X$23211 2416 VIA_via1_4
* cell instance $23212 r0 *1 94.335,90.51
X$23212 2416 VIA_via2_5
* cell instance $23213 r0 *1 93.765,90.51
X$23213 2416 VIA_via1_4
* cell instance $23214 r0 *1 93.765,90.51
X$23214 2416 VIA_via2_5
* cell instance $23215 r0 *1 94.905,90.37
X$23215 2416 VIA_via1_4
* cell instance $23216 r0 *1 94.905,90.51
X$23216 2416 VIA_via2_5
* cell instance $23217 r0 *1 95.855,90.23
X$23217 2417 VIA_via1_4
* cell instance $23218 r0 *1 95.855,90.23
X$23218 2417 VIA_via2_5
* cell instance $23219 r0 *1 95.855,90.23
X$23219 2417 VIA_via3_2
* cell instance $23220 r0 *1 95.855,90.79
X$23220 2417 VIA_via4_0
* cell instance $23221 r0 *1 9.595,94.01
X$23221 2418 VIA_via1_7
* cell instance $23222 r0 *1 10.735,91.49
X$23222 2418 VIA_via2_5
* cell instance $23223 r0 *1 9.785,91.49
X$23223 2418 VIA_via2_5
* cell instance $23224 r0 *1 10.735,90.37
X$23224 2418 VIA_via1_4
* cell instance $23225 r0 *1 13.015,90.37
X$23225 2419 VIA_via1_4
* cell instance $23226 r0 *1 13.015,90.51
X$23226 2419 VIA_via2_5
* cell instance $23227 r0 *1 10.925,90.51
X$23227 2419 VIA_via1_4
* cell instance $23228 r0 *1 10.925,90.51
X$23228 2419 VIA_via2_5
* cell instance $23229 r0 *1 17.195,89.39
X$23229 2420 VIA_via1_7
* cell instance $23230 r0 *1 17.195,90.51
X$23230 2420 VIA_via2_5
* cell instance $23231 r0 *1 19.855,90.37
X$23231 2420 VIA_via1_4
* cell instance $23232 r0 *1 19.855,90.51
X$23232 2420 VIA_via2_5
* cell instance $23233 r0 *1 18.715,90.37
X$23233 2421 VIA_via1_4
* cell instance $23234 r0 *1 18.715,90.37
X$23234 2421 VIA_via2_5
* cell instance $23235 r0 *1 20.425,90.37
X$23235 2421 VIA_via1_4
* cell instance $23236 r0 *1 20.425,90.37
X$23236 2421 VIA_via2_5
* cell instance $23237 r0 *1 84.835,90.37
X$23237 2422 VIA_via1_4
* cell instance $23238 r0 *1 84.835,90.51
X$23238 2422 VIA_via2_5
* cell instance $23239 r0 *1 88.445,90.51
X$23239 2422 VIA_via1_4
* cell instance $23240 r0 *1 88.445,90.51
X$23240 2422 VIA_via2_5
* cell instance $23241 r0 *1 84.075,90.37
X$23241 2423 VIA_via1_4
* cell instance $23242 r0 *1 84.075,90.37
X$23242 2423 VIA_via2_5
* cell instance $23243 r0 *1 86.165,90.37
X$23243 2423 VIA_via1_4
* cell instance $23244 r0 *1 86.165,90.37
X$23244 2423 VIA_via2_5
* cell instance $23245 r0 *1 38.285,90.37
X$23245 2424 VIA_via1_4
* cell instance $23246 r0 *1 38.095,90.37
X$23246 2424 VIA_via1_4
* cell instance $23247 r0 *1 40.755,90.37
X$23247 2425 VIA_via1_4
* cell instance $23248 r0 *1 40.755,90.51
X$23248 2425 VIA_via2_5
* cell instance $23249 r0 *1 43.605,90.51
X$23249 2425 VIA_via1_4
* cell instance $23250 r0 *1 43.605,90.51
X$23250 2425 VIA_via2_5
* cell instance $23251 r0 *1 43.415,92.61
X$23251 2426 VIA_via1_7
* cell instance $23252 r0 *1 43.225,90.37
X$23252 2426 VIA_via2_5
* cell instance $23253 r0 *1 41.705,90.37
X$23253 2426 VIA_via1_4
* cell instance $23254 r0 *1 41.705,90.37
X$23254 2426 VIA_via2_5
* cell instance $23255 r0 *1 48.735,90.79
X$23255 2427 VIA_via1_7
* cell instance $23256 r0 *1 49.875,91.07
X$23256 2427 VIA_via2_5
* cell instance $23257 r0 *1 48.735,91.07
X$23257 2427 VIA_via2_5
* cell instance $23258 r0 *1 49.875,91.63
X$23258 2427 VIA_via1_4
* cell instance $23259 r0 *1 74.385,91.35
X$23259 2428 VIA_via1_7
* cell instance $23260 r0 *1 74.385,90.65
X$23260 2428 VIA_via2_5
* cell instance $23261 r0 *1 75.715,90.65
X$23261 2428 VIA_via1_4
* cell instance $23262 r0 *1 75.715,90.65
X$23262 2428 VIA_via2_5
* cell instance $23263 r0 *1 74.575,91.35
X$23263 2429 VIA_via2_5
* cell instance $23264 r0 *1 74.575,91.63
X$23264 2429 VIA_via1_4
* cell instance $23265 r0 *1 72.295,91.35
X$23265 2429 VIA_via1_4
* cell instance $23266 r0 *1 72.295,91.35
X$23266 2429 VIA_via2_5
* cell instance $23267 r0 *1 50.825,90.65
X$23267 2430 VIA_via2_5
* cell instance $23268 r0 *1 55.195,90.65
X$23268 2430 VIA_via2_5
* cell instance $23269 r0 *1 55.195,90.23
X$23269 2430 VIA_via1_4
* cell instance $23270 r0 *1 50.825,91.63
X$23270 2430 VIA_via1_4
* cell instance $23271 r0 *1 55.005,90.37
X$23271 2431 VIA_via1_4
* cell instance $23272 r0 *1 54.815,90.37
X$23272 2431 VIA_via1_4
* cell instance $23273 r0 *1 9.215,92.33
X$23273 2432 VIA_via2_5
* cell instance $23274 r0 *1 8.645,92.33
X$23274 2432 VIA_via2_5
* cell instance $23275 r0 *1 8.265,92.05
X$23275 2432 VIA_via1_4
* cell instance $23276 r0 *1 8.645,94.43
X$23276 2432 VIA_via1_4
* cell instance $23277 r0 *1 9.215,91.63
X$23277 2432 VIA_via1_4
* cell instance $23278 r0 *1 12.065,92.75
X$23278 2433 VIA_via2_5
* cell instance $23279 r0 *1 11.115,92.75
X$23279 2433 VIA_via2_5
* cell instance $23280 r0 *1 12.635,92.75
X$23280 2433 VIA_via1_4
* cell instance $23281 r0 *1 12.635,92.75
X$23281 2433 VIA_via2_5
* cell instance $23282 r0 *1 11.115,91.63
X$23282 2433 VIA_via1_4
* cell instance $23283 r0 *1 12.065,91.63
X$23283 2433 VIA_via1_4
* cell instance $23284 r0 *1 12.445,93.17
X$23284 2434 VIA_via2_5
* cell instance $23285 r0 *1 14.345,93.17
X$23285 2434 VIA_via2_5
* cell instance $23286 r0 *1 15.865,93.17
X$23286 2434 VIA_via2_5
* cell instance $23287 r0 *1 16.625,93.17
X$23287 2434 VIA_via2_5
* cell instance $23288 r0 *1 14.345,87.57
X$23288 2434 VIA_via1_4
* cell instance $23289 r0 *1 16.625,91.63
X$23289 2434 VIA_via1_4
* cell instance $23290 r0 *1 14.155,93.17
X$23290 2434 VIA_via1_4
* cell instance $23291 r0 *1 15.865,94.43
X$23291 2434 VIA_via1_4
* cell instance $23292 r0 *1 20.235,93.17
X$23292 2434 VIA_via1_4
* cell instance $23293 r0 *1 20.235,93.17
X$23293 2434 VIA_via2_5
* cell instance $23294 r0 *1 14.345,92.05
X$23294 2434 VIA_via1_4
* cell instance $23295 r0 *1 6.935,93.17
X$23295 2434 VIA_via1_4
* cell instance $23296 r0 *1 6.935,93.17
X$23296 2434 VIA_via2_5
* cell instance $23297 r0 *1 11.115,93.17
X$23297 2434 VIA_via1_4
* cell instance $23298 r0 *1 11.115,93.17
X$23298 2434 VIA_via2_5
* cell instance $23299 r0 *1 12.445,94.43
X$23299 2434 VIA_via1_4
* cell instance $23300 r0 *1 15.105,94.43
X$23300 2435 VIA_via1_4
* cell instance $23301 r0 *1 15.865,92.89
X$23301 2435 VIA_via1_4
* cell instance $23302 r0 *1 20.425,92.19
X$23302 2436 VIA_via1_7
* cell instance $23303 r0 *1 19.475,93.17
X$23303 2436 VIA_via1_4
* cell instance $23304 r0 *1 21.375,91.63
X$23304 2437 VIA_via1_4
* cell instance $23305 r0 *1 21.375,91.63
X$23305 2437 VIA_via2_5
* cell instance $23306 r0 *1 20.045,91.63
X$23306 2437 VIA_via1_4
* cell instance $23307 r0 *1 20.045,91.63
X$23307 2437 VIA_via2_5
* cell instance $23308 r0 *1 21.755,92.75
X$23308 2437 VIA_via1_4
* cell instance $23309 r0 *1 20.805,92.05
X$23309 2438 VIA_via2_5
* cell instance $23310 r0 *1 22.515,92.05
X$23310 2438 VIA_via2_5
* cell instance $23311 r0 *1 20.805,91.63
X$23311 2438 VIA_via1_4
* cell instance $23312 r0 *1 22.705,93.17
X$23312 2438 VIA_via1_4
* cell instance $23313 r0 *1 24.985,92.05
X$23313 2438 VIA_via1_4
* cell instance $23314 r0 *1 24.985,92.05
X$23314 2438 VIA_via2_5
* cell instance $23315 r0 *1 23.085,92.61
X$23315 2439 VIA_via1_7
* cell instance $23316 r0 *1 22.705,91.63
X$23316 2439 VIA_via1_4
* cell instance $23317 r0 *1 28.025,91.91
X$23317 2440 VIA_via2_5
* cell instance $23318 r0 *1 27.075,91.63
X$23318 2440 VIA_via1_4
* cell instance $23319 r0 *1 27.075,91.77
X$23319 2440 VIA_via2_5
* cell instance $23320 r0 *1 28.785,91.63
X$23320 2440 VIA_via1_4
* cell instance $23321 r0 *1 28.785,91.77
X$23321 2440 VIA_via2_5
* cell instance $23322 r0 *1 28.025,92.75
X$23322 2440 VIA_via1_4
* cell instance $23323 r0 *1 28.215,94.15
X$23323 2441 VIA_via1_4
* cell instance $23324 r0 *1 28.215,91.63
X$23324 2441 VIA_via1_4
* cell instance $23325 r0 *1 28.975,93.17
X$23325 2441 VIA_via1_4
* cell instance $23326 r0 *1 33.155,92.61
X$23326 2442 VIA_via1_7
* cell instance $23327 r0 *1 32.965,91.63
X$23327 2442 VIA_via1_4
* cell instance $23328 r0 *1 42.275,92.05
X$23328 2443 VIA_via1_4
* cell instance $23329 r0 *1 42.465,93.17
X$23329 2443 VIA_via1_4
* cell instance $23330 r0 *1 42.465,93.17
X$23330 2443 VIA_via2_5
* cell instance $23331 r0 *1 41.705,93.17
X$23331 2443 VIA_via1_4
* cell instance $23332 r0 *1 41.705,93.17
X$23332 2443 VIA_via2_5
* cell instance $23333 r0 *1 50.255,92.05
X$23333 2444 VIA_via1_4
* cell instance $23334 r0 *1 50.635,91.63
X$23334 2444 VIA_via1_4
* cell instance $23335 r0 *1 51.585,92.61
X$23335 2445 VIA_via1_7
* cell instance $23336 r0 *1 51.775,91.7
X$23336 2445 VIA_via1_4
* cell instance $23337 r0 *1 52.915,94.57
X$23337 2446 VIA_via2_5
* cell instance $23338 r0 *1 57.285,94.57
X$23338 2446 VIA_via1_4
* cell instance $23339 r0 *1 57.285,94.57
X$23339 2446 VIA_via2_5
* cell instance $23340 r0 *1 53.105,91.63
X$23340 2446 VIA_via1_4
* cell instance $23341 r0 *1 56.145,92.61
X$23341 2447 VIA_via1_7
* cell instance $23342 r0 *1 55.765,91.63
X$23342 2447 VIA_via1_4
* cell instance $23343 r0 *1 70.015,94.43
X$23343 2448 VIA_via1_4
* cell instance $23344 r0 *1 70.965,92.89
X$23344 2448 VIA_via1_4
* cell instance $23345 r0 *1 69.825,92.19
X$23345 2449 VIA_via1_7
* cell instance $23346 r0 *1 69.825,92.19
X$23346 2449 VIA_via2_5
* cell instance $23347 r0 *1 72.485,92.19
X$23347 2449 VIA_via2_5
* cell instance $23348 r0 *1 71.345,92.19
X$23348 2449 VIA_via2_5
* cell instance $23349 r0 *1 72.485,91.63
X$23349 2449 VIA_via1_4
* cell instance $23350 r0 *1 71.345,93.17
X$23350 2449 VIA_via1_4
* cell instance $23351 r0 *1 77.995,91.77
X$23351 2450 VIA_via1_7
* cell instance $23352 r0 *1 77.995,91.77
X$23352 2450 VIA_via2_5
* cell instance $23353 r0 *1 71.725,90.65
X$23353 2450 VIA_via1_7
* cell instance $23354 r0 *1 71.725,91.77
X$23354 2450 VIA_via2_5
* cell instance $23355 r0 *1 73.815,91.63
X$23355 2450 VIA_via1_4
* cell instance $23356 r0 *1 73.815,91.77
X$23356 2450 VIA_via2_5
* cell instance $23357 r0 *1 76.665,92.47
X$23357 2451 VIA_via2_5
* cell instance $23358 r0 *1 74.195,92.47
X$23358 2451 VIA_via2_5
* cell instance $23359 r0 *1 75.335,92.47
X$23359 2451 VIA_via2_5
* cell instance $23360 r0 *1 75.335,94.15
X$23360 2451 VIA_via2_5
* cell instance $23361 r0 *1 76.665,91.63
X$23361 2451 VIA_via1_4
* cell instance $23362 r0 *1 75.905,94.43
X$23362 2451 VIA_via1_4
* cell instance $23363 r0 *1 75.905,94.43
X$23363 2451 VIA_via2_5
* cell instance $23364 r0 *1 74.765,94.43
X$23364 2451 VIA_via1_4
* cell instance $23365 r0 *1 74.765,94.43
X$23365 2451 VIA_via2_5
* cell instance $23366 r0 *1 75.335,91.63
X$23366 2451 VIA_via1_4
* cell instance $23367 r0 *1 74.005,92.05
X$23367 2451 VIA_via1_4
* cell instance $23368 r0 *1 76.285,95.97
X$23368 2451 VIA_via1_4
* cell instance $23369 r0 *1 78.945,93.87
X$23369 2452 VIA_via2_5
* cell instance $23370 r0 *1 74.765,93.87
X$23370 2452 VIA_via2_5
* cell instance $23371 r0 *1 75.525,93.87
X$23371 2452 VIA_via2_5
* cell instance $23372 r0 *1 76.475,93.87
X$23372 2452 VIA_via2_5
* cell instance $23373 r0 *1 74.385,94.43
X$23373 2452 VIA_via1_4
* cell instance $23374 r0 *1 74.385,94.43
X$23374 2452 VIA_via2_5
* cell instance $23375 r0 *1 75.525,94.43
X$23375 2452 VIA_via1_4
* cell instance $23376 r0 *1 78.945,94.43
X$23376 2452 VIA_via1_4
* cell instance $23377 r0 *1 74.955,91.63
X$23377 2452 VIA_via1_4
* cell instance $23378 r0 *1 76.475,91.63
X$23378 2452 VIA_via1_4
* cell instance $23379 r0 *1 75.715,95.97
X$23379 2452 VIA_via1_4
* cell instance $23380 r0 *1 75.715,95.97
X$23380 2452 VIA_via2_5
* cell instance $23381 r0 *1 77.615,95.97
X$23381 2452 VIA_via1_4
* cell instance $23382 r0 *1 77.615,95.97
X$23382 2452 VIA_via2_5
* cell instance $23383 r0 *1 72.675,94.15
X$23383 2452 VIA_via1_4
* cell instance $23384 r0 *1 72.675,94.15
X$23384 2452 VIA_via2_5
* cell instance $23385 r0 *1 77.235,93.17
X$23385 2453 VIA_via1_4
* cell instance $23386 r0 *1 77.425,92.05
X$23386 2453 VIA_via1_4
* cell instance $23387 r0 *1 78.495,94.71
X$23387 2454 VIA_via5_0
* cell instance $23388 r0 *1 78.495,94.71
X$23388 2454 VIA_via4_0
* cell instance $23389 r0 *1 77.995,92.47
X$23389 2454 VIA_via2_5
* cell instance $23390 r0 *1 78.375,90.37
X$23390 2454 VIA_via1_4
* cell instance $23391 r0 *1 78.495,92.47
X$23391 2454 VIA_via3_2
* cell instance $23392 r0 *1 78.565,92.05
X$23392 2455 VIA_via1_7
* cell instance $23393 r0 *1 78.185,94.43
X$23393 2455 VIA_via1_4
* cell instance $23394 r0 *1 84.075,92.19
X$23394 2456 VIA_via1_7
* cell instance $23395 r0 *1 84.265,93.17
X$23395 2456 VIA_via1_4
* cell instance $23396 r0 *1 84.835,93.17
X$23396 2457 VIA_via1_4
* cell instance $23397 r0 *1 85.025,91.91
X$23397 2457 VIA_via1_4
* cell instance $23398 r0 *1 88.825,91.77
X$23398 2458 VIA_via1_7
* cell instance $23399 r0 *1 89.205,90.79
X$23399 2458 VIA_via1_7
* cell instance $23400 r0 *1 89.965,92.19
X$23400 2459 VIA_via1_7
* cell instance $23401 r0 *1 90.155,93.17
X$23401 2459 VIA_via1_4
* cell instance $23402 r0 *1 5.985,91.63
X$23402 2460 VIA_via1_4
* cell instance $23403 r0 *1 5.985,91.63
X$23403 2460 VIA_via2_5
* cell instance $23404 r0 *1 9.595,91.63
X$23404 2460 VIA_via1_4
* cell instance $23405 r0 *1 9.595,91.63
X$23405 2460 VIA_via2_5
* cell instance $23406 r0 *1 11.495,92.19
X$23406 2461 VIA_via1_7
* cell instance $23407 r0 *1 10.355,92.47
X$23407 2461 VIA_via2_5
* cell instance $23408 r0 *1 11.495,92.47
X$23408 2461 VIA_via2_5
* cell instance $23409 r0 *1 10.355,93.17
X$23409 2461 VIA_via1_4
* cell instance $23410 r0 *1 87.685,91.77
X$23410 2462 VIA_via1_4
* cell instance $23411 r0 *1 87.685,91.77
X$23411 2462 VIA_via2_5
* cell instance $23412 r0 *1 89.585,91.63
X$23412 2462 VIA_via1_4
* cell instance $23413 r0 *1 89.585,91.77
X$23413 2462 VIA_via2_5
* cell instance $23414 r0 *1 12.635,92.05
X$23414 2463 VIA_via2_5
* cell instance $23415 r0 *1 13.585,92.05
X$23415 2463 VIA_via2_5
* cell instance $23416 r0 *1 12.635,91.63
X$23416 2463 VIA_via1_4
* cell instance $23417 r0 *1 13.585,93.17
X$23417 2463 VIA_via1_4
* cell instance $23418 r0 *1 13.965,94.15
X$23418 2463 VIA_via1_4
* cell instance $23419 r0 *1 13.015,91.63
X$23419 2464 VIA_via1_4
* cell instance $23420 r0 *1 13.205,91.63
X$23420 2464 VIA_via1_4
* cell instance $23421 r0 *1 17.195,92.61
X$23421 2465 VIA_via1_7
* cell instance $23422 r0 *1 17.195,91.63
X$23422 2465 VIA_via2_5
* cell instance $23423 r0 *1 15.865,91.63
X$23423 2465 VIA_via1_4
* cell instance $23424 r0 *1 15.865,91.63
X$23424 2465 VIA_via2_5
* cell instance $23425 r0 *1 18.525,92.61
X$23425 2466 VIA_via1_7
* cell instance $23426 r0 *1 18.525,90.37
X$23426 2466 VIA_via1_4
* cell instance $23427 r0 *1 29.165,91.63
X$23427 2467 VIA_via1_4
* cell instance $23428 r0 *1 29.165,91.63
X$23428 2467 VIA_via2_5
* cell instance $23429 r0 *1 31.255,91.63
X$23429 2467 VIA_via1_4
* cell instance $23430 r0 *1 31.255,91.63
X$23430 2467 VIA_via2_5
* cell instance $23431 r0 *1 33.535,92.05
X$23431 2468 VIA_via2_5
* cell instance $23432 r0 *1 31.635,92.05
X$23432 2468 VIA_via1_4
* cell instance $23433 r0 *1 31.635,92.05
X$23433 2468 VIA_via2_5
* cell instance $23434 r0 *1 33.535,88.83
X$23434 2468 VIA_via1_4
* cell instance $23435 r0 *1 42.085,92.61
X$23435 2469 VIA_via1_7
* cell instance $23436 r0 *1 42.085,91.77
X$23436 2469 VIA_via2_5
* cell instance $23437 r0 *1 39.995,91.63
X$23437 2469 VIA_via1_4
* cell instance $23438 r0 *1 39.995,91.77
X$23438 2469 VIA_via2_5
* cell instance $23439 r0 *1 51.395,92.05
X$23439 2470 VIA_via2_5
* cell instance $23440 r0 *1 52.155,92.05
X$23440 2470 VIA_via1_4
* cell instance $23441 r0 *1 52.155,92.05
X$23441 2470 VIA_via2_5
* cell instance $23442 r0 *1 51.395,91.63
X$23442 2470 VIA_via1_4
* cell instance $23443 r0 *1 51.585,91.63
X$23443 2471 VIA_via1_4
* cell instance $23444 r0 *1 51.585,91.77
X$23444 2471 VIA_via2_5
* cell instance $23445 r0 *1 53.295,91.77
X$23445 2471 VIA_via1_4
* cell instance $23446 r0 *1 53.295,91.77
X$23446 2471 VIA_via2_5
* cell instance $23447 r0 *1 70.965,92.33
X$23447 2472 VIA_via2_5
* cell instance $23448 r0 *1 71.535,92.33
X$23448 2472 VIA_via2_5
* cell instance $23449 r0 *1 74.005,92.33
X$23449 2472 VIA_via2_5
* cell instance $23450 r0 *1 74.005,93.03
X$23450 2472 VIA_via1_4
* cell instance $23451 r0 *1 70.965,91.63
X$23451 2472 VIA_via1_4
* cell instance $23452 r0 *1 71.535,88.83
X$23452 2472 VIA_via1_4
* cell instance $23453 r0 *1 69.065,91.63
X$23453 2473 VIA_via1_4
* cell instance $23454 r0 *1 69.065,91.63
X$23454 2473 VIA_via2_5
* cell instance $23455 r0 *1 67.355,91.63
X$23455 2473 VIA_via1_4
* cell instance $23456 r0 *1 67.355,91.63
X$23456 2473 VIA_via2_5
* cell instance $23457 r0 *1 8.265,94.43
X$23457 2474 VIA_via2_5
* cell instance $23458 r0 *1 8.455,93.45
X$23458 2474 VIA_via1_4
* cell instance $23459 r0 *1 7.315,94.43
X$23459 2474 VIA_via1_4
* cell instance $23460 r0 *1 7.315,94.43
X$23460 2474 VIA_via2_5
* cell instance $23461 r0 *1 9.215,94.43
X$23461 2474 VIA_via1_4
* cell instance $23462 r0 *1 9.215,94.43
X$23462 2474 VIA_via2_5
* cell instance $23463 r0 *1 16.815,93.17
X$23463 2475 VIA_via1_4
* cell instance $23464 r0 *1 17.575,93.17
X$23464 2475 VIA_via1_4
* cell instance $23465 r0 *1 18.145,92.05
X$23465 2475 VIA_via1_4
* cell instance $23466 r0 *1 49.495,93.17
X$23466 2476 VIA_via1_4
* cell instance $23467 r0 *1 49.495,93.17
X$23467 2476 VIA_via2_5
* cell instance $23468 r0 *1 50.635,93.17
X$23468 2476 VIA_via1_4
* cell instance $23469 r0 *1 50.635,93.17
X$23469 2476 VIA_via2_5
* cell instance $23470 r0 *1 48.545,93.17
X$23470 2476 VIA_via1_4
* cell instance $23471 r0 *1 48.545,93.17
X$23471 2476 VIA_via2_5
* cell instance $23472 r0 *1 54.245,93.59
X$23472 2477 VIA_via1_7
* cell instance $23473 r0 *1 53.675,94.43
X$23473 2477 VIA_via1_4
* cell instance $23474 r0 *1 71.345,93.45
X$23474 2478 VIA_via2_5
* cell instance $23475 r0 *1 71.915,93.31
X$23475 2478 VIA_via2_5
* cell instance $23476 r0 *1 71.915,91.63
X$23476 2478 VIA_via1_4
* cell instance $23477 r0 *1 70.585,93.17
X$23477 2478 VIA_via1_4
* cell instance $23478 r0 *1 70.585,93.17
X$23478 2478 VIA_via2_5
* cell instance $23479 r0 *1 71.345,94.15
X$23479 2478 VIA_via1_4
* cell instance $23480 r0 *1 70.775,93.17
X$23480 2478 VIA_via1_4
* cell instance $23481 r0 *1 70.775,93.31
X$23481 2478 VIA_via2_5
* cell instance $23482 r0 *1 69.065,93.17
X$23482 2478 VIA_via1_4
* cell instance $23483 r0 *1 69.065,93.17
X$23483 2478 VIA_via2_5
* cell instance $23484 r0 *1 70.585,93.59
X$23484 2479 VIA_via1_7
* cell instance $23485 r0 *1 70.775,94.43
X$23485 2479 VIA_via1_4
* cell instance $23486 r0 *1 71.535,93.59
X$23486 2480 VIA_via1_7
* cell instance $23487 r0 *1 72.295,91.63
X$23487 2480 VIA_via1_4
* cell instance $23488 r0 *1 71.725,94.43
X$23488 2480 VIA_via1_4
* cell instance $23489 r0 *1 72.295,94.43
X$23489 2480 VIA_via1_4
* cell instance $23490 r0 *1 74.385,93.45
X$23490 2481 VIA_via1_4
* cell instance $23491 r0 *1 75.145,95.97
X$23491 2481 VIA_via1_4
* cell instance $23492 r0 *1 73.815,94.43
X$23492 2481 VIA_via1_4
* cell instance $23493 r0 *1 75.715,93.17
X$23493 2482 VIA_via1_7
* cell instance $23494 r0 *1 77.425,93.17
X$23494 2482 VIA_via1_7
* cell instance $23495 r0 *1 71.155,93.59
X$23495 2482 VIA_via2_5
* cell instance $23496 r0 *1 77.425,93.59
X$23496 2482 VIA_via2_5
* cell instance $23497 r0 *1 77.045,93.59
X$23497 2482 VIA_via2_5
* cell instance $23498 r0 *1 75.715,93.59
X$23498 2482 VIA_via2_5
* cell instance $23499 r0 *1 77.045,94.71
X$23499 2482 VIA_via1_4
* cell instance $23500 r0 *1 71.155,94.29
X$23500 2482 VIA_via1_4
* cell instance $23501 r0 *1 84.645,90.79
X$23501 2483 VIA_via1_7
* cell instance $23502 r0 *1 84.075,93.17
X$23502 2483 VIA_via1_4
* cell instance $23503 r0 *1 85.215,93.59
X$23503 2484 VIA_via1_7
* cell instance $23504 r0 *1 84.645,94.43
X$23504 2484 VIA_via1_4
* cell instance $23505 r0 *1 87.495,93.17
X$23505 2485 VIA_via1_4
* cell instance $23506 r0 *1 86.165,93.45
X$23506 2485 VIA_via1_4
* cell instance $23507 r0 *1 88.445,93.59
X$23507 2486 VIA_via1_7
* cell instance $23508 r0 *1 88.255,94.43
X$23508 2486 VIA_via1_4
* cell instance $23509 r0 *1 88.065,93.17
X$23509 2487 VIA_via1_4
* cell instance $23510 r0 *1 88.065,93.17
X$23510 2487 VIA_via2_5
* cell instance $23511 r0 *1 88.825,93.17
X$23511 2487 VIA_via1_4
* cell instance $23512 r0 *1 88.825,93.17
X$23512 2487 VIA_via2_5
* cell instance $23513 r0 *1 13.965,93.59
X$23513 2488 VIA_via1_7
* cell instance $23514 r0 *1 13.965,93.59
X$23514 2488 VIA_via2_5
* cell instance $23515 r0 *1 11.685,93.59
X$23515 2488 VIA_via2_5
* cell instance $23516 r0 *1 11.685,94.43
X$23516 2488 VIA_via1_4
* cell instance $23517 r0 *1 17.765,93.03
X$23517 2489 VIA_via2_5
* cell instance $23518 r0 *1 15.485,93.17
X$23518 2489 VIA_via1_4
* cell instance $23519 r0 *1 15.485,93.03
X$23519 2489 VIA_via2_5
* cell instance $23520 r0 *1 18.145,93.17
X$23520 2489 VIA_via1_4
* cell instance $23521 r0 *1 18.145,93.03
X$23521 2489 VIA_via2_5
* cell instance $23522 r0 *1 17.385,94.15
X$23522 2489 VIA_via1_4
* cell instance $23523 r0 *1 27.455,92.19
X$23523 2490 VIA_via1_7
* cell instance $23524 r0 *1 27.455,93.17
X$23524 2490 VIA_via2_5
* cell instance $23525 r0 *1 25.745,93.17
X$23525 2490 VIA_via1_4
* cell instance $23526 r0 *1 25.745,93.17
X$23526 2490 VIA_via2_5
* cell instance $23527 r0 *1 29.355,93.59
X$23527 2491 VIA_via1_7
* cell instance $23528 r0 *1 29.355,93.59
X$23528 2491 VIA_via2_5
* cell instance $23529 r0 *1 25.935,93.59
X$23529 2491 VIA_via2_5
* cell instance $23530 r0 *1 25.935,94.43
X$23530 2491 VIA_via1_4
* cell instance $23531 r0 *1 30.685,93.59
X$23531 2492 VIA_via1_7
* cell instance $23532 r0 *1 30.685,93.73
X$23532 2492 VIA_via2_5
* cell instance $23533 r0 *1 30.115,93.73
X$23533 2492 VIA_via2_5
* cell instance $23534 r0 *1 30.115,94.43
X$23534 2492 VIA_via1_4
* cell instance $23535 r0 *1 78.565,93.45
X$23535 2493 VIA_via1_7
* cell instance $23536 r0 *1 78.565,93.45
X$23536 2493 VIA_via2_5
* cell instance $23537 r0 *1 77.995,93.45
X$23537 2493 VIA_via2_5
* cell instance $23538 r0 *1 78.185,95.97
X$23538 2493 VIA_via1_4
* cell instance $23539 r0 *1 77.805,95.41
X$23539 2494 VIA_via1_7
* cell instance $23540 r0 *1 78.755,93.59
X$23540 2494 VIA_via2_5
* cell instance $23541 r0 *1 77.805,93.59
X$23541 2494 VIA_via2_5
* cell instance $23542 r0 *1 78.755,93.17
X$23542 2494 VIA_via1_4
* cell instance $23543 r0 *1 32.395,94.15
X$23543 2495 VIA_via1_4
* cell instance $23544 r0 *1 30.305,93.17
X$23544 2495 VIA_via1_4
* cell instance $23545 r0 *1 30.305,93.17
X$23545 2495 VIA_via2_5
* cell instance $23546 r0 *1 32.205,93.17
X$23546 2495 VIA_via1_4
* cell instance $23547 r0 *1 32.205,93.17
X$23547 2495 VIA_via2_5
* cell instance $23548 r0 *1 36.385,93.17
X$23548 2496 VIA_via1_4
* cell instance $23549 r0 *1 36.385,93.17
X$23549 2496 VIA_via2_5
* cell instance $23550 r0 *1 39.995,93.17
X$23550 2496 VIA_via1_4
* cell instance $23551 r0 *1 39.995,93.17
X$23551 2496 VIA_via2_5
* cell instance $23552 r0 *1 39.235,93.31
X$23552 2497 VIA_via2_5
* cell instance $23553 r0 *1 39.235,94.43
X$23553 2497 VIA_via1_4
* cell instance $23554 r0 *1 38.665,93.31
X$23554 2497 VIA_via1_4
* cell instance $23555 r0 *1 38.665,93.31
X$23555 2497 VIA_via2_5
* cell instance $23556 r0 *1 39.615,93.17
X$23556 2497 VIA_via1_4
* cell instance $23557 r0 *1 39.615,93.31
X$23557 2497 VIA_via2_5
* cell instance $23558 r0 *1 75.525,93.17
X$23558 2498 VIA_via1_4
* cell instance $23559 r0 *1 75.525,91.91
X$23559 2498 VIA_via1_4
* cell instance $23560 r0 *1 49.875,93.31
X$23560 2499 VIA_via1_4
* cell instance $23561 r0 *1 49.875,93.31
X$23561 2499 VIA_via2_5
* cell instance $23562 r0 *1 46.265,93.17
X$23562 2499 VIA_via1_4
* cell instance $23563 r0 *1 46.265,93.31
X$23563 2499 VIA_via2_5
* cell instance $23564 r0 *1 73.625,92.19
X$23564 2500 VIA_via1_7
* cell instance $23565 r0 *1 73.625,93.21
X$23565 2500 VIA_via1_7
* cell instance $23566 r0 *1 71.725,92.19
X$23566 2501 VIA_via1_7
* cell instance $23567 r0 *1 71.725,93.17
X$23567 2501 VIA_via2_5
* cell instance $23568 r0 *1 71.155,93.17
X$23568 2501 VIA_via1_4
* cell instance $23569 r0 *1 71.155,93.17
X$23569 2501 VIA_via2_5
* cell instance $23570 r0 *1 55.955,93.17
X$23570 2502 VIA_via2_5
* cell instance $23571 r0 *1 55.955,94.15
X$23571 2502 VIA_via1_4
* cell instance $23572 r0 *1 55.955,94.29
X$23572 2502 VIA_via2_5
* cell instance $23573 r0 *1 56.335,94.43
X$23573 2502 VIA_via1_4
* cell instance $23574 r0 *1 56.335,94.29
X$23574 2502 VIA_via2_5
* cell instance $23575 r0 *1 53.865,93.17
X$23575 2502 VIA_via1_4
* cell instance $23576 r0 *1 53.865,93.17
X$23576 2502 VIA_via2_5
* cell instance $23577 r0 *1 70.205,91.35
X$23577 2503 VIA_via1_7
* cell instance $23578 r0 *1 70.205,93.17
X$23578 2503 VIA_via1_4
* cell instance $23579 r0 *1 68.115,91.91
X$23579 2504 VIA_via1_4
* cell instance $23580 r0 *1 68.115,93.17
X$23580 2504 VIA_via1_4
* cell instance $23581 r0 *1 36.195,94.29
X$23581 2505 VIA_via2_5
* cell instance $23582 r0 *1 32.775,94.29
X$23582 2505 VIA_via2_5
* cell instance $23583 r0 *1 33.725,94.43
X$23583 2505 VIA_via1_4
* cell instance $23584 r0 *1 33.725,94.29
X$23584 2505 VIA_via2_5
* cell instance $23585 r0 *1 32.775,93.17
X$23585 2505 VIA_via1_4
* cell instance $23586 r0 *1 36.195,95.55
X$23586 2505 VIA_via1_4
* cell instance $23587 r0 *1 51.015,94.43
X$23587 2506 VIA_via1_4
* cell instance $23588 r0 *1 51.585,95.55
X$23588 2506 VIA_via1_4
* cell instance $23589 r0 *1 51.205,93.17
X$23589 2506 VIA_via1_4
* cell instance $23590 r0 *1 62.985,94.43
X$23590 2507 VIA_via2_5
* cell instance $23591 r0 *1 59.185,94.43
X$23591 2507 VIA_via1_4
* cell instance $23592 r0 *1 59.185,94.43
X$23592 2507 VIA_via2_5
* cell instance $23593 r0 *1 56.905,94.43
X$23593 2507 VIA_via1_4
* cell instance $23594 r0 *1 56.905,94.43
X$23594 2507 VIA_via2_5
* cell instance $23595 r0 *1 62.985,95.55
X$23595 2507 VIA_via1_4
* cell instance $23596 r0 *1 64.885,94.43
X$23596 2508 VIA_via1_4
* cell instance $23597 r0 *1 64.885,94.43
X$23597 2508 VIA_via2_5
* cell instance $23598 r0 *1 65.455,94.43
X$23598 2508 VIA_via1_4
* cell instance $23599 r0 *1 65.455,94.43
X$23599 2508 VIA_via2_5
* cell instance $23600 r0 *1 65.645,93.31
X$23600 2508 VIA_via1_4
* cell instance $23601 r0 *1 66.025,94.43
X$23601 2508 VIA_via1_4
* cell instance $23602 r0 *1 76.665,93.17
X$23602 2509 VIA_via1_4
* cell instance $23603 r0 *1 76.285,94.15
X$23603 2509 VIA_via1_4
* cell instance $23604 r0 *1 77.425,94.85
X$23604 2510 VIA_via1_7
* cell instance $23605 r0 *1 77.425,94.85
X$23605 2510 VIA_via2_5
* cell instance $23606 r0 *1 78.755,94.85
X$23606 2510 VIA_via2_5
* cell instance $23607 r0 *1 80.085,94.85
X$23607 2510 VIA_via2_5
* cell instance $23608 r0 *1 78.375,93.17
X$23608 2510 VIA_via1_4
* cell instance $23609 r0 *1 80.085,95.97
X$23609 2510 VIA_via1_4
* cell instance $23610 r0 *1 7.695,94.01
X$23610 2511 VIA_via1_7
* cell instance $23611 r0 *1 7.695,94.01
X$23611 2511 VIA_via2_5
* cell instance $23612 r0 *1 6.175,94.01
X$23612 2511 VIA_via2_5
* cell instance $23613 r0 *1 6.175,93.17
X$23613 2511 VIA_via1_4
* cell instance $23614 r0 *1 79.135,96.11
X$23614 2512 VIA_via2_5
* cell instance $23615 r0 *1 81.225,94.29
X$23615 2512 VIA_via2_5
* cell instance $23616 r0 *1 79.135,94.43
X$23616 2512 VIA_via1_4
* cell instance $23617 r0 *1 81.035,95.97
X$23617 2512 VIA_via1_4
* cell instance $23618 r0 *1 81.035,96.11
X$23618 2512 VIA_via2_5
* cell instance $23619 r0 *1 83.315,94.29
X$23619 2512 VIA_via1_4
* cell instance $23620 r0 *1 83.315,94.29
X$23620 2512 VIA_via2_5
* cell instance $23621 r0 *1 79.515,95.97
X$23621 2512 VIA_via1_4
* cell instance $23622 r0 *1 79.515,96.11
X$23622 2512 VIA_via2_5
* cell instance $23623 r0 *1 74.955,93.17
X$23623 2513 VIA_via1_4
* cell instance $23624 r0 *1 74.955,94.15
X$23624 2513 VIA_via1_4
* cell instance $23625 r0 *1 38.095,95.41
X$23625 2514 VIA_via1_7
* cell instance $23626 r0 *1 38.095,94.29
X$23626 2514 VIA_via2_5
* cell instance $23627 r0 *1 36.575,94.43
X$23627 2514 VIA_via1_4
* cell instance $23628 r0 *1 36.575,94.29
X$23628 2514 VIA_via2_5
* cell instance $23629 r0 *1 13.395,95.97
X$23629 2515 VIA_via1_4
* cell instance $23630 r0 *1 13.395,95.97
X$23630 2515 VIA_via2_5
* cell instance $23631 r0 *1 14.095,97.23
X$23631 2515 VIA_via4_0
* cell instance $23632 r0 *1 14.095,97.23
X$23632 2515 VIA_via5_0
* cell instance $23633 r0 *1 14.095,95.97
X$23633 2515 VIA_via3_2
* cell instance $23634 r0 *1 14.655,97.23
X$23634 2516 VIA_via5_0
* cell instance $23635 r0 *1 14.725,95.97
X$23635 2516 VIA_via1_4
* cell instance $23636 r0 *1 14.725,95.97
X$23636 2516 VIA_via2_5
* cell instance $23637 r0 *1 14.935,97.23
X$23637 2516 VIA_via4_0
* cell instance $23638 r0 *1 14.935,95.97
X$23638 2516 VIA_via3_2
* cell instance $23639 r0 *1 29.735,95.97
X$23639 2517 VIA_via1_4
* cell instance $23640 r0 *1 29.735,95.97
X$23640 2517 VIA_via2_5
* cell instance $23641 r0 *1 29.775,95.97
X$23641 2517 VIA_via3_2
* cell instance $23642 r0 *1 29.775,97.79
X$23642 2517 VIA_via4_0
* cell instance $23643 r0 *1 29.775,97.79
X$23643 2517 VIA_via5_0
* cell instance $23644 r0 *1 30.685,96.39
X$23644 2518 VIA_via1_7
* cell instance $23645 r0 *1 30.685,96.39
X$23645 2518 VIA_via2_5
* cell instance $23646 r0 *1 31.455,96.39
X$23646 2518 VIA_via5_0
* cell instance $23647 r0 *1 31.455,96.39
X$23647 2518 VIA_via4_0
* cell instance $23648 r0 *1 31.455,96.39
X$23648 2518 VIA_via3_2
* cell instance $23649 r0 *1 31.255,96.39
X$23649 2519 VIA_via1_7
* cell instance $23650 r0 *1 31.255,96.95
X$23650 2519 VIA_via2_5
* cell instance $23651 r0 *1 32.015,96.95
X$23651 2519 VIA_via4_0
* cell instance $23652 r0 *1 32.015,96.95
X$23652 2519 VIA_via3_2
* cell instance $23653 r0 *1 32.015,96.95
X$23653 2519 VIA_via5_0
* cell instance $23654 r0 *1 31.825,96.39
X$23654 2520 VIA_via1_7
* cell instance $23655 r0 *1 31.825,96.39
X$23655 2520 VIA_via2_5
* cell instance $23656 r0 *1 32.575,96.39
X$23656 2520 VIA_via5_0
* cell instance $23657 r0 *1 32.575,96.39
X$23657 2520 VIA_via4_0
* cell instance $23658 r0 *1 32.575,96.39
X$23658 2520 VIA_via3_2
* cell instance $23659 r0 *1 34.105,94.99
X$23659 2521 VIA_via1_7
* cell instance $23660 r0 *1 33.915,95.97
X$23660 2521 VIA_via1_4
* cell instance $23661 r0 *1 39.235,96.39
X$23661 2522 VIA_via1_7
* cell instance $23662 r0 *1 39.235,96.39
X$23662 2522 VIA_via2_5
* cell instance $23663 r0 *1 37.615,96.39
X$23663 2522 VIA_via5_0
* cell instance $23664 r0 *1 39.015,96.39
X$23664 2522 VIA_via3_2
* cell instance $23665 r0 *1 39.015,96.39
X$23665 2522 VIA_via4_0
* cell instance $23666 r0 *1 38.285,95.97
X$23666 2523 VIA_via1_4
* cell instance $23667 r0 *1 38.285,95.97
X$23667 2523 VIA_via2_5
* cell instance $23668 r0 *1 38.175,95.97
X$23668 2523 VIA_via3_2
* cell instance $23669 r0 *1 38.175,97.23
X$23669 2523 VIA_via4_0
* cell instance $23670 r0 *1 38.175,97.23
X$23670 2523 VIA_via5_0
* cell instance $23671 r0 *1 37.715,94.85
X$23671 2524 VIA_via2_5
* cell instance $23672 r0 *1 38.855,94.85
X$23672 2524 VIA_via2_5
* cell instance $23673 r0 *1 39.805,94.85
X$23673 2524 VIA_via2_5
* cell instance $23674 r0 *1 39.805,94.43
X$23674 2524 VIA_via1_4
* cell instance $23675 r0 *1 37.715,95.97
X$23675 2524 VIA_via1_4
* cell instance $23676 r0 *1 38.855,94.43
X$23676 2524 VIA_via1_4
* cell instance $23677 r0 *1 41.535,94.99
X$23677 2525 VIA_via5_0
* cell instance $23678 r0 *1 42.655,94.99
X$23678 2525 VIA_via4_0
* cell instance $23679 r0 *1 42.655,94.99
X$23679 2525 VIA_via3_2
* cell instance $23680 r0 *1 42.655,94.99
X$23680 2525 VIA_via2_5
* cell instance $23681 r0 *1 42.655,94.99
X$23681 2525 VIA_via1_7
* cell instance $23682 r0 *1 46.015,96.39
X$23682 2526 VIA_via5_0
* cell instance $23683 r0 *1 46.015,96.39
X$23683 2526 VIA_via4_0
* cell instance $23684 r0 *1 46.265,94.43
X$23684 2526 VIA_via1_4
* cell instance $23685 r0 *1 46.265,94.43
X$23685 2526 VIA_via2_5
* cell instance $23686 r0 *1 46.015,94.43
X$23686 2526 VIA_via3_2
* cell instance $23687 r0 *1 52.155,96.39
X$23687 2527 VIA_via1_7
* cell instance $23688 r0 *1 52.155,96.39
X$23688 2527 VIA_via2_5
* cell instance $23689 r0 *1 51.615,96.39
X$23689 2527 VIA_via4_0
* cell instance $23690 r0 *1 51.615,96.39
X$23690 2527 VIA_via3_2
* cell instance $23691 r0 *1 51.615,96.39
X$23691 2527 VIA_via5_0
* cell instance $23692 r0 *1 54.055,96.39
X$23692 2528 VIA_via1_7
* cell instance $23693 r0 *1 54.055,96.39
X$23693 2528 VIA_via2_5
* cell instance $23694 r0 *1 52.735,96.39
X$23694 2528 VIA_via4_0
* cell instance $23695 r0 *1 52.735,96.39
X$23695 2528 VIA_via5_0
* cell instance $23696 r0 *1 52.735,96.39
X$23696 2528 VIA_via3_2
* cell instance $23697 r0 *1 54.415,96.39
X$23697 2529 VIA_via5_0
* cell instance $23698 r0 *1 55.535,96.39
X$23698 2529 VIA_via4_0
* cell instance $23699 r0 *1 55.535,96.39
X$23699 2529 VIA_via3_2
* cell instance $23700 r0 *1 55.575,96.39
X$23700 2529 VIA_via2_5
* cell instance $23701 r0 *1 55.575,96.39
X$23701 2529 VIA_via1_7
* cell instance $23702 r0 *1 57.215,96.95
X$23702 2530 VIA_via5_0
* cell instance $23703 r0 *1 57.215,96.95
X$23703 2530 VIA_via4_0
* cell instance $23704 r0 *1 57.095,95.97
X$23704 2530 VIA_via1_4
* cell instance $23705 r0 *1 57.095,95.97
X$23705 2530 VIA_via2_5
* cell instance $23706 r0 *1 57.215,95.97
X$23706 2530 VIA_via3_2
* cell instance $23707 r0 *1 59.565,94.99
X$23707 2531 VIA_via1_7
* cell instance $23708 r0 *1 60.705,95.97
X$23708 2531 VIA_via1_4
* cell instance $23709 r0 *1 58.805,95.97
X$23709 2532 VIA_via1_4
* cell instance $23710 r0 *1 58.805,95.97
X$23710 2532 VIA_via2_5
* cell instance $23711 r0 *1 60.015,97.23
X$23711 2532 VIA_via4_0
* cell instance $23712 r0 *1 60.015,97.23
X$23712 2532 VIA_via5_0
* cell instance $23713 r0 *1 60.015,95.97
X$23713 2532 VIA_via3_2
* cell instance $23714 r0 *1 63.935,97.23
X$23714 2533 VIA_via5_0
* cell instance $23715 r0 *1 63.935,97.23
X$23715 2533 VIA_via4_0
* cell instance $23716 r0 *1 63.935,95.97
X$23716 2533 VIA_via1_4
* cell instance $23717 r0 *1 63.935,95.97
X$23717 2533 VIA_via3_2
* cell instance $23718 r0 *1 63.935,95.97
X$23718 2533 VIA_via2_5
* cell instance $23719 r0 *1 64.695,94.99
X$23719 2534 VIA_via1_7
* cell instance $23720 r0 *1 64.695,94.99
X$23720 2534 VIA_via2_5
* cell instance $23721 r0 *1 64.495,94.99
X$23721 2534 VIA_via4_0
* cell instance $23722 r0 *1 64.495,94.99
X$23722 2534 VIA_via5_0
* cell instance $23723 r0 *1 64.495,94.99
X$23723 2534 VIA_via3_2
* cell instance $23724 r0 *1 65.055,96.39
X$23724 2535 VIA_via5_0
* cell instance $23725 r0 *1 65.335,96.39
X$23725 2535 VIA_via3_2
* cell instance $23726 r0 *1 65.335,96.39
X$23726 2535 VIA_via4_0
* cell instance $23727 r0 *1 65.455,96.39
X$23727 2535 VIA_via2_5
* cell instance $23728 r0 *1 65.455,96.39
X$23728 2535 VIA_via1_7
* cell instance $23729 r0 *1 65.265,94.99
X$23729 2536 VIA_via1_7
* cell instance $23730 r0 *1 65.075,95.97
X$23730 2536 VIA_via1_4
* cell instance $23731 r0 *1 65.835,94.99
X$23731 2537 VIA_via1_7
* cell instance $23732 r0 *1 65.835,94.99
X$23732 2537 VIA_via2_5
* cell instance $23733 r0 *1 65.615,94.99
X$23733 2537 VIA_via4_0
* cell instance $23734 r0 *1 65.615,94.99
X$23734 2537 VIA_via3_2
* cell instance $23735 r0 *1 65.615,94.99
X$23735 2537 VIA_via5_0
* cell instance $23736 r0 *1 66.595,96.39
X$23736 2538 VIA_via1_7
* cell instance $23737 r0 *1 66.595,96.39
X$23737 2538 VIA_via2_5
* cell instance $23738 r0 *1 66.175,96.39
X$23738 2538 VIA_via4_0
* cell instance $23739 r0 *1 66.175,96.39
X$23739 2538 VIA_via3_2
* cell instance $23740 r0 *1 66.175,96.39
X$23740 2538 VIA_via5_0
* cell instance $23741 r0 *1 67.855,98.07
X$23741 2539 VIA_via5_0
* cell instance $23742 r0 *1 67.855,98.07
X$23742 2539 VIA_via4_0
* cell instance $23743 r0 *1 67.925,95.97
X$23743 2539 VIA_via1_4
* cell instance $23744 r0 *1 67.925,95.97
X$23744 2539 VIA_via2_5
* cell instance $23745 r0 *1 67.855,95.97
X$23745 2539 VIA_via3_2
* cell instance $23746 r0 *1 74.955,96.39
X$23746 2540 VIA_via1_7
* cell instance $23747 r0 *1 74.955,96.39
X$23747 2540 VIA_via2_5
* cell instance $23748 r0 *1 75.135,96.39
X$23748 2540 VIA_via3_2
* cell instance $23749 r0 *1 75.135,96.39
X$23749 2540 VIA_via4_0
* cell instance $23750 r0 *1 75.135,96.39
X$23750 2540 VIA_via5_0
* cell instance $23751 r0 *1 75.525,96.39
X$23751 2541 VIA_via1_7
* cell instance $23752 r0 *1 75.525,96.39
X$23752 2541 VIA_via2_5
* cell instance $23753 r0 *1 75.695,96.39
X$23753 2541 VIA_via4_0
* cell instance $23754 r0 *1 75.695,96.39
X$23754 2541 VIA_via3_2
* cell instance $23755 r0 *1 75.695,96.39
X$23755 2541 VIA_via5_0
* cell instance $23756 r0 *1 76.095,96.39
X$23756 2542 VIA_via1_7
* cell instance $23757 r0 *1 76.095,96.39
X$23757 2542 VIA_via2_5
* cell instance $23758 r0 *1 76.255,96.39
X$23758 2542 VIA_via3_2
* cell instance $23759 r0 *1 76.255,96.39
X$23759 2542 VIA_via4_0
* cell instance $23760 r0 *1 76.255,96.39
X$23760 2542 VIA_via5_0
* cell instance $23761 r0 *1 76.665,96.39
X$23761 2543 VIA_via1_7
* cell instance $23762 r0 *1 76.665,96.39
X$23762 2543 VIA_via2_5
* cell instance $23763 r0 *1 76.815,96.39
X$23763 2543 VIA_via4_0
* cell instance $23764 r0 *1 76.815,96.39
X$23764 2543 VIA_via5_0
* cell instance $23765 r0 *1 76.815,96.39
X$23765 2543 VIA_via3_2
* cell instance $23766 r0 *1 77.235,96.39
X$23766 2544 VIA_via1_7
* cell instance $23767 r0 *1 77.235,96.39
X$23767 2544 VIA_via2_5
* cell instance $23768 r0 *1 77.375,96.39
X$23768 2544 VIA_via3_2
* cell instance $23769 r0 *1 77.375,96.39
X$23769 2544 VIA_via4_0
* cell instance $23770 r0 *1 77.375,96.39
X$23770 2544 VIA_via5_0
* cell instance $23771 r0 *1 78.565,96.39
X$23771 2545 VIA_via1_7
* cell instance $23772 r0 *1 78.565,96.39
X$23772 2545 VIA_via2_5
* cell instance $23773 r0 *1 77.935,96.39
X$23773 2545 VIA_via4_0
* cell instance $23774 r0 *1 77.935,96.39
X$23774 2545 VIA_via5_0
* cell instance $23775 r0 *1 77.935,96.39
X$23775 2545 VIA_via3_2
* cell instance $23776 r0 *1 78.565,94.5
X$23776 2546 VIA_via1_4
* cell instance $23777 r0 *1 80.275,95.97
X$23777 2546 VIA_via1_4
* cell instance $23778 r0 *1 80.275,95.97
X$23778 2546 VIA_via2_5
* cell instance $23779 r0 *1 78.755,95.97
X$23779 2546 VIA_via1_4
* cell instance $23780 r0 *1 78.755,95.97
X$23780 2546 VIA_via2_5
* cell instance $23781 r0 *1 79.055,96.39
X$23781 2547 VIA_via5_0
* cell instance $23782 r0 *1 79.055,96.39
X$23782 2547 VIA_via4_0
* cell instance $23783 r0 *1 79.055,96.39
X$23783 2547 VIA_via3_2
* cell instance $23784 r0 *1 79.135,96.39
X$23784 2547 VIA_via2_5
* cell instance $23785 r0 *1 79.135,96.39
X$23785 2547 VIA_via1_7
* cell instance $23786 r0 *1 79.895,96.39
X$23786 2548 VIA_via1_7
* cell instance $23787 r0 *1 79.895,96.39
X$23787 2548 VIA_via2_5
* cell instance $23788 r0 *1 79.895,96.39
X$23788 2548 VIA_via3_2
* cell instance $23789 r0 *1 79.895,96.39
X$23789 2548 VIA_via4_0
* cell instance $23790 r0 *1 79.615,96.39
X$23790 2548 VIA_via5_0
* cell instance $23791 r0 *1 80.085,93.17
X$23791 2549 VIA_via1_4
* cell instance $23792 r0 *1 79.705,94.57
X$23792 2549 VIA_via1_4
* cell instance $23793 r0 *1 80.655,93.17
X$23793 2550 VIA_via1_4
* cell instance $23794 r0 *1 80.845,95.69
X$23794 2550 VIA_via1_4
* cell instance $23795 r0 *1 83.505,96.39
X$23795 2551 VIA_via1_7
* cell instance $23796 r0 *1 83.505,96.39
X$23796 2551 VIA_via2_5
* cell instance $23797 r0 *1 82.975,96.39
X$23797 2551 VIA_via4_0
* cell instance $23798 r0 *1 82.975,96.39
X$23798 2551 VIA_via3_2
* cell instance $23799 r0 *1 82.975,96.39
X$23799 2551 VIA_via5_0
* cell instance $23800 r0 *1 84.075,96.39
X$23800 2552 VIA_via1_7
* cell instance $23801 r0 *1 84.075,96.39
X$23801 2552 VIA_via2_5
* cell instance $23802 r0 *1 83.535,96.39
X$23802 2552 VIA_via5_0
* cell instance $23803 r0 *1 84.375,96.39
X$23803 2552 VIA_via3_2
* cell instance $23804 r0 *1 84.375,96.39
X$23804 2552 VIA_via4_0
* cell instance $23805 r0 *1 84.645,96.39
X$23805 2553 VIA_via1_7
* cell instance $23806 r0 *1 84.645,96.95
X$23806 2553 VIA_via2_5
* cell instance $23807 r0 *1 84.095,96.95
X$23807 2553 VIA_via4_0
* cell instance $23808 r0 *1 84.095,96.95
X$23808 2553 VIA_via3_2
* cell instance $23809 r0 *1 84.095,96.95
X$23809 2553 VIA_via5_0
* cell instance $23810 r0 *1 85.215,96.39
X$23810 2554 VIA_via3_2
* cell instance $23811 r0 *1 85.215,96.39
X$23811 2554 VIA_via4_0
* cell instance $23812 r0 *1 85.215,96.39
X$23812 2554 VIA_via2_5
* cell instance $23813 r0 *1 85.215,96.39
X$23813 2554 VIA_via1_7
* cell instance $23814 r0 *1 85.215,96.39
X$23814 2554 VIA_via5_0
* cell instance $23815 r0 *1 89.015,96.39
X$23815 2555 VIA_via1_7
* cell instance $23816 r0 *1 89.015,96.39
X$23816 2555 VIA_via2_5
* cell instance $23817 r0 *1 89.135,96.39
X$23817 2555 VIA_via3_2
* cell instance $23818 r0 *1 89.135,96.39
X$23818 2555 VIA_via4_0
* cell instance $23819 r0 *1 89.135,96.39
X$23819 2555 VIA_via5_0
* cell instance $23820 r0 *1 91.865,96.39
X$23820 2556 VIA_via1_7
* cell instance $23821 r0 *1 91.865,96.39
X$23821 2556 VIA_via2_5
* cell instance $23822 r0 *1 91.935,96.39
X$23822 2556 VIA_via3_2
* cell instance $23823 r0 *1 91.935,96.39
X$23823 2556 VIA_via4_0
* cell instance $23824 r0 *1 91.935,96.39
X$23824 2556 VIA_via5_0
* cell instance $23825 r0 *1 41.515,94.99
X$23825 2557 VIA_via1_7
* cell instance $23826 r0 *1 41.515,94.99
X$23826 2557 VIA_via2_5
* cell instance $23827 r0 *1 40.755,94.99
X$23827 2557 VIA_via2_5
* cell instance $23828 r0 *1 40.755,95.97
X$23828 2557 VIA_via1_4
* cell instance $23829 r0 *1 43.035,94.43
X$23829 2558 VIA_via2_5
* cell instance $23830 r0 *1 41.135,94.43
X$23830 2558 VIA_via1_4
* cell instance $23831 r0 *1 41.135,94.43
X$23831 2558 VIA_via2_5
* cell instance $23832 r0 *1 43.035,95.55
X$23832 2558 VIA_via1_4
* cell instance $23833 r0 *1 43.035,93.17
X$23833 2558 VIA_via1_4
* cell instance $23834 r0 *1 51.395,94.99
X$23834 2559 VIA_via1_7
* cell instance $23835 r0 *1 51.395,94.99
X$23835 2559 VIA_via2_5
* cell instance $23836 r0 *1 49.305,94.99
X$23836 2559 VIA_via2_5
* cell instance $23837 r0 *1 49.305,95.97
X$23837 2559 VIA_via1_4
* cell instance $23838 r0 *1 81.035,93.59
X$23838 2560 VIA_via1_7
* cell instance $23839 r0 *1 81.035,94.43
X$23839 2560 VIA_via1_4
* cell instance $23840 r0 *1 66.215,94.99
X$23840 2561 VIA_via1_7
* cell instance $23841 r0 *1 66.215,95.97
X$23841 2561 VIA_via1_4
* cell instance $23842 r0 *1 73.245,92.19
X$23842 2562 VIA_via1_7
* cell instance $23843 r0 *1 73.245,94.43
X$23843 2562 VIA_via2_5
* cell instance $23844 r0 *1 70.395,94.43
X$23844 2562 VIA_via1_4
* cell instance $23845 r0 *1 70.395,94.43
X$23845 2562 VIA_via2_5
* cell instance $23846 r0 *1 78.945,94.99
X$23846 2563 VIA_via1_7
* cell instance $23847 r0 *1 78.945,94.99
X$23847 2563 VIA_via2_5
* cell instance $23848 r0 *1 76.855,94.99
X$23848 2563 VIA_via2_5
* cell instance $23849 r0 *1 76.855,95.97
X$23849 2563 VIA_via1_4
.ENDS smart_fifo

* cell OR2_X1
* pin A1
* pin A2
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR2_X1 1 2 3 5 6
* net 1 A1
* net 2 A2
* net 3 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 7 1 4 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 7 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 4 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.195 NMOS_VTL
M$4 4 1 3 3 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $5 r0 *1 0.36,0.195 NMOS_VTL
M$5 3 2 4 3 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 4 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OR2_X1

* cell OAI22_X1
* pin B2
* pin B1
* pin A1
* pin A2
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT OAI22_X1 1 2 3 4 6 7 8
* net 1 B2
* net 2 B1
* net 3 A1
* net 4 A2
* net 6 NWELL,VDD
* net 7 PWELL,VSS
* net 8 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 10 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 8 2 10 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.565,0.995 PMOS_VTL
M$3 9 3 8 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.755,0.995 PMOS_VTL
M$4 6 4 9 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.185,0.2975 NMOS_VTL
M$5 7 1 5 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.375,0.2975 NMOS_VTL
M$6 5 2 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.565,0.2975 NMOS_VTL
M$7 8 3 5 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.755,0.2975 NMOS_VTL
M$8 5 4 8 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI22_X1

* cell NOR3_X2
* pin A3
* pin A2
* pin A1
* pin NWELL,VDD
* pin ZN
* pin PWELL,VSS
.SUBCKT NOR3_X2 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 NWELL,VDD
* net 5 ZN
* net 6 PWELL,VSS
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 10 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 9 2 10 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 5 3 9 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 8 3 5 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 7 2 8 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 4 1 7 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.21,0.2975 NMOS_VTL
M$7 5 1 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $8 r0 *1 0.4,0.2975 NMOS_VTL
M$8 6 2 5 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.59,0.2975 NMOS_VTL
M$9 5 3 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.78,0.2975 NMOS_VTL
M$10 6 3 5 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.97,0.2975 NMOS_VTL
M$11 5 2 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 1.16,0.2975 NMOS_VTL
M$12 6 1 5 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NOR3_X2

* cell AND4_X1
* pin A1
* pin A2
* pin A3
* pin A4
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND4_X1 1 2 3 4 6 7 8
* net 1 A1
* net 2 A2
* net 3 A3
* net 4 A4
* net 6 NWELL,VDD
* net 7 PWELL,VSS
* net 8 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 5 1 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 6 2 5 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 5 3 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $4 r0 *1 0.74,1.1525 PMOS_VTL
M$4 5 4 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 8 5 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.17,0.195 NMOS_VTL
M$6 10 1 5 7 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $7 r0 *1 0.36,0.195 NMOS_VTL
M$7 11 2 10 7 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $8 r0 *1 0.55,0.195 NMOS_VTL
M$8 9 3 11 7 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $9 r0 *1 0.74,0.195 NMOS_VTL
M$9 7 4 9 7 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $10 r0 *1 0.93,0.2975 NMOS_VTL
M$10 8 5 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AND4_X1

* cell NAND3_X2
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND3_X2 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 6 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 5 2 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 6 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 5 3 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 6 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 5 1 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.21,0.2975 NMOS_VTL
M$7 10 1 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $8 r0 *1 0.4,0.2975 NMOS_VTL
M$8 9 2 10 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.59,0.2975 NMOS_VTL
M$9 6 3 9 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.78,0.2975 NMOS_VTL
M$10 8 3 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.97,0.2975 NMOS_VTL
M$11 7 2 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 1.16,0.2975 NMOS_VTL
M$12 4 1 7 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND3_X2

* cell INV_X8
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT INV_X8 1 2 3 4
* net 1 A
* net 2 PWELL,VSS
* net 3 NWELL,VDD
* net 4 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 3 3 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 3 1 4 3 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 4 1 3 3 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 3 1 4 3 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 4 1 3 3 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 3 1 4 3 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.31,0.995 PMOS_VTL
M$7 4 1 3 3 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.5,0.995 PMOS_VTL
M$8 3 1 4 3 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 0.17,0.2975 NMOS_VTL
M$9 4 1 2 2 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $10 r0 *1 0.36,0.2975 NMOS_VTL
M$10 2 1 4 2 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.55,0.2975 NMOS_VTL
M$11 4 1 2 2 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 0.74,0.2975 NMOS_VTL
M$12 2 1 4 2 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.93,0.2975 NMOS_VTL
M$13 4 1 2 2 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 1.12,0.2975 NMOS_VTL
M$14 2 1 4 2 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 1.31,0.2975 NMOS_VTL
M$15 4 1 2 2 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 1.5,0.2975 NMOS_VTL
M$16 2 1 4 2 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS INV_X8

* cell OAI21_X1
* pin B2
* pin B1
* pin A
* pin NWELL,VDD
* pin ZN
* pin PWELL,VSS
.SUBCKT OAI21_X1 1 2 3 5 6 7
* net 1 B2
* net 2 B1
* net 3 A
* net 5 NWELL,VDD
* net 6 ZN
* net 7 PWELL,VSS
* device instance $1 r0 *1 0.195,0.995 PMOS_VTL
M$1 8 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.385,0.995 PMOS_VTL
M$2 6 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.575,0.995 PMOS_VTL
M$3 5 3 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.195,0.2975 NMOS_VTL
M$4 6 1 4 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.385,0.2975 NMOS_VTL
M$5 4 2 6 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.575,0.2975 NMOS_VTL
M$6 7 3 4 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI21_X1

* cell XNOR2_X1
* pin A
* pin B
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT XNOR2_X1 1 2 4 5 7
* net 1 A
* net 2 B
* net 4 NWELL,VDD
* net 5 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.18,1.1525 PMOS_VTL
M$1 3 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.37,1.1525 PMOS_VTL
M$2 3 2 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.0338625P AD=0.02205P PS=0.775U
+ PD=0.455U
* device instance $3 r0 *1 0.565,0.995 PMOS_VTL
M$3 7 3 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.0338625P AD=0.0441P PS=0.775U PD=0.77U
* device instance $4 r0 *1 0.755,0.995 PMOS_VTL
M$4 8 1 7 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.945,0.995 PMOS_VTL
M$5 4 2 8 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.18,0.195 NMOS_VTL
M$6 9 1 3 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $7 r0 *1 0.37,0.195 NMOS_VTL
M$7 5 2 9 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0224P PS=0.35U PD=0.56U
* device instance $8 r0 *1 0.565,0.2975 NMOS_VTL
M$8 6 3 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.0224P AD=0.02905P PS=0.56U PD=0.555U
* device instance $9 r0 *1 0.755,0.2975 NMOS_VTL
M$9 7 1 6 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.945,0.2975 NMOS_VTL
M$10 6 2 7 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS XNOR2_X1

* cell AOI21_X1
* pin A
* pin B2
* pin B1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT AOI21_X1 1 2 3 4 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 4 PWELL,VSS
* net 6 ZN
* net 7 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 6 2 5 7 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 5 3 6 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 7 1 5 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.21,0.2975 NMOS_VTL
M$4 8 2 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.4,0.2975 NMOS_VTL
M$5 6 3 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.59,0.2975 NMOS_VTL
M$6 4 1 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI21_X1

* cell XOR2_X2
* pin B
* pin A
* pin NWELL,VDD
* pin Z
* pin PWELL,VSS
.SUBCKT XOR2_X2 1 2 4 5 7
* net 1 B
* net 2 A
* net 4 NWELL,VDD
* net 5 Z
* net 7 PWELL,VSS
* device instance $1 r0 *1 0.2,0.995 PMOS_VTL
M$1 8 2 3 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.39,0.995 PMOS_VTL
M$2 4 1 8 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.58,0.995 PMOS_VTL
M$3 6 3 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.77,0.995 PMOS_VTL
M$4 5 2 6 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.96,0.995 PMOS_VTL
M$5 6 1 5 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.15,0.995 PMOS_VTL
M$6 5 1 6 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.34,0.995 PMOS_VTL
M$7 6 2 5 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.53,0.995 PMOS_VTL
M$8 4 3 6 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 0.2,0.2975 NMOS_VTL
M$9 3 2 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $10 r0 *1 0.39,0.2975 NMOS_VTL
M$10 7 1 3 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.58,0.2975 NMOS_VTL
M$11 5 3 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 0.77,0.2975 NMOS_VTL
M$12 10 2 5 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.96,0.2975 NMOS_VTL
M$13 7 1 10 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 1.15,0.2975 NMOS_VTL
M$14 9 1 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 1.34,0.2975 NMOS_VTL
M$15 5 2 9 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 1.53,0.2975 NMOS_VTL
M$16 7 3 5 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS XOR2_X2

* cell XOR2_X1
* pin A
* pin B
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT XOR2_X1 1 3 4 5 6
* net 1 A
* net 3 B
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 Z
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 8 1 2 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 8 3 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.0338625P AD=0.02205P PS=0.775U
+ PD=0.455U
* device instance $3 r0 *1 0.555,0.995 PMOS_VTL
M$3 7 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0338625P AD=0.0441P PS=0.775U PD=0.77U
* device instance $4 r0 *1 0.745,0.995 PMOS_VTL
M$4 6 1 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.935,0.995 PMOS_VTL
M$5 7 3 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.17,0.195 NMOS_VTL
M$6 2 1 4 4 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $7 r0 *1 0.36,0.195 NMOS_VTL
M$7 4 3 2 4 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0224P PS=0.35U PD=0.56U
* device instance $8 r0 *1 0.555,0.2975 NMOS_VTL
M$8 6 2 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.0224P AD=0.02905P PS=0.56U PD=0.555U
* device instance $9 r0 *1 0.745,0.2975 NMOS_VTL
M$9 9 1 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.935,0.2975 NMOS_VTL
M$10 4 3 9 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS XOR2_X1

* cell NOR2_X4
* pin A2
* pin A1
* pin ZN
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT NOR2_X4 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 ZN
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 9 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 3 2 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 8 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 5 1 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 7 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 3 2 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.35,0.995 PMOS_VTL
M$7 6 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.54,0.995 PMOS_VTL
M$8 5 1 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 0.21,0.2975 NMOS_VTL
M$9 3 1 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $10 r0 *1 0.4,0.2975 NMOS_VTL
M$10 4 2 3 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.59,0.2975 NMOS_VTL
M$11 3 2 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 0.78,0.2975 NMOS_VTL
M$12 4 1 3 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.97,0.2975 NMOS_VTL
M$13 3 1 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 1.16,0.2975 NMOS_VTL
M$14 4 2 3 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 1.35,0.2975 NMOS_VTL
M$15 3 2 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 1.54,0.2975 NMOS_VTL
M$16 4 1 3 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NOR2_X4

* cell OR4_X2
* pin A1
* pin A2
* pin A3
* pin A4
* pin NWELL,VDD
* pin ZN
* pin PWELL,VSS
.SUBCKT OR4_X2 1 2 3 4 6 7 8
* net 1 A1
* net 2 A2
* net 3 A3
* net 4 A4
* net 6 NWELL,VDD
* net 7 ZN
* net 8 PWELL,VSS
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 11 1 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 10 2 11 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 9 3 10 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 6 4 9 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 7 5 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 6 5 7 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.17,0.2975 NMOS_VTL
M$7 5 1 8 8 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $8 r0 *1 0.36,0.2975 NMOS_VTL
M$8 8 2 5 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.55,0.2975 NMOS_VTL
M$9 5 3 8 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.74,0.2975 NMOS_VTL
M$10 8 4 5 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.93,0.2975 NMOS_VTL
M$11 7 5 8 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 1.12,0.2975 NMOS_VTL
M$12 8 5 7 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OR4_X2

* cell MUX2_X2
* pin A
* pin B
* pin S
* pin NWELL,VDD
* pin PWELL,VSS
* pin Z
.SUBCKT MUX2_X2 1 2 3 6 7 8
* net 1 A
* net 2 B
* net 3 S
* net 6 NWELL,VDD
* net 7 PWELL,VSS
* net 8 Z
* device instance $1 r0 *1 1.16,0.995 PMOS_VTL
M$1 8 4 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 1.35,0.995 PMOS_VTL
M$2 6 4 8 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.033075P PS=0.77U PD=0.77U
* device instance $3 r0 *1 1.54,1.1525 PMOS_VTL
M$3 9 3 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.033075P PS=0.77U
+ PD=0.84U
* device instance $4 r0 *1 0.215,0.995 PMOS_VTL
M$4 6 1 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $5 r0 *1 0.405,0.995 PMOS_VTL
M$5 5 9 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 0.595,0.995 PMOS_VTL
M$6 4 2 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.045675P PS=0.77U PD=0.775U
* device instance $7 r0 *1 0.79,0.995 PMOS_VTL
M$7 5 3 4 6 PMOS_VTL L=0.05U W=0.63U AS=0.045675P AD=0.0693P PS=0.775U PD=1.48U
* device instance $8 r0 *1 1.54,0.195 NMOS_VTL
M$8 9 3 7 7 NMOS_VTL L=0.05U W=0.21U AS=0.021875P AD=0.02205P PS=0.555U PD=0.63U
* device instance $9 r0 *1 1.16,0.2975 NMOS_VTL
M$9 8 4 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $10 r0 *1 1.35,0.2975 NMOS_VTL
M$10 7 4 8 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.021875P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.215,0.2975 NMOS_VTL
M$11 11 1 4 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $12 r0 *1 0.405,0.2975 NMOS_VTL
M$12 7 9 11 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.595,0.2975 NMOS_VTL
M$13 10 2 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.0300875P PS=0.555U
+ PD=0.56U
* device instance $14 r0 *1 0.79,0.2975 NMOS_VTL
M$14 4 3 10 7 NMOS_VTL L=0.05U W=0.415U AS=0.0300875P AD=0.043575P PS=0.56U
+ PD=1.04U
.ENDS MUX2_X2

* cell NOR4_X1
* pin A4
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NOR4_X1 1 2 3 4 5 6 7
* net 1 A4
* net 2 A3
* net 3 A2
* net 4 A1
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 10 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 9 2 10 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 8 3 9 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 4 8 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 7 1 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.36,0.2975 NMOS_VTL
M$6 5 2 7 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.55,0.2975 NMOS_VTL
M$7 7 3 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.74,0.2975 NMOS_VTL
M$8 5 4 7 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NOR4_X1

* cell NOR3_X1
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NOR3_X1 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 8 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 7 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.2975 NMOS_VTL
M$4 6 1 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.36,0.2975 NMOS_VTL
M$5 4 2 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 3 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NOR3_X1

* cell NAND4_X2
* pin A3
* pin A2
* pin A1
* pin A4
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT NAND4_X2 1 2 3 4 5 6 7
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 A4
* net 5 PWELL,VSS
* net 6 ZN
* net 7 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 6 4 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 7 1 6 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 6 2 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 7 3 6 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 6 3 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 7 2 6 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.35,0.995 PMOS_VTL
M$7 6 1 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.54,0.995 PMOS_VTL
M$8 7 4 6 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 0.21,0.2975 NMOS_VTL
M$9 13 4 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $10 r0 *1 0.4,0.2975 NMOS_VTL
M$10 12 1 13 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.59,0.2975 NMOS_VTL
M$11 11 2 12 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 0.78,0.2975 NMOS_VTL
M$12 6 3 11 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.97,0.2975 NMOS_VTL
M$13 8 3 6 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 1.16,0.2975 NMOS_VTL
M$14 10 2 8 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 1.35,0.2975 NMOS_VTL
M$15 9 1 10 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 1.54,0.2975 NMOS_VTL
M$16 5 4 9 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND4_X2

* cell NAND3_X1
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND3_X1 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 6 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.2975 NMOS_VTL
M$4 8 1 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.36,0.2975 NMOS_VTL
M$5 7 2 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 3 7 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND3_X1

* cell AND3_X1
* pin A1
* pin A2
* pin A3
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND3_X1 1 2 3 5 6 7
* net 1 A1
* net 2 A2
* net 3 A3
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 5 1 4 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 4 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 4 3 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 4 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.195 NMOS_VTL
M$5 8 1 4 6 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $6 r0 *1 0.36,0.195 NMOS_VTL
M$6 9 2 8 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $7 r0 *1 0.55,0.195 NMOS_VTL
M$7 6 3 9 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $8 r0 *1 0.74,0.2975 NMOS_VTL
M$8 7 4 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AND3_X1

* cell DFF_X2
* pin PWELL,VSS
* pin D
* pin CK
* pin QN
* pin Q
* pin NWELL,VDD
.SUBCKT DFF_X2 1 6 8 10 11 16
* net 1 PWELL,VSS
* net 6 D
* net 8 CK
* net 10 QN
* net 11 Q
* net 16 NWELL,VDD
* device instance $1 r0 *1 2.855,0.995 PMOS_VTL
M$1 10 9 16 16 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 3.045,0.995 PMOS_VTL
M$2 16 9 10 16 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 3.235,0.995 PMOS_VTL
M$3 11 2 16 16 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 3.425,0.995 PMOS_VTL
M$4 16 2 11 16 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.2,0.9275 PMOS_VTL
M$5 16 7 3 16 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.014175P PS=0.84U
+ PD=0.455U
* device instance $6 r0 *1 0.39,1.04 PMOS_VTL
M$6 17 4 16 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.0063P PS=0.455U
+ PD=0.23U
* device instance $7 r0 *1 0.58,1.04 PMOS_VTL
M$7 17 7 5 16 PMOS_VTL L=0.05U W=0.09U AS=0.01785P AD=0.0063P PS=0.56U PD=0.23U
* device instance $8 r0 *1 0.77,0.975 PMOS_VTL
M$8 18 3 5 16 PMOS_VTL L=0.05U W=0.42U AS=0.01785P AD=0.0294P PS=0.56U PD=0.56U
* device instance $9 r0 *1 0.96,0.975 PMOS_VTL
M$9 16 6 18 16 PMOS_VTL L=0.05U W=0.42U AS=0.0294P AD=0.025725P PS=0.56U
+ PD=0.56U
* device instance $10 r0 *1 1.15,1.0275 PMOS_VTL
M$10 4 5 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.025725P AD=0.0567P PS=0.56U
+ PD=0.99U
* device instance $11 r0 *1 2.135,0.915 PMOS_VTL
M$11 20 3 9 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.0063P PS=0.455U
+ PD=0.23U
* device instance $12 r0 *1 2.325,0.915 PMOS_VTL
M$12 20 2 16 16 PMOS_VTL L=0.05U W=0.09U AS=0.0252P AD=0.0063P PS=0.77U PD=0.23U
* device instance $13 r0 *1 1.565,1.0275 PMOS_VTL
M$13 16 8 7 16 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $14 r0 *1 1.755,1.0275 PMOS_VTL
M$14 19 5 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $15 r0 *1 1.945,1.0275 PMOS_VTL
M$15 9 7 19 16 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.014175P PS=0.455U
+ PD=0.455U
* device instance $16 r0 *1 2.515,0.995 PMOS_VTL
M$16 2 9 16 16 PMOS_VTL L=0.05U W=0.63U AS=0.0252P AD=0.06615P PS=0.77U PD=1.47U
* device instance $17 r0 *1 2.855,0.2975 NMOS_VTL
M$17 10 9 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $18 r0 *1 3.045,0.2975 NMOS_VTL
M$18 1 9 10 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 3.235,0.2975 NMOS_VTL
M$19 11 2 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $20 r0 *1 3.425,0.2975 NMOS_VTL
M$20 1 2 11 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
* device instance $21 r0 *1 0.39,0.31 NMOS_VTL
M$21 12 4 1 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.0063P PS=0.35U PD=0.23U
* device instance $22 r0 *1 0.58,0.31 NMOS_VTL
M$22 12 3 5 1 NMOS_VTL L=0.05U W=0.09U AS=0.012775P AD=0.0063P PS=0.415U
+ PD=0.23U
* device instance $23 r0 *1 1.15,0.25 NMOS_VTL
M$23 4 5 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.016975P AD=0.02205P PS=0.415U
+ PD=0.63U
* device instance $24 r0 *1 0.77,0.2825 NMOS_VTL
M$24 13 7 5 1 NMOS_VTL L=0.05U W=0.275U AS=0.012775P AD=0.01925P PS=0.415U
+ PD=0.415U
* device instance $25 r0 *1 0.96,0.2825 NMOS_VTL
M$25 1 6 13 1 NMOS_VTL L=0.05U W=0.275U AS=0.01925P AD=0.016975P PS=0.415U
+ PD=0.415U
* device instance $26 r0 *1 0.2,0.37 NMOS_VTL
M$26 1 7 3 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0105P PS=0.63U PD=0.35U
* device instance $27 r0 *1 1.565,0.35 NMOS_VTL
M$27 1 8 7 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $28 r0 *1 1.755,0.35 NMOS_VTL
M$28 14 5 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $29 r0 *1 1.945,0.35 NMOS_VTL
M$29 9 3 14 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0105P PS=0.35U PD=0.35U
* device instance $30 r0 *1 2.135,0.41 NMOS_VTL
M$30 15 7 9 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.0063P PS=0.35U PD=0.23U
* device instance $31 r0 *1 2.325,0.41 NMOS_VTL
M$31 15 2 1 1 NMOS_VTL L=0.05U W=0.09U AS=0.017675P AD=0.0063P PS=0.555U
+ PD=0.23U
* device instance $32 r0 *1 2.515,0.2975 NMOS_VTL
M$32 2 9 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.017675P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS DFF_X2

* cell HA_X1
* pin A
* pin B
* pin S
* pin NWELL,VDD
* pin PWELL,VSS
* pin CO
.SUBCKT HA_X1 1 2 4 5 6 9
* net 1 A
* net 2 B
* net 4 S
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 9 CO
* device instance $1 r0 *1 0.785,1.0275 PMOS_VTL
M$1 10 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.0338625P AD=0.02205P PS=0.775U
+ PD=0.455U
* device instance $2 r0 *1 0.975,1.0275 PMOS_VTL
M$2 7 1 10 5 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.033075P PS=0.455U
+ PD=0.84U
* device instance $3 r0 *1 0.21,0.995 PMOS_VTL
M$3 4 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $4 r0 *1 0.4,0.995 PMOS_VTL
M$4 3 1 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.59,0.995 PMOS_VTL
M$5 5 7 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0338625P PS=0.77U PD=0.775U
* device instance $6 r0 *1 1.345,1.0275 PMOS_VTL
M$6 8 1 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $7 r0 *1 1.535,1.0275 PMOS_VTL
M$7 8 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $8 r0 *1 1.725,0.995 PMOS_VTL
M$8 9 8 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 1.345,0.195 NMOS_VTL
M$9 12 1 8 6 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $10 r0 *1 1.535,0.195 NMOS_VTL
M$10 6 2 12 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
* device instance $11 r0 *1 1.725,0.2975 NMOS_VTL
M$11 9 8 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
* device instance $12 r0 *1 0.785,0.195 NMOS_VTL
M$12 7 2 6 6 NMOS_VTL L=0.05U W=0.21U AS=0.0224P AD=0.0147P PS=0.56U PD=0.35U
* device instance $13 r0 *1 0.975,0.195 NMOS_VTL
M$13 6 1 7 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.02205P PS=0.35U PD=0.63U
* device instance $14 r0 *1 0.21,0.2975 NMOS_VTL
M$14 11 2 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $15 r0 *1 0.4,0.2975 NMOS_VTL
M$15 4 1 11 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 0.59,0.2975 NMOS_VTL
M$16 6 7 4 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.0224P PS=0.555U PD=0.56U
.ENDS HA_X1

* cell FA_X1
* pin PWELL,VSS
* pin B
* pin CO
* pin S
* pin CI
* pin A
* pin NWELL,VDD
.SUBCKT FA_X1 1 2 3 8 11 12 14
* net 1 PWELL,VSS
* net 2 B
* net 3 CO
* net 8 S
* net 11 CI
* net 12 A
* net 14 NWELL,VDD
* device instance $1 r0 *1 0.385,1.0275 PMOS_VTL
M$1 17 2 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $2 r0 *1 0.575,1.0275 PMOS_VTL
M$2 4 12 17 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.765,1.0275 PMOS_VTL
M$3 15 11 4 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02265P PS=0.455U
+ PD=0.535U
* device instance $4 r0 *1 0.96,1.1025 PMOS_VTL
M$4 14 12 15 14 PMOS_VTL L=0.05U W=0.315U AS=0.02265P AD=0.02205P PS=0.535U
+ PD=0.455U
* device instance $5 r0 *1 1.15,1.1025 PMOS_VTL
M$5 15 2 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.033075P PS=0.455U
+ PD=0.84U
* device instance $6 r0 *1 0.195,0.995 PMOS_VTL
M$6 14 4 3 14 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.033075P PS=1.47U
+ PD=0.77U
* device instance $7 r0 *1 1.49,1.1525 PMOS_VTL
M$7 16 2 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $8 r0 *1 1.68,1.1525 PMOS_VTL
M$8 14 11 16 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $9 r0 *1 1.87,1.1525 PMOS_VTL
M$9 16 12 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $10 r0 *1 2.06,1.1525 PMOS_VTL
M$10 7 4 16 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.023625P PS=0.455U
+ PD=0.465U
* device instance $11 r0 *1 2.26,1.1525 PMOS_VTL
M$11 18 11 7 14 PMOS_VTL L=0.05U W=0.315U AS=0.023625P AD=0.02205P PS=0.465U
+ PD=0.455U
* device instance $12 r0 *1 2.45,1.1525 PMOS_VTL
M$12 19 2 18 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $13 r0 *1 2.64,1.1525 PMOS_VTL
M$13 19 12 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $14 r0 *1 2.83,0.995 PMOS_VTL
M$14 8 7 14 14 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U
+ PD=1.47U
* device instance $15 r0 *1 0.385,0.32 NMOS_VTL
M$15 13 2 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.021875P AD=0.0147P PS=0.555U
+ PD=0.35U
* device instance $16 r0 *1 0.575,0.32 NMOS_VTL
M$16 4 12 13 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $17 r0 *1 0.765,0.32 NMOS_VTL
M$17 5 11 4 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.015225P PS=0.35U
+ PD=0.355U
* device instance $18 r0 *1 0.96,0.32 NMOS_VTL
M$18 1 12 5 1 NMOS_VTL L=0.05U W=0.21U AS=0.015225P AD=0.0147P PS=0.355U
+ PD=0.35U
* device instance $19 r0 *1 1.15,0.32 NMOS_VTL
M$19 5 2 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.02205P PS=0.35U PD=0.63U
* device instance $20 r0 *1 0.195,0.2975 NMOS_VTL
M$20 1 4 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.021875P PS=1.04U
+ PD=0.555U
* device instance $21 r0 *1 1.49,0.195 NMOS_VTL
M$21 6 2 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $22 r0 *1 1.68,0.195 NMOS_VTL
M$22 1 11 6 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $23 r0 *1 1.87,0.195 NMOS_VTL
M$23 6 12 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $24 r0 *1 2.06,0.195 NMOS_VTL
M$24 7 4 6 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.01575P PS=0.35U PD=0.36U
* device instance $25 r0 *1 2.26,0.195 NMOS_VTL
M$25 9 11 7 1 NMOS_VTL L=0.05U W=0.21U AS=0.01575P AD=0.0147P PS=0.36U PD=0.35U
* device instance $26 r0 *1 2.45,0.195 NMOS_VTL
M$26 10 2 9 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $27 r0 *1 2.64,0.195 NMOS_VTL
M$27 1 12 10 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
* device instance $28 r0 *1 2.83,0.2975 NMOS_VTL
M$28 8 7 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS FA_X1

* cell BUF_X8
* pin PWELL,VSS
* pin Z
* pin NWELL,VDD
* pin A
.SUBCKT BUF_X8 1 3 4 5
* net 1 PWELL,VSS
* net 3 Z
* net 4 NWELL,VDD
* net 5 A
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 2 5 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 4 5 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 2 5 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 4 5 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 3 2 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 4 2 3 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.31,0.995 PMOS_VTL
M$7 3 2 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.5,0.995 PMOS_VTL
M$8 4 2 3 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $9 r0 *1 1.69,0.995 PMOS_VTL
M$9 3 2 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $10 r0 *1 1.88,0.995 PMOS_VTL
M$10 4 2 3 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $11 r0 *1 2.07,0.995 PMOS_VTL
M$11 3 2 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $12 r0 *1 2.26,0.995 PMOS_VTL
M$12 4 2 3 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $13 r0 *1 0.17,0.2975 NMOS_VTL
M$13 2 5 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $14 r0 *1 0.36,0.2975 NMOS_VTL
M$14 1 5 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 0.55,0.2975 NMOS_VTL
M$15 2 5 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 0.74,0.2975 NMOS_VTL
M$16 1 5 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $17 r0 *1 0.93,0.2975 NMOS_VTL
M$17 3 2 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $18 r0 *1 1.12,0.2975 NMOS_VTL
M$18 1 2 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 1.31,0.2975 NMOS_VTL
M$19 3 2 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $20 r0 *1 1.5,0.2975 NMOS_VTL
M$20 1 2 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $21 r0 *1 1.69,0.2975 NMOS_VTL
M$21 3 2 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $22 r0 *1 1.88,0.2975 NMOS_VTL
M$22 1 2 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $23 r0 *1 2.07,0.2975 NMOS_VTL
M$23 3 2 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $24 r0 *1 2.26,0.2975 NMOS_VTL
M$24 1 2 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS BUF_X8

* cell NAND4_X1
* pin A4
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND4_X1 1 2 3 4 5 6 7
* net 1 A4
* net 2 A3
* net 3 A2
* net 4 A1
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 6 2 7 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 7 3 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 6 4 7 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 10 1 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.36,0.2975 NMOS_VTL
M$6 9 2 10 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.55,0.2975 NMOS_VTL
M$7 8 3 9 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.74,0.2975 NMOS_VTL
M$8 7 4 8 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND4_X1

* cell AND2_X1
* pin A1
* pin A2
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND2_X1 1 2 4 5 6
* net 1 A1
* net 2 A2
* net 4 NWELL,VDD
* net 5 PWELL,VSS
* net 6 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 3 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 3 2 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.195 NMOS_VTL
M$4 7 1 3 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $5 r0 *1 0.36,0.195 NMOS_VTL
M$5 5 2 7 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 3 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AND2_X1

* cell INV_X1
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT INV_X1 1 2 3 4
* net 1 A
* net 2 PWELL,VSS
* net 3 NWELL,VDD
* net 4 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 3 3 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.06615P PS=1.47U PD=1.47U
* device instance $2 r0 *1 0.17,0.2975 NMOS_VTL
M$2 4 1 2 2 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.043575P PS=1.04U
+ PD=1.04U
.ENDS INV_X1

* cell BUF_X16
* pin PWELL,VSS
* pin A
* pin Z
* pin NWELL,VDD
.SUBCKT BUF_X16 1 2 4 5
* net 1 PWELL,VSS
* net 2 A
* net 4 Z
* net 5 NWELL,VDD
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 3 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 5 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.565,0.995 PMOS_VTL
M$3 3 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.755,0.995 PMOS_VTL
M$4 5 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.945,0.995 PMOS_VTL
M$5 3 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.135,0.995 PMOS_VTL
M$6 5 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.325,0.995 PMOS_VTL
M$7 3 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.515,0.995 PMOS_VTL
M$8 5 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $9 r0 *1 1.705,0.995 PMOS_VTL
M$9 4 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $10 r0 *1 1.895,0.995 PMOS_VTL
M$10 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $11 r0 *1 2.085,0.995 PMOS_VTL
M$11 4 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $12 r0 *1 2.275,0.995 PMOS_VTL
M$12 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $13 r0 *1 2.465,0.995 PMOS_VTL
M$13 4 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $14 r0 *1 2.655,0.995 PMOS_VTL
M$14 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $15 r0 *1 2.845,0.995 PMOS_VTL
M$15 4 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $16 r0 *1 3.035,0.995 PMOS_VTL
M$16 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $17 r0 *1 3.225,0.995 PMOS_VTL
M$17 4 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $18 r0 *1 3.415,0.995 PMOS_VTL
M$18 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $19 r0 *1 3.605,0.995 PMOS_VTL
M$19 4 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $20 r0 *1 3.795,0.995 PMOS_VTL
M$20 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $21 r0 *1 3.985,0.995 PMOS_VTL
M$21 4 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $22 r0 *1 4.175,0.995 PMOS_VTL
M$22 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $23 r0 *1 4.365,0.995 PMOS_VTL
M$23 4 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $24 r0 *1 4.555,0.995 PMOS_VTL
M$24 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $25 r0 *1 0.185,0.2975 NMOS_VTL
M$25 3 2 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $26 r0 *1 0.375,0.2975 NMOS_VTL
M$26 1 2 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $27 r0 *1 0.565,0.2975 NMOS_VTL
M$27 3 2 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $28 r0 *1 0.755,0.2975 NMOS_VTL
M$28 1 2 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $29 r0 *1 0.945,0.2975 NMOS_VTL
M$29 3 2 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $30 r0 *1 1.135,0.2975 NMOS_VTL
M$30 1 2 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $31 r0 *1 1.325,0.2975 NMOS_VTL
M$31 3 2 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $32 r0 *1 1.515,0.2975 NMOS_VTL
M$32 1 2 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $33 r0 *1 1.705,0.2975 NMOS_VTL
M$33 4 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $34 r0 *1 1.895,0.2975 NMOS_VTL
M$34 1 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $35 r0 *1 2.085,0.2975 NMOS_VTL
M$35 4 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $36 r0 *1 2.275,0.2975 NMOS_VTL
M$36 1 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $37 r0 *1 2.465,0.2975 NMOS_VTL
M$37 4 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $38 r0 *1 2.655,0.2975 NMOS_VTL
M$38 1 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $39 r0 *1 2.845,0.2975 NMOS_VTL
M$39 4 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $40 r0 *1 3.035,0.2975 NMOS_VTL
M$40 1 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $41 r0 *1 3.225,0.2975 NMOS_VTL
M$41 4 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $42 r0 *1 3.415,0.2975 NMOS_VTL
M$42 1 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $43 r0 *1 3.605,0.2975 NMOS_VTL
M$43 4 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $44 r0 *1 3.795,0.2975 NMOS_VTL
M$44 1 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $45 r0 *1 3.985,0.2975 NMOS_VTL
M$45 4 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $46 r0 *1 4.175,0.2975 NMOS_VTL
M$46 1 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $47 r0 *1 4.365,0.2975 NMOS_VTL
M$47 4 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $48 r0 *1 4.555,0.2975 NMOS_VTL
M$48 1 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS BUF_X16

* cell CLKBUF_X1
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT CLKBUF_X1 1 3 4
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.19,1.1525 PMOS_VTL
M$1 2 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.033075P PS=0.77U
+ PD=0.84U
* device instance $2 r0 *1 0.38,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.19,0.2075 NMOS_VTL
M$3 3 1 2 3 NMOS_VTL L=0.05U W=0.095U AS=0.009975P AD=0.01015P PS=0.4U PD=0.335U
* device instance $4 r0 *1 0.38,0.2575 NMOS_VTL
M$4 5 2 3 3 NMOS_VTL L=0.05U W=0.195U AS=0.01015P AD=0.020475P PS=0.335U PD=0.6U
.ENDS CLKBUF_X1

* cell DFF_X1
* pin PWELL,VSS
* pin QN
* pin Q
* pin D
* pin CK
* pin NWELL,VDD
.SUBCKT DFF_X1 1 8 9 14 15 16
* net 1 PWELL,VSS
* net 8 QN
* net 9 Q
* net 14 D
* net 15 CK
* net 16 NWELL,VDD
* device instance $1 r0 *1 2.85,0.995 PMOS_VTL
M$1 16 6 8 16 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 3.04,0.995 PMOS_VTL
M$2 9 7 16 16 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.185,0.9425 PMOS_VTL
M$3 16 5 2 16 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.014175P PS=0.84U
+ PD=0.455U
* device instance $4 r0 *1 0.375,1.055 PMOS_VTL
M$4 17 3 16 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.0063P PS=0.455U
+ PD=0.23U
* device instance $5 r0 *1 0.565,1.055 PMOS_VTL
M$5 17 5 4 16 PMOS_VTL L=0.05U W=0.09U AS=0.018075P AD=0.0063P PS=0.565U
+ PD=0.23U
* device instance $6 r0 *1 0.76,0.975 PMOS_VTL
M$6 18 2 4 16 PMOS_VTL L=0.05U W=0.42U AS=0.018075P AD=0.0294P PS=0.565U
+ PD=0.56U
* device instance $7 r0 *1 0.95,0.975 PMOS_VTL
M$7 16 14 18 16 PMOS_VTL L=0.05U W=0.42U AS=0.0294P AD=0.025725P PS=0.56U
+ PD=0.56U
* device instance $8 r0 *1 1.14,1.0275 PMOS_VTL
M$8 3 4 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.025725P AD=0.0567P PS=0.56U
+ PD=0.99U
* device instance $9 r0 *1 1.555,1.0275 PMOS_VTL
M$9 16 15 5 16 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $10 r0 *1 1.745,1.0275 PMOS_VTL
M$10 19 4 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $11 r0 *1 1.935,1.0275 PMOS_VTL
M$11 6 5 19 16 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.014175P PS=0.455U
+ PD=0.455U
* device instance $12 r0 *1 2.125,1.14 PMOS_VTL
M$12 20 2 6 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.006525P PS=0.455U
+ PD=0.235U
* device instance $13 r0 *1 2.32,1.14 PMOS_VTL
M$13 20 7 16 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.006525P PS=0.455U
+ PD=0.235U
* device instance $14 r0 *1 2.51,1.0275 PMOS_VTL
M$14 7 6 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.014175P AD=0.033075P PS=0.455U
+ PD=0.84U
* device instance $15 r0 *1 2.85,0.2975 NMOS_VTL
M$15 1 6 8 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $16 r0 *1 3.04,0.2975 NMOS_VTL
M$16 9 7 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
* device instance $17 r0 *1 2.125,0.345 NMOS_VTL
M$17 12 5 6 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.006525P PS=0.35U
+ PD=0.235U
* device instance $18 r0 *1 2.32,0.345 NMOS_VTL
M$18 12 7 1 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.006525P PS=0.35U
+ PD=0.235U
* device instance $19 r0 *1 1.555,0.36 NMOS_VTL
M$19 1 15 5 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $20 r0 *1 1.745,0.36 NMOS_VTL
M$20 13 4 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $21 r0 *1 1.935,0.36 NMOS_VTL
M$21 6 2 13 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0105P PS=0.35U PD=0.35U
* device instance $22 r0 *1 2.51,0.36 NMOS_VTL
M$22 7 6 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0105P AD=0.02205P PS=0.35U PD=0.63U
* device instance $23 r0 *1 0.185,0.285 NMOS_VTL
M$23 1 5 2 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0105P PS=0.63U PD=0.35U
* device instance $24 r0 *1 0.375,0.345 NMOS_VTL
M$24 10 3 1 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.0063P PS=0.35U PD=0.23U
* device instance $25 r0 *1 0.565,0.345 NMOS_VTL
M$25 10 2 4 1 NMOS_VTL L=0.05U W=0.09U AS=0.013P AD=0.0063P PS=0.42U PD=0.23U
* device instance $26 r0 *1 1.14,0.285 NMOS_VTL
M$26 3 4 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.016975P AD=0.02205P PS=0.415U
+ PD=0.63U
* device instance $27 r0 *1 0.76,0.3175 NMOS_VTL
M$27 11 5 4 1 NMOS_VTL L=0.05U W=0.275U AS=0.013P AD=0.01925P PS=0.42U PD=0.415U
* device instance $28 r0 *1 0.95,0.3175 NMOS_VTL
M$28 1 14 11 1 NMOS_VTL L=0.05U W=0.275U AS=0.01925P AD=0.016975P PS=0.415U
+ PD=0.415U
.ENDS DFF_X1

* cell OAI22_X4
* pin PWELL,VSS
* pin B2
* pin B1
* pin A2
* pin ZN
* pin A1
* pin NWELL,VDD
.SUBCKT OAI22_X4 1 3 4 5 6 7 8
* net 1 PWELL,VSS
* net 3 B2
* net 4 B1
* net 5 A2
* net 6 ZN
* net 7 A1
* net 8 NWELL,VDD
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 9 3 8 8 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 6 4 9 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 11 4 6 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 8 3 11 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 10 3 8 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 6 4 10 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.31,0.995 PMOS_VTL
M$7 12 4 6 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.5,0.995 PMOS_VTL
M$8 8 3 12 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $9 r0 *1 1.69,0.995 PMOS_VTL
M$9 13 5 8 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $10 r0 *1 1.88,0.995 PMOS_VTL
M$10 6 7 13 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $11 r0 *1 2.07,0.995 PMOS_VTL
M$11 14 7 6 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $12 r0 *1 2.26,0.995 PMOS_VTL
M$12 8 5 14 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $13 r0 *1 2.45,0.995 PMOS_VTL
M$13 15 5 8 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $14 r0 *1 2.64,0.995 PMOS_VTL
M$14 6 7 15 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $15 r0 *1 2.83,0.995 PMOS_VTL
M$15 16 7 6 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $16 r0 *1 3.02,0.995 PMOS_VTL
M$16 8 5 16 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $17 r0 *1 0.17,0.2975 NMOS_VTL
M$17 1 3 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $18 r0 *1 0.36,0.2975 NMOS_VTL
M$18 2 4 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 0.55,0.2975 NMOS_VTL
M$19 1 4 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $20 r0 *1 0.74,0.2975 NMOS_VTL
M$20 2 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $21 r0 *1 0.93,0.2975 NMOS_VTL
M$21 1 3 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $22 r0 *1 1.12,0.2975 NMOS_VTL
M$22 2 4 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $23 r0 *1 1.31,0.2975 NMOS_VTL
M$23 1 4 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $24 r0 *1 1.5,0.2975 NMOS_VTL
M$24 2 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $25 r0 *1 1.69,0.2975 NMOS_VTL
M$25 6 5 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $26 r0 *1 1.88,0.2975 NMOS_VTL
M$26 2 7 6 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $27 r0 *1 2.07,0.2975 NMOS_VTL
M$27 6 7 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $28 r0 *1 2.26,0.2975 NMOS_VTL
M$28 2 5 6 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $29 r0 *1 2.45,0.2975 NMOS_VTL
M$29 6 5 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $30 r0 *1 2.64,0.2975 NMOS_VTL
M$30 2 7 6 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $31 r0 *1 2.83,0.2975 NMOS_VTL
M$31 6 7 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $32 r0 *1 3.02,0.2975 NMOS_VTL
M$32 2 5 6 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI22_X4

* cell OAI21_X4
* pin A
* pin B2
* pin B1
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT OAI21_X4 1 2 3 5 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 1 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 7 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 5 1 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 11 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 7 3 11 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.31,0.995 PMOS_VTL
M$7 10 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.5,0.995 PMOS_VTL
M$8 5 2 10 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $9 r0 *1 1.69,0.995 PMOS_VTL
M$9 9 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $10 r0 *1 1.88,0.995 PMOS_VTL
M$10 7 3 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $11 r0 *1 2.07,0.995 PMOS_VTL
M$11 8 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $12 r0 *1 2.26,0.995 PMOS_VTL
M$12 5 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $13 r0 *1 0.17,0.2975 NMOS_VTL
M$13 6 1 4 6 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $14 r0 *1 0.36,0.2975 NMOS_VTL
M$14 4 1 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 0.55,0.2975 NMOS_VTL
M$15 6 1 4 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 0.74,0.2975 NMOS_VTL
M$16 4 1 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $17 r0 *1 0.93,0.2975 NMOS_VTL
M$17 7 2 4 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $18 r0 *1 1.12,0.2975 NMOS_VTL
M$18 4 3 7 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 1.31,0.2975 NMOS_VTL
M$19 7 3 4 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $20 r0 *1 1.5,0.2975 NMOS_VTL
M$20 4 2 7 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $21 r0 *1 1.69,0.2975 NMOS_VTL
M$21 7 2 4 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $22 r0 *1 1.88,0.2975 NMOS_VTL
M$22 4 3 7 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $23 r0 *1 2.07,0.2975 NMOS_VTL
M$23 7 3 4 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $24 r0 *1 2.26,0.2975 NMOS_VTL
M$24 4 2 7 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI21_X4

* cell OAI22_X2
* pin B2
* pin B1
* pin A2
* pin A1
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT OAI22_X2 1 2 3 4 6 7 8
* net 1 B2
* net 2 B1
* net 3 A2
* net 4 A1
* net 6 NWELL,VDD
* net 7 PWELL,VSS
* net 8 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 10 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 8 2 10 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 9 2 8 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 6 1 9 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 12 3 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 8 4 12 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.31,0.995 PMOS_VTL
M$7 11 4 8 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.5,0.995 PMOS_VTL
M$8 6 3 11 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 0.17,0.2975 NMOS_VTL
M$9 7 1 5 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $10 r0 *1 0.36,0.2975 NMOS_VTL
M$10 5 2 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.55,0.2975 NMOS_VTL
M$11 7 2 5 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 0.74,0.2975 NMOS_VTL
M$12 5 1 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.93,0.2975 NMOS_VTL
M$13 8 3 5 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 1.12,0.2975 NMOS_VTL
M$14 5 4 8 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 1.31,0.2975 NMOS_VTL
M$15 8 4 5 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 1.5,0.2975 NMOS_VTL
M$16 5 3 8 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI22_X2

* cell OAI221_X1
* pin B2
* pin B1
* pin A
* pin C2
* pin C1
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT OAI221_X1 1 2 3 4 5 7 8 9
* net 1 B2
* net 2 B1
* net 3 A
* net 4 C2
* net 5 C1
* net 7 NWELL,VDD
* net 8 PWELL,VSS
* net 9 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 12 1 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 9 2 12 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 7 3 9 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 11 4 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 9 5 11 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.17,0.2975 NMOS_VTL
M$6 8 1 6 8 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $7 r0 *1 0.36,0.2975 NMOS_VTL
M$7 6 2 8 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.55,0.2975 NMOS_VTL
M$8 10 3 6 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.74,0.2975 NMOS_VTL
M$9 9 4 10 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.93,0.2975 NMOS_VTL
M$10 10 5 9 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI221_X1

* cell OAI33_X1
* pin B3
* pin B2
* pin B1
* pin A1
* pin A2
* pin A3
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OAI33_X1 1 2 3 4 5 6 7 8 10
* net 1 B3
* net 2 B2
* net 3 B1
* net 4 A1
* net 5 A2
* net 6 A3
* net 7 PWELL,VSS
* net 8 NWELL,VDD
* net 10 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 14 1 8 8 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 13 2 14 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.565,0.995 PMOS_VTL
M$3 10 3 13 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.755,0.995 PMOS_VTL
M$4 12 4 10 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.945,0.995 PMOS_VTL
M$5 11 5 12 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.135,0.995 PMOS_VTL
M$6 8 6 11 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.185,0.2975 NMOS_VTL
M$7 9 1 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $8 r0 *1 0.375,0.2975 NMOS_VTL
M$8 7 2 9 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.565,0.2975 NMOS_VTL
M$9 9 3 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.755,0.2975 NMOS_VTL
M$10 10 4 9 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.945,0.2975 NMOS_VTL
M$11 9 5 10 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 1.135,0.2975 NMOS_VTL
M$12 10 6 9 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI33_X1

* cell NOR2_X1
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NOR2_X1 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 6 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 5 2 6 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.185,0.2975 NMOS_VTL
M$3 5 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $4 r0 *1 0.375,0.2975 NMOS_VTL
M$4 3 2 5 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NOR2_X1

* cell NAND2_X4
* pin A2
* pin A1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT NAND2_X4 1 2 4 5 6
* net 1 A2
* net 2 A1
* net 4 PWELL,VSS
* net 5 ZN
* net 6 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 5 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 6 1 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 5 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 6 1 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 5 2 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 6 2 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.35,0.995 PMOS_VTL
M$7 5 2 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.54,0.995 PMOS_VTL
M$8 6 2 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 0.21,0.2975 NMOS_VTL
M$9 4 1 3 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $10 r0 *1 0.4,0.2975 NMOS_VTL
M$10 3 1 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.59,0.2975 NMOS_VTL
M$11 4 1 3 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 0.78,0.2975 NMOS_VTL
M$12 3 1 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.97,0.2975 NMOS_VTL
M$13 5 2 3 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 1.16,0.2975 NMOS_VTL
M$14 3 2 5 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 1.35,0.2975 NMOS_VTL
M$15 5 2 3 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 1.54,0.2975 NMOS_VTL
M$16 3 2 5 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND2_X4

* cell NAND2_X2
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND2_X2 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.195,0.995 PMOS_VTL
M$1 5 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.385,0.995 PMOS_VTL
M$2 4 2 5 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.575,0.995 PMOS_VTL
M$3 5 2 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.765,0.995 PMOS_VTL
M$4 4 1 5 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.195,0.2975 NMOS_VTL
M$5 7 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.385,0.2975 NMOS_VTL
M$6 5 2 7 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.575,0.2975 NMOS_VTL
M$7 6 2 5 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.765,0.2975 NMOS_VTL
M$8 3 1 6 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND2_X2

* cell MUX2_X1
* pin A
* pin S
* pin B
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT MUX2_X1 1 2 3 5 6 8
* net 1 A
* net 2 S
* net 3 B
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 8 Z
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 6 2 4 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 9 1 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 7 2 9 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $4 r0 *1 0.74,1.1525 PMOS_VTL
M$4 10 4 7 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $5 r0 *1 0.93,1.1525 PMOS_VTL
M$5 10 3 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 8 7 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.17,0.195 NMOS_VTL
M$7 5 2 4 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $8 r0 *1 0.36,0.195 NMOS_VTL
M$8 12 1 5 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $9 r0 *1 0.55,0.195 NMOS_VTL
M$9 7 4 12 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $10 r0 *1 0.74,0.195 NMOS_VTL
M$10 11 2 7 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $11 r0 *1 0.93,0.195 NMOS_VTL
M$11 5 3 11 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
* device instance $12 r0 *1 1.12,0.2975 NMOS_VTL
M$12 8 7 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS MUX2_X1

* cell INV_X2
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT INV_X2 1 2 3 4
* net 1 A
* net 2 PWELL,VSS
* net 3 NWELL,VDD
* net 4 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 4 1 3 3 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 3 1 4 3 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.185,0.2975 NMOS_VTL
M$3 4 1 2 2 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $4 r0 *1 0.375,0.2975 NMOS_VTL
M$4 2 1 4 2 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS INV_X2

* cell BUF_X2
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT BUF_X2 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 4 1 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 4 2 5 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.21,0.2975 NMOS_VTL
M$4 3 1 2 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.4,0.2975 NMOS_VTL
M$5 5 2 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.59,0.2975 NMOS_VTL
M$6 3 2 5 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS BUF_X2

* cell CLKBUF_X2
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT CLKBUF_X2 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 4 2 5 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.1875 NMOS_VTL
M$4 3 1 2 3 NMOS_VTL L=0.05U W=0.195U AS=0.020475P AD=0.01365P PS=0.6U PD=0.335U
* device instance $5 r0 *1 0.36,0.1875 NMOS_VTL
M$5 5 2 3 3 NMOS_VTL L=0.05U W=0.195U AS=0.01365P AD=0.01365P PS=0.335U
+ PD=0.335U
* device instance $6 r0 *1 0.55,0.1875 NMOS_VTL
M$6 3 2 5 3 NMOS_VTL L=0.05U W=0.195U AS=0.01365P AD=0.020475P PS=0.335U PD=0.6U
.ENDS CLKBUF_X2

* cell BUF_X32
* pin PWELL,VSS
* pin A
* pin Z
* pin NWELL,VDD
.SUBCKT BUF_X32 1 2 4 5
* net 1 PWELL,VSS
* net 2 A
* net 4 Z
* net 5 NWELL,VDD
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 3 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 3 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 5 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 3 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 5 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.31,0.995 PMOS_VTL
M$7 3 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.5,0.995 PMOS_VTL
M$8 5 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $9 r0 *1 1.69,0.995 PMOS_VTL
M$9 3 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $10 r0 *1 1.88,0.995 PMOS_VTL
M$10 5 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $11 r0 *1 2.07,0.995 PMOS_VTL
M$11 3 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $12 r0 *1 2.26,0.995 PMOS_VTL
M$12 5 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $13 r0 *1 2.45,0.995 PMOS_VTL
M$13 3 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $14 r0 *1 2.64,0.995 PMOS_VTL
M$14 5 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $15 r0 *1 2.83,0.995 PMOS_VTL
M$15 3 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.045675P PS=0.77U PD=0.775U
* device instance $16 r0 *1 3.025,0.995 PMOS_VTL
M$16 5 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.045675P AD=0.0441P PS=0.775U PD=0.77U
* device instance $17 r0 *1 3.215,0.995 PMOS_VTL
M$17 4 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0504P PS=0.77U PD=0.79U
* device instance $18 r0 *1 3.425,0.995 PMOS_VTL
M$18 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0504P AD=0.0441P PS=0.79U PD=0.77U
* device instance $19 r0 *1 3.615,0.995 PMOS_VTL
M$19 4 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $20 r0 *1 3.805,0.995 PMOS_VTL
M$20 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $21 r0 *1 3.995,0.995 PMOS_VTL
M$21 4 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $22 r0 *1 4.185,0.995 PMOS_VTL
M$22 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $23 r0 *1 4.375,0.995 PMOS_VTL
M$23 4 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $24 r0 *1 4.565,0.995 PMOS_VTL
M$24 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $25 r0 *1 4.755,0.995 PMOS_VTL
M$25 4 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $26 r0 *1 4.945,0.995 PMOS_VTL
M$26 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $27 r0 *1 5.135,0.995 PMOS_VTL
M$27 4 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $28 r0 *1 5.325,0.995 PMOS_VTL
M$28 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $29 r0 *1 5.515,0.995 PMOS_VTL
M$29 4 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $30 r0 *1 5.705,0.995 PMOS_VTL
M$30 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $31 r0 *1 5.895,0.995 PMOS_VTL
M$31 4 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $32 r0 *1 6.085,0.995 PMOS_VTL
M$32 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $33 r0 *1 6.275,0.995 PMOS_VTL
M$33 4 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $34 r0 *1 6.465,0.995 PMOS_VTL
M$34 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $35 r0 *1 6.655,0.995 PMOS_VTL
M$35 4 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $36 r0 *1 6.845,0.995 PMOS_VTL
M$36 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $37 r0 *1 7.035,0.995 PMOS_VTL
M$37 4 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $38 r0 *1 7.225,0.995 PMOS_VTL
M$38 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $39 r0 *1 7.415,0.995 PMOS_VTL
M$39 4 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $40 r0 *1 7.605,0.995 PMOS_VTL
M$40 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $41 r0 *1 7.795,0.995 PMOS_VTL
M$41 4 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $42 r0 *1 7.985,0.995 PMOS_VTL
M$42 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $43 r0 *1 8.175,0.995 PMOS_VTL
M$43 4 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $44 r0 *1 8.365,0.995 PMOS_VTL
M$44 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $45 r0 *1 8.555,0.995 PMOS_VTL
M$45 4 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $46 r0 *1 8.745,0.995 PMOS_VTL
M$46 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $47 r0 *1 8.935,0.995 PMOS_VTL
M$47 4 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $48 r0 *1 9.125,0.995 PMOS_VTL
M$48 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $49 r0 *1 0.17,0.2975 NMOS_VTL
M$49 3 2 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $50 r0 *1 0.36,0.2975 NMOS_VTL
M$50 1 2 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $51 r0 *1 0.55,0.2975 NMOS_VTL
M$51 3 2 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $52 r0 *1 0.74,0.2975 NMOS_VTL
M$52 1 2 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $53 r0 *1 0.93,0.2975 NMOS_VTL
M$53 3 2 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $54 r0 *1 1.12,0.2975 NMOS_VTL
M$54 1 2 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $55 r0 *1 1.31,0.2975 NMOS_VTL
M$55 3 2 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $56 r0 *1 1.5,0.2975 NMOS_VTL
M$56 1 2 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $57 r0 *1 1.69,0.2975 NMOS_VTL
M$57 3 2 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $58 r0 *1 1.88,0.2975 NMOS_VTL
M$58 1 2 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $59 r0 *1 2.07,0.2975 NMOS_VTL
M$59 3 2 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $60 r0 *1 2.26,0.2975 NMOS_VTL
M$60 1 2 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $61 r0 *1 2.45,0.2975 NMOS_VTL
M$61 3 2 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $62 r0 *1 2.64,0.2975 NMOS_VTL
M$62 1 2 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $63 r0 *1 2.83,0.2975 NMOS_VTL
M$63 3 2 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.0300875P PS=0.555U
+ PD=0.56U
* device instance $64 r0 *1 3.025,0.2975 NMOS_VTL
M$64 1 2 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.0300875P AD=0.02905P PS=0.56U
+ PD=0.555U
* device instance $65 r0 *1 3.215,0.2975 NMOS_VTL
M$65 4 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.0332P PS=0.555U
+ PD=0.575U
* device instance $66 r0 *1 3.425,0.2975 NMOS_VTL
M$66 1 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.0332P AD=0.02905P PS=0.575U
+ PD=0.555U
* device instance $67 r0 *1 3.615,0.2975 NMOS_VTL
M$67 4 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $68 r0 *1 3.805,0.2975 NMOS_VTL
M$68 1 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $69 r0 *1 3.995,0.2975 NMOS_VTL
M$69 4 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $70 r0 *1 4.185,0.2975 NMOS_VTL
M$70 1 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $71 r0 *1 4.375,0.2975 NMOS_VTL
M$71 4 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $72 r0 *1 4.565,0.2975 NMOS_VTL
M$72 1 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $73 r0 *1 4.755,0.2975 NMOS_VTL
M$73 4 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $74 r0 *1 4.945,0.2975 NMOS_VTL
M$74 1 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $75 r0 *1 5.135,0.2975 NMOS_VTL
M$75 4 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $76 r0 *1 5.325,0.2975 NMOS_VTL
M$76 1 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $77 r0 *1 5.515,0.2975 NMOS_VTL
M$77 4 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $78 r0 *1 5.705,0.2975 NMOS_VTL
M$78 1 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $79 r0 *1 5.895,0.2975 NMOS_VTL
M$79 4 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $80 r0 *1 6.085,0.2975 NMOS_VTL
M$80 1 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $81 r0 *1 6.275,0.2975 NMOS_VTL
M$81 4 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $82 r0 *1 6.465,0.2975 NMOS_VTL
M$82 1 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $83 r0 *1 6.655,0.2975 NMOS_VTL
M$83 4 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $84 r0 *1 6.845,0.2975 NMOS_VTL
M$84 1 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $85 r0 *1 7.035,0.2975 NMOS_VTL
M$85 4 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $86 r0 *1 7.225,0.2975 NMOS_VTL
M$86 1 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $87 r0 *1 7.415,0.2975 NMOS_VTL
M$87 4 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $88 r0 *1 7.605,0.2975 NMOS_VTL
M$88 1 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $89 r0 *1 7.795,0.2975 NMOS_VTL
M$89 4 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $90 r0 *1 7.985,0.2975 NMOS_VTL
M$90 1 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $91 r0 *1 8.175,0.2975 NMOS_VTL
M$91 4 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $92 r0 *1 8.365,0.2975 NMOS_VTL
M$92 1 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $93 r0 *1 8.555,0.2975 NMOS_VTL
M$93 4 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $94 r0 *1 8.745,0.2975 NMOS_VTL
M$94 1 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $95 r0 *1 8.935,0.2975 NMOS_VTL
M$95 4 3 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $96 r0 *1 9.125,0.2975 NMOS_VTL
M$96 1 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS BUF_X32

* cell BUF_X1
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT BUF_X1 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 2 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.033075P PS=0.77U
+ PD=0.84U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.17,0.195 NMOS_VTL
M$3 3 1 2 3 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.021875P PS=0.63U PD=0.555U
* device instance $4 r0 *1 0.36,0.2975 NMOS_VTL
M$4 5 2 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS BUF_X1

* cell CLKBUF_X3
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT CLKBUF_X3 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 4 2 5 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 5 2 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.1875 NMOS_VTL
M$5 3 1 2 3 NMOS_VTL L=0.05U W=0.195U AS=0.020475P AD=0.01365P PS=0.6U PD=0.335U
* device instance $6 r0 *1 0.36,0.1875 NMOS_VTL
M$6 5 2 3 3 NMOS_VTL L=0.05U W=0.195U AS=0.01365P AD=0.01365P PS=0.335U
+ PD=0.335U
* device instance $7 r0 *1 0.55,0.1875 NMOS_VTL
M$7 3 2 5 3 NMOS_VTL L=0.05U W=0.195U AS=0.01365P AD=0.01365P PS=0.335U
+ PD=0.335U
* device instance $8 r0 *1 0.74,0.1875 NMOS_VTL
M$8 5 2 3 3 NMOS_VTL L=0.05U W=0.195U AS=0.01365P AD=0.020475P PS=0.335U PD=0.6U
.ENDS CLKBUF_X3

* cell OAI21_X2
* pin A
* pin B2
* pin B1
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT OAI21_X2 1 2 3 5 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 1 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 8 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 3 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 9 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 5 2 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.17,0.2975 NMOS_VTL
M$7 6 1 4 6 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $8 r0 *1 0.36,0.2975 NMOS_VTL
M$8 4 1 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.55,0.2975 NMOS_VTL
M$9 7 2 4 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.74,0.2975 NMOS_VTL
M$10 4 3 7 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.93,0.2975 NMOS_VTL
M$11 7 3 4 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 1.12,0.2975 NMOS_VTL
M$12 4 2 7 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI21_X2

* cell NAND2_X1
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND2_X1 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 5 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 4 2 5 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.185,0.2975 NMOS_VTL
M$3 6 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $4 r0 *1 0.375,0.2975 NMOS_VTL
M$4 5 2 6 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND2_X1

* cell BUF_X4
* pin A
* pin NWELL,VDD
* pin Z
* pin PWELL,VSS
.SUBCKT BUF_X4 1 3 4 5
* net 1 A
* net 3 NWELL,VDD
* net 4 Z
* net 5 PWELL,VSS
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 2 1 3 3 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 3 1 2 3 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 4 2 3 3 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 3 2 4 3 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 4 2 3 3 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 3 2 4 3 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.17,0.2975 NMOS_VTL
M$7 2 1 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $8 r0 *1 0.36,0.2975 NMOS_VTL
M$8 5 1 2 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.55,0.2975 NMOS_VTL
M$9 4 2 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.74,0.2975 NMOS_VTL
M$10 5 2 4 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.93,0.2975 NMOS_VTL
M$11 4 2 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 1.12,0.2975 NMOS_VTL
M$12 5 2 4 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS BUF_X4

* cell TAPCELL_X1
* pin VSS
* pin VDD
* pin PWELL
* pin NWELL
.SUBCKT TAPCELL_X1 1 2 3 4
* net 1 VSS
* net 2 VDD
* net 3 PWELL
* net 4 NWELL
.ENDS TAPCELL_X1

* cell FILLCELL_X4
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT FILLCELL_X4 1 2
* net 1 PWELL,VSS
* net 2 NWELL,VDD
.ENDS FILLCELL_X4

* cell FILLCELL_X16
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT FILLCELL_X16 1 2
* net 1 PWELL,VSS
* net 2 NWELL,VDD
.ENDS FILLCELL_X16

* cell FILLCELL_X1
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT FILLCELL_X1 1 2
* net 1 PWELL,VSS
* net 2 NWELL,VDD
.ENDS FILLCELL_X1

* cell FILLCELL_X2
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT FILLCELL_X2 1 2
* net 1 PWELL,VSS
* net 2 NWELL,VDD
.ENDS FILLCELL_X2

* cell FILLCELL_X8
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT FILLCELL_X8 1 2
* net 1 PWELL,VSS
* net 2 NWELL,VDD
.ENDS FILLCELL_X8

* cell FILLCELL_X32
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT FILLCELL_X32 1 2
* net 1 PWELL,VSS
* net 2 NWELL,VDD
.ENDS FILLCELL_X32

* cell VIA_via6_0
* pin 
.SUBCKT VIA_via6_0 1
.ENDS VIA_via6_0

* cell VIA_via4_5_960_2800_5_2_600_600
* pin 
.SUBCKT VIA_via4_5_960_2800_5_2_600_600 1
.ENDS VIA_via4_5_960_2800_5_2_600_600

* cell VIA_via5_6_960_2800_5_2_600_600
* pin 
.SUBCKT VIA_via5_6_960_2800_5_2_600_600 1
.ENDS VIA_via5_6_960_2800_5_2_600_600

* cell VIA_via2_3_960_340_1_3_320_320
* pin 
.SUBCKT VIA_via2_3_960_340_1_3_320_320 1
.ENDS VIA_via2_3_960_340_1_3_320_320

* cell VIA_via3_4_960_340_1_3_320_320
* pin 
.SUBCKT VIA_via3_4_960_340_1_3_320_320 1
.ENDS VIA_via3_4_960_340_1_3_320_320

* cell VIA_via5_0
* pin 
.SUBCKT VIA_via5_0 1
.ENDS VIA_via5_0

* cell VIA_via4_0
* pin 
.SUBCKT VIA_via4_0 1
.ENDS VIA_via4_0

* cell VIA_via1_7
* pin 
.SUBCKT VIA_via1_7 1
.ENDS VIA_via1_7

* cell VIA_via3_2
* pin 
.SUBCKT VIA_via3_2 1
.ENDS VIA_via3_2

* cell VIA_via2_5
* pin 
.SUBCKT VIA_via2_5 1
.ENDS VIA_via2_5

* cell VIA_via1_4
* pin 
.SUBCKT VIA_via1_4 1
.ENDS VIA_via1_4

* cell VIA_via1_2_960_340_1_3_300_300
* pin 
.SUBCKT VIA_via1_2_960_340_1_3_300_300 1
.ENDS VIA_via1_2_960_340_1_3_300_300

* cell VIA_via6_7_960_2800_4_1_600_600
* pin 
.SUBCKT VIA_via6_7_960_2800_4_1_600_600 1
.ENDS VIA_via6_7_960_2800_4_1_600_600
