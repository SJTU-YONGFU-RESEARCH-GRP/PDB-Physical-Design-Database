module configurable_carry_select_adder (cin,
    cout,
    a,
    b,
    sum);
 input cin;
 output cout;
 input [63:0] a;
 input [63:0] b;
 output [63:0] sum;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire \first_block.full_adders[0].fa.sum ;
 wire \first_block.full_adders[1].fa.sum ;
 wire \first_block.full_adders[2].fa.sum ;
 wire \first_block.full_adders[3].fa.sum ;
 wire \first_block.full_adders[4].fa.sum ;
 wire \first_block.full_adders[5].fa.sum ;
 wire \first_block.full_adders[6].fa.sum ;
 wire \first_block.full_adders[7].fa.sum ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;

 sky130_fd_sc_hd__inv_1 _408_ (.A(net1),
    .Y(_249_));
 sky130_fd_sc_hd__inv_1 _409_ (.A(net65),
    .Y(_250_));
 sky130_fd_sc_hd__inv_1 _410_ (.A(net129),
    .Y(_251_));
 sky130_fd_sc_hd__inv_1 _411_ (.A(_252_),
    .Y(_253_));
 sky130_fd_sc_hd__inv_1 _412_ (.A(_255_),
    .Y(\first_block.full_adders[1].fa.sum ));
 sky130_fd_sc_hd__inv_1 _413_ (.A(_257_),
    .Y(\first_block.full_adders[2].fa.sum ));
 sky130_fd_sc_hd__inv_1 _414_ (.A(_259_),
    .Y(\first_block.full_adders[3].fa.sum ));
 sky130_fd_sc_hd__inv_1 _415_ (.A(_261_),
    .Y(\first_block.full_adders[4].fa.sum ));
 sky130_fd_sc_hd__inv_1 _416_ (.A(_263_),
    .Y(\first_block.full_adders[5].fa.sum ));
 sky130_fd_sc_hd__inv_1 _417_ (.A(_265_),
    .Y(\first_block.full_adders[6].fa.sum ));
 sky130_fd_sc_hd__inv_1 _418_ (.A(_267_),
    .Y(\first_block.full_adders[7].fa.sum ));
 sky130_fd_sc_hd__inv_1 _419_ (.A(net43),
    .Y(_268_));
 sky130_fd_sc_hd__inv_1 _420_ (.A(net52),
    .Y(_274_));
 sky130_fd_sc_hd__inv_1 _421_ (.A(net8),
    .Y(_280_));
 sky130_fd_sc_hd__inv_1 _422_ (.A(net17),
    .Y(_286_));
 sky130_fd_sc_hd__inv_1 _423_ (.A(net26),
    .Y(_292_));
 sky130_fd_sc_hd__inv_1 _424_ (.A(net35),
    .Y(_298_));
 sky130_fd_sc_hd__inv_1 _425_ (.A(net63),
    .Y(_402_));
 sky130_fd_sc_hd__inv_1 _426_ (.A(net107),
    .Y(_269_));
 sky130_fd_sc_hd__inv_1 _427_ (.A(net116),
    .Y(_275_));
 sky130_fd_sc_hd__inv_1 _428_ (.A(net72),
    .Y(_281_));
 sky130_fd_sc_hd__inv_1 _429_ (.A(net81),
    .Y(_287_));
 sky130_fd_sc_hd__inv_1 _430_ (.A(net90),
    .Y(_293_));
 sky130_fd_sc_hd__inv_1 _431_ (.A(net99),
    .Y(_299_));
 sky130_fd_sc_hd__inv_1 _432_ (.A(net127),
    .Y(_403_));
 sky130_fd_sc_hd__or3_1 _433_ (.A(net58),
    .B(net122),
    .C(_392_),
    .X(_000_));
 sky130_fd_sc_hd__o21a_1 _434_ (.A1(net59),
    .A2(net123),
    .B1(_000_),
    .X(_001_));
 sky130_fd_sc_hd__or2_0 _435_ (.A(net50),
    .B(net114),
    .X(_002_));
 sky130_fd_sc_hd__inv_1 _436_ (.A(_386_),
    .Y(_003_));
 sky130_fd_sc_hd__or2_0 _437_ (.A(net44),
    .B(net108),
    .X(_004_));
 sky130_fd_sc_hd__nand2b_1 _438_ (.A_N(_270_),
    .B(_004_),
    .Y(_005_));
 sky130_fd_sc_hd__nor2_1 _439_ (.A(net46),
    .B(net110),
    .Y(_006_));
 sky130_fd_sc_hd__a21oi_1 _440_ (.A1(_003_),
    .A2(_005_),
    .B1(_006_),
    .Y(_007_));
 sky130_fd_sc_hd__o22a_1 _441_ (.A1(net47),
    .A2(net111),
    .B1(_384_),
    .B2(_007_),
    .X(_008_));
 sky130_fd_sc_hd__nor2_1 _442_ (.A(_382_),
    .B(_008_),
    .Y(_009_));
 sky130_fd_sc_hd__nor2_1 _443_ (.A(net48),
    .B(net112),
    .Y(_010_));
 sky130_fd_sc_hd__o21ba_1 _444_ (.A1(_009_),
    .A2(_010_),
    .B1_N(_380_),
    .X(_011_));
 sky130_fd_sc_hd__nor2_1 _445_ (.A(net49),
    .B(net113),
    .Y(_012_));
 sky130_fd_sc_hd__o21bai_1 _446_ (.A1(_011_),
    .A2(_012_),
    .B1_N(_378_),
    .Y(_013_));
 sky130_fd_sc_hd__a21o_1 _447_ (.A1(_002_),
    .A2(_013_),
    .B1(_376_),
    .X(_014_));
 sky130_fd_sc_hd__inv_1 _448_ (.A(_360_),
    .Y(_015_));
 sky130_fd_sc_hd__nor2_1 _449_ (.A(_342_),
    .B(_344_),
    .Y(_016_));
 sky130_fd_sc_hd__o21ai_0 _450_ (.A1(net18),
    .A2(net82),
    .B1(_290_),
    .Y(_017_));
 sky130_fd_sc_hd__o22ai_1 _451_ (.A1(net20),
    .A2(net84),
    .B1(net21),
    .B2(net85),
    .Y(_018_));
 sky130_fd_sc_hd__nor3_1 _452_ (.A(net19),
    .B(net83),
    .C(_342_),
    .Y(_019_));
 sky130_fd_sc_hd__a211oi_1 _453_ (.A1(_016_),
    .A2(_017_),
    .B1(_018_),
    .C1(_019_),
    .Y(_020_));
 sky130_fd_sc_hd__inv_1 _454_ (.A(_338_),
    .Y(_021_));
 sky130_fd_sc_hd__nor3_1 _455_ (.A(_332_),
    .B(_334_),
    .C(_336_),
    .Y(_022_));
 sky130_fd_sc_hd__o21ai_0 _456_ (.A1(net21),
    .A2(net85),
    .B1(_340_),
    .Y(_023_));
 sky130_fd_sc_hd__nand3_1 _457_ (.A(_021_),
    .B(_022_),
    .C(_023_),
    .Y(_024_));
 sky130_fd_sc_hd__nor2_1 _458_ (.A(net25),
    .B(net89),
    .Y(_025_));
 sky130_fd_sc_hd__nor3_1 _459_ (.A(net24),
    .B(net88),
    .C(_334_),
    .Y(_026_));
 sky130_fd_sc_hd__nor4_1 _460_ (.A(net22),
    .B(net86),
    .C(_334_),
    .D(_336_),
    .Y(_027_));
 sky130_fd_sc_hd__inv_1 _461_ (.A(_332_),
    .Y(_028_));
 sky130_fd_sc_hd__o31ai_2 _462_ (.A1(_025_),
    .A2(_026_),
    .A3(_027_),
    .B1(_028_),
    .Y(_029_));
 sky130_fd_sc_hd__o21a_1 _463_ (.A1(_020_),
    .A2(_024_),
    .B1(_029_),
    .X(_030_));
 sky130_fd_sc_hd__o22ai_1 _464_ (.A1(net15),
    .A2(net79),
    .B1(net16),
    .B2(net80),
    .Y(_031_));
 sky130_fd_sc_hd__nor4_1 _465_ (.A(net11),
    .B(net75),
    .C(_324_),
    .D(_326_),
    .Y(_032_));
 sky130_fd_sc_hd__nor3_1 _466_ (.A(net13),
    .B(net77),
    .C(_324_),
    .Y(_033_));
 sky130_fd_sc_hd__or2_0 _467_ (.A(net14),
    .B(net78),
    .X(_034_));
 sky130_fd_sc_hd__nor4b_1 _468_ (.A(_031_),
    .B(_032_),
    .C(_033_),
    .D_N(_034_),
    .Y(_035_));
 sky130_fd_sc_hd__inv_1 _469_ (.A(_284_),
    .Y(_036_));
 sky130_fd_sc_hd__nor2_1 _470_ (.A(net10),
    .B(net74),
    .Y(_037_));
 sky130_fd_sc_hd__nor2_1 _471_ (.A(net9),
    .B(net73),
    .Y(_038_));
 sky130_fd_sc_hd__nor3_1 _472_ (.A(_324_),
    .B(_326_),
    .C(_328_),
    .Y(_039_));
 sky130_fd_sc_hd__o21ai_0 _473_ (.A1(net10),
    .A2(net74),
    .B1(_330_),
    .Y(_040_));
 sky130_fd_sc_hd__o311ai_0 _474_ (.A1(_036_),
    .A2(_037_),
    .A3(_038_),
    .B1(_039_),
    .C1(_040_),
    .Y(_041_));
 sky130_fd_sc_hd__inv_1 _475_ (.A(_322_),
    .Y(_042_));
 sky130_fd_sc_hd__o21ai_0 _476_ (.A1(net16),
    .A2(net80),
    .B1(_320_),
    .Y(_043_));
 sky130_fd_sc_hd__inv_1 _477_ (.A(_318_),
    .Y(_044_));
 sky130_fd_sc_hd__o211ai_1 _478_ (.A1(_042_),
    .A2(_031_),
    .B1(_043_),
    .C1(_044_),
    .Y(_045_));
 sky130_fd_sc_hd__a21oi_1 _479_ (.A1(_035_),
    .A2(_041_),
    .B1(_045_),
    .Y(_046_));
 sky130_fd_sc_hd__nand2b_1 _480_ (.A_N(_404_),
    .B(_266_),
    .Y(_047_));
 sky130_fd_sc_hd__nand2b_1 _481_ (.A_N(_266_),
    .B(_406_),
    .Y(_048_));
 sky130_fd_sc_hd__nor2_1 _482_ (.A(net64),
    .B(net128),
    .Y(_049_));
 sky130_fd_sc_hd__a21oi_2 _483_ (.A1(_047_),
    .A2(_048_),
    .B1(_049_),
    .Y(_050_));
 sky130_fd_sc_hd__o32a_1 _484_ (.A1(net2),
    .A2(net66),
    .A3(_314_),
    .B1(net67),
    .B2(net3),
    .X(_051_));
 sky130_fd_sc_hd__o22a_1 _485_ (.A1(net4),
    .A2(net68),
    .B1(_312_),
    .B2(_051_),
    .X(_052_));
 sky130_fd_sc_hd__o41ai_4 _486_ (.A1(_312_),
    .A2(_314_),
    .A3(_316_),
    .A4(_050_),
    .B1(_052_),
    .Y(_053_));
 sky130_fd_sc_hd__or3_1 _487_ (.A(net7),
    .B(net71),
    .C(_304_),
    .X(_054_));
 sky130_fd_sc_hd__nor2_1 _488_ (.A(net6),
    .B(net70),
    .Y(_055_));
 sky130_fd_sc_hd__nor2_1 _489_ (.A(net5),
    .B(net69),
    .Y(_056_));
 sky130_fd_sc_hd__nor2_1 _490_ (.A(_055_),
    .B(_056_),
    .Y(_057_));
 sky130_fd_sc_hd__nand2_1 _491_ (.A(_054_),
    .B(_057_),
    .Y(_058_));
 sky130_fd_sc_hd__o21a_1 _492_ (.A1(net5),
    .A2(net69),
    .B1(_310_),
    .X(_059_));
 sky130_fd_sc_hd__nor2_1 _493_ (.A(_308_),
    .B(_059_),
    .Y(_060_));
 sky130_fd_sc_hd__o21ai_0 _494_ (.A1(net6),
    .A2(net70),
    .B1(_054_),
    .Y(_061_));
 sky130_fd_sc_hd__o21ai_0 _495_ (.A1(_304_),
    .A2(_306_),
    .B1(_054_),
    .Y(_062_));
 sky130_fd_sc_hd__o21a_1 _496_ (.A1(_060_),
    .A2(_061_),
    .B1(_062_),
    .X(_063_));
 sky130_fd_sc_hd__o21a_2 _497_ (.A1(_053_),
    .A2(_058_),
    .B1(_063_),
    .X(_064_));
 sky130_fd_sc_hd__nand3_1 _498_ (.A(_030_),
    .B(_046_),
    .C(_064_),
    .Y(_065_));
 sky130_fd_sc_hd__o41a_1 _499_ (.A1(_312_),
    .A2(_314_),
    .A3(_316_),
    .A4(_050_),
    .B1(_052_),
    .X(_066_));
 sky130_fd_sc_hd__nor2_1 _500_ (.A(_304_),
    .B(_306_),
    .Y(_067_));
 sky130_fd_sc_hd__o21ai_0 _501_ (.A1(_055_),
    .A2(_060_),
    .B1(_067_),
    .Y(_068_));
 sky130_fd_sc_hd__a21oi_1 _502_ (.A1(_066_),
    .A2(_057_),
    .B1(_068_),
    .Y(_069_));
 sky130_fd_sc_hd__o311ai_0 _503_ (.A1(_282_),
    .A2(_037_),
    .A3(_038_),
    .B1(_039_),
    .C1(_040_),
    .Y(_070_));
 sky130_fd_sc_hd__a21oi_1 _504_ (.A1(_035_),
    .A2(_070_),
    .B1(_045_),
    .Y(_071_));
 sky130_fd_sc_hd__nand3_1 _505_ (.A(_030_),
    .B(_054_),
    .C(_071_),
    .Y(_072_));
 sky130_fd_sc_hd__o32a_1 _506_ (.A1(net20),
    .A2(net84),
    .A3(_340_),
    .B1(net85),
    .B2(net21),
    .X(_073_));
 sky130_fd_sc_hd__nor2_1 _507_ (.A(net19),
    .B(net83),
    .Y(_074_));
 sky130_fd_sc_hd__nor3_1 _508_ (.A(net18),
    .B(net82),
    .C(_344_),
    .Y(_075_));
 sky130_fd_sc_hd__nor2b_1 _509_ (.A(_344_),
    .B_N(_288_),
    .Y(_076_));
 sky130_fd_sc_hd__nor2_1 _510_ (.A(_340_),
    .B(_342_),
    .Y(_077_));
 sky130_fd_sc_hd__o31ai_1 _511_ (.A1(_074_),
    .A2(_075_),
    .A3(_076_),
    .B1(_077_),
    .Y(_078_));
 sky130_fd_sc_hd__a21oi_1 _512_ (.A1(_073_),
    .A2(_078_),
    .B1(_338_),
    .Y(_079_));
 sky130_fd_sc_hd__nand2_2 _513_ (.A(_022_),
    .B(_079_),
    .Y(_080_));
 sky130_fd_sc_hd__a2bb2oi_2 _514_ (.A1_N(_069_),
    .A2_N(_072_),
    .B1(_080_),
    .B2(_030_),
    .Y(_081_));
 sky130_fd_sc_hd__inv_1 _515_ (.A(_071_),
    .Y(_082_));
 sky130_fd_sc_hd__o211ai_2 _516_ (.A1(_053_),
    .A2(_058_),
    .B1(_063_),
    .C1(_046_),
    .Y(_083_));
 sky130_fd_sc_hd__o2111ai_4 _517_ (.A1(_064_),
    .A2(_082_),
    .B1(_080_),
    .C1(_083_),
    .D1(_029_),
    .Y(_084_));
 sky130_fd_sc_hd__nor2_1 _518_ (.A(net32),
    .B(net96),
    .Y(_085_));
 sky130_fd_sc_hd__nor2_1 _519_ (.A(net31),
    .B(net95),
    .Y(_086_));
 sky130_fd_sc_hd__nor2_1 _520_ (.A(net33),
    .B(net97),
    .Y(_087_));
 sky130_fd_sc_hd__nor2_1 _521_ (.A(net30),
    .B(net94),
    .Y(_088_));
 sky130_fd_sc_hd__nor4_1 _522_ (.A(_085_),
    .B(_086_),
    .C(_087_),
    .D(_088_),
    .Y(_089_));
 sky130_fd_sc_hd__nor2_1 _523_ (.A(net29),
    .B(net93),
    .Y(_090_));
 sky130_fd_sc_hd__inv_1 _524_ (.A(_358_),
    .Y(_091_));
 sky130_fd_sc_hd__o21bai_1 _525_ (.A1(net27),
    .A2(net91),
    .B1_N(_294_),
    .Y(_092_));
 sky130_fd_sc_hd__nor2_1 _526_ (.A(net28),
    .B(net92),
    .Y(_093_));
 sky130_fd_sc_hd__a21oi_1 _527_ (.A1(_091_),
    .A2(_092_),
    .B1(_093_),
    .Y(_094_));
 sky130_fd_sc_hd__nor2_1 _528_ (.A(_356_),
    .B(_094_),
    .Y(_095_));
 sky130_fd_sc_hd__o21bai_1 _529_ (.A1(_090_),
    .A2(_095_),
    .B1_N(_354_),
    .Y(_096_));
 sky130_fd_sc_hd__o21a_1 _530_ (.A1(net31),
    .A2(net95),
    .B1(_352_),
    .X(_097_));
 sky130_fd_sc_hd__nor2_1 _531_ (.A(_350_),
    .B(_097_),
    .Y(_098_));
 sky130_fd_sc_hd__o21bai_1 _532_ (.A1(_085_),
    .A2(_098_),
    .B1_N(_348_),
    .Y(_099_));
 sky130_fd_sc_hd__inv_1 _533_ (.A(_087_),
    .Y(_100_));
 sky130_fd_sc_hd__a21o_1 _534_ (.A1(_099_),
    .A2(_100_),
    .B1(_346_),
    .X(_101_));
 sky130_fd_sc_hd__a21o_1 _535_ (.A1(_089_),
    .A2(_096_),
    .B1(_101_),
    .X(_102_));
 sky130_fd_sc_hd__a31o_1 _536_ (.A1(_065_),
    .A2(_081_),
    .A3(_084_),
    .B1(_102_),
    .X(_103_));
 sky130_fd_sc_hd__o21ai_0 _537_ (.A1(net27),
    .A2(net91),
    .B1(_296_),
    .Y(_104_));
 sky130_fd_sc_hd__a21oi_1 _538_ (.A1(_091_),
    .A2(_104_),
    .B1(_093_),
    .Y(_105_));
 sky130_fd_sc_hd__nor2_1 _539_ (.A(_356_),
    .B(_105_),
    .Y(_106_));
 sky130_fd_sc_hd__o21bai_1 _540_ (.A1(_090_),
    .A2(_106_),
    .B1_N(_354_),
    .Y(_107_));
 sky130_fd_sc_hd__a21oi_1 _541_ (.A1(_089_),
    .A2(_107_),
    .B1(_101_),
    .Y(_108_));
 sky130_fd_sc_hd__nand4_2 _542_ (.A(_065_),
    .B(_081_),
    .C(_084_),
    .D(_108_),
    .Y(_109_));
 sky130_fd_sc_hd__or2_0 _543_ (.A(net41),
    .B(net105),
    .X(_110_));
 sky130_fd_sc_hd__or2_0 _544_ (.A(net40),
    .B(net104),
    .X(_111_));
 sky130_fd_sc_hd__nand2_1 _545_ (.A(_110_),
    .B(_111_),
    .Y(_112_));
 sky130_fd_sc_hd__inv_1 _546_ (.A(_368_),
    .Y(_113_));
 sky130_fd_sc_hd__inv_1 _547_ (.A(_372_),
    .Y(_114_));
 sky130_fd_sc_hd__o21ai_0 _548_ (.A1(net36),
    .A2(net100),
    .B1(_302_),
    .Y(_115_));
 sky130_fd_sc_hd__nor2_1 _549_ (.A(net37),
    .B(net101),
    .Y(_116_));
 sky130_fd_sc_hd__a21oi_1 _550_ (.A1(_114_),
    .A2(_115_),
    .B1(_116_),
    .Y(_117_));
 sky130_fd_sc_hd__or2_0 _551_ (.A(net38),
    .B(net102),
    .X(_118_));
 sky130_fd_sc_hd__o21ai_0 _552_ (.A1(_370_),
    .A2(_117_),
    .B1(_118_),
    .Y(_119_));
 sky130_fd_sc_hd__nor2_1 _553_ (.A(net39),
    .B(net103),
    .Y(_120_));
 sky130_fd_sc_hd__a21oi_1 _554_ (.A1(_113_),
    .A2(_119_),
    .B1(_120_),
    .Y(_121_));
 sky130_fd_sc_hd__nor2_1 _555_ (.A(_366_),
    .B(_121_),
    .Y(_122_));
 sky130_fd_sc_hd__a21oi_1 _556_ (.A1(_364_),
    .A2(_110_),
    .B1(_362_),
    .Y(_123_));
 sky130_fd_sc_hd__o21a_1 _557_ (.A1(_112_),
    .A2(_122_),
    .B1(_123_),
    .X(_124_));
 sky130_fd_sc_hd__nor2_1 _558_ (.A(net42),
    .B(net106),
    .Y(_125_));
 sky130_fd_sc_hd__a211o_1 _559_ (.A1(_103_),
    .A2(_109_),
    .B1(_124_),
    .C1(_125_),
    .X(_126_));
 sky130_fd_sc_hd__o21bai_1 _560_ (.A1(net36),
    .A2(net100),
    .B1_N(_300_),
    .Y(_127_));
 sky130_fd_sc_hd__a21oi_1 _561_ (.A1(_114_),
    .A2(_127_),
    .B1(_116_),
    .Y(_128_));
 sky130_fd_sc_hd__o21ai_0 _562_ (.A1(_370_),
    .A2(_128_),
    .B1(_118_),
    .Y(_129_));
 sky130_fd_sc_hd__a21oi_1 _563_ (.A1(_113_),
    .A2(_129_),
    .B1(_120_),
    .Y(_130_));
 sky130_fd_sc_hd__o21bai_1 _564_ (.A1(_366_),
    .A2(_130_),
    .B1_N(_112_),
    .Y(_131_));
 sky130_fd_sc_hd__a21oi_1 _565_ (.A1(_123_),
    .A2(_131_),
    .B1(_125_),
    .Y(_132_));
 sky130_fd_sc_hd__nand3_2 _566_ (.A(_103_),
    .B(_109_),
    .C(_132_),
    .Y(_133_));
 sky130_fd_sc_hd__and3_1 _567_ (.A(_015_),
    .B(_126_),
    .C(_133_),
    .X(_134_));
 sky130_fd_sc_hd__buf_6 _568_ (.A(_134_),
    .X(_135_));
 sky130_fd_sc_hd__o21ai_0 _569_ (.A1(net44),
    .A2(net108),
    .B1(_272_),
    .Y(_136_));
 sky130_fd_sc_hd__a21oi_1 _570_ (.A1(_003_),
    .A2(_136_),
    .B1(_006_),
    .Y(_137_));
 sky130_fd_sc_hd__o22a_1 _571_ (.A1(net47),
    .A2(net111),
    .B1(_384_),
    .B2(_137_),
    .X(_138_));
 sky130_fd_sc_hd__nor2_1 _572_ (.A(_382_),
    .B(_138_),
    .Y(_139_));
 sky130_fd_sc_hd__o21ba_1 _573_ (.A1(_010_),
    .A2(_139_),
    .B1_N(_380_),
    .X(_140_));
 sky130_fd_sc_hd__o21bai_1 _574_ (.A1(_012_),
    .A2(_140_),
    .B1_N(_378_),
    .Y(_141_));
 sky130_fd_sc_hd__a21oi_2 _575_ (.A1(_002_),
    .A2(_141_),
    .B1(_376_),
    .Y(_142_));
 sky130_fd_sc_hd__nor2_1 _576_ (.A(_360_),
    .B(_374_),
    .Y(_143_));
 sky130_fd_sc_hd__nor3_1 _577_ (.A(net51),
    .B(net115),
    .C(_374_),
    .Y(_144_));
 sky130_fd_sc_hd__a41oi_4 _578_ (.A1(_126_),
    .A2(_133_),
    .A3(_142_),
    .A4(_143_),
    .B1(_144_),
    .Y(_145_));
 sky130_fd_sc_hd__o31ai_4 _579_ (.A1(_374_),
    .A2(_014_),
    .A3(_135_),
    .B1(_145_),
    .Y(_146_));
 sky130_fd_sc_hd__nor2_1 _580_ (.A(net55),
    .B(net119),
    .Y(_147_));
 sky130_fd_sc_hd__or2_0 _581_ (.A(net54),
    .B(net118),
    .X(_148_));
 sky130_fd_sc_hd__o21ai_0 _582_ (.A1(net53),
    .A2(net117),
    .B1(_278_),
    .Y(_149_));
 sky130_fd_sc_hd__nand2b_1 _583_ (.A_N(_400_),
    .B(_149_),
    .Y(_150_));
 sky130_fd_sc_hd__a21oi_1 _584_ (.A1(_148_),
    .A2(_150_),
    .B1(_398_),
    .Y(_151_));
 sky130_fd_sc_hd__nor2_1 _585_ (.A(_147_),
    .B(_151_),
    .Y(_152_));
 sky130_fd_sc_hd__nor2_1 _586_ (.A(_396_),
    .B(_152_),
    .Y(_153_));
 sky130_fd_sc_hd__nor2_1 _587_ (.A(net53),
    .B(net117),
    .Y(_154_));
 sky130_fd_sc_hd__o21bai_1 _588_ (.A1(_276_),
    .A2(_154_),
    .B1_N(_400_),
    .Y(_155_));
 sky130_fd_sc_hd__a21oi_1 _589_ (.A1(_148_),
    .A2(_155_),
    .B1(_398_),
    .Y(_156_));
 sky130_fd_sc_hd__nor2_1 _590_ (.A(_147_),
    .B(_156_),
    .Y(_157_));
 sky130_fd_sc_hd__nor2_1 _591_ (.A(_396_),
    .B(_157_),
    .Y(_158_));
 sky130_fd_sc_hd__o311a_1 _592_ (.A1(_374_),
    .A2(_014_),
    .A3(_135_),
    .B1(_145_),
    .C1(_158_),
    .X(_159_));
 sky130_fd_sc_hd__nor2_1 _593_ (.A(net57),
    .B(net121),
    .Y(_160_));
 sky130_fd_sc_hd__a211oi_2 _594_ (.A1(_146_),
    .A2(_153_),
    .B1(_159_),
    .C1(_160_),
    .Y(_161_));
 sky130_fd_sc_hd__or3_1 _595_ (.A(_390_),
    .B(_392_),
    .C(_394_),
    .X(_162_));
 sky130_fd_sc_hd__o22ai_1 _596_ (.A1(_390_),
    .A2(_001_),
    .B1(_161_),
    .B2(_162_),
    .Y(_163_));
 sky130_fd_sc_hd__nor2_1 _597_ (.A(net60),
    .B(net124),
    .Y(_164_));
 sky130_fd_sc_hd__o21bai_1 _598_ (.A1(_163_),
    .A2(_164_),
    .B1_N(_388_),
    .Y(net130));
 sky130_fd_sc_hd__nor2_1 _599_ (.A(_316_),
    .B(_050_),
    .Y(_165_));
 sky130_fd_sc_hd__xnor2_1 _600_ (.A(_315_),
    .B(_165_),
    .Y(net132));
 sky130_fd_sc_hd__nor2_1 _601_ (.A(net2),
    .B(net66),
    .Y(_166_));
 sky130_fd_sc_hd__o21bai_1 _602_ (.A1(_166_),
    .A2(_165_),
    .B1_N(_314_),
    .Y(_167_));
 sky130_fd_sc_hd__xor2_1 _603_ (.A(_313_),
    .B(_167_),
    .X(net133));
 sky130_fd_sc_hd__or2_0 _604_ (.A(net3),
    .B(net67),
    .X(_168_));
 sky130_fd_sc_hd__a21oi_1 _605_ (.A1(_168_),
    .A2(_167_),
    .B1(_312_),
    .Y(_169_));
 sky130_fd_sc_hd__xnor2_1 _606_ (.A(_311_),
    .B(_169_),
    .Y(net134));
 sky130_fd_sc_hd__nor2_1 _607_ (.A(_310_),
    .B(_066_),
    .Y(_170_));
 sky130_fd_sc_hd__xnor2_1 _608_ (.A(_309_),
    .B(_170_),
    .Y(net135));
 sky130_fd_sc_hd__o21ai_1 _609_ (.A1(_056_),
    .A2(_053_),
    .B1(_060_),
    .Y(_171_));
 sky130_fd_sc_hd__xor2_1 _610_ (.A(_307_),
    .B(_171_),
    .X(net136));
 sky130_fd_sc_hd__inv_1 _611_ (.A(_055_),
    .Y(_172_));
 sky130_fd_sc_hd__a21oi_1 _612_ (.A1(_172_),
    .A2(_171_),
    .B1(_306_),
    .Y(_173_));
 sky130_fd_sc_hd__xnor2_1 _613_ (.A(_305_),
    .B(_173_),
    .Y(net137));
 sky130_fd_sc_hd__xnor2_1 _614_ (.A(_283_),
    .B(_064_),
    .Y(net138));
 sky130_fd_sc_hd__nor2_1 _615_ (.A(_282_),
    .B(_064_),
    .Y(_174_));
 sky130_fd_sc_hd__a21oi_1 _616_ (.A1(_284_),
    .A2(_064_),
    .B1(_174_),
    .Y(_175_));
 sky130_fd_sc_hd__xnor2_1 _617_ (.A(_331_),
    .B(_175_),
    .Y(net139));
 sky130_fd_sc_hd__o21ba_1 _618_ (.A1(_038_),
    .A2(_175_),
    .B1_N(_330_),
    .X(_176_));
 sky130_fd_sc_hd__xnor2_1 _619_ (.A(_329_),
    .B(_176_),
    .Y(net140));
 sky130_fd_sc_hd__o21bai_2 _620_ (.A1(_037_),
    .A2(_176_),
    .B1_N(_328_),
    .Y(_177_));
 sky130_fd_sc_hd__xor2_1 _621_ (.A(_327_),
    .B(_177_),
    .X(net141));
 sky130_fd_sc_hd__or2_0 _622_ (.A(net11),
    .B(net75),
    .X(_178_));
 sky130_fd_sc_hd__a21oi_1 _623_ (.A1(_178_),
    .A2(_177_),
    .B1(_326_),
    .Y(_179_));
 sky130_fd_sc_hd__xnor2_1 _624_ (.A(_325_),
    .B(_179_),
    .Y(net143));
 sky130_fd_sc_hd__nor2_1 _625_ (.A(_032_),
    .B(_033_),
    .Y(_180_));
 sky130_fd_sc_hd__o31a_1 _626_ (.A1(_324_),
    .A2(_326_),
    .A3(_177_),
    .B1(_180_),
    .X(_181_));
 sky130_fd_sc_hd__xor2_1 _627_ (.A(_323_),
    .B(_181_),
    .X(net144));
 sky130_fd_sc_hd__a21oi_1 _628_ (.A1(_034_),
    .A2(_181_),
    .B1(_322_),
    .Y(_182_));
 sky130_fd_sc_hd__xnor2_1 _629_ (.A(_321_),
    .B(_182_),
    .Y(net145));
 sky130_fd_sc_hd__nor2_1 _630_ (.A(net15),
    .B(net79),
    .Y(_183_));
 sky130_fd_sc_hd__o21bai_1 _631_ (.A1(_183_),
    .A2(_182_),
    .B1_N(_320_),
    .Y(_184_));
 sky130_fd_sc_hd__xor2_1 _632_ (.A(_319_),
    .B(_184_),
    .X(net146));
 sky130_fd_sc_hd__o21a_1 _633_ (.A1(_064_),
    .A2(_082_),
    .B1(_083_),
    .X(_185_));
 sky130_fd_sc_hd__xor2_1 _634_ (.A(_289_),
    .B(_185_),
    .X(net147));
 sky130_fd_sc_hd__inv_1 _635_ (.A(_288_),
    .Y(_186_));
 sky130_fd_sc_hd__mux2i_2 _636_ (.A0(_290_),
    .A1(_186_),
    .S(_185_),
    .Y(_187_));
 sky130_fd_sc_hd__xnor2_1 _637_ (.A(_345_),
    .B(_187_),
    .Y(net148));
 sky130_fd_sc_hd__nor2_1 _638_ (.A(net18),
    .B(net82),
    .Y(_188_));
 sky130_fd_sc_hd__nor2_1 _639_ (.A(_188_),
    .B(_187_),
    .Y(_189_));
 sky130_fd_sc_hd__nor2_1 _640_ (.A(_344_),
    .B(_189_),
    .Y(_190_));
 sky130_fd_sc_hd__xnor2_1 _641_ (.A(_343_),
    .B(_190_),
    .Y(net149));
 sky130_fd_sc_hd__nor2_1 _642_ (.A(_074_),
    .B(_190_),
    .Y(_191_));
 sky130_fd_sc_hd__nor2_1 _643_ (.A(_342_),
    .B(_191_),
    .Y(_192_));
 sky130_fd_sc_hd__xnor2_1 _644_ (.A(_341_),
    .B(_192_),
    .Y(net150));
 sky130_fd_sc_hd__o22a_1 _645_ (.A1(net20),
    .A2(net84),
    .B1(_342_),
    .B2(_191_),
    .X(_193_));
 sky130_fd_sc_hd__nor2_1 _646_ (.A(_340_),
    .B(_193_),
    .Y(_194_));
 sky130_fd_sc_hd__xnor2_1 _647_ (.A(_339_),
    .B(_194_),
    .Y(net151));
 sky130_fd_sc_hd__nand2_1 _648_ (.A(_021_),
    .B(_023_),
    .Y(_195_));
 sky130_fd_sc_hd__nand2_1 _649_ (.A(_079_),
    .B(_185_),
    .Y(_196_));
 sky130_fd_sc_hd__o31a_1 _650_ (.A1(_020_),
    .A2(_195_),
    .A3(_185_),
    .B1(_196_),
    .X(_197_));
 sky130_fd_sc_hd__xor2_1 _651_ (.A(_337_),
    .B(_197_),
    .X(net152));
 sky130_fd_sc_hd__or2_0 _652_ (.A(net22),
    .B(net86),
    .X(_198_));
 sky130_fd_sc_hd__a21oi_1 _653_ (.A1(_198_),
    .A2(_197_),
    .B1(_336_),
    .Y(_199_));
 sky130_fd_sc_hd__xnor2_1 _654_ (.A(_335_),
    .B(_199_),
    .Y(net154));
 sky130_fd_sc_hd__nor2_1 _655_ (.A(net24),
    .B(net88),
    .Y(_200_));
 sky130_fd_sc_hd__nor2_1 _656_ (.A(_200_),
    .B(_199_),
    .Y(_201_));
 sky130_fd_sc_hd__nor2_1 _657_ (.A(_334_),
    .B(_201_),
    .Y(_202_));
 sky130_fd_sc_hd__xnor2_1 _658_ (.A(_333_),
    .B(_202_),
    .Y(net155));
 sky130_fd_sc_hd__and3_1 _659_ (.A(_065_),
    .B(_081_),
    .C(_084_),
    .X(_203_));
 sky130_fd_sc_hd__xnor2_1 _660_ (.A(_295_),
    .B(_203_),
    .Y(net156));
 sky130_fd_sc_hd__and3_1 _661_ (.A(_030_),
    .B(_046_),
    .C(_064_),
    .X(_204_));
 sky130_fd_sc_hd__o2bb2ai_1 _662_ (.A1_N(_030_),
    .A2_N(_080_),
    .B1(_072_),
    .B2(_069_),
    .Y(_205_));
 sky130_fd_sc_hd__nor4b_1 _663_ (.A(_296_),
    .B(_204_),
    .C(_205_),
    .D_N(_084_),
    .Y(_206_));
 sky130_fd_sc_hd__inv_1 _664_ (.A(_294_),
    .Y(_207_));
 sky130_fd_sc_hd__a31oi_1 _665_ (.A1(_065_),
    .A2(_081_),
    .A3(_084_),
    .B1(_207_),
    .Y(_208_));
 sky130_fd_sc_hd__or2_0 _666_ (.A(_206_),
    .B(_208_),
    .X(_209_));
 sky130_fd_sc_hd__xnor2_1 _667_ (.A(_359_),
    .B(_209_),
    .Y(net157));
 sky130_fd_sc_hd__nor2_1 _668_ (.A(net27),
    .B(net91),
    .Y(_210_));
 sky130_fd_sc_hd__o31a_1 _669_ (.A1(_210_),
    .A2(_206_),
    .A3(_208_),
    .B1(_091_),
    .X(_211_));
 sky130_fd_sc_hd__xnor2_1 _670_ (.A(_357_),
    .B(_211_),
    .Y(net158));
 sky130_fd_sc_hd__o21ba_1 _671_ (.A1(_093_),
    .A2(_211_),
    .B1_N(_356_),
    .X(_212_));
 sky130_fd_sc_hd__xnor2_1 _672_ (.A(_355_),
    .B(_212_),
    .Y(net159));
 sky130_fd_sc_hd__o21bai_2 _673_ (.A1(_090_),
    .A2(_212_),
    .B1_N(_354_),
    .Y(_213_));
 sky130_fd_sc_hd__xor2_1 _674_ (.A(_353_),
    .B(_213_),
    .X(net160));
 sky130_fd_sc_hd__or2_0 _675_ (.A(net30),
    .B(net94),
    .X(_214_));
 sky130_fd_sc_hd__a21oi_1 _676_ (.A1(_214_),
    .A2(_213_),
    .B1(_352_),
    .Y(_215_));
 sky130_fd_sc_hd__xnor2_1 _677_ (.A(_351_),
    .B(_215_),
    .Y(net161));
 sky130_fd_sc_hd__o21bai_1 _678_ (.A1(_086_),
    .A2(_215_),
    .B1_N(_350_),
    .Y(_216_));
 sky130_fd_sc_hd__xor2_1 _679_ (.A(_349_),
    .B(_216_),
    .X(net162));
 sky130_fd_sc_hd__nor3_1 _680_ (.A(_085_),
    .B(_086_),
    .C(_088_),
    .Y(_217_));
 sky130_fd_sc_hd__a21oi_1 _681_ (.A1(_217_),
    .A2(_213_),
    .B1(_099_),
    .Y(_218_));
 sky130_fd_sc_hd__xnor2_1 _682_ (.A(_347_),
    .B(_218_),
    .Y(net163));
 sky130_fd_sc_hd__and2_0 _683_ (.A(_103_),
    .B(_109_),
    .X(_219_));
 sky130_fd_sc_hd__clkbuf_2 _684_ (.A(_219_),
    .X(_220_));
 sky130_fd_sc_hd__xor2_1 _685_ (.A(_301_),
    .B(_220_),
    .X(net165));
 sky130_fd_sc_hd__nand3_1 _686_ (.A(_300_),
    .B(_103_),
    .C(_109_),
    .Y(_221_));
 sky130_fd_sc_hd__o21ai_1 _687_ (.A1(_302_),
    .A2(_220_),
    .B1(_221_),
    .Y(_222_));
 sky130_fd_sc_hd__xnor2_1 _688_ (.A(_373_),
    .B(_222_),
    .Y(net166));
 sky130_fd_sc_hd__nor2_1 _689_ (.A(net36),
    .B(net100),
    .Y(_223_));
 sky130_fd_sc_hd__o21a_1 _690_ (.A1(_223_),
    .A2(_222_),
    .B1(_114_),
    .X(_224_));
 sky130_fd_sc_hd__xnor2_1 _691_ (.A(_371_),
    .B(_224_),
    .Y(net167));
 sky130_fd_sc_hd__o21bai_1 _692_ (.A1(_116_),
    .A2(_224_),
    .B1_N(_370_),
    .Y(_225_));
 sky130_fd_sc_hd__xor2_1 _693_ (.A(_369_),
    .B(_225_),
    .X(net168));
 sky130_fd_sc_hd__a21oi_1 _694_ (.A1(_118_),
    .A2(_225_),
    .B1(_368_),
    .Y(_226_));
 sky130_fd_sc_hd__xnor2_1 _695_ (.A(_367_),
    .B(_226_),
    .Y(net169));
 sky130_fd_sc_hd__nor2_1 _696_ (.A(_366_),
    .B(_130_),
    .Y(_227_));
 sky130_fd_sc_hd__mux2i_2 _697_ (.A0(_122_),
    .A1(_227_),
    .S(_220_),
    .Y(_228_));
 sky130_fd_sc_hd__xor2_1 _698_ (.A(_365_),
    .B(_228_),
    .X(net170));
 sky130_fd_sc_hd__a21oi_1 _699_ (.A1(_111_),
    .A2(_228_),
    .B1(_364_),
    .Y(_229_));
 sky130_fd_sc_hd__xnor2_1 _700_ (.A(_363_),
    .B(_229_),
    .Y(net171));
 sky130_fd_sc_hd__nor2b_1 _701_ (.A(_220_),
    .B_N(_124_),
    .Y(_230_));
 sky130_fd_sc_hd__a31oi_1 _702_ (.A1(_220_),
    .A2(_123_),
    .A3(_131_),
    .B1(_230_),
    .Y(_231_));
 sky130_fd_sc_hd__xor2_1 _703_ (.A(_361_),
    .B(_231_),
    .X(net172));
 sky130_fd_sc_hd__xnor2_1 _704_ (.A(_271_),
    .B(_135_),
    .Y(net173));
 sky130_fd_sc_hd__nand4_1 _705_ (.A(_272_),
    .B(_015_),
    .C(_126_),
    .D(_133_),
    .Y(_232_));
 sky130_fd_sc_hd__o21ai_1 _706_ (.A1(_270_),
    .A2(_135_),
    .B1(_232_),
    .Y(_233_));
 sky130_fd_sc_hd__xor2_1 _707_ (.A(_387_),
    .B(_233_),
    .X(net174));
 sky130_fd_sc_hd__a21oi_1 _708_ (.A1(_004_),
    .A2(_233_),
    .B1(_386_),
    .Y(_234_));
 sky130_fd_sc_hd__xnor2_1 _709_ (.A(_385_),
    .B(_234_),
    .Y(net176));
 sky130_fd_sc_hd__o21bai_1 _710_ (.A1(_006_),
    .A2(_234_),
    .B1_N(_384_),
    .Y(_235_));
 sky130_fd_sc_hd__xor2_1 _711_ (.A(_383_),
    .B(_235_),
    .X(net177));
 sky130_fd_sc_hd__mux2i_1 _712_ (.A0(_009_),
    .A1(_139_),
    .S(_135_),
    .Y(_236_));
 sky130_fd_sc_hd__xor2_1 _713_ (.A(_381_),
    .B(_236_),
    .X(net178));
 sky130_fd_sc_hd__mux2i_1 _714_ (.A0(_011_),
    .A1(_140_),
    .S(_135_),
    .Y(_237_));
 sky130_fd_sc_hd__xor2_1 _715_ (.A(_379_),
    .B(_237_),
    .X(net179));
 sky130_fd_sc_hd__mux2i_1 _716_ (.A0(_013_),
    .A1(_141_),
    .S(_135_),
    .Y(_238_));
 sky130_fd_sc_hd__xnor2_1 _717_ (.A(_377_),
    .B(_238_),
    .Y(net180));
 sky130_fd_sc_hd__nor2_1 _718_ (.A(_014_),
    .B(_135_),
    .Y(_239_));
 sky130_fd_sc_hd__a21o_1 _719_ (.A1(_135_),
    .A2(_142_),
    .B1(_239_),
    .X(_240_));
 sky130_fd_sc_hd__xnor2_1 _720_ (.A(_375_),
    .B(_240_),
    .Y(net181));
 sky130_fd_sc_hd__xnor2_1 _721_ (.A(_277_),
    .B(_146_),
    .Y(net182));
 sky130_fd_sc_hd__nor2_1 _722_ (.A(_276_),
    .B(_146_),
    .Y(_241_));
 sky130_fd_sc_hd__a21oi_1 _723_ (.A1(_278_),
    .A2(_146_),
    .B1(_241_),
    .Y(_242_));
 sky130_fd_sc_hd__xnor2_1 _724_ (.A(_401_),
    .B(_242_),
    .Y(net183));
 sky130_fd_sc_hd__mux2_1 _725_ (.A0(_155_),
    .A1(_150_),
    .S(_146_),
    .X(_243_));
 sky130_fd_sc_hd__xor2_1 _726_ (.A(_399_),
    .B(_243_),
    .X(net184));
 sky130_fd_sc_hd__a21oi_1 _727_ (.A1(_148_),
    .A2(_243_),
    .B1(_398_),
    .Y(_244_));
 sky130_fd_sc_hd__xnor2_1 _728_ (.A(_397_),
    .B(_244_),
    .Y(net185));
 sky130_fd_sc_hd__a21oi_1 _729_ (.A1(_146_),
    .A2(_153_),
    .B1(_159_),
    .Y(_245_));
 sky130_fd_sc_hd__xor2_1 _730_ (.A(_395_),
    .B(_245_),
    .X(net187));
 sky130_fd_sc_hd__nor2_1 _731_ (.A(_394_),
    .B(_161_),
    .Y(_246_));
 sky130_fd_sc_hd__xnor2_1 _732_ (.A(_393_),
    .B(_246_),
    .Y(net188));
 sky130_fd_sc_hd__o31ai_1 _733_ (.A1(_392_),
    .A2(_394_),
    .A3(_161_),
    .B1(_000_),
    .Y(_247_));
 sky130_fd_sc_hd__xnor2_1 _734_ (.A(_391_),
    .B(_247_),
    .Y(net189));
 sky130_fd_sc_hd__xnor2_1 _735_ (.A(_389_),
    .B(_163_),
    .Y(net190));
 sky130_fd_sc_hd__xor2_1 _736_ (.A(_266_),
    .B(_405_),
    .X(net193));
 sky130_fd_sc_hd__nand2_1 _737_ (.A(_047_),
    .B(_048_),
    .Y(_248_));
 sky130_fd_sc_hd__xor2_1 _738_ (.A(_317_),
    .B(_248_),
    .X(net194));
 sky130_fd_sc_hd__fa_1 _739_ (.A(_249_),
    .B(_250_),
    .CIN(_251_),
    .COUT(_252_),
    .SUM(\first_block.full_adders[0].fa.sum ));
 sky130_fd_sc_hd__fa_1 _740_ (.A(net12),
    .B(net76),
    .CIN(_253_),
    .COUT(_254_),
    .SUM(_255_));
 sky130_fd_sc_hd__fa_1 _741_ (.A(net23),
    .B(net87),
    .CIN(_254_),
    .COUT(_256_),
    .SUM(_257_));
 sky130_fd_sc_hd__fa_1 _742_ (.A(net34),
    .B(net98),
    .CIN(_256_),
    .COUT(_258_),
    .SUM(_259_));
 sky130_fd_sc_hd__fa_1 _743_ (.A(net45),
    .B(net109),
    .CIN(_258_),
    .COUT(_260_),
    .SUM(_261_));
 sky130_fd_sc_hd__fa_1 _744_ (.A(net56),
    .B(net120),
    .CIN(_260_),
    .COUT(_262_),
    .SUM(_263_));
 sky130_fd_sc_hd__fa_1 _745_ (.A(net61),
    .B(net125),
    .CIN(_262_),
    .COUT(_264_),
    .SUM(_265_));
 sky130_fd_sc_hd__fa_1 _746_ (.A(net62),
    .B(net126),
    .CIN(_264_),
    .COUT(_266_),
    .SUM(_267_));
 sky130_fd_sc_hd__ha_1 _747_ (.A(_268_),
    .B(_269_),
    .COUT(_270_),
    .SUM(_271_));
 sky130_fd_sc_hd__ha_1 _748_ (.A(net43),
    .B(net107),
    .COUT(_272_),
    .SUM(_273_));
 sky130_fd_sc_hd__ha_1 _749_ (.A(_274_),
    .B(_275_),
    .COUT(_276_),
    .SUM(_277_));
 sky130_fd_sc_hd__ha_1 _750_ (.A(net52),
    .B(net116),
    .COUT(_278_),
    .SUM(_279_));
 sky130_fd_sc_hd__ha_1 _751_ (.A(_280_),
    .B(_281_),
    .COUT(_282_),
    .SUM(_283_));
 sky130_fd_sc_hd__ha_1 _752_ (.A(net8),
    .B(net72),
    .COUT(_284_),
    .SUM(_285_));
 sky130_fd_sc_hd__ha_1 _753_ (.A(_286_),
    .B(_287_),
    .COUT(_288_),
    .SUM(_289_));
 sky130_fd_sc_hd__ha_1 _754_ (.A(net17),
    .B(net81),
    .COUT(_290_),
    .SUM(_291_));
 sky130_fd_sc_hd__ha_1 _755_ (.A(_292_),
    .B(_293_),
    .COUT(_294_),
    .SUM(_295_));
 sky130_fd_sc_hd__ha_1 _756_ (.A(net26),
    .B(net90),
    .COUT(_296_),
    .SUM(_297_));
 sky130_fd_sc_hd__ha_1 _757_ (.A(_298_),
    .B(_299_),
    .COUT(_300_),
    .SUM(_301_));
 sky130_fd_sc_hd__ha_1 _758_ (.A(net35),
    .B(net99),
    .COUT(_302_),
    .SUM(_303_));
 sky130_fd_sc_hd__ha_1 _759_ (.A(net7),
    .B(net71),
    .COUT(_304_),
    .SUM(_305_));
 sky130_fd_sc_hd__ha_1 _760_ (.A(net6),
    .B(net70),
    .COUT(_306_),
    .SUM(_307_));
 sky130_fd_sc_hd__ha_1 _761_ (.A(net5),
    .B(net69),
    .COUT(_308_),
    .SUM(_309_));
 sky130_fd_sc_hd__ha_1 _762_ (.A(net4),
    .B(net68),
    .COUT(_310_),
    .SUM(_311_));
 sky130_fd_sc_hd__ha_1 _763_ (.A(net3),
    .B(net67),
    .COUT(_312_),
    .SUM(_313_));
 sky130_fd_sc_hd__ha_1 _764_ (.A(net2),
    .B(net66),
    .COUT(_314_),
    .SUM(_315_));
 sky130_fd_sc_hd__ha_1 _765_ (.A(net64),
    .B(net128),
    .COUT(_316_),
    .SUM(_317_));
 sky130_fd_sc_hd__ha_1 _766_ (.A(net16),
    .B(net80),
    .COUT(_318_),
    .SUM(_319_));
 sky130_fd_sc_hd__ha_1 _767_ (.A(net15),
    .B(net79),
    .COUT(_320_),
    .SUM(_321_));
 sky130_fd_sc_hd__ha_1 _768_ (.A(net14),
    .B(net78),
    .COUT(_322_),
    .SUM(_323_));
 sky130_fd_sc_hd__ha_1 _769_ (.A(net13),
    .B(net77),
    .COUT(_324_),
    .SUM(_325_));
 sky130_fd_sc_hd__ha_1 _770_ (.A(net11),
    .B(net75),
    .COUT(_326_),
    .SUM(_327_));
 sky130_fd_sc_hd__ha_1 _771_ (.A(net10),
    .B(net74),
    .COUT(_328_),
    .SUM(_329_));
 sky130_fd_sc_hd__ha_1 _772_ (.A(net9),
    .B(net73),
    .COUT(_330_),
    .SUM(_331_));
 sky130_fd_sc_hd__ha_1 _773_ (.A(net25),
    .B(net89),
    .COUT(_332_),
    .SUM(_333_));
 sky130_fd_sc_hd__ha_1 _774_ (.A(net24),
    .B(net88),
    .COUT(_334_),
    .SUM(_335_));
 sky130_fd_sc_hd__ha_1 _775_ (.A(net22),
    .B(net86),
    .COUT(_336_),
    .SUM(_337_));
 sky130_fd_sc_hd__ha_1 _776_ (.A(net21),
    .B(net85),
    .COUT(_338_),
    .SUM(_339_));
 sky130_fd_sc_hd__ha_1 _777_ (.A(net20),
    .B(net84),
    .COUT(_340_),
    .SUM(_341_));
 sky130_fd_sc_hd__ha_1 _778_ (.A(net19),
    .B(net83),
    .COUT(_342_),
    .SUM(_343_));
 sky130_fd_sc_hd__ha_1 _779_ (.A(net18),
    .B(net82),
    .COUT(_344_),
    .SUM(_345_));
 sky130_fd_sc_hd__ha_1 _780_ (.A(net33),
    .B(net97),
    .COUT(_346_),
    .SUM(_347_));
 sky130_fd_sc_hd__ha_1 _781_ (.A(net32),
    .B(net96),
    .COUT(_348_),
    .SUM(_349_));
 sky130_fd_sc_hd__ha_1 _782_ (.A(net31),
    .B(net95),
    .COUT(_350_),
    .SUM(_351_));
 sky130_fd_sc_hd__ha_1 _783_ (.A(net30),
    .B(net94),
    .COUT(_352_),
    .SUM(_353_));
 sky130_fd_sc_hd__ha_1 _784_ (.A(net29),
    .B(net93),
    .COUT(_354_),
    .SUM(_355_));
 sky130_fd_sc_hd__ha_1 _785_ (.A(net28),
    .B(net92),
    .COUT(_356_),
    .SUM(_357_));
 sky130_fd_sc_hd__ha_1 _786_ (.A(net27),
    .B(net91),
    .COUT(_358_),
    .SUM(_359_));
 sky130_fd_sc_hd__ha_1 _787_ (.A(net42),
    .B(net106),
    .COUT(_360_),
    .SUM(_361_));
 sky130_fd_sc_hd__ha_1 _788_ (.A(net41),
    .B(net105),
    .COUT(_362_),
    .SUM(_363_));
 sky130_fd_sc_hd__ha_1 _789_ (.A(net40),
    .B(net104),
    .COUT(_364_),
    .SUM(_365_));
 sky130_fd_sc_hd__ha_1 _790_ (.A(net39),
    .B(net103),
    .COUT(_366_),
    .SUM(_367_));
 sky130_fd_sc_hd__ha_1 _791_ (.A(net38),
    .B(net102),
    .COUT(_368_),
    .SUM(_369_));
 sky130_fd_sc_hd__ha_1 _792_ (.A(net37),
    .B(net101),
    .COUT(_370_),
    .SUM(_371_));
 sky130_fd_sc_hd__ha_1 _793_ (.A(net36),
    .B(net100),
    .COUT(_372_),
    .SUM(_373_));
 sky130_fd_sc_hd__ha_1 _794_ (.A(net51),
    .B(net115),
    .COUT(_374_),
    .SUM(_375_));
 sky130_fd_sc_hd__ha_1 _795_ (.A(net50),
    .B(net114),
    .COUT(_376_),
    .SUM(_377_));
 sky130_fd_sc_hd__ha_1 _796_ (.A(net49),
    .B(net113),
    .COUT(_378_),
    .SUM(_379_));
 sky130_fd_sc_hd__ha_1 _797_ (.A(net48),
    .B(net112),
    .COUT(_380_),
    .SUM(_381_));
 sky130_fd_sc_hd__ha_1 _798_ (.A(net47),
    .B(net111),
    .COUT(_382_),
    .SUM(_383_));
 sky130_fd_sc_hd__ha_1 _799_ (.A(net46),
    .B(net110),
    .COUT(_384_),
    .SUM(_385_));
 sky130_fd_sc_hd__ha_1 _800_ (.A(net44),
    .B(net108),
    .COUT(_386_),
    .SUM(_387_));
 sky130_fd_sc_hd__ha_1 _801_ (.A(net60),
    .B(net124),
    .COUT(_388_),
    .SUM(_389_));
 sky130_fd_sc_hd__ha_1 _802_ (.A(net59),
    .B(net123),
    .COUT(_390_),
    .SUM(_391_));
 sky130_fd_sc_hd__ha_1 _803_ (.A(net58),
    .B(net122),
    .COUT(_392_),
    .SUM(_393_));
 sky130_fd_sc_hd__ha_1 _804_ (.A(net57),
    .B(net121),
    .COUT(_394_),
    .SUM(_395_));
 sky130_fd_sc_hd__ha_1 _805_ (.A(net55),
    .B(net119),
    .COUT(_396_),
    .SUM(_397_));
 sky130_fd_sc_hd__ha_1 _806_ (.A(net54),
    .B(net118),
    .COUT(_398_),
    .SUM(_399_));
 sky130_fd_sc_hd__ha_1 _807_ (.A(net53),
    .B(net117),
    .COUT(_400_),
    .SUM(_401_));
 sky130_fd_sc_hd__ha_1 _808_ (.A(_402_),
    .B(_403_),
    .COUT(_404_),
    .SUM(_405_));
 sky130_fd_sc_hd__ha_1 _809_ (.A(net63),
    .B(net127),
    .COUT(_406_),
    .SUM(_407_));
 sky130_fd_sc_hd__clkbuf_1 _810_ (.A(\first_block.full_adders[0].fa.sum ),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 _811_ (.A(\first_block.full_adders[1].fa.sum ),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 _812_ (.A(\first_block.full_adders[2].fa.sum ),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 _813_ (.A(\first_block.full_adders[3].fa.sum ),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 _814_ (.A(\first_block.full_adders[4].fa.sum ),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 _815_ (.A(\first_block.full_adders[5].fa.sum ),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 _816_ (.A(\first_block.full_adders[6].fa.sum ),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 _817_ (.A(\first_block.full_adders[7].fa.sum ),
    .X(net192));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_71 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(a[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(a[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(a[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(a[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(a[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(a[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(a[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(a[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(a[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(a[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(a[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(a[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(a[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(a[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(a[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(a[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(a[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(a[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(a[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(a[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(a[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(a[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(a[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(a[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(a[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(a[32]),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(a[33]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(a[34]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(a[35]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(a[36]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(a[37]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(a[38]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(a[39]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(a[3]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(a[40]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(a[41]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(a[42]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(a[43]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(a[44]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(a[45]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(a[46]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(a[47]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(a[48]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(a[49]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(a[4]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(a[50]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(a[51]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(a[52]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(a[53]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(a[54]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(a[55]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(a[56]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(a[57]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(a[58]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(a[59]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(a[5]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(a[60]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(a[61]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(a[62]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(a[63]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(a[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(a[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(a[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(a[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(b[0]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(b[10]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(b[11]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(b[12]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(b[13]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(b[14]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(b[15]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(b[16]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(b[17]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(b[18]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(b[19]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(b[1]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(b[20]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(b[21]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(b[22]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input80 (.A(b[23]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(b[24]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(b[25]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(b[26]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(b[27]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(b[28]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(b[29]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(b[2]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(b[30]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(b[31]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 input90 (.A(b[32]),
    .X(net90));
 sky130_fd_sc_hd__dlymetal6s2s_1 input91 (.A(b[33]),
    .X(net91));
 sky130_fd_sc_hd__dlymetal6s2s_1 input92 (.A(b[34]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(b[35]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 input94 (.A(b[36]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 input95 (.A(b[37]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 input96 (.A(b[38]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(b[39]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 input98 (.A(b[3]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 input99 (.A(b[40]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(b[41]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 input101 (.A(b[42]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 input102 (.A(b[43]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 input103 (.A(b[44]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 input104 (.A(b[45]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 input105 (.A(b[46]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 input106 (.A(b[47]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 input107 (.A(b[48]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 input108 (.A(b[49]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 input109 (.A(b[4]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 input110 (.A(b[50]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_1 input111 (.A(b[51]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 input112 (.A(b[52]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 input113 (.A(b[53]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 input114 (.A(b[54]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 input115 (.A(b[55]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_1 input116 (.A(b[56]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 input117 (.A(b[57]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_1 input118 (.A(b[58]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 input119 (.A(b[59]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 input120 (.A(b[5]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 input121 (.A(b[60]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 input122 (.A(b[61]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(b[62]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 input124 (.A(b[63]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 input125 (.A(b[6]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 input126 (.A(b[7]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 input127 (.A(b[8]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 input128 (.A(b[9]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 input129 (.A(cin),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 output130 (.A(net130),
    .X(cout));
 sky130_fd_sc_hd__clkbuf_1 output131 (.A(net131),
    .X(sum[0]));
 sky130_fd_sc_hd__clkbuf_1 output132 (.A(net132),
    .X(sum[10]));
 sky130_fd_sc_hd__clkbuf_1 output133 (.A(net133),
    .X(sum[11]));
 sky130_fd_sc_hd__clkbuf_1 output134 (.A(net134),
    .X(sum[12]));
 sky130_fd_sc_hd__clkbuf_1 output135 (.A(net135),
    .X(sum[13]));
 sky130_fd_sc_hd__clkbuf_1 output136 (.A(net136),
    .X(sum[14]));
 sky130_fd_sc_hd__clkbuf_1 output137 (.A(net137),
    .X(sum[15]));
 sky130_fd_sc_hd__clkbuf_1 output138 (.A(net138),
    .X(sum[16]));
 sky130_fd_sc_hd__clkbuf_1 output139 (.A(net139),
    .X(sum[17]));
 sky130_fd_sc_hd__clkbuf_1 output140 (.A(net140),
    .X(sum[18]));
 sky130_fd_sc_hd__clkbuf_1 output141 (.A(net141),
    .X(sum[19]));
 sky130_fd_sc_hd__clkbuf_1 output142 (.A(net142),
    .X(sum[1]));
 sky130_fd_sc_hd__clkbuf_1 output143 (.A(net143),
    .X(sum[20]));
 sky130_fd_sc_hd__clkbuf_1 output144 (.A(net144),
    .X(sum[21]));
 sky130_fd_sc_hd__clkbuf_1 output145 (.A(net145),
    .X(sum[22]));
 sky130_fd_sc_hd__clkbuf_1 output146 (.A(net146),
    .X(sum[23]));
 sky130_fd_sc_hd__clkbuf_1 output147 (.A(net147),
    .X(sum[24]));
 sky130_fd_sc_hd__clkbuf_1 output148 (.A(net148),
    .X(sum[25]));
 sky130_fd_sc_hd__clkbuf_1 output149 (.A(net149),
    .X(sum[26]));
 sky130_fd_sc_hd__clkbuf_1 output150 (.A(net150),
    .X(sum[27]));
 sky130_fd_sc_hd__clkbuf_1 output151 (.A(net151),
    .X(sum[28]));
 sky130_fd_sc_hd__clkbuf_1 output152 (.A(net152),
    .X(sum[29]));
 sky130_fd_sc_hd__clkbuf_1 output153 (.A(net153),
    .X(sum[2]));
 sky130_fd_sc_hd__clkbuf_1 output154 (.A(net154),
    .X(sum[30]));
 sky130_fd_sc_hd__clkbuf_1 output155 (.A(net155),
    .X(sum[31]));
 sky130_fd_sc_hd__clkbuf_1 output156 (.A(net156),
    .X(sum[32]));
 sky130_fd_sc_hd__clkbuf_1 output157 (.A(net157),
    .X(sum[33]));
 sky130_fd_sc_hd__clkbuf_1 output158 (.A(net158),
    .X(sum[34]));
 sky130_fd_sc_hd__clkbuf_1 output159 (.A(net159),
    .X(sum[35]));
 sky130_fd_sc_hd__clkbuf_1 output160 (.A(net160),
    .X(sum[36]));
 sky130_fd_sc_hd__clkbuf_1 output161 (.A(net161),
    .X(sum[37]));
 sky130_fd_sc_hd__clkbuf_1 output162 (.A(net162),
    .X(sum[38]));
 sky130_fd_sc_hd__clkbuf_1 output163 (.A(net163),
    .X(sum[39]));
 sky130_fd_sc_hd__clkbuf_1 output164 (.A(net164),
    .X(sum[3]));
 sky130_fd_sc_hd__clkbuf_1 output165 (.A(net165),
    .X(sum[40]));
 sky130_fd_sc_hd__clkbuf_1 output166 (.A(net166),
    .X(sum[41]));
 sky130_fd_sc_hd__clkbuf_1 output167 (.A(net167),
    .X(sum[42]));
 sky130_fd_sc_hd__clkbuf_1 output168 (.A(net168),
    .X(sum[43]));
 sky130_fd_sc_hd__clkbuf_1 output169 (.A(net169),
    .X(sum[44]));
 sky130_fd_sc_hd__clkbuf_1 output170 (.A(net170),
    .X(sum[45]));
 sky130_fd_sc_hd__clkbuf_1 output171 (.A(net171),
    .X(sum[46]));
 sky130_fd_sc_hd__clkbuf_1 output172 (.A(net172),
    .X(sum[47]));
 sky130_fd_sc_hd__clkbuf_1 output173 (.A(net173),
    .X(sum[48]));
 sky130_fd_sc_hd__clkbuf_1 output174 (.A(net174),
    .X(sum[49]));
 sky130_fd_sc_hd__clkbuf_1 output175 (.A(net175),
    .X(sum[4]));
 sky130_fd_sc_hd__clkbuf_1 output176 (.A(net176),
    .X(sum[50]));
 sky130_fd_sc_hd__clkbuf_1 output177 (.A(net177),
    .X(sum[51]));
 sky130_fd_sc_hd__clkbuf_1 output178 (.A(net178),
    .X(sum[52]));
 sky130_fd_sc_hd__clkbuf_1 output179 (.A(net179),
    .X(sum[53]));
 sky130_fd_sc_hd__clkbuf_1 output180 (.A(net180),
    .X(sum[54]));
 sky130_fd_sc_hd__clkbuf_1 output181 (.A(net181),
    .X(sum[55]));
 sky130_fd_sc_hd__clkbuf_1 output182 (.A(net182),
    .X(sum[56]));
 sky130_fd_sc_hd__clkbuf_1 output183 (.A(net183),
    .X(sum[57]));
 sky130_fd_sc_hd__clkbuf_1 output184 (.A(net184),
    .X(sum[58]));
 sky130_fd_sc_hd__clkbuf_1 output185 (.A(net185),
    .X(sum[59]));
 sky130_fd_sc_hd__clkbuf_1 output186 (.A(net186),
    .X(sum[5]));
 sky130_fd_sc_hd__clkbuf_1 output187 (.A(net187),
    .X(sum[60]));
 sky130_fd_sc_hd__clkbuf_1 output188 (.A(net188),
    .X(sum[61]));
 sky130_fd_sc_hd__clkbuf_1 output189 (.A(net189),
    .X(sum[62]));
 sky130_fd_sc_hd__clkbuf_1 output190 (.A(net190),
    .X(sum[63]));
 sky130_fd_sc_hd__clkbuf_1 output191 (.A(net191),
    .X(sum[6]));
 sky130_fd_sc_hd__clkbuf_1 output192 (.A(net192),
    .X(sum[7]));
 sky130_fd_sc_hd__clkbuf_1 output193 (.A(net193),
    .X(sum[8]));
 sky130_fd_sc_hd__clkbuf_1 output194 (.A(net194),
    .X(sum[9]));
 sky130_fd_sc_hd__fill_1 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_90 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_81 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_147 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_120 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_22 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_21 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_72 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_163 ();
endmodule
