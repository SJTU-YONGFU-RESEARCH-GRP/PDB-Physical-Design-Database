module loadable_updown_counter (clk,
    enable,
    load_en,
    overflow,
    rst_n,
    underflow,
    up_down,
    count,
    load_val);
 input clk;
 input enable;
 input load_en;
 output overflow;
 input rst_n;
 output underflow;
 input up_down;
 output [7:0] count;
 input [7:0] load_val;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 BUF_X2 _112_ (.A(net9),
    .Z(_043_));
 INV_X4 _113_ (.A(_043_),
    .ZN(_099_));
 BUF_X2 _114_ (.A(rst_n),
    .Z(_044_));
 CLKBUF_X2 _115_ (.A(net10),
    .Z(_045_));
 BUF_X4 _116_ (.A(load_en),
    .Z(_046_));
 MUX2_X1 _117_ (.A(_095_),
    .B(net1),
    .S(_046_),
    .Z(_047_));
 BUF_X1 _118_ (.A(enable),
    .Z(_048_));
 CLKBUF_X3 _119_ (.A(_048_),
    .Z(_049_));
 MUX2_X1 _120_ (.A(_045_),
    .B(_047_),
    .S(_049_),
    .Z(_050_));
 AND2_X1 _121_ (.A1(_044_),
    .A2(_050_),
    .ZN(_000_));
 NAND2_X1 _122_ (.A1(_046_),
    .A2(net2),
    .ZN(_051_));
 OAI21_X1 _123_ (.A(_051_),
    .B1(_098_),
    .B2(_046_),
    .ZN(_052_));
 MUX2_X1 _124_ (.A(net11),
    .B(_052_),
    .S(_049_),
    .Z(_053_));
 AND2_X1 _125_ (.A1(_044_),
    .A2(_053_),
    .ZN(_001_));
 BUF_X2 _126_ (.A(_103_),
    .Z(_054_));
 XNOR2_X1 _127_ (.A(_054_),
    .B(_097_),
    .ZN(_055_));
 INV_X2 _128_ (.A(_046_),
    .ZN(_056_));
 MUX2_X1 _129_ (.A(net3),
    .B(_055_),
    .S(_056_),
    .Z(_057_));
 MUX2_X1 _130_ (.A(net12),
    .B(_057_),
    .S(_048_),
    .Z(_058_));
 AND2_X1 _131_ (.A1(_044_),
    .A2(_058_),
    .ZN(_002_));
 OAI21_X1 _132_ (.A(_044_),
    .B1(net13),
    .B2(_049_),
    .ZN(_059_));
 AND2_X1 _133_ (.A1(_046_),
    .A2(net4),
    .ZN(_060_));
 INV_X1 _134_ (.A(_107_),
    .ZN(_061_));
 BUF_X4 _135_ (.A(_102_),
    .Z(_062_));
 INV_X1 _136_ (.A(_062_),
    .ZN(_063_));
 AOI21_X1 _137_ (.A(_100_),
    .B1(_101_),
    .B2(_045_),
    .ZN(_064_));
 INV_X1 _138_ (.A(_054_),
    .ZN(_065_));
 OAI21_X1 _139_ (.A(_063_),
    .B1(_064_),
    .B2(_065_),
    .ZN(_066_));
 XNOR2_X1 _140_ (.A(_061_),
    .B(_066_),
    .ZN(_067_));
 AOI21_X1 _141_ (.A(_060_),
    .B1(_067_),
    .B2(_056_),
    .ZN(_068_));
 AOI21_X1 _142_ (.A(_059_),
    .B1(_068_),
    .B2(_049_),
    .ZN(_003_));
 OAI21_X1 _143_ (.A(_044_),
    .B1(net14),
    .B2(_049_),
    .ZN(_069_));
 INV_X1 _144_ (.A(_106_),
    .ZN(_070_));
 BUF_X4 _145_ (.A(_105_),
    .Z(_071_));
 NOR2_X1 _146_ (.A1(_046_),
    .A2(_071_),
    .ZN(_072_));
 INV_X1 _147_ (.A(_097_),
    .ZN(_073_));
 AOI21_X2 _148_ (.A(_062_),
    .B1(_073_),
    .B2(_054_),
    .ZN(_074_));
 OAI211_X2 _149_ (.A(_070_),
    .B(_072_),
    .C1(_074_),
    .C2(_061_),
    .ZN(_075_));
 NAND2_X1 _150_ (.A1(_056_),
    .A2(_071_),
    .ZN(_076_));
 OAI21_X1 _151_ (.A(_063_),
    .B1(_097_),
    .B2(_065_),
    .ZN(_077_));
 AOI21_X1 _152_ (.A(_106_),
    .B1(_077_),
    .B2(_107_),
    .ZN(_078_));
 OAI221_X1 _153_ (.A(_075_),
    .B1(_076_),
    .B2(_078_),
    .C1(_056_),
    .C2(net5),
    .ZN(_079_));
 AOI21_X1 _154_ (.A(_069_),
    .B1(_079_),
    .B2(_049_),
    .ZN(_004_));
 OAI21_X1 _155_ (.A(_044_),
    .B1(net15),
    .B2(_049_),
    .ZN(_080_));
 AND2_X1 _156_ (.A1(_046_),
    .A2(net6),
    .ZN(_081_));
 AOI21_X1 _157_ (.A(_104_),
    .B1(_106_),
    .B2(_071_),
    .ZN(_082_));
 AOI211_X2 _158_ (.A(_100_),
    .B(_062_),
    .C1(_045_),
    .C2(_101_),
    .ZN(_083_));
 OAI211_X2 _159_ (.A(_107_),
    .B(_071_),
    .C1(_062_),
    .C2(_054_),
    .ZN(_084_));
 OAI21_X2 _160_ (.A(_082_),
    .B1(_083_),
    .B2(_084_),
    .ZN(_085_));
 XOR2_X1 _161_ (.A(_109_),
    .B(_085_),
    .Z(_086_));
 AOI21_X1 _162_ (.A(_081_),
    .B1(_086_),
    .B2(_056_),
    .ZN(_087_));
 AOI21_X1 _163_ (.A(_080_),
    .B1(_087_),
    .B2(_049_),
    .ZN(_005_));
 BUF_X2 _164_ (.A(_111_),
    .Z(_088_));
 NAND2_X1 _165_ (.A1(_056_),
    .A2(_048_),
    .ZN(_008_));
 OR3_X1 _166_ (.A1(_088_),
    .A2(_108_),
    .A3(_008_),
    .ZN(_009_));
 OAI21_X1 _167_ (.A(_109_),
    .B1(_104_),
    .B2(_071_),
    .ZN(_010_));
 INV_X1 _168_ (.A(_010_),
    .ZN(_011_));
 NOR2_X1 _169_ (.A1(_104_),
    .A2(_106_),
    .ZN(_012_));
 OAI21_X1 _170_ (.A(_012_),
    .B1(_074_),
    .B2(_061_),
    .ZN(_013_));
 AOI21_X1 _171_ (.A(_009_),
    .B1(_011_),
    .B2(_013_),
    .ZN(_014_));
 AND2_X1 _172_ (.A1(_056_),
    .A2(_048_),
    .ZN(_015_));
 AND4_X1 _173_ (.A1(_088_),
    .A2(_015_),
    .A3(_013_),
    .A4(_011_),
    .ZN(_016_));
 NAND2_X1 _174_ (.A1(_046_),
    .A2(_048_),
    .ZN(_017_));
 NAND2_X1 _175_ (.A1(_088_),
    .A2(_108_),
    .ZN(_018_));
 OAI22_X1 _176_ (.A1(net7),
    .A2(_017_),
    .B1(_008_),
    .B2(_018_),
    .ZN(_019_));
 OAI21_X1 _177_ (.A(_044_),
    .B1(net16),
    .B2(_049_),
    .ZN(_020_));
 NOR4_X1 _178_ (.A1(_014_),
    .A2(_016_),
    .A3(_019_),
    .A4(_020_),
    .ZN(_006_));
 INV_X1 _179_ (.A(net17),
    .ZN(_021_));
 INV_X1 _180_ (.A(net8),
    .ZN(_022_));
 OAI22_X1 _181_ (.A1(_049_),
    .A2(_021_),
    .B1(_022_),
    .B2(_017_),
    .ZN(_023_));
 NAND2_X1 _182_ (.A1(_044_),
    .A2(_023_),
    .ZN(_024_));
 AND3_X1 _183_ (.A1(_021_),
    .A2(_044_),
    .A3(_015_),
    .ZN(_025_));
 AOI21_X1 _184_ (.A(_110_),
    .B1(_108_),
    .B2(_088_),
    .ZN(_026_));
 OR2_X1 _185_ (.A1(_099_),
    .A2(_026_),
    .ZN(_027_));
 NAND2_X1 _186_ (.A1(_099_),
    .A2(_026_),
    .ZN(_028_));
 INV_X1 _187_ (.A(_110_),
    .ZN(_029_));
 OAI21_X1 _188_ (.A(_088_),
    .B1(_108_),
    .B2(_109_),
    .ZN(_030_));
 NAND2_X1 _189_ (.A1(_029_),
    .A2(_030_),
    .ZN(_031_));
 OAI221_X2 _190_ (.A(_027_),
    .B1(_028_),
    .B2(_085_),
    .C1(_031_),
    .C2(_043_),
    .ZN(_032_));
 AND4_X1 _191_ (.A1(_043_),
    .A2(_109_),
    .A3(_088_),
    .A4(_085_),
    .ZN(_033_));
 OAI21_X1 _192_ (.A(_025_),
    .B1(_032_),
    .B2(_033_),
    .ZN(_034_));
 NAND3_X1 _193_ (.A1(_056_),
    .A2(net17),
    .A3(_044_),
    .ZN(_035_));
 OR3_X1 _194_ (.A1(_033_),
    .A2(_032_),
    .A3(_035_),
    .ZN(_036_));
 NAND3_X1 _195_ (.A1(_024_),
    .A2(_034_),
    .A3(_036_),
    .ZN(_007_));
 NAND4_X1 _196_ (.A1(net15),
    .A2(net14),
    .A3(net16),
    .A4(net17),
    .ZN(_037_));
 NAND2_X1 _197_ (.A1(net11),
    .A2(_043_),
    .ZN(_038_));
 NAND3_X1 _198_ (.A1(_045_),
    .A2(net12),
    .A3(net13),
    .ZN(_039_));
 NOR4_X2 _199_ (.A1(_008_),
    .A2(_037_),
    .A3(_038_),
    .A4(_039_),
    .ZN(net18));
 NOR4_X1 _200_ (.A1(net15),
    .A2(net14),
    .A3(net16),
    .A4(net17),
    .ZN(_040_));
 NOR2_X1 _201_ (.A1(net11),
    .A2(_043_),
    .ZN(_041_));
 NAND3_X1 _202_ (.A1(_015_),
    .A2(_040_),
    .A3(_041_),
    .ZN(_042_));
 NOR4_X1 _203_ (.A1(_045_),
    .A2(net12),
    .A3(net13),
    .A4(_042_),
    .ZN(net19));
 FA_X1 _204_ (.A(_095_),
    .B(_096_),
    .CI(net9),
    .CO(_097_),
    .S(_098_));
 HA_X1 _205_ (.A(net11),
    .B(_099_),
    .CO(_100_),
    .S(_101_));
 HA_X1 _206_ (.A(net12),
    .B(_099_),
    .CO(_102_),
    .S(_103_));
 HA_X1 _207_ (.A(net14),
    .B(_099_),
    .CO(_104_),
    .S(_105_));
 HA_X1 _208_ (.A(net13),
    .B(_099_),
    .CO(_106_),
    .S(_107_));
 HA_X1 _209_ (.A(net15),
    .B(_099_),
    .CO(_108_),
    .S(_109_));
 HA_X1 _210_ (.A(net16),
    .B(_099_),
    .CO(_110_),
    .S(_111_));
 DFF_X1 \count[0]$_SDFFE_PN0P_  (.D(_000_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net10),
    .QN(_095_));
 DFF_X2 \count[1]$_SDFFE_PN0P_  (.D(_001_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net11),
    .QN(_096_));
 DFF_X2 \count[2]$_SDFFE_PN0P_  (.D(_002_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net12),
    .QN(_094_));
 DFF_X2 \count[3]$_SDFFE_PN0P_  (.D(_003_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net13),
    .QN(_093_));
 DFF_X2 \count[4]$_SDFFE_PN0P_  (.D(_004_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net14),
    .QN(_092_));
 DFF_X2 \count[5]$_SDFFE_PN0P_  (.D(_005_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net15),
    .QN(_091_));
 DFF_X2 \count[6]$_SDFFE_PN0P_  (.D(_006_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net16),
    .QN(_090_));
 DFF_X2 \count[7]$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net17),
    .QN(_089_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_81 ();
 BUF_X1 input1 (.A(load_val[0]),
    .Z(net1));
 BUF_X1 input2 (.A(load_val[1]),
    .Z(net2));
 BUF_X1 input3 (.A(load_val[2]),
    .Z(net3));
 BUF_X1 input4 (.A(load_val[3]),
    .Z(net4));
 BUF_X1 input5 (.A(load_val[4]),
    .Z(net5));
 BUF_X1 input6 (.A(load_val[5]),
    .Z(net6));
 BUF_X1 input7 (.A(load_val[6]),
    .Z(net7));
 BUF_X1 input8 (.A(load_val[7]),
    .Z(net8));
 BUF_X1 input9 (.A(up_down),
    .Z(net9));
 BUF_X1 output10 (.A(net10),
    .Z(count[0]));
 BUF_X1 output11 (.A(net11),
    .Z(count[1]));
 BUF_X1 output12 (.A(net12),
    .Z(count[2]));
 BUF_X1 output13 (.A(net13),
    .Z(count[3]));
 BUF_X1 output14 (.A(net14),
    .Z(count[4]));
 BUF_X1 output15 (.A(net15),
    .Z(count[5]));
 BUF_X1 output16 (.A(net16),
    .Z(count[6]));
 BUF_X1 output17 (.A(net17),
    .Z(count[7]));
 BUF_X1 output18 (.A(net18),
    .Z(overflow));
 BUF_X1 output19 (.A(net19),
    .Z(underflow));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 CLKBUF_X1 clkload0 (.A(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X16 FILLER_0_97 ();
 FILLCELL_X8 FILLER_0_113 ();
 FILLCELL_X2 FILLER_0_121 ();
 FILLCELL_X1 FILLER_0_123 ();
 FILLCELL_X8 FILLER_0_139 ();
 FILLCELL_X4 FILLER_0_147 ();
 FILLCELL_X4 FILLER_0_166 ();
 FILLCELL_X32 FILLER_0_177 ();
 FILLCELL_X32 FILLER_0_209 ();
 FILLCELL_X32 FILLER_0_241 ();
 FILLCELL_X16 FILLER_0_273 ();
 FILLCELL_X8 FILLER_0_289 ();
 FILLCELL_X4 FILLER_0_297 ();
 FILLCELL_X1 FILLER_0_301 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X16 FILLER_1_97 ();
 FILLCELL_X4 FILLER_1_113 ();
 FILLCELL_X2 FILLER_1_121 ();
 FILLCELL_X1 FILLER_1_123 ();
 FILLCELL_X1 FILLER_1_131 ();
 FILLCELL_X8 FILLER_1_136 ();
 FILLCELL_X2 FILLER_1_144 ();
 FILLCELL_X32 FILLER_1_166 ();
 FILLCELL_X32 FILLER_1_198 ();
 FILLCELL_X32 FILLER_1_230 ();
 FILLCELL_X32 FILLER_1_262 ();
 FILLCELL_X8 FILLER_1_294 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X16 FILLER_2_97 ();
 FILLCELL_X1 FILLER_2_113 ();
 FILLCELL_X2 FILLER_2_142 ();
 FILLCELL_X2 FILLER_2_148 ();
 FILLCELL_X1 FILLER_2_150 ();
 FILLCELL_X32 FILLER_2_158 ();
 FILLCELL_X32 FILLER_2_190 ();
 FILLCELL_X32 FILLER_2_222 ();
 FILLCELL_X32 FILLER_2_254 ();
 FILLCELL_X16 FILLER_2_286 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X8 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_156 ();
 FILLCELL_X32 FILLER_3_188 ();
 FILLCELL_X32 FILLER_3_220 ();
 FILLCELL_X32 FILLER_3_252 ();
 FILLCELL_X16 FILLER_3_284 ();
 FILLCELL_X2 FILLER_3_300 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X16 FILLER_4_129 ();
 FILLCELL_X8 FILLER_4_145 ();
 FILLCELL_X2 FILLER_4_153 ();
 FILLCELL_X32 FILLER_4_159 ();
 FILLCELL_X32 FILLER_4_191 ();
 FILLCELL_X32 FILLER_4_223 ();
 FILLCELL_X32 FILLER_4_255 ();
 FILLCELL_X8 FILLER_4_287 ();
 FILLCELL_X4 FILLER_4_295 ();
 FILLCELL_X2 FILLER_4_299 ();
 FILLCELL_X1 FILLER_4_301 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X4 FILLER_5_129 ();
 FILLCELL_X1 FILLER_5_133 ();
 FILLCELL_X32 FILLER_5_138 ();
 FILLCELL_X32 FILLER_5_170 ();
 FILLCELL_X32 FILLER_5_202 ();
 FILLCELL_X32 FILLER_5_234 ();
 FILLCELL_X32 FILLER_5_266 ();
 FILLCELL_X4 FILLER_5_298 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X16 FILLER_6_129 ();
 FILLCELL_X8 FILLER_6_145 ();
 FILLCELL_X4 FILLER_6_153 ();
 FILLCELL_X1 FILLER_6_157 ();
 FILLCELL_X32 FILLER_6_168 ();
 FILLCELL_X32 FILLER_6_200 ();
 FILLCELL_X32 FILLER_6_232 ();
 FILLCELL_X32 FILLER_6_264 ();
 FILLCELL_X4 FILLER_6_296 ();
 FILLCELL_X2 FILLER_6_300 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X16 FILLER_7_97 ();
 FILLCELL_X8 FILLER_7_113 ();
 FILLCELL_X2 FILLER_7_121 ();
 FILLCELL_X1 FILLER_7_123 ();
 FILLCELL_X2 FILLER_7_147 ();
 FILLCELL_X1 FILLER_7_149 ();
 FILLCELL_X2 FILLER_7_155 ();
 FILLCELL_X4 FILLER_7_161 ();
 FILLCELL_X2 FILLER_7_165 ();
 FILLCELL_X1 FILLER_7_167 ();
 FILLCELL_X32 FILLER_7_185 ();
 FILLCELL_X32 FILLER_7_217 ();
 FILLCELL_X32 FILLER_7_249 ();
 FILLCELL_X16 FILLER_7_281 ();
 FILLCELL_X4 FILLER_7_297 ();
 FILLCELL_X1 FILLER_7_301 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X16 FILLER_8_97 ();
 FILLCELL_X8 FILLER_8_113 ();
 FILLCELL_X1 FILLER_8_121 ();
 FILLCELL_X2 FILLER_8_129 ();
 FILLCELL_X1 FILLER_8_131 ();
 FILLCELL_X2 FILLER_8_139 ();
 FILLCELL_X2 FILLER_8_147 ();
 FILLCELL_X1 FILLER_8_149 ();
 FILLCELL_X1 FILLER_8_154 ();
 FILLCELL_X8 FILLER_8_157 ();
 FILLCELL_X1 FILLER_8_165 ();
 FILLCELL_X32 FILLER_8_179 ();
 FILLCELL_X32 FILLER_8_211 ();
 FILLCELL_X32 FILLER_8_243 ();
 FILLCELL_X16 FILLER_8_275 ();
 FILLCELL_X8 FILLER_8_291 ();
 FILLCELL_X2 FILLER_8_299 ();
 FILLCELL_X1 FILLER_8_301 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X16 FILLER_9_97 ();
 FILLCELL_X8 FILLER_9_113 ();
 FILLCELL_X2 FILLER_9_121 ();
 FILLCELL_X1 FILLER_9_123 ();
 FILLCELL_X4 FILLER_9_128 ();
 FILLCELL_X2 FILLER_9_132 ();
 FILLCELL_X8 FILLER_9_139 ();
 FILLCELL_X8 FILLER_9_159 ();
 FILLCELL_X4 FILLER_9_167 ();
 FILLCELL_X2 FILLER_9_171 ();
 FILLCELL_X1 FILLER_9_173 ();
 FILLCELL_X32 FILLER_9_179 ();
 FILLCELL_X32 FILLER_9_211 ();
 FILLCELL_X32 FILLER_9_243 ();
 FILLCELL_X16 FILLER_9_275 ();
 FILLCELL_X8 FILLER_9_291 ();
 FILLCELL_X2 FILLER_9_299 ();
 FILLCELL_X1 FILLER_9_301 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X16 FILLER_10_97 ();
 FILLCELL_X8 FILLER_10_113 ();
 FILLCELL_X1 FILLER_10_121 ();
 FILLCELL_X2 FILLER_10_126 ();
 FILLCELL_X8 FILLER_10_137 ();
 FILLCELL_X1 FILLER_10_145 ();
 FILLCELL_X32 FILLER_10_159 ();
 FILLCELL_X32 FILLER_10_191 ();
 FILLCELL_X32 FILLER_10_223 ();
 FILLCELL_X32 FILLER_10_255 ();
 FILLCELL_X8 FILLER_10_287 ();
 FILLCELL_X4 FILLER_10_295 ();
 FILLCELL_X2 FILLER_10_299 ();
 FILLCELL_X1 FILLER_10_301 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X8 FILLER_11_97 ();
 FILLCELL_X4 FILLER_11_105 ();
 FILLCELL_X2 FILLER_11_109 ();
 FILLCELL_X4 FILLER_11_130 ();
 FILLCELL_X2 FILLER_11_134 ();
 FILLCELL_X4 FILLER_11_139 ();
 FILLCELL_X2 FILLER_11_143 ();
 FILLCELL_X1 FILLER_11_145 ();
 FILLCELL_X4 FILLER_11_149 ();
 FILLCELL_X2 FILLER_11_155 ();
 FILLCELL_X4 FILLER_11_166 ();
 FILLCELL_X2 FILLER_11_170 ();
 FILLCELL_X32 FILLER_11_179 ();
 FILLCELL_X32 FILLER_11_211 ();
 FILLCELL_X32 FILLER_11_243 ();
 FILLCELL_X16 FILLER_11_275 ();
 FILLCELL_X8 FILLER_11_291 ();
 FILLCELL_X2 FILLER_11_299 ();
 FILLCELL_X1 FILLER_11_301 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X8 FILLER_12_129 ();
 FILLCELL_X2 FILLER_12_137 ();
 FILLCELL_X2 FILLER_12_169 ();
 FILLCELL_X32 FILLER_12_178 ();
 FILLCELL_X32 FILLER_12_210 ();
 FILLCELL_X32 FILLER_12_242 ();
 FILLCELL_X16 FILLER_12_274 ();
 FILLCELL_X8 FILLER_12_290 ();
 FILLCELL_X4 FILLER_12_298 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X16 FILLER_13_129 ();
 FILLCELL_X8 FILLER_13_148 ();
 FILLCELL_X2 FILLER_13_156 ();
 FILLCELL_X4 FILLER_13_165 ();
 FILLCELL_X32 FILLER_13_183 ();
 FILLCELL_X32 FILLER_13_215 ();
 FILLCELL_X32 FILLER_13_247 ();
 FILLCELL_X16 FILLER_13_279 ();
 FILLCELL_X4 FILLER_13_295 ();
 FILLCELL_X2 FILLER_13_299 ();
 FILLCELL_X1 FILLER_13_301 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X16 FILLER_14_97 ();
 FILLCELL_X4 FILLER_14_113 ();
 FILLCELL_X1 FILLER_14_117 ();
 FILLCELL_X1 FILLER_14_122 ();
 FILLCELL_X8 FILLER_14_138 ();
 FILLCELL_X8 FILLER_14_152 ();
 FILLCELL_X2 FILLER_14_160 ();
 FILLCELL_X32 FILLER_14_172 ();
 FILLCELL_X32 FILLER_14_204 ();
 FILLCELL_X32 FILLER_14_236 ();
 FILLCELL_X32 FILLER_14_268 ();
 FILLCELL_X2 FILLER_14_300 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X16 FILLER_15_97 ();
 FILLCELL_X4 FILLER_15_113 ();
 FILLCELL_X2 FILLER_15_117 ();
 FILLCELL_X8 FILLER_15_138 ();
 FILLCELL_X4 FILLER_15_146 ();
 FILLCELL_X2 FILLER_15_150 ();
 FILLCELL_X1 FILLER_15_152 ();
 FILLCELL_X4 FILLER_15_156 ();
 FILLCELL_X1 FILLER_15_160 ();
 FILLCELL_X32 FILLER_15_163 ();
 FILLCELL_X32 FILLER_15_195 ();
 FILLCELL_X32 FILLER_15_227 ();
 FILLCELL_X32 FILLER_15_259 ();
 FILLCELL_X8 FILLER_15_291 ();
 FILLCELL_X2 FILLER_15_299 ();
 FILLCELL_X1 FILLER_15_301 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X1 FILLER_16_129 ();
 FILLCELL_X8 FILLER_16_134 ();
 FILLCELL_X1 FILLER_16_142 ();
 FILLCELL_X1 FILLER_16_152 ();
 FILLCELL_X16 FILLER_16_156 ();
 FILLCELL_X8 FILLER_16_172 ();
 FILLCELL_X4 FILLER_16_180 ();
 FILLCELL_X32 FILLER_16_188 ();
 FILLCELL_X32 FILLER_16_220 ();
 FILLCELL_X32 FILLER_16_252 ();
 FILLCELL_X16 FILLER_16_284 ();
 FILLCELL_X2 FILLER_16_300 ();
 FILLCELL_X16 FILLER_17_1 ();
 FILLCELL_X8 FILLER_17_17 ();
 FILLCELL_X2 FILLER_17_25 ();
 FILLCELL_X32 FILLER_17_30 ();
 FILLCELL_X32 FILLER_17_62 ();
 FILLCELL_X8 FILLER_17_94 ();
 FILLCELL_X2 FILLER_17_102 ();
 FILLCELL_X1 FILLER_17_104 ();
 FILLCELL_X16 FILLER_17_108 ();
 FILLCELL_X1 FILLER_17_124 ();
 FILLCELL_X4 FILLER_17_129 ();
 FILLCELL_X8 FILLER_17_170 ();
 FILLCELL_X2 FILLER_17_178 ();
 FILLCELL_X32 FILLER_17_198 ();
 FILLCELL_X32 FILLER_17_230 ();
 FILLCELL_X32 FILLER_17_262 ();
 FILLCELL_X8 FILLER_17_294 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X16 FILLER_18_97 ();
 FILLCELL_X2 FILLER_18_113 ();
 FILLCELL_X1 FILLER_18_124 ();
 FILLCELL_X16 FILLER_18_132 ();
 FILLCELL_X2 FILLER_18_148 ();
 FILLCELL_X1 FILLER_18_158 ();
 FILLCELL_X1 FILLER_18_163 ();
 FILLCELL_X1 FILLER_18_174 ();
 FILLCELL_X32 FILLER_18_193 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X8 FILLER_18_257 ();
 FILLCELL_X32 FILLER_18_268 ();
 FILLCELL_X2 FILLER_18_300 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X16 FILLER_19_97 ();
 FILLCELL_X1 FILLER_19_113 ();
 FILLCELL_X8 FILLER_19_126 ();
 FILLCELL_X4 FILLER_19_134 ();
 FILLCELL_X2 FILLER_19_138 ();
 FILLCELL_X16 FILLER_19_162 ();
 FILLCELL_X2 FILLER_19_178 ();
 FILLCELL_X1 FILLER_19_183 ();
 FILLCELL_X32 FILLER_19_186 ();
 FILLCELL_X32 FILLER_19_218 ();
 FILLCELL_X32 FILLER_19_250 ();
 FILLCELL_X16 FILLER_19_282 ();
 FILLCELL_X4 FILLER_19_298 ();
 FILLCELL_X4 FILLER_20_1 ();
 FILLCELL_X1 FILLER_20_5 ();
 FILLCELL_X32 FILLER_20_9 ();
 FILLCELL_X32 FILLER_20_41 ();
 FILLCELL_X32 FILLER_20_73 ();
 FILLCELL_X4 FILLER_20_105 ();
 FILLCELL_X2 FILLER_20_109 ();
 FILLCELL_X32 FILLER_20_130 ();
 FILLCELL_X32 FILLER_20_162 ();
 FILLCELL_X32 FILLER_20_194 ();
 FILLCELL_X32 FILLER_20_226 ();
 FILLCELL_X4 FILLER_20_258 ();
 FILLCELL_X1 FILLER_20_262 ();
 FILLCELL_X32 FILLER_20_266 ();
 FILLCELL_X4 FILLER_20_298 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X8 FILLER_21_129 ();
 FILLCELL_X2 FILLER_21_137 ();
 FILLCELL_X1 FILLER_21_139 ();
 FILLCELL_X32 FILLER_21_159 ();
 FILLCELL_X32 FILLER_21_191 ();
 FILLCELL_X32 FILLER_21_223 ();
 FILLCELL_X32 FILLER_21_255 ();
 FILLCELL_X8 FILLER_21_287 ();
 FILLCELL_X4 FILLER_21_295 ();
 FILLCELL_X2 FILLER_21_299 ();
 FILLCELL_X1 FILLER_21_301 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X16 FILLER_22_129 ();
 FILLCELL_X4 FILLER_22_145 ();
 FILLCELL_X32 FILLER_22_168 ();
 FILLCELL_X32 FILLER_22_200 ();
 FILLCELL_X32 FILLER_22_232 ();
 FILLCELL_X32 FILLER_22_264 ();
 FILLCELL_X4 FILLER_22_296 ();
 FILLCELL_X2 FILLER_22_300 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X16 FILLER_23_97 ();
 FILLCELL_X8 FILLER_23_113 ();
 FILLCELL_X2 FILLER_23_121 ();
 FILLCELL_X32 FILLER_23_125 ();
 FILLCELL_X32 FILLER_23_157 ();
 FILLCELL_X32 FILLER_23_189 ();
 FILLCELL_X32 FILLER_23_221 ();
 FILLCELL_X32 FILLER_23_253 ();
 FILLCELL_X16 FILLER_23_285 ();
 FILLCELL_X1 FILLER_23_301 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X32 FILLER_24_193 ();
 FILLCELL_X32 FILLER_24_225 ();
 FILLCELL_X32 FILLER_24_257 ();
 FILLCELL_X8 FILLER_24_289 ();
 FILLCELL_X4 FILLER_24_297 ();
 FILLCELL_X1 FILLER_24_301 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X32 FILLER_25_193 ();
 FILLCELL_X32 FILLER_25_225 ();
 FILLCELL_X32 FILLER_25_257 ();
 FILLCELL_X8 FILLER_25_289 ();
 FILLCELL_X4 FILLER_25_297 ();
 FILLCELL_X1 FILLER_25_301 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X32 FILLER_26_193 ();
 FILLCELL_X32 FILLER_26_225 ();
 FILLCELL_X32 FILLER_26_257 ();
 FILLCELL_X8 FILLER_26_289 ();
 FILLCELL_X4 FILLER_26_297 ();
 FILLCELL_X1 FILLER_26_301 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X32 FILLER_27_225 ();
 FILLCELL_X32 FILLER_27_257 ();
 FILLCELL_X8 FILLER_27_289 ();
 FILLCELL_X4 FILLER_27_297 ();
 FILLCELL_X1 FILLER_27_301 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X32 FILLER_28_225 ();
 FILLCELL_X32 FILLER_28_257 ();
 FILLCELL_X8 FILLER_28_289 ();
 FILLCELL_X4 FILLER_28_297 ();
 FILLCELL_X1 FILLER_28_301 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X32 FILLER_29_225 ();
 FILLCELL_X32 FILLER_29_257 ();
 FILLCELL_X8 FILLER_29_289 ();
 FILLCELL_X4 FILLER_29_297 ();
 FILLCELL_X1 FILLER_29_301 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X32 FILLER_30_225 ();
 FILLCELL_X32 FILLER_30_257 ();
 FILLCELL_X8 FILLER_30_289 ();
 FILLCELL_X4 FILLER_30_297 ();
 FILLCELL_X1 FILLER_30_301 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X32 FILLER_31_193 ();
 FILLCELL_X32 FILLER_31_225 ();
 FILLCELL_X32 FILLER_31_257 ();
 FILLCELL_X8 FILLER_31_289 ();
 FILLCELL_X4 FILLER_31_297 ();
 FILLCELL_X1 FILLER_31_301 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X32 FILLER_32_257 ();
 FILLCELL_X8 FILLER_32_289 ();
 FILLCELL_X4 FILLER_32_297 ();
 FILLCELL_X1 FILLER_32_301 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_225 ();
 FILLCELL_X32 FILLER_33_257 ();
 FILLCELL_X8 FILLER_33_289 ();
 FILLCELL_X4 FILLER_33_297 ();
 FILLCELL_X1 FILLER_33_301 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X32 FILLER_34_161 ();
 FILLCELL_X32 FILLER_34_193 ();
 FILLCELL_X32 FILLER_34_225 ();
 FILLCELL_X32 FILLER_34_257 ();
 FILLCELL_X8 FILLER_34_289 ();
 FILLCELL_X4 FILLER_34_297 ();
 FILLCELL_X1 FILLER_34_301 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X32 FILLER_35_161 ();
 FILLCELL_X32 FILLER_35_193 ();
 FILLCELL_X32 FILLER_35_225 ();
 FILLCELL_X32 FILLER_35_257 ();
 FILLCELL_X8 FILLER_35_289 ();
 FILLCELL_X4 FILLER_35_297 ();
 FILLCELL_X1 FILLER_35_301 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X32 FILLER_36_193 ();
 FILLCELL_X32 FILLER_36_225 ();
 FILLCELL_X32 FILLER_36_257 ();
 FILLCELL_X8 FILLER_36_289 ();
 FILLCELL_X4 FILLER_36_297 ();
 FILLCELL_X1 FILLER_36_301 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X32 FILLER_37_193 ();
 FILLCELL_X32 FILLER_37_225 ();
 FILLCELL_X32 FILLER_37_257 ();
 FILLCELL_X8 FILLER_37_289 ();
 FILLCELL_X4 FILLER_37_297 ();
 FILLCELL_X1 FILLER_37_301 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X32 FILLER_38_193 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X32 FILLER_38_257 ();
 FILLCELL_X8 FILLER_38_289 ();
 FILLCELL_X4 FILLER_38_297 ();
 FILLCELL_X1 FILLER_38_301 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X8 FILLER_39_129 ();
 FILLCELL_X4 FILLER_39_137 ();
 FILLCELL_X1 FILLER_39_141 ();
 FILLCELL_X4 FILLER_39_145 ();
 FILLCELL_X2 FILLER_39_149 ();
 FILLCELL_X1 FILLER_39_151 ();
 FILLCELL_X16 FILLER_39_155 ();
 FILLCELL_X32 FILLER_39_174 ();
 FILLCELL_X32 FILLER_39_206 ();
 FILLCELL_X32 FILLER_39_238 ();
 FILLCELL_X32 FILLER_39_270 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X16 FILLER_40_97 ();
 FILLCELL_X8 FILLER_40_113 ();
 FILLCELL_X2 FILLER_40_121 ();
 FILLCELL_X16 FILLER_40_126 ();
 FILLCELL_X8 FILLER_40_142 ();
 FILLCELL_X1 FILLER_40_150 ();
 FILLCELL_X16 FILLER_40_154 ();
 FILLCELL_X8 FILLER_40_170 ();
 FILLCELL_X1 FILLER_40_178 ();
 FILLCELL_X32 FILLER_40_182 ();
 FILLCELL_X32 FILLER_40_214 ();
 FILLCELL_X32 FILLER_40_246 ();
 FILLCELL_X16 FILLER_40_278 ();
 FILLCELL_X8 FILLER_40_294 ();
endmodule
