module async_fifo (almost_empty,
    almost_full,
    empty,
    full,
    pointer_wraparound_flag,
    rd_clk,
    rd_en,
    rd_rst_n,
    sync_error_flag,
    wr_clk,
    wr_en,
    wr_rst_n,
    rd_count,
    rd_data,
    wr_count,
    wr_data);
 output almost_empty;
 output almost_full;
 output empty;
 output full;
 output pointer_wraparound_flag;
 input rd_clk;
 input rd_en;
 input rd_rst_n;
 output sync_error_flag;
 input wr_clk;
 input wr_en;
 input wr_rst_n;
 output [4:0] rd_count;
 output [7:0] rd_data;
 output [4:0] wr_count;
 input [7:0] wr_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire \mem[0][0] ;
 wire \mem[0][1] ;
 wire \mem[0][2] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[10][0] ;
 wire \mem[10][1] ;
 wire \mem[10][2] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[11][0] ;
 wire \mem[11][1] ;
 wire \mem[11][2] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[12][0] ;
 wire \mem[12][1] ;
 wire \mem[12][2] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[13][0] ;
 wire \mem[13][1] ;
 wire \mem[13][2] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[14][0] ;
 wire \mem[14][1] ;
 wire \mem[14][2] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[15][0] ;
 wire \mem[15][1] ;
 wire \mem[15][2] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[1][0] ;
 wire \mem[1][1] ;
 wire \mem[1][2] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[2][0] ;
 wire \mem[2][1] ;
 wire \mem[2][2] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[3][0] ;
 wire \mem[3][1] ;
 wire \mem[3][2] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[4][0] ;
 wire \mem[4][1] ;
 wire \mem[4][2] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[5][0] ;
 wire \mem[5][1] ;
 wire \mem[5][2] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[6][0] ;
 wire \mem[6][1] ;
 wire \mem[6][2] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[7][0] ;
 wire \mem[7][1] ;
 wire \mem[7][2] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[8][0] ;
 wire \mem[8][1] ;
 wire \mem[8][2] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[9][0] ;
 wire \mem[9][1] ;
 wire \mem[9][2] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \rd_ptr_bin[0] ;
 wire \rd_ptr_bin[1] ;
 wire \rd_ptr_bin[2] ;
 wire \rd_ptr_bin[3] ;
 wire \rd_ptr_bin[4] ;
 wire \rd_ptr_gray[0] ;
 wire \rd_ptr_gray[1] ;
 wire \rd_ptr_gray[2] ;
 wire \rd_ptr_gray[3] ;
 wire \rd_ptr_gray_sync1[0] ;
 wire \rd_ptr_gray_sync1[1] ;
 wire \rd_ptr_gray_sync1[2] ;
 wire \rd_ptr_gray_sync1[3] ;
 wire \rd_ptr_gray_sync1[4] ;
 wire \rd_ptr_gray_sync2[0] ;
 wire \rd_ptr_gray_sync2[1] ;
 wire \rd_ptr_gray_sync2[2] ;
 wire \rd_ptr_gray_sync2[3] ;
 wire \rd_ptr_gray_sync2[4] ;
 wire \rd_ptr_sync[0] ;
 wire \rd_ptr_sync[1] ;
 wire \rd_ptr_sync[2] ;
 wire \rd_ptr_sync[3] ;
 wire \rd_ptr_sync[4] ;
 wire \wr_ptr_bin[0] ;
 wire \wr_ptr_bin[1] ;
 wire \wr_ptr_bin[2] ;
 wire \wr_ptr_bin[3] ;
 wire \wr_ptr_bin[4] ;
 wire \wr_ptr_gray[0] ;
 wire \wr_ptr_gray[1] ;
 wire \wr_ptr_gray[2] ;
 wire \wr_ptr_gray[3] ;
 wire \wr_ptr_gray_sync1[0] ;
 wire \wr_ptr_gray_sync1[1] ;
 wire \wr_ptr_gray_sync1[2] ;
 wire \wr_ptr_gray_sync1[3] ;
 wire \wr_ptr_gray_sync1[4] ;
 wire \wr_ptr_gray_sync2[0] ;
 wire \wr_ptr_gray_sync2[1] ;
 wire \wr_ptr_gray_sync2[2] ;
 wire \wr_ptr_gray_sync2[3] ;
 wire \wr_ptr_gray_sync2[4] ;
 wire \wr_ptr_sync[0] ;
 wire \wr_ptr_sync[1] ;
 wire \wr_ptr_sync[2] ;
 wire \wr_ptr_sync[3] ;
 wire \wr_ptr_sync[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;

 sky130_fd_sc_hd__inv_1 _338_ (.A(_306_),
    .Y(net20));
 sky130_fd_sc_hd__nand2_1 _339_ (.A(_299_),
    .B(_301_),
    .Y(_057_));
 sky130_fd_sc_hd__nand3_1 _340_ (.A(_296_),
    .B(_304_),
    .C(_306_),
    .Y(_058_));
 sky130_fd_sc_hd__nor2_1 _341_ (.A(_057_),
    .B(_058_),
    .Y(_000_));
 sky130_fd_sc_hd__a21o_1 _342_ (.A1(_304_),
    .A2(_290_),
    .B1(_303_),
    .X(_059_));
 sky130_fd_sc_hd__a21oi_1 _343_ (.A1(_296_),
    .A2(_059_),
    .B1(_295_),
    .Y(_060_));
 sky130_fd_sc_hd__xnor2_1 _344_ (.A(_299_),
    .B(_060_),
    .Y(net24));
 sky130_fd_sc_hd__xor2_1 _345_ (.A(_304_),
    .B(_290_),
    .X(net22));
 sky130_fd_sc_hd__nor2b_1 _346_ (.A(_308_),
    .B_N(_301_),
    .Y(_061_));
 sky130_fd_sc_hd__o21a_1 _347_ (.A1(_300_),
    .A2(_061_),
    .B1(_304_),
    .X(_062_));
 sky130_fd_sc_hd__o21ai_0 _348_ (.A1(_303_),
    .A2(_062_),
    .B1(_296_),
    .Y(_063_));
 sky130_fd_sc_hd__or3_1 _349_ (.A(_296_),
    .B(_303_),
    .C(_062_),
    .X(_064_));
 sky130_fd_sc_hd__and2_0 _350_ (.A(_063_),
    .B(_064_),
    .X(net23));
 sky130_fd_sc_hd__inv_1 _351_ (.A(_313_),
    .Y(net34));
 sky130_fd_sc_hd__inv_1 _352_ (.A(_319_),
    .Y(_065_));
 sky130_fd_sc_hd__nor2b_1 _353_ (.A(_314_),
    .B_N(_310_),
    .Y(_066_));
 sky130_fd_sc_hd__o21ai_0 _354_ (.A1(_316_),
    .A2(_066_),
    .B1(_320_),
    .Y(_067_));
 sky130_fd_sc_hd__a21boi_0 _355_ (.A1(_065_),
    .A2(_067_),
    .B1_N(_324_),
    .Y(_068_));
 sky130_fd_sc_hd__nor3b_1 _356_ (.A(_324_),
    .B(_319_),
    .C_N(_067_),
    .Y(_069_));
 sky130_fd_sc_hd__nor2_1 _357_ (.A(_068_),
    .B(_069_),
    .Y(net37));
 sky130_fd_sc_hd__a21o_1 _358_ (.A1(_320_),
    .A2(_293_),
    .B1(_319_),
    .X(_070_));
 sky130_fd_sc_hd__a21oi_1 _359_ (.A1(_324_),
    .A2(_070_),
    .B1(_323_),
    .Y(_071_));
 sky130_fd_sc_hd__xor2_1 _360_ (.A(_328_),
    .B(_071_),
    .X(_072_));
 sky130_fd_sc_hd__inv_1 _361_ (.A(_072_),
    .Y(net38));
 sky130_fd_sc_hd__nor4_1 _362_ (.A(\rd_ptr_sync[1] ),
    .B(\rd_ptr_sync[0] ),
    .C(\rd_ptr_sync[3] ),
    .D(\rd_ptr_sync[2] ),
    .Y(_073_));
 sky130_fd_sc_hd__clkbuf_4 _363_ (.A(\wr_ptr_bin[3] ),
    .X(_074_));
 sky130_fd_sc_hd__clkbuf_4 _364_ (.A(\wr_ptr_bin[2] ),
    .X(_075_));
 sky130_fd_sc_hd__or2_0 _365_ (.A(_074_),
    .B(_075_),
    .X(_076_));
 sky130_fd_sc_hd__buf_4 _366_ (.A(_076_),
    .X(_077_));
 sky130_fd_sc_hd__nand2_1 _367_ (.A(\wr_ptr_bin[4] ),
    .B(_330_),
    .Y(_078_));
 sky130_fd_sc_hd__nor3_1 _368_ (.A(_073_),
    .B(_077_),
    .C(_078_),
    .Y(_010_));
 sky130_fd_sc_hd__nand3_1 _369_ (.A(_310_),
    .B(_324_),
    .C(_320_),
    .Y(_079_));
 sky130_fd_sc_hd__nor3_1 _370_ (.A(net34),
    .B(_328_),
    .C(_079_),
    .Y(_001_));
 sky130_fd_sc_hd__inv_1 _371_ (.A(_075_),
    .Y(_321_));
 sky130_fd_sc_hd__nand2_4 _372_ (.A(_074_),
    .B(_321_),
    .Y(_080_));
 sky130_fd_sc_hd__nor2b_1 _373_ (.A(net18),
    .B_N(net13),
    .Y(_081_));
 sky130_fd_sc_hd__clkbuf_8 _374_ (.A(_081_),
    .X(_082_));
 sky130_fd_sc_hd__nand2_4 _375_ (.A(_331_),
    .B(_082_),
    .Y(_083_));
 sky130_fd_sc_hd__nor2_4 _376_ (.A(_080_),
    .B(_083_),
    .Y(_012_));
 sky130_fd_sc_hd__nand2_8 _377_ (.A(_333_),
    .B(_082_),
    .Y(_084_));
 sky130_fd_sc_hd__nor2_4 _378_ (.A(_080_),
    .B(_084_),
    .Y(_026_));
 sky130_fd_sc_hd__nand2_4 _379_ (.A(_330_),
    .B(_082_),
    .Y(_085_));
 sky130_fd_sc_hd__nor2_4 _380_ (.A(_080_),
    .B(_085_),
    .Y(_025_));
 sky130_fd_sc_hd__inv_1 _381_ (.A(_074_),
    .Y(_325_));
 sky130_fd_sc_hd__nand2_4 _382_ (.A(_325_),
    .B(_075_),
    .Y(_086_));
 sky130_fd_sc_hd__nand2_8 _383_ (.A(_335_),
    .B(_082_),
    .Y(_087_));
 sky130_fd_sc_hd__nor2_4 _384_ (.A(_086_),
    .B(_087_),
    .Y(_024_));
 sky130_fd_sc_hd__nand2_4 _385_ (.A(_074_),
    .B(_075_),
    .Y(_088_));
 sky130_fd_sc_hd__nor2_4 _386_ (.A(_087_),
    .B(_088_),
    .Y(_017_));
 sky130_fd_sc_hd__nor2_4 _387_ (.A(_083_),
    .B(_086_),
    .Y(_023_));
 sky130_fd_sc_hd__nor2_4 _388_ (.A(_083_),
    .B(_088_),
    .Y(_016_));
 sky130_fd_sc_hd__nor2_4 _389_ (.A(_084_),
    .B(_086_),
    .Y(_022_));
 sky130_fd_sc_hd__clkbuf_4 _390_ (.A(\rd_ptr_bin[2] ),
    .X(_089_));
 sky130_fd_sc_hd__inv_1 _391_ (.A(_089_),
    .Y(_302_));
 sky130_fd_sc_hd__buf_2 _392_ (.A(\rd_ptr_bin[3] ),
    .X(_090_));
 sky130_fd_sc_hd__inv_1 _393_ (.A(_090_),
    .Y(_294_));
 sky130_fd_sc_hd__nor2_4 _394_ (.A(_085_),
    .B(_086_),
    .Y(_021_));
 sky130_fd_sc_hd__nor2_4 _395_ (.A(_077_),
    .B(_087_),
    .Y(_020_));
 sky130_fd_sc_hd__nor2_4 _396_ (.A(_077_),
    .B(_083_),
    .Y(_019_));
 sky130_fd_sc_hd__nor2_4 _397_ (.A(_077_),
    .B(_084_),
    .Y(_018_));
 sky130_fd_sc_hd__nor2_4 _398_ (.A(_077_),
    .B(_085_),
    .Y(_011_));
 sky130_fd_sc_hd__nor2_4 _399_ (.A(_084_),
    .B(_088_),
    .Y(_015_));
 sky130_fd_sc_hd__nor2_4 _400_ (.A(_085_),
    .B(_088_),
    .Y(_014_));
 sky130_fd_sc_hd__xor2_1 _401_ (.A(\wr_ptr_gray_sync2[4] ),
    .B(\wr_ptr_gray_sync2[3] ),
    .X(_005_));
 sky130_fd_sc_hd__xnor2_1 _402_ (.A(\wr_ptr_gray_sync2[2] ),
    .B(_005_),
    .Y(_091_));
 sky130_fd_sc_hd__inv_1 _403_ (.A(_091_),
    .Y(_004_));
 sky130_fd_sc_hd__xnor2_1 _404_ (.A(\wr_ptr_gray_sync2[1] ),
    .B(_091_),
    .Y(_003_));
 sky130_fd_sc_hd__xor2_1 _405_ (.A(\wr_ptr_gray_sync2[0] ),
    .B(_003_),
    .X(_002_));
 sky130_fd_sc_hd__xor2_1 _406_ (.A(\rd_ptr_gray_sync2[4] ),
    .B(\rd_ptr_gray_sync2[3] ),
    .X(_009_));
 sky130_fd_sc_hd__xnor2_1 _407_ (.A(\rd_ptr_gray_sync2[2] ),
    .B(_009_),
    .Y(_092_));
 sky130_fd_sc_hd__inv_1 _408_ (.A(_092_),
    .Y(_008_));
 sky130_fd_sc_hd__xnor2_1 _409_ (.A(\rd_ptr_gray_sync2[1] ),
    .B(_092_),
    .Y(_007_));
 sky130_fd_sc_hd__xor2_1 _410_ (.A(\rd_ptr_gray_sync2[0] ),
    .B(_007_),
    .X(_006_));
 sky130_fd_sc_hd__nor2_4 _411_ (.A(_080_),
    .B(_087_),
    .Y(_013_));
 sky130_fd_sc_hd__buf_2 _412_ (.A(\rd_ptr_bin[1] ),
    .X(_093_));
 sky130_fd_sc_hd__buf_4 _413_ (.A(_093_),
    .X(_094_));
 sky130_fd_sc_hd__inv_1 _414_ (.A(_094_),
    .Y(_288_));
 sky130_fd_sc_hd__clkbuf_4 _415_ (.A(\rd_ptr_bin[0] ),
    .X(_095_));
 sky130_fd_sc_hd__inv_1 _416_ (.A(_095_),
    .Y(_029_));
 sky130_fd_sc_hd__inv_1 _417_ (.A(\rd_ptr_sync[0] ),
    .Y(_311_));
 sky130_fd_sc_hd__inv_1 _418_ (.A(\rd_ptr_sync[1] ),
    .Y(_291_));
 sky130_fd_sc_hd__inv_1 _419_ (.A(\rd_ptr_sync[2] ),
    .Y(_318_));
 sky130_fd_sc_hd__inv_1 _420_ (.A(\rd_ptr_sync[3] ),
    .Y(_322_));
 sky130_fd_sc_hd__inv_1 _421_ (.A(\wr_ptr_bin[0] ),
    .Y(_027_));
 sky130_fd_sc_hd__inv_1 _422_ (.A(\wr_ptr_sync[4] ),
    .Y(_297_));
 sky130_fd_sc_hd__inv_1 _423_ (.A(_308_),
    .Y(_289_));
 sky130_fd_sc_hd__inv_1 _424_ (.A(\wr_ptr_sync[0] ),
    .Y(_307_));
 sky130_fd_sc_hd__inv_1 _425_ (.A(_314_),
    .Y(_292_));
 sky130_fd_sc_hd__inv_1 _426_ (.A(\wr_ptr_bin[4] ),
    .Y(_326_));
 sky130_fd_sc_hd__inv_1 _427_ (.A(\wr_ptr_bin[1] ),
    .Y(_317_));
 sky130_fd_sc_hd__nand2b_1 _428_ (.A_N(net17),
    .B(net2),
    .Y(_096_));
 sky130_fd_sc_hd__buf_2 _429_ (.A(_096_),
    .X(_097_));
 sky130_fd_sc_hd__clkbuf_4 _430_ (.A(_097_),
    .X(_098_));
 sky130_fd_sc_hd__nand2_1 _431_ (.A(net25),
    .B(_098_),
    .Y(_099_));
 sky130_fd_sc_hd__nor2b_1 _432_ (.A(_089_),
    .B_N(_095_),
    .Y(_100_));
 sky130_fd_sc_hd__clkbuf_4 _433_ (.A(_100_),
    .X(_101_));
 sky130_fd_sc_hd__buf_2 _434_ (.A(_101_),
    .X(_102_));
 sky130_fd_sc_hd__buf_4 _435_ (.A(_094_),
    .X(_103_));
 sky130_fd_sc_hd__mux2i_1 _436_ (.A0(\mem[9][0] ),
    .A1(\mem[11][0] ),
    .S(_103_),
    .Y(_104_));
 sky130_fd_sc_hd__nand2_1 _437_ (.A(_102_),
    .B(_104_),
    .Y(_105_));
 sky130_fd_sc_hd__and2_0 _438_ (.A(_095_),
    .B(_089_),
    .X(_106_));
 sky130_fd_sc_hd__clkbuf_2 _439_ (.A(_106_),
    .X(_107_));
 sky130_fd_sc_hd__buf_6 _440_ (.A(_107_),
    .X(_108_));
 sky130_fd_sc_hd__buf_4 _441_ (.A(_093_),
    .X(_109_));
 sky130_fd_sc_hd__mux2i_2 _442_ (.A0(\mem[13][0] ),
    .A1(\mem[15][0] ),
    .S(_109_),
    .Y(_110_));
 sky130_fd_sc_hd__nor2b_1 _443_ (.A(_095_),
    .B_N(_089_),
    .Y(_111_));
 sky130_fd_sc_hd__clkbuf_2 _444_ (.A(_111_),
    .X(_112_));
 sky130_fd_sc_hd__clkbuf_4 _445_ (.A(_112_),
    .X(_113_));
 sky130_fd_sc_hd__buf_6 _446_ (.A(_093_),
    .X(_114_));
 sky130_fd_sc_hd__mux2i_1 _447_ (.A0(\mem[12][0] ),
    .A1(\mem[14][0] ),
    .S(_114_),
    .Y(_115_));
 sky130_fd_sc_hd__a22oi_2 _448_ (.A1(_108_),
    .A2(_110_),
    .B1(_113_),
    .B2(_115_),
    .Y(_116_));
 sky130_fd_sc_hd__nor2_4 _449_ (.A(_294_),
    .B(_097_),
    .Y(_117_));
 sky130_fd_sc_hd__nor2_2 _450_ (.A(_095_),
    .B(_089_),
    .Y(_118_));
 sky130_fd_sc_hd__buf_2 _451_ (.A(_118_),
    .X(_119_));
 sky130_fd_sc_hd__mux2i_1 _452_ (.A0(\mem[8][0] ),
    .A1(\mem[10][0] ),
    .S(_103_),
    .Y(_120_));
 sky130_fd_sc_hd__nand2_1 _453_ (.A(_119_),
    .B(_120_),
    .Y(_121_));
 sky130_fd_sc_hd__nand4_1 _454_ (.A(_105_),
    .B(_116_),
    .C(_117_),
    .D(_121_),
    .Y(_122_));
 sky130_fd_sc_hd__mux2i_1 _455_ (.A0(\mem[5][0] ),
    .A1(\mem[7][0] ),
    .S(_114_),
    .Y(_123_));
 sky130_fd_sc_hd__buf_6 _456_ (.A(_094_),
    .X(_124_));
 sky130_fd_sc_hd__mux2i_1 _457_ (.A0(\mem[1][0] ),
    .A1(\mem[3][0] ),
    .S(_124_),
    .Y(_125_));
 sky130_fd_sc_hd__a22oi_1 _458_ (.A1(_108_),
    .A2(_123_),
    .B1(_125_),
    .B2(_102_),
    .Y(_126_));
 sky130_fd_sc_hd__nor2_4 _459_ (.A(_090_),
    .B(_097_),
    .Y(_127_));
 sky130_fd_sc_hd__mux2i_1 _460_ (.A0(\mem[4][0] ),
    .A1(\mem[6][0] ),
    .S(_114_),
    .Y(_128_));
 sky130_fd_sc_hd__buf_6 _461_ (.A(_094_),
    .X(_129_));
 sky130_fd_sc_hd__mux2i_1 _462_ (.A0(\mem[0][0] ),
    .A1(\mem[2][0] ),
    .S(_129_),
    .Y(_130_));
 sky130_fd_sc_hd__a22oi_1 _463_ (.A1(_113_),
    .A2(_128_),
    .B1(_130_),
    .B2(_119_),
    .Y(_131_));
 sky130_fd_sc_hd__nand3_1 _464_ (.A(_126_),
    .B(_127_),
    .C(_131_),
    .Y(_132_));
 sky130_fd_sc_hd__nand3_1 _465_ (.A(_099_),
    .B(_122_),
    .C(_132_),
    .Y(_031_));
 sky130_fd_sc_hd__nand2_1 _466_ (.A(net26),
    .B(_098_),
    .Y(_133_));
 sky130_fd_sc_hd__mux2i_1 _467_ (.A0(\mem[9][1] ),
    .A1(\mem[11][1] ),
    .S(_103_),
    .Y(_134_));
 sky130_fd_sc_hd__nand2_1 _468_ (.A(_102_),
    .B(_134_),
    .Y(_135_));
 sky130_fd_sc_hd__mux2i_1 _469_ (.A0(\mem[13][1] ),
    .A1(\mem[15][1] ),
    .S(_109_),
    .Y(_136_));
 sky130_fd_sc_hd__buf_4 _470_ (.A(_093_),
    .X(_137_));
 sky130_fd_sc_hd__mux2i_1 _471_ (.A0(\mem[12][1] ),
    .A1(\mem[14][1] ),
    .S(_137_),
    .Y(_138_));
 sky130_fd_sc_hd__a22oi_1 _472_ (.A1(_108_),
    .A2(_136_),
    .B1(_138_),
    .B2(_113_),
    .Y(_139_));
 sky130_fd_sc_hd__mux2i_1 _473_ (.A0(\mem[8][1] ),
    .A1(\mem[10][1] ),
    .S(_124_),
    .Y(_140_));
 sky130_fd_sc_hd__nand2_1 _474_ (.A(_119_),
    .B(_140_),
    .Y(_141_));
 sky130_fd_sc_hd__nand4_1 _475_ (.A(_117_),
    .B(_135_),
    .C(_139_),
    .D(_141_),
    .Y(_142_));
 sky130_fd_sc_hd__mux2i_1 _476_ (.A0(\mem[0][1] ),
    .A1(\mem[2][1] ),
    .S(_114_),
    .Y(_143_));
 sky130_fd_sc_hd__mux2i_1 _477_ (.A0(\mem[1][1] ),
    .A1(\mem[3][1] ),
    .S(_124_),
    .Y(_144_));
 sky130_fd_sc_hd__a22oi_1 _478_ (.A1(_118_),
    .A2(_143_),
    .B1(_144_),
    .B2(_102_),
    .Y(_145_));
 sky130_fd_sc_hd__mux2i_1 _479_ (.A0(\mem[4][1] ),
    .A1(\mem[6][1] ),
    .S(_109_),
    .Y(_146_));
 sky130_fd_sc_hd__mux2i_1 _480_ (.A0(\mem[5][1] ),
    .A1(\mem[7][1] ),
    .S(_129_),
    .Y(_147_));
 sky130_fd_sc_hd__a22oi_1 _481_ (.A1(_113_),
    .A2(_146_),
    .B1(_147_),
    .B2(_108_),
    .Y(_148_));
 sky130_fd_sc_hd__nand3_1 _482_ (.A(_127_),
    .B(_145_),
    .C(_148_),
    .Y(_149_));
 sky130_fd_sc_hd__nand3_1 _483_ (.A(_133_),
    .B(_142_),
    .C(_149_),
    .Y(_032_));
 sky130_fd_sc_hd__nand2_1 _484_ (.A(net27),
    .B(_098_),
    .Y(_150_));
 sky130_fd_sc_hd__mux2i_1 _485_ (.A0(\mem[9][2] ),
    .A1(\mem[11][2] ),
    .S(_103_),
    .Y(_151_));
 sky130_fd_sc_hd__nand2_1 _486_ (.A(_102_),
    .B(_151_),
    .Y(_152_));
 sky130_fd_sc_hd__mux2i_1 _487_ (.A0(\mem[13][2] ),
    .A1(\mem[15][2] ),
    .S(_109_),
    .Y(_153_));
 sky130_fd_sc_hd__mux2i_1 _488_ (.A0(\mem[12][2] ),
    .A1(\mem[14][2] ),
    .S(_137_),
    .Y(_154_));
 sky130_fd_sc_hd__a22oi_1 _489_ (.A1(_107_),
    .A2(_153_),
    .B1(_154_),
    .B2(_113_),
    .Y(_155_));
 sky130_fd_sc_hd__mux2i_2 _490_ (.A0(\mem[8][2] ),
    .A1(\mem[10][2] ),
    .S(_124_),
    .Y(_156_));
 sky130_fd_sc_hd__nand2_1 _491_ (.A(_119_),
    .B(_156_),
    .Y(_157_));
 sky130_fd_sc_hd__nand4_1 _492_ (.A(_117_),
    .B(_152_),
    .C(_155_),
    .D(_157_),
    .Y(_158_));
 sky130_fd_sc_hd__mux2i_1 _493_ (.A0(\mem[5][2] ),
    .A1(\mem[7][2] ),
    .S(_114_),
    .Y(_159_));
 sky130_fd_sc_hd__mux2i_1 _494_ (.A0(\mem[1][2] ),
    .A1(\mem[3][2] ),
    .S(_124_),
    .Y(_160_));
 sky130_fd_sc_hd__a22oi_1 _495_ (.A1(_108_),
    .A2(_159_),
    .B1(_160_),
    .B2(_101_),
    .Y(_161_));
 sky130_fd_sc_hd__mux2i_1 _496_ (.A0(\mem[4][2] ),
    .A1(\mem[6][2] ),
    .S(_109_),
    .Y(_162_));
 sky130_fd_sc_hd__mux2i_1 _497_ (.A0(\mem[0][2] ),
    .A1(\mem[2][2] ),
    .S(_129_),
    .Y(_163_));
 sky130_fd_sc_hd__a22oi_1 _498_ (.A1(_112_),
    .A2(_162_),
    .B1(_163_),
    .B2(_119_),
    .Y(_164_));
 sky130_fd_sc_hd__nand3_1 _499_ (.A(_127_),
    .B(_161_),
    .C(_164_),
    .Y(_165_));
 sky130_fd_sc_hd__nand3_1 _500_ (.A(_150_),
    .B(_158_),
    .C(_165_),
    .Y(_033_));
 sky130_fd_sc_hd__nand2_1 _501_ (.A(net28),
    .B(_098_),
    .Y(_166_));
 sky130_fd_sc_hd__mux2i_1 _502_ (.A0(\mem[9][3] ),
    .A1(\mem[11][3] ),
    .S(_103_),
    .Y(_167_));
 sky130_fd_sc_hd__nand2_1 _503_ (.A(_102_),
    .B(_167_),
    .Y(_168_));
 sky130_fd_sc_hd__mux2i_1 _504_ (.A0(\mem[13][3] ),
    .A1(\mem[15][3] ),
    .S(_094_),
    .Y(_169_));
 sky130_fd_sc_hd__mux2i_1 _505_ (.A0(\mem[12][3] ),
    .A1(\mem[14][3] ),
    .S(_137_),
    .Y(_170_));
 sky130_fd_sc_hd__a22oi_1 _506_ (.A1(_107_),
    .A2(_169_),
    .B1(_170_),
    .B2(_113_),
    .Y(_171_));
 sky130_fd_sc_hd__mux2i_1 _507_ (.A0(\mem[8][3] ),
    .A1(\mem[10][3] ),
    .S(_124_),
    .Y(_172_));
 sky130_fd_sc_hd__nand2_1 _508_ (.A(_119_),
    .B(_172_),
    .Y(_173_));
 sky130_fd_sc_hd__nand4_1 _509_ (.A(_117_),
    .B(_168_),
    .C(_171_),
    .D(_173_),
    .Y(_174_));
 sky130_fd_sc_hd__mux2i_1 _510_ (.A0(\mem[5][3] ),
    .A1(\mem[7][3] ),
    .S(_114_),
    .Y(_175_));
 sky130_fd_sc_hd__mux2i_1 _511_ (.A0(\mem[1][3] ),
    .A1(\mem[3][3] ),
    .S(_129_),
    .Y(_176_));
 sky130_fd_sc_hd__a22oi_2 _512_ (.A1(_108_),
    .A2(_175_),
    .B1(_176_),
    .B2(_101_),
    .Y(_177_));
 sky130_fd_sc_hd__mux2i_1 _513_ (.A0(\mem[4][3] ),
    .A1(\mem[6][3] ),
    .S(_109_),
    .Y(_178_));
 sky130_fd_sc_hd__mux2i_1 _514_ (.A0(\mem[0][3] ),
    .A1(\mem[2][3] ),
    .S(_129_),
    .Y(_179_));
 sky130_fd_sc_hd__a22oi_1 _515_ (.A1(_112_),
    .A2(_178_),
    .B1(_179_),
    .B2(_118_),
    .Y(_180_));
 sky130_fd_sc_hd__nand3_2 _516_ (.A(_127_),
    .B(_177_),
    .C(_180_),
    .Y(_181_));
 sky130_fd_sc_hd__nand3_1 _517_ (.A(_166_),
    .B(_174_),
    .C(_181_),
    .Y(_034_));
 sky130_fd_sc_hd__nand2_1 _518_ (.A(net29),
    .B(_098_),
    .Y(_182_));
 sky130_fd_sc_hd__mux2i_1 _519_ (.A0(\mem[9][4] ),
    .A1(\mem[11][4] ),
    .S(_103_),
    .Y(_183_));
 sky130_fd_sc_hd__nand2_1 _520_ (.A(_102_),
    .B(_183_),
    .Y(_184_));
 sky130_fd_sc_hd__mux2i_1 _521_ (.A0(\mem[13][4] ),
    .A1(\mem[15][4] ),
    .S(_094_),
    .Y(_185_));
 sky130_fd_sc_hd__mux2i_1 _522_ (.A0(\mem[12][4] ),
    .A1(\mem[14][4] ),
    .S(_137_),
    .Y(_186_));
 sky130_fd_sc_hd__a22oi_1 _523_ (.A1(_107_),
    .A2(_185_),
    .B1(_186_),
    .B2(_113_),
    .Y(_187_));
 sky130_fd_sc_hd__mux2i_1 _524_ (.A0(\mem[8][4] ),
    .A1(\mem[10][4] ),
    .S(_124_),
    .Y(_188_));
 sky130_fd_sc_hd__nand2_1 _525_ (.A(_119_),
    .B(_188_),
    .Y(_189_));
 sky130_fd_sc_hd__nand4_1 _526_ (.A(_117_),
    .B(_184_),
    .C(_187_),
    .D(_189_),
    .Y(_190_));
 sky130_fd_sc_hd__mux2i_1 _527_ (.A0(\mem[5][4] ),
    .A1(\mem[7][4] ),
    .S(_114_),
    .Y(_191_));
 sky130_fd_sc_hd__mux2i_1 _528_ (.A0(\mem[1][4] ),
    .A1(\mem[3][4] ),
    .S(_129_),
    .Y(_192_));
 sky130_fd_sc_hd__a22oi_2 _529_ (.A1(_108_),
    .A2(_191_),
    .B1(_192_),
    .B2(_101_),
    .Y(_193_));
 sky130_fd_sc_hd__mux2i_1 _530_ (.A0(\mem[4][4] ),
    .A1(\mem[6][4] ),
    .S(_109_),
    .Y(_194_));
 sky130_fd_sc_hd__mux2i_1 _531_ (.A0(\mem[0][4] ),
    .A1(\mem[2][4] ),
    .S(_129_),
    .Y(_195_));
 sky130_fd_sc_hd__a22oi_1 _532_ (.A1(_112_),
    .A2(_194_),
    .B1(_195_),
    .B2(_118_),
    .Y(_196_));
 sky130_fd_sc_hd__nand3_2 _533_ (.A(_127_),
    .B(_193_),
    .C(_196_),
    .Y(_197_));
 sky130_fd_sc_hd__nand3_1 _534_ (.A(_182_),
    .B(_190_),
    .C(_197_),
    .Y(_035_));
 sky130_fd_sc_hd__nand2_1 _535_ (.A(net30),
    .B(_098_),
    .Y(_198_));
 sky130_fd_sc_hd__mux2i_1 _536_ (.A0(\mem[9][5] ),
    .A1(\mem[11][5] ),
    .S(_103_),
    .Y(_199_));
 sky130_fd_sc_hd__nand2_1 _537_ (.A(_102_),
    .B(_199_),
    .Y(_200_));
 sky130_fd_sc_hd__mux2i_1 _538_ (.A0(\mem[13][5] ),
    .A1(\mem[15][5] ),
    .S(_094_),
    .Y(_201_));
 sky130_fd_sc_hd__mux2i_1 _539_ (.A0(\mem[12][5] ),
    .A1(\mem[14][5] ),
    .S(_137_),
    .Y(_202_));
 sky130_fd_sc_hd__a22oi_1 _540_ (.A1(_107_),
    .A2(_201_),
    .B1(_202_),
    .B2(_113_),
    .Y(_203_));
 sky130_fd_sc_hd__mux2i_1 _541_ (.A0(\mem[8][5] ),
    .A1(\mem[10][5] ),
    .S(_124_),
    .Y(_204_));
 sky130_fd_sc_hd__nand2_1 _542_ (.A(_119_),
    .B(_204_),
    .Y(_205_));
 sky130_fd_sc_hd__nand4_1 _543_ (.A(_117_),
    .B(_200_),
    .C(_203_),
    .D(_205_),
    .Y(_206_));
 sky130_fd_sc_hd__mux2i_1 _544_ (.A0(\mem[0][5] ),
    .A1(\mem[2][5] ),
    .S(_114_),
    .Y(_207_));
 sky130_fd_sc_hd__mux2i_1 _545_ (.A0(\mem[1][5] ),
    .A1(\mem[3][5] ),
    .S(_129_),
    .Y(_208_));
 sky130_fd_sc_hd__a22oi_1 _546_ (.A1(_118_),
    .A2(_207_),
    .B1(_208_),
    .B2(_101_),
    .Y(_209_));
 sky130_fd_sc_hd__mux2i_2 _547_ (.A0(\mem[4][5] ),
    .A1(\mem[6][5] ),
    .S(_109_),
    .Y(_210_));
 sky130_fd_sc_hd__mux2i_1 _548_ (.A0(\mem[5][5] ),
    .A1(\mem[7][5] ),
    .S(_137_),
    .Y(_211_));
 sky130_fd_sc_hd__a22oi_1 _549_ (.A1(_112_),
    .A2(_210_),
    .B1(_211_),
    .B2(_108_),
    .Y(_212_));
 sky130_fd_sc_hd__nand3_1 _550_ (.A(_127_),
    .B(_209_),
    .C(_212_),
    .Y(_213_));
 sky130_fd_sc_hd__nand3_1 _551_ (.A(_198_),
    .B(_206_),
    .C(_213_),
    .Y(_036_));
 sky130_fd_sc_hd__nand2_1 _552_ (.A(net31),
    .B(_098_),
    .Y(_214_));
 sky130_fd_sc_hd__mux2i_1 _553_ (.A0(\mem[9][6] ),
    .A1(\mem[11][6] ),
    .S(_103_),
    .Y(_215_));
 sky130_fd_sc_hd__nand2_1 _554_ (.A(_102_),
    .B(_215_),
    .Y(_216_));
 sky130_fd_sc_hd__mux2i_1 _555_ (.A0(\mem[13][6] ),
    .A1(\mem[15][6] ),
    .S(_094_),
    .Y(_217_));
 sky130_fd_sc_hd__mux2i_1 _556_ (.A0(\mem[12][6] ),
    .A1(\mem[14][6] ),
    .S(_137_),
    .Y(_218_));
 sky130_fd_sc_hd__a22oi_1 _557_ (.A1(_107_),
    .A2(_217_),
    .B1(_218_),
    .B2(_113_),
    .Y(_219_));
 sky130_fd_sc_hd__mux2i_1 _558_ (.A0(\mem[8][6] ),
    .A1(\mem[10][6] ),
    .S(_124_),
    .Y(_220_));
 sky130_fd_sc_hd__nand2_1 _559_ (.A(_119_),
    .B(_220_),
    .Y(_221_));
 sky130_fd_sc_hd__nand4_1 _560_ (.A(_117_),
    .B(_216_),
    .C(_219_),
    .D(_221_),
    .Y(_222_));
 sky130_fd_sc_hd__mux2i_1 _561_ (.A0(\mem[0][6] ),
    .A1(\mem[2][6] ),
    .S(_114_),
    .Y(_223_));
 sky130_fd_sc_hd__mux2i_1 _562_ (.A0(\mem[1][6] ),
    .A1(\mem[3][6] ),
    .S(_129_),
    .Y(_224_));
 sky130_fd_sc_hd__a22oi_1 _563_ (.A1(_118_),
    .A2(_223_),
    .B1(_224_),
    .B2(_101_),
    .Y(_225_));
 sky130_fd_sc_hd__mux2i_1 _564_ (.A0(\mem[4][6] ),
    .A1(\mem[6][6] ),
    .S(_109_),
    .Y(_226_));
 sky130_fd_sc_hd__mux2i_1 _565_ (.A0(\mem[5][6] ),
    .A1(\mem[7][6] ),
    .S(_137_),
    .Y(_227_));
 sky130_fd_sc_hd__a22oi_1 _566_ (.A1(_112_),
    .A2(_226_),
    .B1(_227_),
    .B2(_108_),
    .Y(_228_));
 sky130_fd_sc_hd__nand3_1 _567_ (.A(_127_),
    .B(_225_),
    .C(_228_),
    .Y(_229_));
 sky130_fd_sc_hd__nand3_1 _568_ (.A(_214_),
    .B(_222_),
    .C(_229_),
    .Y(_037_));
 sky130_fd_sc_hd__nand2_1 _569_ (.A(net32),
    .B(_098_),
    .Y(_230_));
 sky130_fd_sc_hd__mux2i_1 _570_ (.A0(\mem[9][7] ),
    .A1(\mem[11][7] ),
    .S(_103_),
    .Y(_231_));
 sky130_fd_sc_hd__nand2_1 _571_ (.A(_102_),
    .B(_231_),
    .Y(_232_));
 sky130_fd_sc_hd__mux2i_1 _572_ (.A0(\mem[13][7] ),
    .A1(\mem[15][7] ),
    .S(_094_),
    .Y(_233_));
 sky130_fd_sc_hd__mux2i_1 _573_ (.A0(\mem[12][7] ),
    .A1(\mem[14][7] ),
    .S(_137_),
    .Y(_234_));
 sky130_fd_sc_hd__a22oi_1 _574_ (.A1(_107_),
    .A2(_233_),
    .B1(_234_),
    .B2(_113_),
    .Y(_235_));
 sky130_fd_sc_hd__mux2i_2 _575_ (.A0(\mem[8][7] ),
    .A1(\mem[10][7] ),
    .S(_124_),
    .Y(_236_));
 sky130_fd_sc_hd__nand2_1 _576_ (.A(_119_),
    .B(_236_),
    .Y(_237_));
 sky130_fd_sc_hd__nand4_1 _577_ (.A(_117_),
    .B(_232_),
    .C(_235_),
    .D(_237_),
    .Y(_238_));
 sky130_fd_sc_hd__mux2i_1 _578_ (.A0(\mem[5][7] ),
    .A1(\mem[7][7] ),
    .S(_114_),
    .Y(_239_));
 sky130_fd_sc_hd__mux2i_1 _579_ (.A0(\mem[1][7] ),
    .A1(\mem[3][7] ),
    .S(_129_),
    .Y(_240_));
 sky130_fd_sc_hd__a22oi_1 _580_ (.A1(_108_),
    .A2(_239_),
    .B1(_240_),
    .B2(_101_),
    .Y(_241_));
 sky130_fd_sc_hd__mux2i_1 _581_ (.A0(\mem[4][7] ),
    .A1(\mem[6][7] ),
    .S(_109_),
    .Y(_242_));
 sky130_fd_sc_hd__mux2i_1 _582_ (.A0(\mem[0][7] ),
    .A1(\mem[2][7] ),
    .S(_137_),
    .Y(_243_));
 sky130_fd_sc_hd__a22oi_1 _583_ (.A1(_112_),
    .A2(_242_),
    .B1(_243_),
    .B2(_118_),
    .Y(_244_));
 sky130_fd_sc_hd__nand3_1 _584_ (.A(_127_),
    .B(_241_),
    .C(_244_),
    .Y(_245_));
 sky130_fd_sc_hd__nand3_1 _585_ (.A(_230_),
    .B(_238_),
    .C(_245_),
    .Y(_038_));
 sky130_fd_sc_hd__nor2b_1 _586_ (.A(net17),
    .B_N(net2),
    .Y(_246_));
 sky130_fd_sc_hd__clkbuf_2 _587_ (.A(_246_),
    .X(_247_));
 sky130_fd_sc_hd__xnor2_1 _588_ (.A(_029_),
    .B(_247_),
    .Y(_039_));
 sky130_fd_sc_hd__nand2_1 _589_ (.A(_030_),
    .B(_247_),
    .Y(_248_));
 sky130_fd_sc_hd__o21ai_0 _590_ (.A1(_288_),
    .A2(_247_),
    .B1(_248_),
    .Y(_040_));
 sky130_fd_sc_hd__nand2_1 _591_ (.A(_329_),
    .B(_247_),
    .Y(_249_));
 sky130_fd_sc_hd__xnor2_1 _592_ (.A(_089_),
    .B(_249_),
    .Y(_041_));
 sky130_fd_sc_hd__nand4_1 _593_ (.A(_095_),
    .B(_103_),
    .C(_089_),
    .D(_247_),
    .Y(_250_));
 sky130_fd_sc_hd__xnor2_1 _594_ (.A(_090_),
    .B(_250_),
    .Y(_042_));
 sky130_fd_sc_hd__xor2_1 _595_ (.A(_095_),
    .B(_030_),
    .X(_251_));
 sky130_fd_sc_hd__nand2_1 _596_ (.A(\rd_ptr_gray[0] ),
    .B(_098_),
    .Y(_252_));
 sky130_fd_sc_hd__o21ai_0 _597_ (.A1(_097_),
    .A2(_251_),
    .B1(_252_),
    .Y(_043_));
 sky130_fd_sc_hd__xnor2_1 _598_ (.A(_329_),
    .B(_030_),
    .Y(_253_));
 sky130_fd_sc_hd__xnor2_1 _599_ (.A(_302_),
    .B(_253_),
    .Y(_254_));
 sky130_fd_sc_hd__nand2_1 _600_ (.A(\rd_ptr_gray[1] ),
    .B(_098_),
    .Y(_255_));
 sky130_fd_sc_hd__o21ai_0 _601_ (.A1(_097_),
    .A2(_254_),
    .B1(_255_),
    .Y(_044_));
 sky130_fd_sc_hd__xnor2_1 _602_ (.A(_090_),
    .B(_329_),
    .Y(_256_));
 sky130_fd_sc_hd__o21ai_0 _603_ (.A1(_029_),
    .A2(_288_),
    .B1(_089_),
    .Y(_257_));
 sky130_fd_sc_hd__xnor2_1 _604_ (.A(_256_),
    .B(_257_),
    .Y(_258_));
 sky130_fd_sc_hd__nand2_1 _605_ (.A(\rd_ptr_gray[2] ),
    .B(_097_),
    .Y(_259_));
 sky130_fd_sc_hd__o21ai_0 _606_ (.A1(_097_),
    .A2(_258_),
    .B1(_259_),
    .Y(_045_));
 sky130_fd_sc_hd__a31oi_1 _607_ (.A1(_095_),
    .A2(_094_),
    .A3(_089_),
    .B1(_090_),
    .Y(_260_));
 sky130_fd_sc_hd__nand4b_1 _608_ (.A_N(_329_),
    .B(_090_),
    .C(_093_),
    .D(_095_),
    .Y(_261_));
 sky130_fd_sc_hd__a21bo_1 _609_ (.A1(_095_),
    .A2(_093_),
    .B1_N(_329_),
    .X(_262_));
 sky130_fd_sc_hd__a21oi_1 _610_ (.A1(_261_),
    .A2(_262_),
    .B1(_302_),
    .Y(_263_));
 sky130_fd_sc_hd__o21ai_0 _611_ (.A1(_260_),
    .A2(_263_),
    .B1(\rd_ptr_bin[4] ),
    .Y(_264_));
 sky130_fd_sc_hd__or3_1 _612_ (.A(\rd_ptr_bin[4] ),
    .B(_260_),
    .C(_263_),
    .X(_265_));
 sky130_fd_sc_hd__nor2_1 _613_ (.A(\rd_ptr_gray[3] ),
    .B(_247_),
    .Y(_266_));
 sky130_fd_sc_hd__a31oi_1 _614_ (.A1(_247_),
    .A2(_264_),
    .A3(_265_),
    .B1(_266_),
    .Y(_046_));
 sky130_fd_sc_hd__nand3_1 _615_ (.A(_089_),
    .B(_329_),
    .C(_117_),
    .Y(_267_));
 sky130_fd_sc_hd__xnor2_1 _616_ (.A(\rd_ptr_bin[4] ),
    .B(_267_),
    .Y(_047_));
 sky130_fd_sc_hd__xnor2_1 _617_ (.A(_027_),
    .B(_082_),
    .Y(_048_));
 sky130_fd_sc_hd__nand2_1 _618_ (.A(_028_),
    .B(_082_),
    .Y(_268_));
 sky130_fd_sc_hd__o21ai_0 _619_ (.A1(_317_),
    .A2(_082_),
    .B1(_268_),
    .Y(_049_));
 sky130_fd_sc_hd__xnor2_1 _620_ (.A(_075_),
    .B(_087_),
    .Y(_050_));
 sky130_fd_sc_hd__and2_0 _621_ (.A(\wr_ptr_bin[1] ),
    .B(\wr_ptr_bin[0] ),
    .X(_269_));
 sky130_fd_sc_hd__nand3_1 _622_ (.A(_075_),
    .B(_082_),
    .C(_269_),
    .Y(_270_));
 sky130_fd_sc_hd__xnor2_1 _623_ (.A(_074_),
    .B(_270_),
    .Y(_051_));
 sky130_fd_sc_hd__nand2b_2 _624_ (.A_N(net18),
    .B(net13),
    .Y(_271_));
 sky130_fd_sc_hd__xor2_1 _625_ (.A(\wr_ptr_bin[0] ),
    .B(_028_),
    .X(_272_));
 sky130_fd_sc_hd__nand2_1 _626_ (.A(\wr_ptr_gray[0] ),
    .B(_271_),
    .Y(_273_));
 sky130_fd_sc_hd__o21ai_0 _627_ (.A1(_271_),
    .A2(_272_),
    .B1(_273_),
    .Y(_052_));
 sky130_fd_sc_hd__xnor2_1 _628_ (.A(_335_),
    .B(_028_),
    .Y(_274_));
 sky130_fd_sc_hd__xnor2_1 _629_ (.A(_321_),
    .B(_274_),
    .Y(_275_));
 sky130_fd_sc_hd__nand2_1 _630_ (.A(\wr_ptr_gray[1] ),
    .B(_271_),
    .Y(_276_));
 sky130_fd_sc_hd__o21ai_0 _631_ (.A1(_271_),
    .A2(_275_),
    .B1(_276_),
    .Y(_053_));
 sky130_fd_sc_hd__xnor2_1 _632_ (.A(_074_),
    .B(_335_),
    .Y(_277_));
 sky130_fd_sc_hd__o21ai_0 _633_ (.A1(_317_),
    .A2(_027_),
    .B1(_075_),
    .Y(_278_));
 sky130_fd_sc_hd__xnor2_1 _634_ (.A(_277_),
    .B(_278_),
    .Y(_279_));
 sky130_fd_sc_hd__nand2_1 _635_ (.A(\wr_ptr_gray[2] ),
    .B(_271_),
    .Y(_280_));
 sky130_fd_sc_hd__o21ai_0 _636_ (.A1(_271_),
    .A2(_279_),
    .B1(_280_),
    .Y(_054_));
 sky130_fd_sc_hd__a21boi_0 _637_ (.A1(_075_),
    .A2(_335_),
    .B1_N(_074_),
    .Y(_281_));
 sky130_fd_sc_hd__nand4_1 _638_ (.A(_074_),
    .B(_075_),
    .C(\wr_ptr_bin[1] ),
    .D(\wr_ptr_bin[0] ),
    .Y(_282_));
 sky130_fd_sc_hd__o221ai_2 _639_ (.A1(_269_),
    .A2(_281_),
    .B1(_282_),
    .B2(_335_),
    .C1(_077_),
    .Y(_283_));
 sky130_fd_sc_hd__xnor2_1 _640_ (.A(_326_),
    .B(_283_),
    .Y(_284_));
 sky130_fd_sc_hd__nand2_1 _641_ (.A(\wr_ptr_gray[3] ),
    .B(_271_),
    .Y(_285_));
 sky130_fd_sc_hd__o21ai_0 _642_ (.A1(_271_),
    .A2(_284_),
    .B1(_285_),
    .Y(_055_));
 sky130_fd_sc_hd__xnor2_1 _643_ (.A(_326_),
    .B(_017_),
    .Y(_056_));
 sky130_fd_sc_hd__nor2b_1 _644_ (.A(_306_),
    .B_N(net21),
    .Y(_286_));
 sky130_fd_sc_hd__a2111oi_0 _645_ (.A1(_063_),
    .A2(_064_),
    .B1(_286_),
    .C1(net22),
    .D1(net24),
    .Y(net15));
 sky130_fd_sc_hd__xor2_1 _646_ (.A(_320_),
    .B(_293_),
    .X(net36));
 sky130_fd_sc_hd__nand2_1 _647_ (.A(net35),
    .B(net36),
    .Y(_287_));
 sky130_fd_sc_hd__o31ai_1 _648_ (.A1(_068_),
    .A2(_069_),
    .A3(_287_),
    .B1(_072_),
    .Y(net16));
 sky130_fd_sc_hd__fa_1 _649_ (.A(_288_),
    .B(\wr_ptr_sync[1] ),
    .CIN(_289_),
    .COUT(_290_),
    .SUM(net21));
 sky130_fd_sc_hd__fa_1 _650_ (.A(_291_),
    .B(\wr_ptr_bin[1] ),
    .CIN(_292_),
    .COUT(_293_),
    .SUM(net35));
 sky130_fd_sc_hd__ha_1 _651_ (.A(_294_),
    .B(\wr_ptr_sync[3] ),
    .COUT(_295_),
    .SUM(_296_));
 sky130_fd_sc_hd__ha_1 _652_ (.A(\rd_ptr_bin[4] ),
    .B(_297_),
    .COUT(_298_),
    .SUM(_299_));
 sky130_fd_sc_hd__ha_1 _653_ (.A(_288_),
    .B(\wr_ptr_sync[1] ),
    .COUT(_300_),
    .SUM(_301_));
 sky130_fd_sc_hd__ha_1 _654_ (.A(_302_),
    .B(\wr_ptr_sync[2] ),
    .COUT(_303_),
    .SUM(_304_));
 sky130_fd_sc_hd__ha_1 _655_ (.A(_029_),
    .B(\wr_ptr_sync[0] ),
    .COUT(_305_),
    .SUM(_306_));
 sky130_fd_sc_hd__ha_1 _656_ (.A(\rd_ptr_bin[0] ),
    .B(_307_),
    .COUT(_308_),
    .SUM(_309_));
 sky130_fd_sc_hd__ha_1 _657_ (.A(_311_),
    .B(\wr_ptr_bin[0] ),
    .COUT(_312_),
    .SUM(_313_));
 sky130_fd_sc_hd__ha_1 _658_ (.A(\rd_ptr_sync[0] ),
    .B(_027_),
    .COUT(_314_),
    .SUM(_315_));
 sky130_fd_sc_hd__ha_1 _659_ (.A(_291_),
    .B(\wr_ptr_bin[1] ),
    .COUT(_316_),
    .SUM(_310_));
 sky130_fd_sc_hd__ha_1 _660_ (.A(_318_),
    .B(\wr_ptr_bin[2] ),
    .COUT(_319_),
    .SUM(_320_));
 sky130_fd_sc_hd__ha_1 _661_ (.A(_322_),
    .B(\wr_ptr_bin[3] ),
    .COUT(_323_),
    .SUM(_324_));
 sky130_fd_sc_hd__ha_1 _662_ (.A(\rd_ptr_sync[4] ),
    .B(_326_),
    .COUT(_327_),
    .SUM(_328_));
 sky130_fd_sc_hd__ha_1 _663_ (.A(\rd_ptr_bin[0] ),
    .B(\rd_ptr_bin[1] ),
    .COUT(_329_),
    .SUM(_030_));
 sky130_fd_sc_hd__ha_1 _664_ (.A(_027_),
    .B(_317_),
    .COUT(_330_),
    .SUM(_028_));
 sky130_fd_sc_hd__ha_1 _665_ (.A(_027_),
    .B(\wr_ptr_bin[1] ),
    .COUT(_331_),
    .SUM(_332_));
 sky130_fd_sc_hd__ha_1 _666_ (.A(\wr_ptr_bin[0] ),
    .B(_317_),
    .COUT(_333_),
    .SUM(_334_));
 sky130_fd_sc_hd__ha_2 _667_ (.A(\wr_ptr_bin[0] ),
    .B(\wr_ptr_bin[1] ),
    .COUT(_335_),
    .SUM(_336_));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__dfstp_1 \empty_reg$_DFF_PN1_  (.D(_000_),
    .Q(net17),
    .SET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \full_reg$_DFF_PN0_  (.D(_001_),
    .Q(net18),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][0]$_DFFE_PP_  (.D(net5),
    .DE(_011_),
    .Q(\mem[0][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][1]$_DFFE_PP_  (.D(net6),
    .DE(_011_),
    .Q(\mem[0][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][2]$_DFFE_PP_  (.D(net7),
    .DE(_011_),
    .Q(\mem[0][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][3]$_DFFE_PP_  (.D(net8),
    .DE(_011_),
    .Q(\mem[0][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][4]$_DFFE_PP_  (.D(net9),
    .DE(_011_),
    .Q(\mem[0][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][5]$_DFFE_PP_  (.D(net10),
    .DE(_011_),
    .Q(\mem[0][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][6]$_DFFE_PP_  (.D(net11),
    .DE(_011_),
    .Q(\mem[0][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][7]$_DFFE_PP_  (.D(net12),
    .DE(_011_),
    .Q(\mem[0][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][0]$_DFFE_PP_  (.D(net5),
    .DE(_012_),
    .Q(\mem[10][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][1]$_DFFE_PP_  (.D(net6),
    .DE(_012_),
    .Q(\mem[10][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][2]$_DFFE_PP_  (.D(net7),
    .DE(_012_),
    .Q(\mem[10][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][3]$_DFFE_PP_  (.D(net8),
    .DE(_012_),
    .Q(\mem[10][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][4]$_DFFE_PP_  (.D(net9),
    .DE(_012_),
    .Q(\mem[10][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][5]$_DFFE_PP_  (.D(net10),
    .DE(_012_),
    .Q(\mem[10][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][6]$_DFFE_PP_  (.D(net11),
    .DE(_012_),
    .Q(\mem[10][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][7]$_DFFE_PP_  (.D(net12),
    .DE(_012_),
    .Q(\mem[10][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][0]$_DFFE_PP_  (.D(net5),
    .DE(_013_),
    .Q(\mem[11][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][1]$_DFFE_PP_  (.D(net6),
    .DE(_013_),
    .Q(\mem[11][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][2]$_DFFE_PP_  (.D(net7),
    .DE(_013_),
    .Q(\mem[11][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][3]$_DFFE_PP_  (.D(net8),
    .DE(_013_),
    .Q(\mem[11][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][4]$_DFFE_PP_  (.D(net9),
    .DE(_013_),
    .Q(\mem[11][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][5]$_DFFE_PP_  (.D(net10),
    .DE(_013_),
    .Q(\mem[11][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][6]$_DFFE_PP_  (.D(net11),
    .DE(_013_),
    .Q(\mem[11][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][7]$_DFFE_PP_  (.D(net12),
    .DE(_013_),
    .Q(\mem[11][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][0]$_DFFE_PP_  (.D(net5),
    .DE(_014_),
    .Q(\mem[12][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][1]$_DFFE_PP_  (.D(net6),
    .DE(_014_),
    .Q(\mem[12][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][2]$_DFFE_PP_  (.D(net7),
    .DE(_014_),
    .Q(\mem[12][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][3]$_DFFE_PP_  (.D(net8),
    .DE(_014_),
    .Q(\mem[12][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][4]$_DFFE_PP_  (.D(net9),
    .DE(_014_),
    .Q(\mem[12][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][5]$_DFFE_PP_  (.D(net10),
    .DE(_014_),
    .Q(\mem[12][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][6]$_DFFE_PP_  (.D(net11),
    .DE(_014_),
    .Q(\mem[12][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][7]$_DFFE_PP_  (.D(net12),
    .DE(_014_),
    .Q(\mem[12][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][0]$_DFFE_PP_  (.D(net5),
    .DE(_015_),
    .Q(\mem[13][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][1]$_DFFE_PP_  (.D(net6),
    .DE(_015_),
    .Q(\mem[13][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][2]$_DFFE_PP_  (.D(net7),
    .DE(_015_),
    .Q(\mem[13][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][3]$_DFFE_PP_  (.D(net8),
    .DE(_015_),
    .Q(\mem[13][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][4]$_DFFE_PP_  (.D(net9),
    .DE(_015_),
    .Q(\mem[13][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][5]$_DFFE_PP_  (.D(net10),
    .DE(_015_),
    .Q(\mem[13][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][6]$_DFFE_PP_  (.D(net11),
    .DE(_015_),
    .Q(\mem[13][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][7]$_DFFE_PP_  (.D(net12),
    .DE(_015_),
    .Q(\mem[13][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][0]$_DFFE_PP_  (.D(net5),
    .DE(_016_),
    .Q(\mem[14][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][1]$_DFFE_PP_  (.D(net6),
    .DE(_016_),
    .Q(\mem[14][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][2]$_DFFE_PP_  (.D(net7),
    .DE(_016_),
    .Q(\mem[14][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][3]$_DFFE_PP_  (.D(net8),
    .DE(_016_),
    .Q(\mem[14][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][4]$_DFFE_PP_  (.D(net9),
    .DE(_016_),
    .Q(\mem[14][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][5]$_DFFE_PP_  (.D(net10),
    .DE(_016_),
    .Q(\mem[14][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][6]$_DFFE_PP_  (.D(net11),
    .DE(_016_),
    .Q(\mem[14][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][7]$_DFFE_PP_  (.D(net12),
    .DE(_016_),
    .Q(\mem[14][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][0]$_DFFE_PP_  (.D(net5),
    .DE(_017_),
    .Q(\mem[15][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][1]$_DFFE_PP_  (.D(net6),
    .DE(_017_),
    .Q(\mem[15][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][2]$_DFFE_PP_  (.D(net7),
    .DE(_017_),
    .Q(\mem[15][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][3]$_DFFE_PP_  (.D(net8),
    .DE(_017_),
    .Q(\mem[15][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][4]$_DFFE_PP_  (.D(net9),
    .DE(_017_),
    .Q(\mem[15][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][5]$_DFFE_PP_  (.D(net10),
    .DE(_017_),
    .Q(\mem[15][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][6]$_DFFE_PP_  (.D(net11),
    .DE(_017_),
    .Q(\mem[15][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][7]$_DFFE_PP_  (.D(net12),
    .DE(_017_),
    .Q(\mem[15][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][0]$_DFFE_PP_  (.D(net5),
    .DE(_018_),
    .Q(\mem[1][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][1]$_DFFE_PP_  (.D(net6),
    .DE(_018_),
    .Q(\mem[1][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][2]$_DFFE_PP_  (.D(net7),
    .DE(_018_),
    .Q(\mem[1][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][3]$_DFFE_PP_  (.D(net8),
    .DE(_018_),
    .Q(\mem[1][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][4]$_DFFE_PP_  (.D(net9),
    .DE(_018_),
    .Q(\mem[1][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][5]$_DFFE_PP_  (.D(net10),
    .DE(_018_),
    .Q(\mem[1][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][6]$_DFFE_PP_  (.D(net11),
    .DE(_018_),
    .Q(\mem[1][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][7]$_DFFE_PP_  (.D(net12),
    .DE(_018_),
    .Q(\mem[1][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][0]$_DFFE_PP_  (.D(net5),
    .DE(_019_),
    .Q(\mem[2][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][1]$_DFFE_PP_  (.D(net6),
    .DE(_019_),
    .Q(\mem[2][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][2]$_DFFE_PP_  (.D(net7),
    .DE(_019_),
    .Q(\mem[2][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][3]$_DFFE_PP_  (.D(net8),
    .DE(_019_),
    .Q(\mem[2][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][4]$_DFFE_PP_  (.D(net9),
    .DE(_019_),
    .Q(\mem[2][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][5]$_DFFE_PP_  (.D(net10),
    .DE(_019_),
    .Q(\mem[2][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][6]$_DFFE_PP_  (.D(net11),
    .DE(_019_),
    .Q(\mem[2][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][7]$_DFFE_PP_  (.D(net12),
    .DE(_019_),
    .Q(\mem[2][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][0]$_DFFE_PP_  (.D(net5),
    .DE(_020_),
    .Q(\mem[3][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][1]$_DFFE_PP_  (.D(net6),
    .DE(_020_),
    .Q(\mem[3][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][2]$_DFFE_PP_  (.D(net7),
    .DE(_020_),
    .Q(\mem[3][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][3]$_DFFE_PP_  (.D(net8),
    .DE(_020_),
    .Q(\mem[3][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][4]$_DFFE_PP_  (.D(net9),
    .DE(_020_),
    .Q(\mem[3][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][5]$_DFFE_PP_  (.D(net10),
    .DE(_020_),
    .Q(\mem[3][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][6]$_DFFE_PP_  (.D(net11),
    .DE(_020_),
    .Q(\mem[3][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][7]$_DFFE_PP_  (.D(net12),
    .DE(_020_),
    .Q(\mem[3][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][0]$_DFFE_PP_  (.D(net5),
    .DE(_021_),
    .Q(\mem[4][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][1]$_DFFE_PP_  (.D(net6),
    .DE(_021_),
    .Q(\mem[4][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][2]$_DFFE_PP_  (.D(net7),
    .DE(_021_),
    .Q(\mem[4][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][3]$_DFFE_PP_  (.D(net8),
    .DE(_021_),
    .Q(\mem[4][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][4]$_DFFE_PP_  (.D(net9),
    .DE(_021_),
    .Q(\mem[4][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][5]$_DFFE_PP_  (.D(net10),
    .DE(_021_),
    .Q(\mem[4][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][6]$_DFFE_PP_  (.D(net11),
    .DE(_021_),
    .Q(\mem[4][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][7]$_DFFE_PP_  (.D(net12),
    .DE(_021_),
    .Q(\mem[4][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][0]$_DFFE_PP_  (.D(net5),
    .DE(_022_),
    .Q(\mem[5][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][1]$_DFFE_PP_  (.D(net6),
    .DE(_022_),
    .Q(\mem[5][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][2]$_DFFE_PP_  (.D(net7),
    .DE(_022_),
    .Q(\mem[5][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][3]$_DFFE_PP_  (.D(net8),
    .DE(_022_),
    .Q(\mem[5][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][4]$_DFFE_PP_  (.D(net9),
    .DE(_022_),
    .Q(\mem[5][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][5]$_DFFE_PP_  (.D(net10),
    .DE(_022_),
    .Q(\mem[5][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][6]$_DFFE_PP_  (.D(net11),
    .DE(_022_),
    .Q(\mem[5][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][7]$_DFFE_PP_  (.D(net12),
    .DE(_022_),
    .Q(\mem[5][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][0]$_DFFE_PP_  (.D(net5),
    .DE(_023_),
    .Q(\mem[6][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][1]$_DFFE_PP_  (.D(net6),
    .DE(_023_),
    .Q(\mem[6][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][2]$_DFFE_PP_  (.D(net7),
    .DE(_023_),
    .Q(\mem[6][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][3]$_DFFE_PP_  (.D(net8),
    .DE(_023_),
    .Q(\mem[6][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][4]$_DFFE_PP_  (.D(net9),
    .DE(_023_),
    .Q(\mem[6][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][5]$_DFFE_PP_  (.D(net10),
    .DE(_023_),
    .Q(\mem[6][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][6]$_DFFE_PP_  (.D(net11),
    .DE(_023_),
    .Q(\mem[6][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][7]$_DFFE_PP_  (.D(net12),
    .DE(_023_),
    .Q(\mem[6][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][0]$_DFFE_PP_  (.D(net5),
    .DE(_024_),
    .Q(\mem[7][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][1]$_DFFE_PP_  (.D(net6),
    .DE(_024_),
    .Q(\mem[7][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][2]$_DFFE_PP_  (.D(net7),
    .DE(_024_),
    .Q(\mem[7][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][3]$_DFFE_PP_  (.D(net8),
    .DE(_024_),
    .Q(\mem[7][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][4]$_DFFE_PP_  (.D(net9),
    .DE(_024_),
    .Q(\mem[7][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][5]$_DFFE_PP_  (.D(net10),
    .DE(_024_),
    .Q(\mem[7][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][6]$_DFFE_PP_  (.D(net11),
    .DE(_024_),
    .Q(\mem[7][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][7]$_DFFE_PP_  (.D(net12),
    .DE(_024_),
    .Q(\mem[7][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][0]$_DFFE_PP_  (.D(net5),
    .DE(_025_),
    .Q(\mem[8][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][1]$_DFFE_PP_  (.D(net6),
    .DE(_025_),
    .Q(\mem[8][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][2]$_DFFE_PP_  (.D(net7),
    .DE(_025_),
    .Q(\mem[8][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][3]$_DFFE_PP_  (.D(net8),
    .DE(_025_),
    .Q(\mem[8][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][4]$_DFFE_PP_  (.D(net9),
    .DE(_025_),
    .Q(\mem[8][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][5]$_DFFE_PP_  (.D(net10),
    .DE(_025_),
    .Q(\mem[8][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][6]$_DFFE_PP_  (.D(net11),
    .DE(_025_),
    .Q(\mem[8][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][7]$_DFFE_PP_  (.D(net12),
    .DE(_025_),
    .Q(\mem[8][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][0]$_DFFE_PP_  (.D(net5),
    .DE(_026_),
    .Q(\mem[9][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][1]$_DFFE_PP_  (.D(net6),
    .DE(_026_),
    .Q(\mem[9][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][2]$_DFFE_PP_  (.D(net7),
    .DE(_026_),
    .Q(\mem[9][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][3]$_DFFE_PP_  (.D(net8),
    .DE(_026_),
    .Q(\mem[9][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][4]$_DFFE_PP_  (.D(net9),
    .DE(_026_),
    .Q(\mem[9][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][5]$_DFFE_PP_  (.D(net10),
    .DE(_026_),
    .Q(\mem[9][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][6]$_DFFE_PP_  (.D(net11),
    .DE(_026_),
    .Q(\mem[9][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][7]$_DFFE_PP_  (.D(net12),
    .DE(_026_),
    .Q(\mem[9][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \pointer_wraparound_error$_DFF_PN0_  (.D(_010_),
    .Q(net19),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_reg[0]$_DFFE_PN0P_  (.D(_031_),
    .Q(net25),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_reg[1]$_DFFE_PN0P_  (.D(_032_),
    .Q(net26),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_reg[2]$_DFFE_PN0P_  (.D(_033_),
    .Q(net27),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_reg[3]$_DFFE_PN0P_  (.D(_034_),
    .Q(net28),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_reg[4]$_DFFE_PN0P_  (.D(_035_),
    .Q(net29),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_reg[5]$_DFFE_PN0P_  (.D(_036_),
    .Q(net30),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_reg[6]$_DFFE_PN0P_  (.D(_037_),
    .Q(net31),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_reg[7]$_DFFE_PN0P_  (.D(_038_),
    .Q(net32),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_bin[0]$_DFFE_PN0P_  (.D(_039_),
    .Q(\rd_ptr_bin[0] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_bin[1]$_DFFE_PN0P_  (.D(_040_),
    .Q(\rd_ptr_bin[1] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_bin[2]$_DFFE_PN0P_  (.D(_041_),
    .Q(\rd_ptr_bin[2] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_bin[3]$_DFFE_PN0P_  (.D(_042_),
    .Q(\rd_ptr_bin[3] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray[0]$_DFFE_PN0P_  (.D(_043_),
    .Q(\rd_ptr_gray[0] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray[1]$_DFFE_PN0P_  (.D(_044_),
    .Q(\rd_ptr_gray[1] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray[2]$_DFFE_PN0P_  (.D(_045_),
    .Q(\rd_ptr_gray[2] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray[3]$_DFFE_PN0P_  (.D(_046_),
    .Q(\rd_ptr_gray[3] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_2 \rd_ptr_gray[4]$_DFFE_PN0P_  (.D(_047_),
    .Q(\rd_ptr_bin[4] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync1[0]$_DFF_PN0_  (.D(\rd_ptr_gray[0] ),
    .Q(\rd_ptr_gray_sync1[0] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync1[1]$_DFF_PN0_  (.D(\rd_ptr_gray[1] ),
    .Q(\rd_ptr_gray_sync1[1] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync1[2]$_DFF_PN0_  (.D(\rd_ptr_gray[2] ),
    .Q(\rd_ptr_gray_sync1[2] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync1[3]$_DFF_PN0_  (.D(\rd_ptr_gray[3] ),
    .Q(\rd_ptr_gray_sync1[3] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync1[4]$_DFF_PN0_  (.D(\rd_ptr_bin[4] ),
    .Q(\rd_ptr_gray_sync1[4] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync2[0]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[0] ),
    .Q(\rd_ptr_gray_sync2[0] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync2[1]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[1] ),
    .Q(\rd_ptr_gray_sync2[1] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync2[2]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[2] ),
    .Q(\rd_ptr_gray_sync2[2] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync2[3]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[3] ),
    .Q(\rd_ptr_gray_sync2[3] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync2[4]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[4] ),
    .Q(\rd_ptr_gray_sync2[4] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_sync[0]$_DFF_PN0_  (.D(_006_),
    .Q(\rd_ptr_sync[0] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_sync[1]$_DFF_PN0_  (.D(_007_),
    .Q(\rd_ptr_sync[1] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_sync[2]$_DFF_PN0_  (.D(_008_),
    .Q(\rd_ptr_sync[2] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_sync[3]$_DFF_PN0_  (.D(_009_),
    .Q(\rd_ptr_sync[3] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_sync[4]$_DFF_PN0_  (.D(\rd_ptr_gray_sync2[4] ),
    .Q(\rd_ptr_sync[4] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \sync_error$_DFF_PN0_  (.D(net39),
    .Q(net33),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_2 \wr_ptr_bin[0]$_DFFE_PN0P_  (.D(_048_),
    .Q(\wr_ptr_bin[0] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_2 \wr_ptr_bin[1]$_DFFE_PN0P_  (.D(_049_),
    .Q(\wr_ptr_bin[1] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_bin[2]$_DFFE_PN0P_  (.D(_050_),
    .Q(\wr_ptr_bin[2] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_bin[3]$_DFFE_PN0P_  (.D(_051_),
    .Q(\wr_ptr_bin[3] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray[0]$_DFFE_PN0P_  (.D(_052_),
    .Q(\wr_ptr_gray[0] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray[1]$_DFFE_PN0P_  (.D(_053_),
    .Q(\wr_ptr_gray[1] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray[2]$_DFFE_PN0P_  (.D(_054_),
    .Q(\wr_ptr_gray[2] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray[3]$_DFFE_PN0P_  (.D(_055_),
    .Q(\wr_ptr_gray[3] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray[4]$_DFFE_PN0P_  (.D(_056_),
    .Q(\wr_ptr_bin[4] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync1[0]$_DFF_PN0_  (.D(\wr_ptr_gray[0] ),
    .Q(\wr_ptr_gray_sync1[0] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync1[1]$_DFF_PN0_  (.D(\wr_ptr_gray[1] ),
    .Q(\wr_ptr_gray_sync1[1] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync1[2]$_DFF_PN0_  (.D(\wr_ptr_gray[2] ),
    .Q(\wr_ptr_gray_sync1[2] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync1[3]$_DFF_PN0_  (.D(\wr_ptr_gray[3] ),
    .Q(\wr_ptr_gray_sync1[3] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync1[4]$_DFF_PN0_  (.D(\wr_ptr_bin[4] ),
    .Q(\wr_ptr_gray_sync1[4] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync2[0]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[0] ),
    .Q(\wr_ptr_gray_sync2[0] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync2[1]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[1] ),
    .Q(\wr_ptr_gray_sync2[1] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync2[2]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[2] ),
    .Q(\wr_ptr_gray_sync2[2] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync2[3]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[3] ),
    .Q(\wr_ptr_gray_sync2[3] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync2[4]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[4] ),
    .Q(\wr_ptr_gray_sync2[4] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_sync[0]$_DFF_PN0_  (.D(_002_),
    .Q(\wr_ptr_sync[0] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_sync[1]$_DFF_PN0_  (.D(_003_),
    .Q(\wr_ptr_sync[1] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_sync[2]$_DFF_PN0_  (.D(_004_),
    .Q(\wr_ptr_sync[2] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_sync[3]$_DFF_PN0_  (.D(_005_),
    .Q(\wr_ptr_sync[3] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_sync[4]$_DFF_PN0_  (.D(\wr_ptr_gray_sync2[4] ),
    .Q(\wr_ptr_sync[4] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_175 ();
 sky130_fd_sc_hd__buf_8 input1 (.A(rd_clk),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(rd_en),
    .X(net2));
 sky130_fd_sc_hd__buf_12 input3 (.A(rd_rst_n),
    .X(net3));
 sky130_fd_sc_hd__buf_16 input4 (.A(wr_clk),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(wr_data[0]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input6 (.A(wr_data[1]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input7 (.A(wr_data[2]),
    .X(net7));
 sky130_fd_sc_hd__buf_6 input8 (.A(wr_data[3]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input9 (.A(wr_data[4]),
    .X(net9));
 sky130_fd_sc_hd__buf_4 input10 (.A(wr_data[5]),
    .X(net10));
 sky130_fd_sc_hd__buf_4 input11 (.A(wr_data[6]),
    .X(net11));
 sky130_fd_sc_hd__buf_4 input12 (.A(wr_data[7]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(wr_en),
    .X(net13));
 sky130_fd_sc_hd__buf_16 input14 (.A(wr_rst_n),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net15),
    .X(almost_empty));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net16),
    .X(almost_full));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net17),
    .X(empty));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net18),
    .X(full));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net19),
    .X(pointer_wraparound_flag));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net20),
    .X(rd_count[0]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net21),
    .X(rd_count[1]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net22),
    .X(rd_count[2]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net23),
    .X(rd_count[3]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net24),
    .X(rd_count[4]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net25),
    .X(rd_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net26),
    .X(rd_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net27),
    .X(rd_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net28),
    .X(rd_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(net29),
    .X(rd_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output30 (.A(net30),
    .X(rd_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(net31),
    .X(rd_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output32 (.A(net32),
    .X(rd_data[7]));
 sky130_fd_sc_hd__clkbuf_1 output33 (.A(net33),
    .X(sync_error_flag));
 sky130_fd_sc_hd__clkbuf_1 output34 (.A(net34),
    .X(wr_count[0]));
 sky130_fd_sc_hd__clkbuf_1 output35 (.A(net35),
    .X(wr_count[1]));
 sky130_fd_sc_hd__clkbuf_1 output36 (.A(net36),
    .X(wr_count[2]));
 sky130_fd_sc_hd__clkbuf_1 output37 (.A(net37),
    .X(wr_count[3]));
 sky130_fd_sc_hd__clkbuf_1 output38 (.A(net38),
    .X(wr_count[4]));
 sky130_fd_sc_hd__conb_1 \sync_error$_DFF_PN0__39  (.HI(net39));
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_173 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_34 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_240 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_143 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_74 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_126 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_94 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_224 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_53 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_253 ();
endmodule
