module multi_phase_pwm_controller (clk,
    enable,
    rst_n,
    deadtime,
    duty,
    pwm_n_out,
    pwm_p_out);
 input clk;
 input enable;
 input rst_n;
 input [5:0] deadtime;
 input [7:0] duty;
 output [2:0] pwm_n_out;
 output [2:0] pwm_p_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire _433_;
 wire _434_;
 wire _435_;
 wire _436_;
 wire _437_;
 wire _438_;
 wire _439_;
 wire _440_;
 wire _441_;
 wire _442_;
 wire _443_;
 wire _444_;
 wire _445_;
 wire _446_;
 wire _447_;
 wire _448_;
 wire _449_;
 wire _450_;
 wire _451_;
 wire _452_;
 wire _453_;
 wire _454_;
 wire _455_;
 wire _456_;
 wire _457_;
 wire _458_;
 wire _459_;
 wire _460_;
 wire _461_;
 wire _462_;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 sky130_fd_sc_hd__inv_1 _463_ (.A(net13),
    .Y(_448_));
 sky130_fd_sc_hd__inv_1 _464_ (.A(_294_),
    .Y(_214_));
 sky130_fd_sc_hd__inv_2 _465_ (.A(net14),
    .Y(_445_));
 sky130_fd_sc_hd__buf_4 _466_ (.A(\counter[4] ),
    .X(_014_));
 sky130_fd_sc_hd__clkinv_4 _467_ (.A(_014_),
    .Y(_237_));
 sky130_fd_sc_hd__inv_2 _468_ (.A(\counter[6] ),
    .Y(_229_));
 sky130_fd_sc_hd__clkbuf_4 _469_ (.A(\counter[2] ),
    .X(_015_));
 sky130_fd_sc_hd__inv_1 _470_ (.A(_015_),
    .Y(_245_));
 sky130_fd_sc_hd__a211oi_2 _471_ (.A1(\counter[0] ),
    .A2(_378_),
    .B1(_015_),
    .C1(_014_),
    .Y(_016_));
 sky130_fd_sc_hd__clkbuf_4 _472_ (.A(\counter[3] ),
    .X(_017_));
 sky130_fd_sc_hd__o21ai_1 _473_ (.A1(_014_),
    .A2(_017_),
    .B1(\counter[5] ),
    .Y(_018_));
 sky130_fd_sc_hd__o21ai_1 _474_ (.A1(_016_),
    .A2(_018_),
    .B1(_229_),
    .Y(_019_));
 sky130_fd_sc_hd__xnor2_2 _475_ (.A(\counter[7] ),
    .B(_019_),
    .Y(_310_));
 sky130_fd_sc_hd__o21a_1 _476_ (.A1(_015_),
    .A2(_328_),
    .B1(_017_),
    .X(_020_));
 sky130_fd_sc_hd__o21ai_1 _477_ (.A1(_014_),
    .A2(_020_),
    .B1(\counter[5] ),
    .Y(_021_));
 sky130_fd_sc_hd__xnor2_2 _478_ (.A(\counter[6] ),
    .B(_021_),
    .Y(_313_));
 sky130_fd_sc_hd__clkinv_4 _479_ (.A(_017_),
    .Y(_241_));
 sky130_fd_sc_hd__a21oi_2 _480_ (.A1(\counter[0] ),
    .A2(_378_),
    .B1(_015_),
    .Y(_022_));
 sky130_fd_sc_hd__clkinv_4 _481_ (.A(\counter[5] ),
    .Y(_233_));
 sky130_fd_sc_hd__o211ai_2 _482_ (.A1(_241_),
    .A2(_022_),
    .B1(_233_),
    .C1(_237_),
    .Y(_023_));
 sky130_fd_sc_hd__o21ai_4 _483_ (.A1(_016_),
    .A2(_018_),
    .B1(_023_),
    .Y(_316_));
 sky130_fd_sc_hd__xnor2_4 _484_ (.A(_237_),
    .B(_020_),
    .Y(_319_));
 sky130_fd_sc_hd__xnor2_4 _485_ (.A(_241_),
    .B(_022_),
    .Y(_322_));
 sky130_fd_sc_hd__xor2_2 _486_ (.A(_015_),
    .B(_328_),
    .X(_325_));
 sky130_fd_sc_hd__inv_1 _487_ (.A(\counter[7] ),
    .Y(_225_));
 sky130_fd_sc_hd__nor2_1 _488_ (.A(_017_),
    .B(_380_),
    .Y(_024_));
 sky130_fd_sc_hd__nor2_2 _489_ (.A(_237_),
    .B(_024_),
    .Y(_025_));
 sky130_fd_sc_hd__o21ai_0 _490_ (.A1(\counter[5] ),
    .A2(_025_),
    .B1(\counter[6] ),
    .Y(_026_));
 sky130_fd_sc_hd__xnor2_1 _491_ (.A(_225_),
    .B(_026_),
    .Y(_027_));
 sky130_fd_sc_hd__inv_1 _492_ (.A(_027_),
    .Y(_363_));
 sky130_fd_sc_hd__a21o_2 _493_ (.A1(_015_),
    .A2(\counter[1] ),
    .B1(_017_),
    .X(_028_));
 sky130_fd_sc_hd__a21oi_2 _494_ (.A1(_014_),
    .A2(_028_),
    .B1(\counter[5] ),
    .Y(_029_));
 sky130_fd_sc_hd__xnor2_4 _495_ (.A(_229_),
    .B(_029_),
    .Y(_366_));
 sky130_fd_sc_hd__xnor2_4 _496_ (.A(_233_),
    .B(_025_),
    .Y(_369_));
 sky130_fd_sc_hd__xnor2_4 _497_ (.A(_014_),
    .B(_028_),
    .Y(_372_));
 sky130_fd_sc_hd__xor2_4 _498_ (.A(_017_),
    .B(_380_),
    .X(_375_));
 sky130_fd_sc_hd__inv_1 _499_ (.A(\counter[0] ),
    .Y(_297_));
 sky130_fd_sc_hd__inv_1 _500_ (.A(net6),
    .Y(_252_));
 sky130_fd_sc_hd__inv_1 _501_ (.A(net5),
    .Y(_257_));
 sky130_fd_sc_hd__inv_1 _502_ (.A(net4),
    .Y(_262_));
 sky130_fd_sc_hd__inv_1 _503_ (.A(net3),
    .Y(_220_));
 sky130_fd_sc_hd__inv_1 _504_ (.A(\counter[1] ),
    .Y(_288_));
 sky130_fd_sc_hd__clkbuf_4 _505_ (.A(_254_),
    .X(_030_));
 sky130_fd_sc_hd__nand2_1 _506_ (.A(net13),
    .B(_445_),
    .Y(_031_));
 sky130_fd_sc_hd__clkinvlp_4 _507_ (.A(_259_),
    .Y(_032_));
 sky130_fd_sc_hd__clkinvlp_4 _508_ (.A(_264_),
    .Y(_033_));
 sky130_fd_sc_hd__a21o_1 _509_ (.A1(_033_),
    .A2(_223_),
    .B1(_265_),
    .X(_034_));
 sky130_fd_sc_hd__nor2_1 _510_ (.A(_259_),
    .B(_264_),
    .Y(_035_));
 sky130_fd_sc_hd__inv_1 _511_ (.A(_268_),
    .Y(_036_));
 sky130_fd_sc_hd__nand2b_1 _512_ (.A_N(_249_),
    .B(_217_),
    .Y(_037_));
 sky130_fd_sc_hd__a21oi_2 _513_ (.A1(_036_),
    .A2(_037_),
    .B1(_222_),
    .Y(_038_));
 sky130_fd_sc_hd__a22oi_2 _514_ (.A1(_032_),
    .A2(_034_),
    .B1(_035_),
    .B2(_038_),
    .Y(_039_));
 sky130_fd_sc_hd__or3_1 _515_ (.A(_260_),
    .B(_445_),
    .C(_255_),
    .X(_040_));
 sky130_fd_sc_hd__a221o_1 _516_ (.A1(_032_),
    .A2(_034_),
    .B1(_035_),
    .B2(_038_),
    .C1(_040_),
    .X(_041_));
 sky130_fd_sc_hd__inv_1 _517_ (.A(_030_),
    .Y(_042_));
 sky130_fd_sc_hd__a21oi_1 _518_ (.A1(_042_),
    .A2(_260_),
    .B1(_255_),
    .Y(_043_));
 sky130_fd_sc_hd__o21ai_0 _519_ (.A1(_042_),
    .A2(_255_),
    .B1(net13),
    .Y(_044_));
 sky130_fd_sc_hd__a2bb2oi_1 _520_ (.A1_N(_031_),
    .A2_N(_043_),
    .B1(_044_),
    .B2(net14),
    .Y(_045_));
 sky130_fd_sc_hd__o311ai_4 _521_ (.A1(_030_),
    .A2(_031_),
    .A3(_039_),
    .B1(_041_),
    .C1(_045_),
    .Y(_270_));
 sky130_fd_sc_hd__inv_1 _522_ (.A(_329_),
    .Y(_330_));
 sky130_fd_sc_hd__inv_1 _523_ (.A(_221_),
    .Y(_046_));
 sky130_fd_sc_hd__nor2b_1 _524_ (.A(_294_),
    .B_N(_249_),
    .Y(_047_));
 sky130_fd_sc_hd__o21ai_1 _525_ (.A1(_267_),
    .A2(_047_),
    .B1(_222_),
    .Y(_048_));
 sky130_fd_sc_hd__a21oi_1 _526_ (.A1(_046_),
    .A2(_048_),
    .B1(_033_),
    .Y(_049_));
 sky130_fd_sc_hd__o21ai_1 _527_ (.A1(_263_),
    .A2(_049_),
    .B1(_259_),
    .Y(_050_));
 sky130_fd_sc_hd__nor3_1 _528_ (.A(net13),
    .B(_253_),
    .C(_258_),
    .Y(_051_));
 sky130_fd_sc_hd__nor3_1 _529_ (.A(net13),
    .B(_030_),
    .C(_253_),
    .Y(_052_));
 sky130_fd_sc_hd__a21oi_1 _530_ (.A1(_050_),
    .A2(_051_),
    .B1(_052_),
    .Y(_053_));
 sky130_fd_sc_hd__xnor2_2 _531_ (.A(net14),
    .B(_053_),
    .Y(_226_));
 sky130_fd_sc_hd__a21oi_1 _532_ (.A1(_222_),
    .A2(_215_),
    .B1(_221_),
    .Y(_054_));
 sky130_fd_sc_hd__nor2_1 _533_ (.A(_033_),
    .B(_054_),
    .Y(_055_));
 sky130_fd_sc_hd__nor2_1 _534_ (.A(_263_),
    .B(_055_),
    .Y(_056_));
 sky130_fd_sc_hd__o21bai_1 _535_ (.A1(_032_),
    .A2(_056_),
    .B1_N(_258_),
    .Y(_057_));
 sky130_fd_sc_hd__a21oi_1 _536_ (.A1(_030_),
    .A2(_057_),
    .B1(_253_),
    .Y(_058_));
 sky130_fd_sc_hd__xnor2_1 _537_ (.A(_448_),
    .B(_058_),
    .Y(_230_));
 sky130_fd_sc_hd__nor2b_1 _538_ (.A(_258_),
    .B_N(_050_),
    .Y(_059_));
 sky130_fd_sc_hd__xnor2_2 _539_ (.A(_030_),
    .B(_059_),
    .Y(_234_));
 sky130_fd_sc_hd__xnor2_2 _540_ (.A(_259_),
    .B(_056_),
    .Y(_238_));
 sky130_fd_sc_hd__and3_1 _541_ (.A(_033_),
    .B(_046_),
    .C(_048_),
    .X(_060_));
 sky130_fd_sc_hd__nor2_1 _542_ (.A(_049_),
    .B(_060_),
    .Y(_242_));
 sky130_fd_sc_hd__xor2_2 _543_ (.A(_222_),
    .B(_215_),
    .X(_246_));
 sky130_fd_sc_hd__inv_1 _544_ (.A(_260_),
    .Y(_061_));
 sky130_fd_sc_hd__nor2b_1 _545_ (.A(_222_),
    .B_N(_218_),
    .Y(_062_));
 sky130_fd_sc_hd__o21a_1 _546_ (.A1(_223_),
    .A2(_062_),
    .B1(_033_),
    .X(_063_));
 sky130_fd_sc_hd__o21ai_0 _547_ (.A1(_265_),
    .A2(_063_),
    .B1(_032_),
    .Y(_064_));
 sky130_fd_sc_hd__a21oi_1 _548_ (.A1(_061_),
    .A2(_064_),
    .B1(_030_),
    .Y(_065_));
 sky130_fd_sc_hd__nor2_1 _549_ (.A(_255_),
    .B(_065_),
    .Y(_066_));
 sky130_fd_sc_hd__xnor2_2 _550_ (.A(net13),
    .B(_066_),
    .Y(_273_));
 sky130_fd_sc_hd__nand2_1 _551_ (.A(_061_),
    .B(_039_),
    .Y(_067_));
 sky130_fd_sc_hd__xnor2_2 _552_ (.A(_030_),
    .B(_067_),
    .Y(_276_));
 sky130_fd_sc_hd__nor2_1 _553_ (.A(_265_),
    .B(_063_),
    .Y(_068_));
 sky130_fd_sc_hd__xnor2_2 _554_ (.A(_032_),
    .B(_068_),
    .Y(_279_));
 sky130_fd_sc_hd__nor2_1 _555_ (.A(_223_),
    .B(_038_),
    .Y(_069_));
 sky130_fd_sc_hd__xnor2_2 _556_ (.A(_033_),
    .B(_069_),
    .Y(_282_));
 sky130_fd_sc_hd__xnor2_2 _557_ (.A(_222_),
    .B(_218_),
    .Y(_285_));
 sky130_fd_sc_hd__clkinvlp_4 _558_ (.A(net2),
    .Y(_213_));
 sky130_fd_sc_hd__inv_1 _559_ (.A(net8),
    .Y(_420_));
 sky130_fd_sc_hd__inv_1 _560_ (.A(net7),
    .Y(_293_));
 sky130_fd_sc_hd__inv_1 _561_ (.A(net12),
    .Y(_451_));
 sky130_fd_sc_hd__inv_1 _562_ (.A(net11),
    .Y(_454_));
 sky130_fd_sc_hd__inv_1 _563_ (.A(net10),
    .Y(_457_));
 sky130_fd_sc_hd__inv_1 _564_ (.A(net9),
    .Y(_460_));
 sky130_fd_sc_hd__nand2_1 _565_ (.A(\counter[6] ),
    .B(\counter[7] ),
    .Y(_070_));
 sky130_fd_sc_hd__nand2_1 _566_ (.A(\counter[5] ),
    .B(_014_),
    .Y(_071_));
 sky130_fd_sc_hd__clkbuf_4 _567_ (.A(enable),
    .X(_072_));
 sky130_fd_sc_hd__nand4_4 _568_ (.A(_072_),
    .B(_017_),
    .C(_015_),
    .D(_328_),
    .Y(_073_));
 sky130_fd_sc_hd__o31ai_4 _569_ (.A1(_070_),
    .A2(_071_),
    .A3(_073_),
    .B1(net15),
    .Y(_074_));
 sky130_fd_sc_hd__xnor2_1 _570_ (.A(_072_),
    .B(\counter[0] ),
    .Y(_075_));
 sky130_fd_sc_hd__nor2_1 _571_ (.A(_074_),
    .B(_075_),
    .Y(_000_));
 sky130_fd_sc_hd__mux2i_1 _572_ (.A0(\counter[1] ),
    .A1(_329_),
    .S(_072_),
    .Y(_076_));
 sky130_fd_sc_hd__nor2_1 _573_ (.A(_074_),
    .B(_076_),
    .Y(_001_));
 sky130_fd_sc_hd__nand2_1 _574_ (.A(_072_),
    .B(_328_),
    .Y(_077_));
 sky130_fd_sc_hd__xnor2_1 _575_ (.A(_015_),
    .B(_077_),
    .Y(_078_));
 sky130_fd_sc_hd__and2_0 _576_ (.A(net15),
    .B(_078_),
    .X(_002_));
 sky130_fd_sc_hd__nand3_1 _577_ (.A(_072_),
    .B(\counter[0] ),
    .C(_380_),
    .Y(_079_));
 sky130_fd_sc_hd__xnor2_1 _578_ (.A(_241_),
    .B(_079_),
    .Y(_080_));
 sky130_fd_sc_hd__nor2_1 _579_ (.A(_074_),
    .B(_080_),
    .Y(_003_));
 sky130_fd_sc_hd__xnor2_1 _580_ (.A(_014_),
    .B(_073_),
    .Y(_081_));
 sky130_fd_sc_hd__and2_0 _581_ (.A(net15),
    .B(_081_),
    .X(_004_));
 sky130_fd_sc_hd__nor3_1 _582_ (.A(_237_),
    .B(_241_),
    .C(_079_),
    .Y(_082_));
 sky130_fd_sc_hd__xnor2_1 _583_ (.A(\counter[5] ),
    .B(_082_),
    .Y(_083_));
 sky130_fd_sc_hd__nor2_1 _584_ (.A(_074_),
    .B(_083_),
    .Y(_005_));
 sky130_fd_sc_hd__o21ai_0 _585_ (.A1(_071_),
    .A2(_073_),
    .B1(\counter[6] ),
    .Y(_084_));
 sky130_fd_sc_hd__or3_1 _586_ (.A(\counter[6] ),
    .B(_071_),
    .C(_073_),
    .X(_085_));
 sky130_fd_sc_hd__a21boi_0 _587_ (.A1(_084_),
    .A2(_085_),
    .B1_N(net15),
    .Y(_006_));
 sky130_fd_sc_hd__nor4_1 _588_ (.A(_229_),
    .B(_241_),
    .C(_071_),
    .D(_079_),
    .Y(_086_));
 sky130_fd_sc_hd__xnor2_1 _589_ (.A(\counter[7] ),
    .B(_086_),
    .Y(_087_));
 sky130_fd_sc_hd__nor2_1 _590_ (.A(_074_),
    .B(_087_),
    .Y(_007_));
 sky130_fd_sc_hd__nand4_2 _591_ (.A(_228_),
    .B(_232_),
    .C(_236_),
    .D(_240_),
    .Y(_088_));
 sky130_fd_sc_hd__nand2_1 _592_ (.A(_244_),
    .B(_248_),
    .Y(_089_));
 sky130_fd_sc_hd__o21bai_1 _593_ (.A1(_335_),
    .A2(_251_),
    .B1_N(_384_),
    .Y(_090_));
 sky130_fd_sc_hd__a21o_1 _594_ (.A1(_248_),
    .A2(_090_),
    .B1(_247_),
    .X(_091_));
 sky130_fd_sc_hd__a21oi_1 _595_ (.A1(_244_),
    .A2(_091_),
    .B1(_243_),
    .Y(_092_));
 sky130_fd_sc_hd__a21o_1 _596_ (.A1(_239_),
    .A2(_236_),
    .B1(_235_),
    .X(_093_));
 sky130_fd_sc_hd__a21o_1 _597_ (.A1(_232_),
    .A2(_093_),
    .B1(_231_),
    .X(_094_));
 sky130_fd_sc_hd__a21oi_1 _598_ (.A1(_228_),
    .A2(_094_),
    .B1(_227_),
    .Y(_095_));
 sky130_fd_sc_hd__o21ai_0 _599_ (.A1(_088_),
    .A2(_092_),
    .B1(_095_),
    .Y(_096_));
 sky130_fd_sc_hd__o41ai_1 _600_ (.A1(_251_),
    .A2(_334_),
    .A3(_088_),
    .A4(_089_),
    .B1(_096_),
    .Y(_097_));
 sky130_fd_sc_hd__nor2b_1 _601_ (.A(_300_),
    .B_N(_290_),
    .Y(_098_));
 sky130_fd_sc_hd__o21ai_0 _602_ (.A1(_289_),
    .A2(_098_),
    .B1(_287_),
    .Y(_099_));
 sky130_fd_sc_hd__nand2b_1 _603_ (.A_N(_286_),
    .B(_099_),
    .Y(_100_));
 sky130_fd_sc_hd__a21oi_1 _604_ (.A1(_284_),
    .A2(_100_),
    .B1(_283_),
    .Y(_101_));
 sky130_fd_sc_hd__nand4_1 _605_ (.A(_272_),
    .B(_275_),
    .C(_278_),
    .D(_281_),
    .Y(_102_));
 sky130_fd_sc_hd__nand4b_1 _606_ (.A_N(_299_),
    .B(_287_),
    .C(_284_),
    .D(_290_),
    .Y(_103_));
 sky130_fd_sc_hd__nand2b_1 _607_ (.A_N(_102_),
    .B(_103_),
    .Y(_104_));
 sky130_fd_sc_hd__nor2b_1 _608_ (.A(_361_),
    .B_N(_405_),
    .Y(_105_));
 sky130_fd_sc_hd__o21ai_0 _609_ (.A1(_404_),
    .A2(_105_),
    .B1(_309_),
    .Y(_106_));
 sky130_fd_sc_hd__nor2_1 _610_ (.A(_306_),
    .B(_308_),
    .Y(_107_));
 sky130_fd_sc_hd__o21ai_0 _611_ (.A1(_307_),
    .A2(_306_),
    .B1(_305_),
    .Y(_108_));
 sky130_fd_sc_hd__a21oi_1 _612_ (.A1(_106_),
    .A2(_107_),
    .B1(_108_),
    .Y(_109_));
 sky130_fd_sc_hd__and4b_1 _613_ (.A_N(_360_),
    .B(_305_),
    .C(_309_),
    .D(_307_),
    .X(_110_));
 sky130_fd_sc_hd__nor2_1 _614_ (.A(_303_),
    .B(_302_),
    .Y(_111_));
 sky130_fd_sc_hd__a31oi_1 _615_ (.A1(_405_),
    .A2(_303_),
    .A3(_110_),
    .B1(_111_),
    .Y(_112_));
 sky130_fd_sc_hd__o31a_1 _616_ (.A1(_304_),
    .A2(_302_),
    .A3(_109_),
    .B1(_112_),
    .X(_113_));
 sky130_fd_sc_hd__a21o_1 _617_ (.A1(_280_),
    .A2(_278_),
    .B1(_277_),
    .X(_114_));
 sky130_fd_sc_hd__a21oi_1 _618_ (.A1(_275_),
    .A2(_114_),
    .B1(_274_),
    .Y(_115_));
 sky130_fd_sc_hd__nor2b_1 _619_ (.A(_115_),
    .B_N(_272_),
    .Y(_116_));
 sky130_fd_sc_hd__o22ai_1 _620_ (.A1(_102_),
    .A2(_103_),
    .B1(_116_),
    .B2(_271_),
    .Y(_117_));
 sky130_fd_sc_hd__o221ai_1 _621_ (.A1(_101_),
    .A2(_104_),
    .B1(_113_),
    .B2(_070_),
    .C1(_117_),
    .Y(_118_));
 sky130_fd_sc_hd__nand2_2 _622_ (.A(net15),
    .B(_072_),
    .Y(_119_));
 sky130_fd_sc_hd__a21oi_1 _623_ (.A1(_097_),
    .A2(_118_),
    .B1(_119_),
    .Y(_008_));
 sky130_fd_sc_hd__nand4_1 _624_ (.A(_312_),
    .B(_315_),
    .C(_318_),
    .D(_321_),
    .Y(_120_));
 sky130_fd_sc_hd__nand4_1 _625_ (.A(_334_),
    .B(_324_),
    .C(_327_),
    .D(_332_),
    .Y(_121_));
 sky130_fd_sc_hd__nor2_1 _626_ (.A(_120_),
    .B(_121_),
    .Y(_122_));
 sky130_fd_sc_hd__nor2b_1 _627_ (.A(_333_),
    .B_N(_332_),
    .Y(_123_));
 sky130_fd_sc_hd__o21ai_0 _628_ (.A1(_331_),
    .A2(_123_),
    .B1(_327_),
    .Y(_124_));
 sky130_fd_sc_hd__nand2b_1 _629_ (.A_N(_326_),
    .B(_124_),
    .Y(_125_));
 sky130_fd_sc_hd__a21oi_1 _630_ (.A1(_324_),
    .A2(_125_),
    .B1(_323_),
    .Y(_126_));
 sky130_fd_sc_hd__a21o_1 _631_ (.A1(_320_),
    .A2(_318_),
    .B1(_317_),
    .X(_127_));
 sky130_fd_sc_hd__a21oi_1 _632_ (.A1(_315_),
    .A2(_127_),
    .B1(_314_),
    .Y(_128_));
 sky130_fd_sc_hd__nor2b_1 _633_ (.A(_128_),
    .B_N(_312_),
    .Y(_129_));
 sky130_fd_sc_hd__o22ai_1 _634_ (.A1(_120_),
    .A2(_121_),
    .B1(_129_),
    .B2(_311_),
    .Y(_130_));
 sky130_fd_sc_hd__o31ai_1 _635_ (.A1(_120_),
    .A2(_122_),
    .A3(_126_),
    .B1(_130_),
    .Y(_131_));
 sky130_fd_sc_hd__nand4_1 _636_ (.A(_344_),
    .B(_340_),
    .C(_342_),
    .D(_346_),
    .Y(_132_));
 sky130_fd_sc_hd__nand3_1 _637_ (.A(_299_),
    .B(_348_),
    .C(_338_),
    .Y(_133_));
 sky130_fd_sc_hd__inv_1 _638_ (.A(_298_),
    .Y(_134_));
 sky130_fd_sc_hd__a21oi_1 _639_ (.A1(_348_),
    .A2(_134_),
    .B1(_347_),
    .Y(_135_));
 sky130_fd_sc_hd__a21o_1 _640_ (.A1(_342_),
    .A2(_343_),
    .B1(_341_),
    .X(_136_));
 sky130_fd_sc_hd__and4_1 _641_ (.A(_344_),
    .B(_340_),
    .C(_342_),
    .D(_345_),
    .X(_137_));
 sky130_fd_sc_hd__a2111oi_0 _642_ (.A1(_340_),
    .A2(_136_),
    .B1(_137_),
    .C1(_337_),
    .D1(_339_),
    .Y(_138_));
 sky130_fd_sc_hd__o21ai_0 _643_ (.A1(_132_),
    .A2(_135_),
    .B1(_138_),
    .Y(_139_));
 sky130_fd_sc_hd__o221a_1 _644_ (.A1(_338_),
    .A2(_337_),
    .B1(_132_),
    .B2(_133_),
    .C1(_139_),
    .X(_140_));
 sky130_fd_sc_hd__nor2b_1 _645_ (.A(_359_),
    .B_N(_358_),
    .Y(_141_));
 sky130_fd_sc_hd__nand3_1 _646_ (.A(_354_),
    .B(_352_),
    .C(_356_),
    .Y(_142_));
 sky130_fd_sc_hd__o21bai_1 _647_ (.A1(_357_),
    .A2(_141_),
    .B1_N(_142_),
    .Y(_143_));
 sky130_fd_sc_hd__a21o_1 _648_ (.A1(_354_),
    .A2(_355_),
    .B1(_353_),
    .X(_144_));
 sky130_fd_sc_hd__nand2_1 _649_ (.A(_352_),
    .B(_144_),
    .Y(_145_));
 sky130_fd_sc_hd__nor2_1 _650_ (.A(_351_),
    .B(_349_),
    .Y(_146_));
 sky130_fd_sc_hd__nand3_1 _651_ (.A(_360_),
    .B(_350_),
    .C(_358_),
    .Y(_147_));
 sky130_fd_sc_hd__o22ai_1 _652_ (.A1(_350_),
    .A2(_349_),
    .B1(_142_),
    .B2(_147_),
    .Y(_148_));
 sky130_fd_sc_hd__a31oi_1 _653_ (.A1(_143_),
    .A2(_145_),
    .A3(_146_),
    .B1(_148_),
    .Y(_149_));
 sky130_fd_sc_hd__nor2_1 _654_ (.A(_313_),
    .B(_149_),
    .Y(_150_));
 sky130_fd_sc_hd__a211oi_1 _655_ (.A1(_270_),
    .A2(_140_),
    .B1(_150_),
    .C1(_310_),
    .Y(_151_));
 sky130_fd_sc_hd__nor3b_1 _656_ (.A(_270_),
    .B(_140_),
    .C_N(_310_),
    .Y(_152_));
 sky130_fd_sc_hd__o311a_1 _657_ (.A1(_131_),
    .A2(_151_),
    .A3(_152_),
    .B1(_072_),
    .C1(net15),
    .X(_009_));
 sky130_fd_sc_hd__nand4_1 _658_ (.A(_365_),
    .B(_368_),
    .C(_371_),
    .D(_374_),
    .Y(_153_));
 sky130_fd_sc_hd__or4bb_1 _659_ (.A(_334_),
    .B(_385_),
    .C_N(_383_),
    .D_N(_377_),
    .X(_154_));
 sky130_fd_sc_hd__o21bai_1 _660_ (.A1(_335_),
    .A2(_385_),
    .B1_N(_250_),
    .Y(_155_));
 sky130_fd_sc_hd__a21o_1 _661_ (.A1(_383_),
    .A2(_155_),
    .B1(_382_),
    .X(_156_));
 sky130_fd_sc_hd__a21oi_1 _662_ (.A1(_377_),
    .A2(_156_),
    .B1(_376_),
    .Y(_157_));
 sky130_fd_sc_hd__a21o_1 _663_ (.A1(_373_),
    .A2(_371_),
    .B1(_370_),
    .X(_158_));
 sky130_fd_sc_hd__a21o_1 _664_ (.A1(_368_),
    .A2(_158_),
    .B1(_367_),
    .X(_159_));
 sky130_fd_sc_hd__a21oi_1 _665_ (.A1(_365_),
    .A2(_159_),
    .B1(_364_),
    .Y(_160_));
 sky130_fd_sc_hd__o21ai_0 _666_ (.A1(_153_),
    .A2(_157_),
    .B1(_160_),
    .Y(_161_));
 sky130_fd_sc_hd__o21ai_0 _667_ (.A1(_153_),
    .A2(_154_),
    .B1(_161_),
    .Y(_162_));
 sky130_fd_sc_hd__nand4_1 _668_ (.A(_393_),
    .B(_389_),
    .C(_391_),
    .D(_395_),
    .Y(_163_));
 sky130_fd_sc_hd__or4b_1 _669_ (.A(_290_),
    .B(_163_),
    .C(_299_),
    .D_N(_387_),
    .X(_164_));
 sky130_fd_sc_hd__nor2_1 _670_ (.A(_290_),
    .B(_300_),
    .Y(_165_));
 sky130_fd_sc_hd__nor2_1 _671_ (.A(_291_),
    .B(_165_),
    .Y(_166_));
 sky130_fd_sc_hd__a211oi_1 _672_ (.A1(_393_),
    .A2(_394_),
    .B1(_392_),
    .C1(_390_),
    .Y(_167_));
 sky130_fd_sc_hd__o21ai_0 _673_ (.A1(_390_),
    .A2(_391_),
    .B1(_389_),
    .Y(_168_));
 sky130_fd_sc_hd__inv_1 _674_ (.A(_388_),
    .Y(_169_));
 sky130_fd_sc_hd__o221ai_1 _675_ (.A1(_163_),
    .A2(_166_),
    .B1(_167_),
    .B2(_168_),
    .C1(_169_),
    .Y(_170_));
 sky130_fd_sc_hd__a21o_1 _676_ (.A1(_387_),
    .A2(_170_),
    .B1(_386_),
    .X(_171_));
 sky130_fd_sc_hd__a211o_1 _677_ (.A1(_164_),
    .A2(_171_),
    .B1(_027_),
    .C1(_270_),
    .X(_172_));
 sky130_fd_sc_hd__nand3b_1 _678_ (.A_N(_405_),
    .B(_403_),
    .C(_401_),
    .Y(_173_));
 sky130_fd_sc_hd__a21o_1 _679_ (.A1(_403_),
    .A2(_406_),
    .B1(_402_),
    .X(_174_));
 sky130_fd_sc_hd__a211o_1 _680_ (.A1(_398_),
    .A2(_397_),
    .B1(_396_),
    .C1(_400_),
    .X(_175_));
 sky130_fd_sc_hd__a21oi_1 _681_ (.A1(_401_),
    .A2(_174_),
    .B1(_175_),
    .Y(_176_));
 sky130_fd_sc_hd__o21ai_0 _682_ (.A1(_361_),
    .A2(_173_),
    .B1(_176_),
    .Y(_177_));
 sky130_fd_sc_hd__nand3b_1 _683_ (.A_N(_360_),
    .B(_397_),
    .C(_399_),
    .Y(_178_));
 sky130_fd_sc_hd__o21a_1 _684_ (.A1(_398_),
    .A2(_399_),
    .B1(_397_),
    .X(_179_));
 sky130_fd_sc_hd__o22a_1 _685_ (.A1(_173_),
    .A2(_178_),
    .B1(_179_),
    .B2(_396_),
    .X(_180_));
 sky130_fd_sc_hd__a21oi_1 _686_ (.A1(_177_),
    .A2(_180_),
    .B1(_366_),
    .Y(_181_));
 sky130_fd_sc_hd__a311o_1 _687_ (.A1(_270_),
    .A2(_164_),
    .A3(_171_),
    .B1(_181_),
    .C1(_363_),
    .X(_182_));
 sky130_fd_sc_hd__a31oi_1 _688_ (.A1(_162_),
    .A2(_172_),
    .A3(_182_),
    .B1(_119_),
    .Y(_010_));
 sky130_fd_sc_hd__nor2b_1 _689_ (.A(_441_),
    .B_N(_422_),
    .Y(_183_));
 sky130_fd_sc_hd__o21ai_0 _690_ (.A1(_421_),
    .A2(_183_),
    .B1(_462_),
    .Y(_184_));
 sky130_fd_sc_hd__nand2b_1 _691_ (.A_N(_461_),
    .B(_184_),
    .Y(_185_));
 sky130_fd_sc_hd__a21oi_1 _692_ (.A1(_459_),
    .A2(_185_),
    .B1(_458_),
    .Y(_186_));
 sky130_fd_sc_hd__nand2_1 _693_ (.A(_453_),
    .B(_456_),
    .Y(_187_));
 sky130_fd_sc_hd__a21oi_1 _694_ (.A1(_455_),
    .A2(_453_),
    .B1(_452_),
    .Y(_188_));
 sky130_fd_sc_hd__o21ai_0 _695_ (.A1(_186_),
    .A2(_187_),
    .B1(_188_),
    .Y(_189_));
 sky130_fd_sc_hd__a211o_1 _696_ (.A1(_447_),
    .A2(_449_),
    .B1(_119_),
    .C1(_446_),
    .X(_190_));
 sky130_fd_sc_hd__a31oi_1 _697_ (.A1(_447_),
    .A2(_450_),
    .A3(_189_),
    .B1(_190_),
    .Y(_011_));
 sky130_fd_sc_hd__nand4_1 _698_ (.A(_426_),
    .B(_430_),
    .C(_432_),
    .D(_428_),
    .Y(_191_));
 sky130_fd_sc_hd__nand4_1 _699_ (.A(_440_),
    .B(_434_),
    .C(_436_),
    .D(_438_),
    .Y(_192_));
 sky130_fd_sc_hd__nor2_1 _700_ (.A(_191_),
    .B(_192_),
    .Y(_193_));
 sky130_fd_sc_hd__nor2b_1 _701_ (.A(_439_),
    .B_N(_438_),
    .Y(_194_));
 sky130_fd_sc_hd__o21ai_0 _702_ (.A1(_437_),
    .A2(_194_),
    .B1(_436_),
    .Y(_195_));
 sky130_fd_sc_hd__nand2b_1 _703_ (.A_N(_435_),
    .B(_195_),
    .Y(_196_));
 sky130_fd_sc_hd__a21oi_1 _704_ (.A1(_434_),
    .A2(_196_),
    .B1(_433_),
    .Y(_197_));
 sky130_fd_sc_hd__a21o_1 _705_ (.A1(_430_),
    .A2(_431_),
    .B1(_429_),
    .X(_198_));
 sky130_fd_sc_hd__a21o_1 _706_ (.A1(_428_),
    .A2(_198_),
    .B1(_427_),
    .X(_199_));
 sky130_fd_sc_hd__a21oi_1 _707_ (.A1(_426_),
    .A2(_199_),
    .B1(_425_),
    .Y(_200_));
 sky130_fd_sc_hd__o21ai_0 _708_ (.A1(_191_),
    .A2(_197_),
    .B1(_200_),
    .Y(_201_));
 sky130_fd_sc_hd__nor3b_1 _709_ (.A(_119_),
    .B(_193_),
    .C_N(_201_),
    .Y(_012_));
 sky130_fd_sc_hd__nand4_2 _710_ (.A(_409_),
    .B(_411_),
    .C(_413_),
    .D(_415_),
    .Y(_202_));
 sky130_fd_sc_hd__nand2_1 _711_ (.A(_417_),
    .B(_419_),
    .Y(_203_));
 sky130_fd_sc_hd__nor4_1 _712_ (.A(_422_),
    .B(_440_),
    .C(_202_),
    .D(_203_),
    .Y(_204_));
 sky130_fd_sc_hd__nor2_1 _713_ (.A(_422_),
    .B(_443_),
    .Y(_205_));
 sky130_fd_sc_hd__o21ai_0 _714_ (.A1(_423_),
    .A2(_205_),
    .B1(_419_),
    .Y(_206_));
 sky130_fd_sc_hd__nand2b_1 _715_ (.A_N(_418_),
    .B(_206_),
    .Y(_207_));
 sky130_fd_sc_hd__a21oi_1 _716_ (.A1(_417_),
    .A2(_207_),
    .B1(_416_),
    .Y(_208_));
 sky130_fd_sc_hd__a21o_1 _717_ (.A1(_414_),
    .A2(_413_),
    .B1(_412_),
    .X(_209_));
 sky130_fd_sc_hd__a21o_1 _718_ (.A1(_411_),
    .A2(_209_),
    .B1(_410_),
    .X(_210_));
 sky130_fd_sc_hd__a21oi_1 _719_ (.A1(_409_),
    .A2(_210_),
    .B1(_408_),
    .Y(_211_));
 sky130_fd_sc_hd__o21ai_0 _720_ (.A1(_202_),
    .A2(_208_),
    .B1(_211_),
    .Y(_212_));
 sky130_fd_sc_hd__nor3b_1 _721_ (.A(_119_),
    .B(_204_),
    .C_N(_212_),
    .Y(_013_));
 sky130_fd_sc_hd__fa_1 _722_ (.A(_213_),
    .B(net8),
    .CIN(_214_),
    .COUT(_215_),
    .SUM(_216_));
 sky130_fd_sc_hd__fa_1 _723_ (.A(net2),
    .B(net8),
    .CIN(_217_),
    .COUT(_218_),
    .SUM(_219_));
 sky130_fd_sc_hd__ha_2 _724_ (.A(_220_),
    .B(net9),
    .COUT(_221_),
    .SUM(_222_));
 sky130_fd_sc_hd__ha_1 _725_ (.A(net3),
    .B(net9),
    .COUT(_223_),
    .SUM(_224_));
 sky130_fd_sc_hd__ha_1 _726_ (.A(_225_),
    .B(_226_),
    .COUT(_227_),
    .SUM(_228_));
 sky130_fd_sc_hd__ha_1 _727_ (.A(_229_),
    .B(_230_),
    .COUT(_231_),
    .SUM(_232_));
 sky130_fd_sc_hd__ha_1 _728_ (.A(_233_),
    .B(_234_),
    .COUT(_235_),
    .SUM(_236_));
 sky130_fd_sc_hd__ha_1 _729_ (.A(_237_),
    .B(_238_),
    .COUT(_239_),
    .SUM(_240_));
 sky130_fd_sc_hd__ha_1 _730_ (.A(_241_),
    .B(_242_),
    .COUT(_243_),
    .SUM(_244_));
 sky130_fd_sc_hd__ha_1 _731_ (.A(_245_),
    .B(_246_),
    .COUT(_247_),
    .SUM(_248_));
 sky130_fd_sc_hd__ha_1 _732_ (.A(_216_),
    .B(\counter[1] ),
    .COUT(_250_),
    .SUM(_251_));
 sky130_fd_sc_hd__ha_1 _733_ (.A(_252_),
    .B(net12),
    .COUT(_253_),
    .SUM(_254_));
 sky130_fd_sc_hd__ha_1 _734_ (.A(net6),
    .B(net12),
    .COUT(_255_),
    .SUM(_256_));
 sky130_fd_sc_hd__ha_2 _735_ (.A(_257_),
    .B(net11),
    .COUT(_258_),
    .SUM(_259_));
 sky130_fd_sc_hd__ha_1 _736_ (.A(net5),
    .B(net11),
    .COUT(_260_),
    .SUM(_261_));
 sky130_fd_sc_hd__ha_1 _737_ (.A(_262_),
    .B(net10),
    .COUT(_263_),
    .SUM(_264_));
 sky130_fd_sc_hd__ha_1 _738_ (.A(net4),
    .B(net10),
    .COUT(_265_),
    .SUM(_266_));
 sky130_fd_sc_hd__ha_1 _739_ (.A(_213_),
    .B(net8),
    .COUT(_267_),
    .SUM(_249_));
 sky130_fd_sc_hd__ha_1 _740_ (.A(net2),
    .B(net8),
    .COUT(_268_),
    .SUM(_269_));
 sky130_fd_sc_hd__ha_1 _741_ (.A(_225_),
    .B(_270_),
    .COUT(_271_),
    .SUM(_272_));
 sky130_fd_sc_hd__ha_1 _742_ (.A(_229_),
    .B(_273_),
    .COUT(_274_),
    .SUM(_275_));
 sky130_fd_sc_hd__ha_1 _743_ (.A(_233_),
    .B(_276_),
    .COUT(_277_),
    .SUM(_278_));
 sky130_fd_sc_hd__ha_1 _744_ (.A(_237_),
    .B(_279_),
    .COUT(_280_),
    .SUM(_281_));
 sky130_fd_sc_hd__ha_1 _745_ (.A(_241_),
    .B(_282_),
    .COUT(_283_),
    .SUM(_284_));
 sky130_fd_sc_hd__ha_1 _746_ (.A(_245_),
    .B(_285_),
    .COUT(_286_),
    .SUM(_287_));
 sky130_fd_sc_hd__ha_1 _747_ (.A(_288_),
    .B(_219_),
    .COUT(_289_),
    .SUM(_290_));
 sky130_fd_sc_hd__ha_1 _748_ (.A(\counter[1] ),
    .B(_219_),
    .COUT(_291_),
    .SUM(_292_));
 sky130_fd_sc_hd__ha_1 _749_ (.A(net1),
    .B(_293_),
    .COUT(_294_),
    .SUM(_295_));
 sky130_fd_sc_hd__ha_1 _750_ (.A(net1),
    .B(net7),
    .COUT(_217_),
    .SUM(_296_));
 sky130_fd_sc_hd__ha_1 _751_ (.A(_297_),
    .B(_295_),
    .COUT(_298_),
    .SUM(_299_));
 sky130_fd_sc_hd__ha_1 _752_ (.A(\counter[0] ),
    .B(_295_),
    .COUT(_300_),
    .SUM(_301_));
 sky130_fd_sc_hd__ha_1 _753_ (.A(_233_),
    .B(_252_),
    .COUT(_302_),
    .SUM(_303_));
 sky130_fd_sc_hd__ha_1 _754_ (.A(_237_),
    .B(_257_),
    .COUT(_304_),
    .SUM(_305_));
 sky130_fd_sc_hd__ha_1 _755_ (.A(_241_),
    .B(_262_),
    .COUT(_306_),
    .SUM(_307_));
 sky130_fd_sc_hd__ha_1 _756_ (.A(_245_),
    .B(_220_),
    .COUT(_308_),
    .SUM(_309_));
 sky130_fd_sc_hd__ha_1 _757_ (.A(_226_),
    .B(_310_),
    .COUT(_311_),
    .SUM(_312_));
 sky130_fd_sc_hd__ha_1 _758_ (.A(_230_),
    .B(_313_),
    .COUT(_314_),
    .SUM(_315_));
 sky130_fd_sc_hd__ha_1 _759_ (.A(_234_),
    .B(_316_),
    .COUT(_317_),
    .SUM(_318_));
 sky130_fd_sc_hd__ha_1 _760_ (.A(_238_),
    .B(_319_),
    .COUT(_320_),
    .SUM(_321_));
 sky130_fd_sc_hd__ha_1 _761_ (.A(_242_),
    .B(_322_),
    .COUT(_323_),
    .SUM(_324_));
 sky130_fd_sc_hd__ha_1 _762_ (.A(_246_),
    .B(_325_),
    .COUT(_326_),
    .SUM(_327_));
 sky130_fd_sc_hd__ha_2 _763_ (.A(\counter[0] ),
    .B(\counter[1] ),
    .COUT(_328_),
    .SUM(_329_));
 sky130_fd_sc_hd__ha_1 _764_ (.A(_216_),
    .B(_330_),
    .COUT(_331_),
    .SUM(_332_));
 sky130_fd_sc_hd__ha_1 _765_ (.A(_297_),
    .B(_295_),
    .COUT(_333_),
    .SUM(_334_));
 sky130_fd_sc_hd__ha_1 _766_ (.A(\counter[0] ),
    .B(_295_),
    .COUT(_335_),
    .SUM(_336_));
 sky130_fd_sc_hd__ha_1 _767_ (.A(_273_),
    .B(_313_),
    .COUT(_337_),
    .SUM(_338_));
 sky130_fd_sc_hd__ha_1 _768_ (.A(_276_),
    .B(_316_),
    .COUT(_339_),
    .SUM(_340_));
 sky130_fd_sc_hd__ha_1 _769_ (.A(_279_),
    .B(_319_),
    .COUT(_341_),
    .SUM(_342_));
 sky130_fd_sc_hd__ha_1 _770_ (.A(_282_),
    .B(_322_),
    .COUT(_343_),
    .SUM(_344_));
 sky130_fd_sc_hd__ha_1 _771_ (.A(_285_),
    .B(_325_),
    .COUT(_345_),
    .SUM(_346_));
 sky130_fd_sc_hd__ha_1 _772_ (.A(_219_),
    .B(_330_),
    .COUT(_347_),
    .SUM(_348_));
 sky130_fd_sc_hd__ha_1 _773_ (.A(_252_),
    .B(_316_),
    .COUT(_349_),
    .SUM(_350_));
 sky130_fd_sc_hd__ha_1 _774_ (.A(_257_),
    .B(_319_),
    .COUT(_351_),
    .SUM(_352_));
 sky130_fd_sc_hd__ha_1 _775_ (.A(_262_),
    .B(_322_),
    .COUT(_353_),
    .SUM(_354_));
 sky130_fd_sc_hd__ha_1 _776_ (.A(_220_),
    .B(_325_),
    .COUT(_355_),
    .SUM(_356_));
 sky130_fd_sc_hd__ha_1 _777_ (.A(_213_),
    .B(_330_),
    .COUT(_357_),
    .SUM(_358_));
 sky130_fd_sc_hd__ha_1 _778_ (.A(_297_),
    .B(net1),
    .COUT(_359_),
    .SUM(_360_));
 sky130_fd_sc_hd__ha_1 _779_ (.A(\counter[0] ),
    .B(net1),
    .COUT(_361_),
    .SUM(_362_));
 sky130_fd_sc_hd__ha_1 _780_ (.A(_363_),
    .B(_226_),
    .COUT(_364_),
    .SUM(_365_));
 sky130_fd_sc_hd__ha_1 _781_ (.A(_366_),
    .B(_230_),
    .COUT(_367_),
    .SUM(_368_));
 sky130_fd_sc_hd__ha_1 _782_ (.A(_369_),
    .B(_234_),
    .COUT(_370_),
    .SUM(_371_));
 sky130_fd_sc_hd__ha_1 _783_ (.A(_372_),
    .B(_238_),
    .COUT(_373_),
    .SUM(_374_));
 sky130_fd_sc_hd__ha_1 _784_ (.A(_375_),
    .B(_242_),
    .COUT(_376_),
    .SUM(_377_));
 sky130_fd_sc_hd__ha_2 _785_ (.A(\counter[1] ),
    .B(_245_),
    .COUT(_378_),
    .SUM(_379_));
 sky130_fd_sc_hd__ha_2 _786_ (.A(\counter[1] ),
    .B(\counter[2] ),
    .COUT(_380_),
    .SUM(_381_));
 sky130_fd_sc_hd__ha_1 _787_ (.A(_379_),
    .B(_246_),
    .COUT(_382_),
    .SUM(_383_));
 sky130_fd_sc_hd__ha_1 _788_ (.A(_288_),
    .B(_216_),
    .COUT(_384_),
    .SUM(_385_));
 sky130_fd_sc_hd__ha_1 _789_ (.A(_366_),
    .B(_273_),
    .COUT(_386_),
    .SUM(_387_));
 sky130_fd_sc_hd__ha_1 _790_ (.A(_369_),
    .B(_276_),
    .COUT(_388_),
    .SUM(_389_));
 sky130_fd_sc_hd__ha_1 _791_ (.A(_372_),
    .B(_279_),
    .COUT(_390_),
    .SUM(_391_));
 sky130_fd_sc_hd__ha_1 _792_ (.A(_375_),
    .B(_282_),
    .COUT(_392_),
    .SUM(_393_));
 sky130_fd_sc_hd__ha_1 _793_ (.A(_379_),
    .B(_285_),
    .COUT(_394_),
    .SUM(_395_));
 sky130_fd_sc_hd__ha_1 _794_ (.A(_252_),
    .B(_369_),
    .COUT(_396_),
    .SUM(_397_));
 sky130_fd_sc_hd__ha_1 _795_ (.A(_257_),
    .B(_372_),
    .COUT(_398_),
    .SUM(_399_));
 sky130_fd_sc_hd__ha_1 _796_ (.A(_262_),
    .B(_375_),
    .COUT(_400_),
    .SUM(_401_));
 sky130_fd_sc_hd__ha_1 _797_ (.A(_220_),
    .B(_379_),
    .COUT(_402_),
    .SUM(_403_));
 sky130_fd_sc_hd__ha_1 _798_ (.A(_288_),
    .B(_213_),
    .COUT(_404_),
    .SUM(_405_));
 sky130_fd_sc_hd__ha_1 _799_ (.A(\counter[1] ),
    .B(_213_),
    .COUT(_406_),
    .SUM(_407_));
 sky130_fd_sc_hd__ha_1 _800_ (.A(_363_),
    .B(net14),
    .COUT(_408_),
    .SUM(_409_));
 sky130_fd_sc_hd__ha_1 _801_ (.A(_366_),
    .B(net13),
    .COUT(_410_),
    .SUM(_411_));
 sky130_fd_sc_hd__ha_1 _802_ (.A(net12),
    .B(_369_),
    .COUT(_412_),
    .SUM(_413_));
 sky130_fd_sc_hd__ha_1 _803_ (.A(net11),
    .B(_372_),
    .COUT(_414_),
    .SUM(_415_));
 sky130_fd_sc_hd__ha_1 _804_ (.A(net10),
    .B(_375_),
    .COUT(_416_),
    .SUM(_417_));
 sky130_fd_sc_hd__ha_1 _805_ (.A(net9),
    .B(_379_),
    .COUT(_418_),
    .SUM(_419_));
 sky130_fd_sc_hd__ha_1 _806_ (.A(\counter[1] ),
    .B(_420_),
    .COUT(_421_),
    .SUM(_422_));
 sky130_fd_sc_hd__ha_1 _807_ (.A(\counter[1] ),
    .B(net8),
    .COUT(_423_),
    .SUM(_424_));
 sky130_fd_sc_hd__ha_1 _808_ (.A(net14),
    .B(_310_),
    .COUT(_425_),
    .SUM(_426_));
 sky130_fd_sc_hd__ha_1 _809_ (.A(net13),
    .B(_313_),
    .COUT(_427_),
    .SUM(_428_));
 sky130_fd_sc_hd__ha_1 _810_ (.A(net12),
    .B(_316_),
    .COUT(_429_),
    .SUM(_430_));
 sky130_fd_sc_hd__ha_1 _811_ (.A(net11),
    .B(_319_),
    .COUT(_431_),
    .SUM(_432_));
 sky130_fd_sc_hd__ha_1 _812_ (.A(net10),
    .B(_322_),
    .COUT(_433_),
    .SUM(_434_));
 sky130_fd_sc_hd__ha_1 _813_ (.A(net9),
    .B(_325_),
    .COUT(_435_),
    .SUM(_436_));
 sky130_fd_sc_hd__ha_1 _814_ (.A(net8),
    .B(_330_),
    .COUT(_437_),
    .SUM(_438_));
 sky130_fd_sc_hd__ha_1 _815_ (.A(_297_),
    .B(_293_),
    .COUT(_439_),
    .SUM(_440_));
 sky130_fd_sc_hd__ha_1 _816_ (.A(_297_),
    .B(net7),
    .COUT(_441_),
    .SUM(_442_));
 sky130_fd_sc_hd__ha_1 _817_ (.A(\counter[0] ),
    .B(_293_),
    .COUT(_443_),
    .SUM(_444_));
 sky130_fd_sc_hd__ha_1 _818_ (.A(\counter[7] ),
    .B(_445_),
    .COUT(_446_),
    .SUM(_447_));
 sky130_fd_sc_hd__ha_1 _819_ (.A(\counter[6] ),
    .B(_448_),
    .COUT(_449_),
    .SUM(_450_));
 sky130_fd_sc_hd__ha_1 _820_ (.A(\counter[5] ),
    .B(_451_),
    .COUT(_452_),
    .SUM(_453_));
 sky130_fd_sc_hd__ha_1 _821_ (.A(\counter[4] ),
    .B(_454_),
    .COUT(_455_),
    .SUM(_456_));
 sky130_fd_sc_hd__ha_1 _822_ (.A(\counter[3] ),
    .B(_457_),
    .COUT(_458_),
    .SUM(_459_));
 sky130_fd_sc_hd__ha_1 _823_ (.A(\counter[2] ),
    .B(_460_),
    .COUT(_461_),
    .SUM(_462_));
 sky130_fd_sc_hd__dfxtp_4 \counter[0]$_SDFFE_PN0P_  (.D(_000_),
    .Q(\counter[0] ),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_4 \counter[1]$_SDFFE_PN0P_  (.D(_001_),
    .Q(\counter[1] ),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \counter[2]$_SDFFE_PN0P_  (.D(_002_),
    .Q(\counter[2] ),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \counter[3]$_SDFFE_PN0P_  (.D(_003_),
    .Q(\counter[3] ),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \counter[4]$_SDFFE_PN0P_  (.D(_004_),
    .Q(\counter[4] ),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_2 \counter[5]$_SDFFE_PN0P_  (.D(_005_),
    .Q(\counter[5] ),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_2 \counter[6]$_SDFFE_PN0P_  (.D(_006_),
    .Q(\counter[6] ),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_2 \counter[7]$_SDFFE_PN0P_  (.D(_007_),
    .Q(\counter[7] ),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \pwm_n_reg[0]$_SDFF_PN0_  (.D(_008_),
    .Q(net16),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \pwm_n_reg[1]$_SDFF_PN0_  (.D(_009_),
    .Q(net17),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \pwm_n_reg[2]$_SDFF_PN0_  (.D(_010_),
    .Q(net18),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \pwm_p_reg[0]$_SDFF_PN0_  (.D(_011_),
    .Q(net19),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \pwm_p_reg[1]$_SDFF_PN0_  (.D(_012_),
    .Q(net20),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \pwm_p_reg[2]$_SDFF_PN0_  (.D(_013_),
    .Q(net21),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_71 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(deadtime[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(deadtime[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(deadtime[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(deadtime[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(deadtime[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(deadtime[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(duty[0]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(duty[1]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(duty[2]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(duty[3]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(duty[4]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(duty[5]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(duty[6]),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input14 (.A(duty[7]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input15 (.A(rst_n),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net16),
    .X(pwm_n_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net17),
    .X(pwm_n_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net18),
    .X(pwm_n_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net19),
    .X(pwm_p_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net20),
    .X(pwm_p_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net21),
    .X(pwm_p_out[2]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload0 (.A(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_114 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_54 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_143 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_162 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_87 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_13 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_62 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_53 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_122 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_92 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_162 ();
endmodule
