module multi_ported_fifo (almost_empty,
    almost_full,
    clk,
    empty,
    full,
    rst_n,
    data_count,
    rd_data,
    rd_en,
    rd_valid,
    wr_data,
    wr_en,
    wr_ready);
 output almost_empty;
 output almost_full;
 input clk;
 output empty;
 output full;
 input rst_n;
 output [4:0] data_count;
 output [63:0] rd_data;
 input [1:0] rd_en;
 output [1:0] rd_valid;
 input [63:0] wr_data;
 input [1:0] wr_en;
 output [1:0] wr_ready;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire net166;
 wire _0714_;
 wire _0715_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire \mem[0][0] ;
 wire \mem[0][10] ;
 wire \mem[0][11] ;
 wire \mem[0][12] ;
 wire \mem[0][13] ;
 wire \mem[0][14] ;
 wire \mem[0][15] ;
 wire \mem[0][16] ;
 wire \mem[0][17] ;
 wire \mem[0][18] ;
 wire \mem[0][19] ;
 wire \mem[0][1] ;
 wire \mem[0][20] ;
 wire \mem[0][21] ;
 wire \mem[0][22] ;
 wire \mem[0][23] ;
 wire \mem[0][24] ;
 wire \mem[0][25] ;
 wire \mem[0][26] ;
 wire \mem[0][27] ;
 wire \mem[0][28] ;
 wire \mem[0][29] ;
 wire \mem[0][2] ;
 wire \mem[0][30] ;
 wire \mem[0][31] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[0][8] ;
 wire \mem[0][9] ;
 wire \mem[10][0] ;
 wire \mem[10][10] ;
 wire \mem[10][11] ;
 wire \mem[10][12] ;
 wire \mem[10][13] ;
 wire \mem[10][14] ;
 wire \mem[10][15] ;
 wire \mem[10][16] ;
 wire \mem[10][17] ;
 wire \mem[10][18] ;
 wire \mem[10][19] ;
 wire \mem[10][1] ;
 wire \mem[10][20] ;
 wire \mem[10][21] ;
 wire \mem[10][22] ;
 wire \mem[10][23] ;
 wire \mem[10][24] ;
 wire \mem[10][25] ;
 wire \mem[10][26] ;
 wire \mem[10][27] ;
 wire \mem[10][28] ;
 wire \mem[10][29] ;
 wire \mem[10][2] ;
 wire \mem[10][30] ;
 wire \mem[10][31] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[10][8] ;
 wire \mem[10][9] ;
 wire \mem[11][0] ;
 wire \mem[11][10] ;
 wire \mem[11][11] ;
 wire \mem[11][12] ;
 wire \mem[11][13] ;
 wire \mem[11][14] ;
 wire \mem[11][15] ;
 wire \mem[11][16] ;
 wire \mem[11][17] ;
 wire \mem[11][18] ;
 wire \mem[11][19] ;
 wire \mem[11][1] ;
 wire \mem[11][20] ;
 wire \mem[11][21] ;
 wire \mem[11][22] ;
 wire \mem[11][23] ;
 wire \mem[11][24] ;
 wire \mem[11][25] ;
 wire \mem[11][26] ;
 wire \mem[11][27] ;
 wire \mem[11][28] ;
 wire \mem[11][29] ;
 wire \mem[11][2] ;
 wire \mem[11][30] ;
 wire \mem[11][31] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[11][8] ;
 wire \mem[11][9] ;
 wire \mem[12][0] ;
 wire \mem[12][10] ;
 wire \mem[12][11] ;
 wire \mem[12][12] ;
 wire \mem[12][13] ;
 wire \mem[12][14] ;
 wire \mem[12][15] ;
 wire \mem[12][16] ;
 wire \mem[12][17] ;
 wire \mem[12][18] ;
 wire \mem[12][19] ;
 wire \mem[12][1] ;
 wire \mem[12][20] ;
 wire \mem[12][21] ;
 wire \mem[12][22] ;
 wire \mem[12][23] ;
 wire \mem[12][24] ;
 wire \mem[12][25] ;
 wire \mem[12][26] ;
 wire \mem[12][27] ;
 wire \mem[12][28] ;
 wire \mem[12][29] ;
 wire \mem[12][2] ;
 wire \mem[12][30] ;
 wire \mem[12][31] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[12][8] ;
 wire \mem[12][9] ;
 wire \mem[13][0] ;
 wire \mem[13][10] ;
 wire \mem[13][11] ;
 wire \mem[13][12] ;
 wire \mem[13][13] ;
 wire \mem[13][14] ;
 wire \mem[13][15] ;
 wire \mem[13][16] ;
 wire \mem[13][17] ;
 wire \mem[13][18] ;
 wire \mem[13][19] ;
 wire \mem[13][1] ;
 wire \mem[13][20] ;
 wire \mem[13][21] ;
 wire \mem[13][22] ;
 wire \mem[13][23] ;
 wire \mem[13][24] ;
 wire \mem[13][25] ;
 wire \mem[13][26] ;
 wire \mem[13][27] ;
 wire \mem[13][28] ;
 wire \mem[13][29] ;
 wire \mem[13][2] ;
 wire \mem[13][30] ;
 wire \mem[13][31] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[13][8] ;
 wire \mem[13][9] ;
 wire \mem[14][0] ;
 wire \mem[14][10] ;
 wire \mem[14][11] ;
 wire \mem[14][12] ;
 wire \mem[14][13] ;
 wire \mem[14][14] ;
 wire \mem[14][15] ;
 wire \mem[14][16] ;
 wire \mem[14][17] ;
 wire \mem[14][18] ;
 wire \mem[14][19] ;
 wire \mem[14][1] ;
 wire \mem[14][20] ;
 wire \mem[14][21] ;
 wire \mem[14][22] ;
 wire \mem[14][23] ;
 wire \mem[14][24] ;
 wire \mem[14][25] ;
 wire \mem[14][26] ;
 wire \mem[14][27] ;
 wire \mem[14][28] ;
 wire \mem[14][29] ;
 wire \mem[14][2] ;
 wire \mem[14][30] ;
 wire \mem[14][31] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[14][8] ;
 wire \mem[14][9] ;
 wire \mem[15][0] ;
 wire \mem[15][10] ;
 wire \mem[15][11] ;
 wire \mem[15][12] ;
 wire \mem[15][13] ;
 wire \mem[15][14] ;
 wire \mem[15][15] ;
 wire \mem[15][16] ;
 wire \mem[15][17] ;
 wire \mem[15][18] ;
 wire \mem[15][19] ;
 wire \mem[15][1] ;
 wire \mem[15][20] ;
 wire \mem[15][21] ;
 wire \mem[15][22] ;
 wire \mem[15][23] ;
 wire \mem[15][24] ;
 wire \mem[15][25] ;
 wire \mem[15][26] ;
 wire \mem[15][27] ;
 wire \mem[15][28] ;
 wire \mem[15][29] ;
 wire \mem[15][2] ;
 wire \mem[15][30] ;
 wire \mem[15][31] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[15][8] ;
 wire \mem[15][9] ;
 wire \mem[1][0] ;
 wire \mem[1][10] ;
 wire \mem[1][11] ;
 wire \mem[1][12] ;
 wire \mem[1][13] ;
 wire \mem[1][14] ;
 wire \mem[1][15] ;
 wire \mem[1][16] ;
 wire \mem[1][17] ;
 wire \mem[1][18] ;
 wire \mem[1][19] ;
 wire \mem[1][1] ;
 wire \mem[1][20] ;
 wire \mem[1][21] ;
 wire \mem[1][22] ;
 wire \mem[1][23] ;
 wire \mem[1][24] ;
 wire \mem[1][25] ;
 wire \mem[1][26] ;
 wire \mem[1][27] ;
 wire \mem[1][28] ;
 wire \mem[1][29] ;
 wire \mem[1][2] ;
 wire \mem[1][30] ;
 wire \mem[1][31] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[1][8] ;
 wire \mem[1][9] ;
 wire \mem[2][0] ;
 wire \mem[2][10] ;
 wire \mem[2][11] ;
 wire \mem[2][12] ;
 wire \mem[2][13] ;
 wire \mem[2][14] ;
 wire \mem[2][15] ;
 wire \mem[2][16] ;
 wire \mem[2][17] ;
 wire \mem[2][18] ;
 wire \mem[2][19] ;
 wire \mem[2][1] ;
 wire \mem[2][20] ;
 wire \mem[2][21] ;
 wire \mem[2][22] ;
 wire \mem[2][23] ;
 wire \mem[2][24] ;
 wire \mem[2][25] ;
 wire \mem[2][26] ;
 wire \mem[2][27] ;
 wire \mem[2][28] ;
 wire \mem[2][29] ;
 wire \mem[2][2] ;
 wire \mem[2][30] ;
 wire \mem[2][31] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[2][8] ;
 wire \mem[2][9] ;
 wire \mem[3][0] ;
 wire \mem[3][10] ;
 wire \mem[3][11] ;
 wire \mem[3][12] ;
 wire \mem[3][13] ;
 wire \mem[3][14] ;
 wire \mem[3][15] ;
 wire \mem[3][16] ;
 wire \mem[3][17] ;
 wire \mem[3][18] ;
 wire \mem[3][19] ;
 wire \mem[3][1] ;
 wire \mem[3][20] ;
 wire \mem[3][21] ;
 wire \mem[3][22] ;
 wire \mem[3][23] ;
 wire \mem[3][24] ;
 wire \mem[3][25] ;
 wire \mem[3][26] ;
 wire \mem[3][27] ;
 wire \mem[3][28] ;
 wire \mem[3][29] ;
 wire \mem[3][2] ;
 wire \mem[3][30] ;
 wire \mem[3][31] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[3][8] ;
 wire \mem[3][9] ;
 wire \mem[4][0] ;
 wire \mem[4][10] ;
 wire \mem[4][11] ;
 wire \mem[4][12] ;
 wire \mem[4][13] ;
 wire \mem[4][14] ;
 wire \mem[4][15] ;
 wire \mem[4][16] ;
 wire \mem[4][17] ;
 wire \mem[4][18] ;
 wire \mem[4][19] ;
 wire \mem[4][1] ;
 wire \mem[4][20] ;
 wire \mem[4][21] ;
 wire \mem[4][22] ;
 wire \mem[4][23] ;
 wire \mem[4][24] ;
 wire \mem[4][25] ;
 wire \mem[4][26] ;
 wire \mem[4][27] ;
 wire \mem[4][28] ;
 wire \mem[4][29] ;
 wire \mem[4][2] ;
 wire \mem[4][30] ;
 wire \mem[4][31] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[4][8] ;
 wire \mem[4][9] ;
 wire \mem[5][0] ;
 wire \mem[5][10] ;
 wire \mem[5][11] ;
 wire \mem[5][12] ;
 wire \mem[5][13] ;
 wire \mem[5][14] ;
 wire \mem[5][15] ;
 wire \mem[5][16] ;
 wire \mem[5][17] ;
 wire \mem[5][18] ;
 wire \mem[5][19] ;
 wire \mem[5][1] ;
 wire \mem[5][20] ;
 wire \mem[5][21] ;
 wire \mem[5][22] ;
 wire \mem[5][23] ;
 wire \mem[5][24] ;
 wire \mem[5][25] ;
 wire \mem[5][26] ;
 wire \mem[5][27] ;
 wire \mem[5][28] ;
 wire \mem[5][29] ;
 wire \mem[5][2] ;
 wire \mem[5][30] ;
 wire \mem[5][31] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[5][8] ;
 wire \mem[5][9] ;
 wire \mem[6][0] ;
 wire \mem[6][10] ;
 wire \mem[6][11] ;
 wire \mem[6][12] ;
 wire \mem[6][13] ;
 wire \mem[6][14] ;
 wire \mem[6][15] ;
 wire \mem[6][16] ;
 wire \mem[6][17] ;
 wire \mem[6][18] ;
 wire \mem[6][19] ;
 wire \mem[6][1] ;
 wire \mem[6][20] ;
 wire \mem[6][21] ;
 wire \mem[6][22] ;
 wire \mem[6][23] ;
 wire \mem[6][24] ;
 wire \mem[6][25] ;
 wire \mem[6][26] ;
 wire \mem[6][27] ;
 wire \mem[6][28] ;
 wire \mem[6][29] ;
 wire \mem[6][2] ;
 wire \mem[6][30] ;
 wire \mem[6][31] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[6][8] ;
 wire \mem[6][9] ;
 wire \mem[7][0] ;
 wire \mem[7][10] ;
 wire \mem[7][11] ;
 wire \mem[7][12] ;
 wire \mem[7][13] ;
 wire \mem[7][14] ;
 wire \mem[7][15] ;
 wire \mem[7][16] ;
 wire \mem[7][17] ;
 wire \mem[7][18] ;
 wire \mem[7][19] ;
 wire \mem[7][1] ;
 wire \mem[7][20] ;
 wire \mem[7][21] ;
 wire \mem[7][22] ;
 wire \mem[7][23] ;
 wire \mem[7][24] ;
 wire \mem[7][25] ;
 wire \mem[7][26] ;
 wire \mem[7][27] ;
 wire \mem[7][28] ;
 wire \mem[7][29] ;
 wire \mem[7][2] ;
 wire \mem[7][30] ;
 wire \mem[7][31] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[7][8] ;
 wire \mem[7][9] ;
 wire \mem[8][0] ;
 wire \mem[8][10] ;
 wire \mem[8][11] ;
 wire \mem[8][12] ;
 wire \mem[8][13] ;
 wire \mem[8][14] ;
 wire \mem[8][15] ;
 wire \mem[8][16] ;
 wire \mem[8][17] ;
 wire \mem[8][18] ;
 wire \mem[8][19] ;
 wire \mem[8][1] ;
 wire \mem[8][20] ;
 wire \mem[8][21] ;
 wire \mem[8][22] ;
 wire \mem[8][23] ;
 wire \mem[8][24] ;
 wire \mem[8][25] ;
 wire \mem[8][26] ;
 wire \mem[8][27] ;
 wire \mem[8][28] ;
 wire \mem[8][29] ;
 wire \mem[8][2] ;
 wire \mem[8][30] ;
 wire \mem[8][31] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[8][8] ;
 wire \mem[8][9] ;
 wire \mem[9][0] ;
 wire \mem[9][10] ;
 wire \mem[9][11] ;
 wire \mem[9][12] ;
 wire \mem[9][13] ;
 wire \mem[9][14] ;
 wire \mem[9][15] ;
 wire \mem[9][16] ;
 wire \mem[9][17] ;
 wire \mem[9][18] ;
 wire \mem[9][19] ;
 wire \mem[9][1] ;
 wire \mem[9][20] ;
 wire \mem[9][21] ;
 wire \mem[9][22] ;
 wire \mem[9][23] ;
 wire \mem[9][24] ;
 wire \mem[9][25] ;
 wire \mem[9][26] ;
 wire \mem[9][27] ;
 wire \mem[9][28] ;
 wire \mem[9][29] ;
 wire \mem[9][2] ;
 wire \mem[9][30] ;
 wire \mem[9][31] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \mem[9][8] ;
 wire \mem[9][9] ;
 wire \next_count[0] ;
 wire \next_count[1] ;
 wire \next_count[2] ;
 wire \next_count[3] ;
 wire \next_count[4] ;
 wire \rd_ptr[0] ;
 wire \rd_ptr[1] ;
 wire \rd_ptr[2] ;
 wire \rd_ptr[3] ;
 wire \wr_ptr[0] ;
 wire \wr_ptr[1] ;
 wire \wr_ptr[2] ;
 wire \wr_ptr[3] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net163;
 wire net164;
 wire net165;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;

 sky130_fd_sc_hd__inv_1 _2568_ (.A(_2512_),
    .Y(net77));
 sky130_fd_sc_hd__buf_6 _2569_ (.A(net71),
    .X(_0607_));
 sky130_fd_sc_hd__inv_1 _2570_ (.A(_0607_),
    .Y(_2514_));
 sky130_fd_sc_hd__nand2_2 _2571_ (.A(net67),
    .B(_2512_),
    .Y(_0608_));
 sky130_fd_sc_hd__clkbuf_4 _2572_ (.A(net72),
    .X(_0609_));
 sky130_fd_sc_hd__nor4_1 _2573_ (.A(_0609_),
    .B(_0607_),
    .C(net73),
    .D(_2548_),
    .Y(_0610_));
 sky130_fd_sc_hd__clkinv_4 _2574_ (.A(net75),
    .Y(_2510_));
 sky130_fd_sc_hd__a21oi_2 _2575_ (.A1(_2561_),
    .A2(_0610_),
    .B1(_2510_),
    .Y(_0611_));
 sky130_fd_sc_hd__nor2_1 _2576_ (.A(_0608_),
    .B(_0611_),
    .Y(_0612_));
 sky130_fd_sc_hd__inv_2 _2577_ (.A(_0612_),
    .Y(_2526_));
 sky130_fd_sc_hd__buf_2 _2578_ (.A(\wr_ptr[1] ),
    .X(_0613_));
 sky130_fd_sc_hd__inv_1 _2579_ (.A(_0613_),
    .Y(_2501_));
 sky130_fd_sc_hd__and2_0 _2580_ (.A(net67),
    .B(_2512_),
    .X(_0614_));
 sky130_fd_sc_hd__clkbuf_2 _2581_ (.A(_0614_),
    .X(_0615_));
 sky130_fd_sc_hd__nand2b_1 _2582_ (.A_N(net168),
    .B(_2552_),
    .Y(_0616_));
 sky130_fd_sc_hd__nand2_1 _2583_ (.A(net73),
    .B(_2565_),
    .Y(_0617_));
 sky130_fd_sc_hd__nand2_1 _2584_ (.A(_0609_),
    .B(_0607_),
    .Y(_0618_));
 sky130_fd_sc_hd__a21oi_2 _2585_ (.A1(_0616_),
    .A2(_0617_),
    .B1(_0618_),
    .Y(_0619_));
 sky130_fd_sc_hd__nand3_1 _2586_ (.A(_2510_),
    .B(net68),
    .C(_2512_),
    .Y(_0620_));
 sky130_fd_sc_hd__a21oi_1 _2587_ (.A1(_0615_),
    .A2(_0619_),
    .B1(_0620_),
    .Y(_2519_));
 sky130_fd_sc_hd__inv_1 _2588_ (.A(_2519_),
    .Y(_2525_));
 sky130_fd_sc_hd__clkbuf_4 _2589_ (.A(\wr_ptr[3] ),
    .X(_0621_));
 sky130_fd_sc_hd__clkbuf_4 _2590_ (.A(\wr_ptr[2] ),
    .X(_0622_));
 sky130_fd_sc_hd__or2_4 _2591_ (.A(_0621_),
    .B(_0622_),
    .X(_0623_));
 sky130_fd_sc_hd__clkbuf_8 _2592_ (.A(_0612_),
    .X(_2520_));
 sky130_fd_sc_hd__nand2_4 _2593_ (.A(_2504_),
    .B(_2520_),
    .Y(_0624_));
 sky130_fd_sc_hd__and3_1 _2594_ (.A(_2510_),
    .B(net68),
    .C(_2512_),
    .X(_0625_));
 sky130_fd_sc_hd__clkbuf_2 _2595_ (.A(_0625_),
    .X(_0626_));
 sky130_fd_sc_hd__nor3_1 _2596_ (.A(_0621_),
    .B(\wr_ptr[0] ),
    .C(_0615_),
    .Y(_0627_));
 sky130_fd_sc_hd__nand2_1 _2597_ (.A(\wr_ptr[2] ),
    .B(_0613_),
    .Y(_0628_));
 sky130_fd_sc_hd__nand2_1 _2598_ (.A(_0621_),
    .B(\wr_ptr[0] ),
    .Y(_0629_));
 sky130_fd_sc_hd__nor4_1 _2599_ (.A(_0608_),
    .B(_0619_),
    .C(_0628_),
    .D(_0629_),
    .Y(_0630_));
 sky130_fd_sc_hd__nor2b_1 _2600_ (.A(\wr_ptr[3] ),
    .B_N(\wr_ptr[0] ),
    .Y(_0631_));
 sky130_fd_sc_hd__nand2_1 _2601_ (.A(_0628_),
    .B(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__nor3_1 _2602_ (.A(_0608_),
    .B(_0619_),
    .C(_0632_),
    .Y(_0633_));
 sky130_fd_sc_hd__or3_1 _2603_ (.A(_0627_),
    .B(_0630_),
    .C(_0633_),
    .X(_0634_));
 sky130_fd_sc_hd__nand2b_1 _2604_ (.A_N(\wr_ptr[2] ),
    .B(_2508_),
    .Y(_0635_));
 sky130_fd_sc_hd__nand2b_1 _2605_ (.A_N(_2508_),
    .B(\wr_ptr[2] ),
    .Y(_0636_));
 sky130_fd_sc_hd__nand3_1 _2606_ (.A(_2503_),
    .B(_0635_),
    .C(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__nand2b_1 _2607_ (.A_N(_0622_),
    .B(_0613_),
    .Y(_0638_));
 sky130_fd_sc_hd__mux2i_1 _2608_ (.A0(_0637_),
    .A1(_0638_),
    .S(_2526_),
    .Y(_0639_));
 sky130_fd_sc_hd__and3_1 _2609_ (.A(_0626_),
    .B(_0634_),
    .C(_0639_),
    .X(_0640_));
 sky130_fd_sc_hd__buf_4 _2610_ (.A(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__buf_6 _2611_ (.A(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__o21bai_4 _2612_ (.A1(_0623_),
    .A2(_0624_),
    .B1_N(_0642_),
    .Y(_0007_));
 sky130_fd_sc_hd__nand2_1 _2613_ (.A(\wr_ptr[0] ),
    .B(_0608_),
    .Y(_0643_));
 sky130_fd_sc_hd__inv_1 _2614_ (.A(\wr_ptr[0] ),
    .Y(_2500_));
 sky130_fd_sc_hd__a21o_1 _2615_ (.A1(_0616_),
    .A2(_0617_),
    .B1(_0618_),
    .X(_0644_));
 sky130_fd_sc_hd__nand3_2 _2616_ (.A(_2500_),
    .B(_0615_),
    .C(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hd__a211o_4 _2617_ (.A1(_0643_),
    .A2(_0645_),
    .B1(_0621_),
    .C1(_0620_),
    .X(_0646_));
 sky130_fd_sc_hd__nor2_1 _2618_ (.A(\wr_ptr[2] ),
    .B(_2508_),
    .Y(_0647_));
 sky130_fd_sc_hd__and2_0 _2619_ (.A(\wr_ptr[2] ),
    .B(_2508_),
    .X(_0648_));
 sky130_fd_sc_hd__inv_1 _2620_ (.A(_2503_),
    .Y(_0649_));
 sky130_fd_sc_hd__a21o_1 _2621_ (.A1(_2561_),
    .A2(_0610_),
    .B1(_2510_),
    .X(_0650_));
 sky130_fd_sc_hd__o2111ai_2 _2622_ (.A1(_0647_),
    .A2(_0648_),
    .B1(_0649_),
    .C1(_0615_),
    .D1(_0650_),
    .Y(_0651_));
 sky130_fd_sc_hd__o31a_2 _2623_ (.A1(_0622_),
    .A2(_0613_),
    .A3(_2520_),
    .B1(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__nand2_4 _2624_ (.A(_2506_),
    .B(_2520_),
    .Y(_0653_));
 sky130_fd_sc_hd__o22ai_4 _2625_ (.A1(_0646_),
    .A2(_0652_),
    .B1(_0653_),
    .B2(_0623_),
    .Y(_0008_));
 sky130_fd_sc_hd__nand2_4 _2626_ (.A(_2508_),
    .B(_2520_),
    .Y(_0654_));
 sky130_fd_sc_hd__nand2_4 _2627_ (.A(_0621_),
    .B(_0622_),
    .Y(_0655_));
 sky130_fd_sc_hd__nand2_1 _2628_ (.A(_0621_),
    .B(_0626_),
    .Y(_0656_));
 sky130_fd_sc_hd__a21oi_4 _2629_ (.A1(_0643_),
    .A2(_0645_),
    .B1(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__nor2_1 _2630_ (.A(_0649_),
    .B(_0635_),
    .Y(_0658_));
 sky130_fd_sc_hd__nor2_1 _2631_ (.A(_0649_),
    .B(_0636_),
    .Y(_0659_));
 sky130_fd_sc_hd__o211ai_2 _2632_ (.A1(_0658_),
    .A2(_0659_),
    .B1(_0615_),
    .C1(_0650_),
    .Y(_0660_));
 sky130_fd_sc_hd__o21ai_4 _2633_ (.A1(_2520_),
    .A2(_0628_),
    .B1(_0660_),
    .Y(_0661_));
 sky130_fd_sc_hd__nand2_8 _2634_ (.A(_0657_),
    .B(_0661_),
    .Y(_0662_));
 sky130_fd_sc_hd__buf_6 _2635_ (.A(_0662_),
    .X(_0663_));
 sky130_fd_sc_hd__o21ai_4 _2636_ (.A1(_0654_),
    .A2(_0655_),
    .B1(_0663_),
    .Y(_0009_));
 sky130_fd_sc_hd__nand3_1 _2637_ (.A(_0621_),
    .B(_2500_),
    .C(_0608_),
    .Y(_0664_));
 sky130_fd_sc_hd__and2_0 _2638_ (.A(\wr_ptr[2] ),
    .B(\wr_ptr[1] ),
    .X(_0665_));
 sky130_fd_sc_hd__nand4_1 _2639_ (.A(_0615_),
    .B(_0644_),
    .C(_0665_),
    .D(_0631_),
    .Y(_0666_));
 sky130_fd_sc_hd__or4_1 _2640_ (.A(_0608_),
    .B(_0619_),
    .C(_0665_),
    .D(_0629_),
    .X(_0667_));
 sky130_fd_sc_hd__nand3_1 _2641_ (.A(_0664_),
    .B(_0666_),
    .C(_0667_),
    .Y(_0668_));
 sky130_fd_sc_hd__and3_1 _2642_ (.A(_0626_),
    .B(_0661_),
    .C(_0668_),
    .X(_0669_));
 sky130_fd_sc_hd__buf_6 _2643_ (.A(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__buf_6 _2644_ (.A(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__o21bai_4 _2645_ (.A1(_0624_),
    .A2(_0655_),
    .B1_N(_0671_),
    .Y(_0010_));
 sky130_fd_sc_hd__nand2_1 _2646_ (.A(_0622_),
    .B(_2501_),
    .Y(_0672_));
 sky130_fd_sc_hd__a2111o_1 _2647_ (.A1(_0635_),
    .A2(_0636_),
    .B1(_2503_),
    .C1(_0608_),
    .D1(_0611_),
    .X(_0673_));
 sky130_fd_sc_hd__o21ai_1 _2648_ (.A1(_2520_),
    .A2(_0672_),
    .B1(_0673_),
    .Y(_0674_));
 sky130_fd_sc_hd__and2_0 _2649_ (.A(_0657_),
    .B(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__buf_6 _2650_ (.A(_0675_),
    .X(_0676_));
 sky130_fd_sc_hd__buf_6 _2651_ (.A(_0676_),
    .X(_0677_));
 sky130_fd_sc_hd__o21bai_4 _2652_ (.A1(_0653_),
    .A2(_0655_),
    .B1_N(_0677_),
    .Y(_0011_));
 sky130_fd_sc_hd__nand2_4 _2653_ (.A(_2502_),
    .B(_2520_),
    .Y(_0678_));
 sky130_fd_sc_hd__and3_1 _2654_ (.A(_0626_),
    .B(_0668_),
    .C(_0674_),
    .X(_0679_));
 sky130_fd_sc_hd__buf_6 _2655_ (.A(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__buf_6 _2656_ (.A(_0680_),
    .X(_0681_));
 sky130_fd_sc_hd__o21bai_4 _2657_ (.A1(_0655_),
    .A2(_0678_),
    .B1_N(_0681_),
    .Y(_0012_));
 sky130_fd_sc_hd__nand2b_4 _2658_ (.A_N(_0622_),
    .B(_0621_),
    .Y(_0682_));
 sky130_fd_sc_hd__and3_1 _2659_ (.A(_0626_),
    .B(_0639_),
    .C(_0668_),
    .X(_0683_));
 sky130_fd_sc_hd__buf_6 _2660_ (.A(_0683_),
    .X(_0684_));
 sky130_fd_sc_hd__buf_6 _2661_ (.A(_0684_),
    .X(_0685_));
 sky130_fd_sc_hd__o21bai_4 _2662_ (.A1(_0624_),
    .A2(_0682_),
    .B1_N(_0685_),
    .Y(_0014_));
 sky130_fd_sc_hd__nand2b_4 _2663_ (.A_N(_0621_),
    .B(_0622_),
    .Y(_0686_));
 sky130_fd_sc_hd__nor2b_1 _2664_ (.A(_0646_),
    .B_N(_0661_),
    .Y(_0687_));
 sky130_fd_sc_hd__buf_4 _2665_ (.A(_0687_),
    .X(_0688_));
 sky130_fd_sc_hd__buf_6 _2666_ (.A(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__o21bai_4 _2667_ (.A1(_0654_),
    .A2(_0686_),
    .B1_N(_0689_),
    .Y(_0002_));
 sky130_fd_sc_hd__and2_0 _2668_ (.A(_0639_),
    .B(_0657_),
    .X(_0690_));
 sky130_fd_sc_hd__buf_6 _2669_ (.A(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__buf_6 _2670_ (.A(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__o21bai_4 _2671_ (.A1(_0654_),
    .A2(_0682_),
    .B1_N(_0692_),
    .Y(_0013_));
 sky130_fd_sc_hd__o31ai_1 _2672_ (.A1(_0622_),
    .A2(_0613_),
    .A3(_2520_),
    .B1(_0651_),
    .Y(_0693_));
 sky130_fd_sc_hd__and3_1 _2673_ (.A(_0626_),
    .B(_0634_),
    .C(_0693_),
    .X(_0694_));
 sky130_fd_sc_hd__buf_4 _2674_ (.A(_0694_),
    .X(_0695_));
 sky130_fd_sc_hd__buf_6 _2675_ (.A(_0695_),
    .X(_0696_));
 sky130_fd_sc_hd__o21bai_4 _2676_ (.A1(_0623_),
    .A2(_0678_),
    .B1_N(_0696_),
    .Y(_0015_));
 sky130_fd_sc_hd__and3_1 _2677_ (.A(_0626_),
    .B(_0634_),
    .C(_0661_),
    .X(_0697_));
 sky130_fd_sc_hd__buf_4 _2678_ (.A(_0697_),
    .X(_0698_));
 sky130_fd_sc_hd__buf_6 _2679_ (.A(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__o21bai_4 _2680_ (.A1(_0624_),
    .A2(_0686_),
    .B1_N(_0699_),
    .Y(_0003_));
 sky130_fd_sc_hd__o21a_1 _2681_ (.A1(_2520_),
    .A2(_0672_),
    .B1(_0673_),
    .X(_0700_));
 sky130_fd_sc_hd__o22ai_4 _2682_ (.A1(_0646_),
    .A2(_0700_),
    .B1(_0686_),
    .B2(_0653_),
    .Y(_0004_));
 sky130_fd_sc_hd__and3_1 _2683_ (.A(_0626_),
    .B(_0634_),
    .C(_0674_),
    .X(_0701_));
 sky130_fd_sc_hd__buf_4 _2684_ (.A(_0701_),
    .X(_0702_));
 sky130_fd_sc_hd__buf_6 _2685_ (.A(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__o21bai_4 _2686_ (.A1(_0678_),
    .A2(_0686_),
    .B1_N(_0703_),
    .Y(_0005_));
 sky130_fd_sc_hd__mux2_2 _2687_ (.A0(_0637_),
    .A1(_0638_),
    .S(_2526_),
    .X(_0704_));
 sky130_fd_sc_hd__o22ai_4 _2688_ (.A1(_0704_),
    .A2(_0646_),
    .B1(_0654_),
    .B2(_0623_),
    .Y(_0006_));
 sky130_fd_sc_hd__and3_1 _2689_ (.A(_0626_),
    .B(_0693_),
    .C(_0668_),
    .X(_0705_));
 sky130_fd_sc_hd__buf_4 _2690_ (.A(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__buf_6 _2691_ (.A(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__o21bai_4 _2692_ (.A1(_0678_),
    .A2(_0682_),
    .B1_N(_0707_),
    .Y(_0001_));
 sky130_fd_sc_hd__and2_0 _2693_ (.A(_0693_),
    .B(_0657_),
    .X(_0708_));
 sky130_fd_sc_hd__buf_6 _2694_ (.A(_0708_),
    .X(_0709_));
 sky130_fd_sc_hd__buf_6 _2695_ (.A(_0709_),
    .X(_0710_));
 sky130_fd_sc_hd__o21bai_4 _2696_ (.A1(_0653_),
    .A2(_0682_),
    .B1_N(_0710_),
    .Y(_0000_));
 sky130_fd_sc_hd__clkbuf_4 _2697_ (.A(rd_en[0]),
    .X(_0711_));
 sky130_fd_sc_hd__or4b_4 _2698_ (.A(net72),
    .B(_0607_),
    .C(net73),
    .D_N(_2557_),
    .X(_0712_));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net219),
    .X(net166));
 sky130_fd_sc_hd__nand2_8 _2700_ (.A(_0711_),
    .B(_0712_),
    .Y(_0714_));
 sky130_fd_sc_hd__inv_2 _2701_ (.A(_0714_),
    .Y(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0997_));
 sky130_fd_sc_hd__clkbuf_16 _2703_ (.A(_0715_),
    .X(_0529_));
 sky130_fd_sc_hd__inv_1 _2704_ (.A(_2559_),
    .Y(_0717_));
 sky130_fd_sc_hd__or4bb_1 _2705_ (.A(net72),
    .B(net73),
    .C_N(_2559_),
    .D_N(_2515_),
    .X(_0718_));
 sky130_fd_sc_hd__or4bb_4 _2706_ (.A(net72),
    .B(net168),
    .C_N(_2516_),
    .D_N(_2548_),
    .X(_0719_));
 sky130_fd_sc_hd__o2111ai_4 _2707_ (.A1(_0717_),
    .A2(_2557_),
    .B1(_0718_),
    .C1(net2),
    .D1(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__inv_4 _2708_ (.A(_0720_),
    .Y(_0721_));
 sky130_fd_sc_hd__buf_6 _2709_ (.A(_0721_),
    .X(_2537_));
 sky130_fd_sc_hd__buf_6 _2710_ (.A(\rd_ptr[1] ),
    .X(_0722_));
 sky130_fd_sc_hd__inv_1 _2711_ (.A(_0722_),
    .Y(_2492_));
 sky130_fd_sc_hd__clkbuf_2 _2712_ (.A(net3),
    .X(_0723_));
 sky130_fd_sc_hd__buf_2 _2713_ (.A(net28),
    .X(_0724_));
 sky130_fd_sc_hd__mux2_1 _2714_ (.A0(_0723_),
    .A1(_0724_),
    .S(_0696_),
    .X(_0016_));
 sky130_fd_sc_hd__buf_2 _2715_ (.A(net14),
    .X(_0725_));
 sky130_fd_sc_hd__buf_2 _2716_ (.A(net29),
    .X(_0726_));
 sky130_fd_sc_hd__mux2_1 _2717_ (.A0(_0725_),
    .A1(_0726_),
    .S(_0696_),
    .X(_0027_));
 sky130_fd_sc_hd__buf_2 _2718_ (.A(net25),
    .X(_0727_));
 sky130_fd_sc_hd__buf_2 _2719_ (.A(net30),
    .X(_0728_));
 sky130_fd_sc_hd__mux2_1 _2720_ (.A0(_0727_),
    .A1(_0728_),
    .S(_0696_),
    .X(_0038_));
 sky130_fd_sc_hd__clkbuf_2 _2721_ (.A(net36),
    .X(_0729_));
 sky130_fd_sc_hd__buf_2 _2722_ (.A(net31),
    .X(_0730_));
 sky130_fd_sc_hd__mux2_1 _2723_ (.A0(_0729_),
    .A1(_0730_),
    .S(_0696_),
    .X(_0041_));
 sky130_fd_sc_hd__buf_2 _2724_ (.A(net47),
    .X(_0731_));
 sky130_fd_sc_hd__buf_2 _2725_ (.A(net32),
    .X(_0732_));
 sky130_fd_sc_hd__mux2_1 _2726_ (.A0(_0731_),
    .A1(_0732_),
    .S(_0696_),
    .X(_0042_));
 sky130_fd_sc_hd__buf_2 _2727_ (.A(net58),
    .X(_0733_));
 sky130_fd_sc_hd__buf_2 _2728_ (.A(net33),
    .X(_0734_));
 sky130_fd_sc_hd__mux2_1 _2729_ (.A0(_0733_),
    .A1(_0734_),
    .S(_0696_),
    .X(_0043_));
 sky130_fd_sc_hd__clkbuf_2 _2730_ (.A(net63),
    .X(_0735_));
 sky130_fd_sc_hd__buf_2 _2731_ (.A(net34),
    .X(_0736_));
 sky130_fd_sc_hd__mux2_1 _2732_ (.A0(_0735_),
    .A1(_0736_),
    .S(_0696_),
    .X(_0044_));
 sky130_fd_sc_hd__clkbuf_2 _2733_ (.A(net64),
    .X(_0737_));
 sky130_fd_sc_hd__clkbuf_2 _2734_ (.A(net35),
    .X(_0738_));
 sky130_fd_sc_hd__mux2_1 _2735_ (.A0(_0737_),
    .A1(_0738_),
    .S(_0696_),
    .X(_0045_));
 sky130_fd_sc_hd__clkbuf_2 _2736_ (.A(net65),
    .X(_0739_));
 sky130_fd_sc_hd__buf_2 _2737_ (.A(net37),
    .X(_0740_));
 sky130_fd_sc_hd__mux2_1 _2738_ (.A0(_0739_),
    .A1(_0740_),
    .S(_0696_),
    .X(_0046_));
 sky130_fd_sc_hd__buf_2 _2739_ (.A(net66),
    .X(_0741_));
 sky130_fd_sc_hd__buf_2 _2740_ (.A(net38),
    .X(_0742_));
 sky130_fd_sc_hd__buf_6 _2741_ (.A(_0695_),
    .X(_0743_));
 sky130_fd_sc_hd__mux2_1 _2742_ (.A0(_0741_),
    .A1(_0742_),
    .S(_0743_),
    .X(_0047_));
 sky130_fd_sc_hd__clkbuf_2 _2743_ (.A(net4),
    .X(_0744_));
 sky130_fd_sc_hd__buf_2 _2744_ (.A(net39),
    .X(_0745_));
 sky130_fd_sc_hd__mux2_1 _2745_ (.A0(_0744_),
    .A1(_0745_),
    .S(_0743_),
    .X(_0017_));
 sky130_fd_sc_hd__buf_2 _2746_ (.A(net5),
    .X(_0746_));
 sky130_fd_sc_hd__buf_2 _2747_ (.A(net40),
    .X(_0747_));
 sky130_fd_sc_hd__mux2_1 _2748_ (.A0(_0746_),
    .A1(_0747_),
    .S(_0743_),
    .X(_0018_));
 sky130_fd_sc_hd__buf_2 _2749_ (.A(net6),
    .X(_0748_));
 sky130_fd_sc_hd__buf_2 _2750_ (.A(net41),
    .X(_0749_));
 sky130_fd_sc_hd__mux2_1 _2751_ (.A0(_0748_),
    .A1(_0749_),
    .S(_0743_),
    .X(_0019_));
 sky130_fd_sc_hd__buf_2 _2752_ (.A(net7),
    .X(_0750_));
 sky130_fd_sc_hd__buf_2 _2753_ (.A(net42),
    .X(_0751_));
 sky130_fd_sc_hd__mux2_1 _2754_ (.A0(_0750_),
    .A1(_0751_),
    .S(_0743_),
    .X(_0020_));
 sky130_fd_sc_hd__buf_2 _2755_ (.A(net8),
    .X(_0752_));
 sky130_fd_sc_hd__buf_2 _2756_ (.A(net43),
    .X(_0753_));
 sky130_fd_sc_hd__mux2_1 _2757_ (.A0(_0752_),
    .A1(_0753_),
    .S(_0743_),
    .X(_0021_));
 sky130_fd_sc_hd__buf_2 _2758_ (.A(net9),
    .X(_0754_));
 sky130_fd_sc_hd__buf_2 _2759_ (.A(net44),
    .X(_0755_));
 sky130_fd_sc_hd__mux2_1 _2760_ (.A0(_0754_),
    .A1(_0755_),
    .S(_0743_),
    .X(_0022_));
 sky130_fd_sc_hd__buf_2 _2761_ (.A(net10),
    .X(_0756_));
 sky130_fd_sc_hd__buf_2 _2762_ (.A(net45),
    .X(_0757_));
 sky130_fd_sc_hd__mux2_1 _2763_ (.A0(_0756_),
    .A1(_0757_),
    .S(_0743_),
    .X(_0023_));
 sky130_fd_sc_hd__buf_2 _2764_ (.A(net11),
    .X(_0758_));
 sky130_fd_sc_hd__buf_2 _2765_ (.A(net46),
    .X(_0759_));
 sky130_fd_sc_hd__mux2_1 _2766_ (.A0(_0758_),
    .A1(_0759_),
    .S(_0743_),
    .X(_0024_));
 sky130_fd_sc_hd__clkbuf_2 _2767_ (.A(net12),
    .X(_0760_));
 sky130_fd_sc_hd__buf_2 _2768_ (.A(net48),
    .X(_0761_));
 sky130_fd_sc_hd__mux2_1 _2769_ (.A0(_0760_),
    .A1(_0761_),
    .S(_0743_),
    .X(_0025_));
 sky130_fd_sc_hd__buf_2 _2770_ (.A(net13),
    .X(_0762_));
 sky130_fd_sc_hd__buf_2 _2771_ (.A(net49),
    .X(_0763_));
 sky130_fd_sc_hd__buf_4 _2772_ (.A(_0695_),
    .X(_0764_));
 sky130_fd_sc_hd__mux2_1 _2773_ (.A0(_0762_),
    .A1(_0763_),
    .S(_0764_),
    .X(_0026_));
 sky130_fd_sc_hd__buf_2 _2774_ (.A(net15),
    .X(_0765_));
 sky130_fd_sc_hd__buf_2 _2775_ (.A(net50),
    .X(_0766_));
 sky130_fd_sc_hd__mux2_1 _2776_ (.A0(_0765_),
    .A1(_0766_),
    .S(_0764_),
    .X(_0028_));
 sky130_fd_sc_hd__buf_2 _2777_ (.A(net16),
    .X(_0767_));
 sky130_fd_sc_hd__buf_2 _2778_ (.A(net51),
    .X(_0768_));
 sky130_fd_sc_hd__mux2_1 _2779_ (.A0(_0767_),
    .A1(_0768_),
    .S(_0764_),
    .X(_0029_));
 sky130_fd_sc_hd__buf_2 _2780_ (.A(net17),
    .X(_0769_));
 sky130_fd_sc_hd__buf_2 _2781_ (.A(net52),
    .X(_0770_));
 sky130_fd_sc_hd__mux2_1 _2782_ (.A0(_0769_),
    .A1(_0770_),
    .S(_0764_),
    .X(_0030_));
 sky130_fd_sc_hd__buf_2 _2783_ (.A(net18),
    .X(_0771_));
 sky130_fd_sc_hd__buf_2 _2784_ (.A(net53),
    .X(_0772_));
 sky130_fd_sc_hd__mux2_1 _2785_ (.A0(_0771_),
    .A1(_0772_),
    .S(_0764_),
    .X(_0031_));
 sky130_fd_sc_hd__clkbuf_2 _2786_ (.A(net19),
    .X(_0773_));
 sky130_fd_sc_hd__clkbuf_2 _2787_ (.A(net54),
    .X(_0774_));
 sky130_fd_sc_hd__mux2_1 _2788_ (.A0(_0773_),
    .A1(_0774_),
    .S(_0764_),
    .X(_0032_));
 sky130_fd_sc_hd__buf_2 _2789_ (.A(net20),
    .X(_0775_));
 sky130_fd_sc_hd__clkbuf_4 _2790_ (.A(net55),
    .X(_0776_));
 sky130_fd_sc_hd__mux2_1 _2791_ (.A0(_0775_),
    .A1(_0776_),
    .S(_0764_),
    .X(_0033_));
 sky130_fd_sc_hd__buf_2 _2792_ (.A(net21),
    .X(_0777_));
 sky130_fd_sc_hd__buf_2 _2793_ (.A(net56),
    .X(_0778_));
 sky130_fd_sc_hd__mux2_1 _2794_ (.A0(_0777_),
    .A1(_0778_),
    .S(_0764_),
    .X(_0034_));
 sky130_fd_sc_hd__buf_2 _2795_ (.A(net22),
    .X(_0779_));
 sky130_fd_sc_hd__buf_2 _2796_ (.A(net57),
    .X(_0780_));
 sky130_fd_sc_hd__mux2_1 _2797_ (.A0(_0779_),
    .A1(_0780_),
    .S(_0764_),
    .X(_0035_));
 sky130_fd_sc_hd__buf_2 _2798_ (.A(net23),
    .X(_0781_));
 sky130_fd_sc_hd__buf_2 _2799_ (.A(net59),
    .X(_0782_));
 sky130_fd_sc_hd__mux2_1 _2800_ (.A0(_0781_),
    .A1(_0782_),
    .S(_0764_),
    .X(_0036_));
 sky130_fd_sc_hd__buf_2 _2801_ (.A(net24),
    .X(_0783_));
 sky130_fd_sc_hd__buf_2 _2802_ (.A(net60),
    .X(_0784_));
 sky130_fd_sc_hd__mux2_1 _2803_ (.A0(_0783_),
    .A1(_0784_),
    .S(_0695_),
    .X(_0037_));
 sky130_fd_sc_hd__buf_2 _2804_ (.A(net26),
    .X(_0785_));
 sky130_fd_sc_hd__buf_2 _2805_ (.A(net61),
    .X(_0786_));
 sky130_fd_sc_hd__mux2_1 _2806_ (.A0(_0785_),
    .A1(_0786_),
    .S(_0695_),
    .X(_0039_));
 sky130_fd_sc_hd__buf_2 _2807_ (.A(net27),
    .X(_0787_));
 sky130_fd_sc_hd__buf_2 _2808_ (.A(net62),
    .X(_0788_));
 sky130_fd_sc_hd__mux2_1 _2809_ (.A0(_0787_),
    .A1(_0788_),
    .S(_0695_),
    .X(_0040_));
 sky130_fd_sc_hd__nor2_4 _2810_ (.A(_0646_),
    .B(_0652_),
    .Y(_0789_));
 sky130_fd_sc_hd__buf_6 _2811_ (.A(_0789_),
    .X(_0790_));
 sky130_fd_sc_hd__mux2_1 _2812_ (.A0(_0723_),
    .A1(_0724_),
    .S(_0790_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _2813_ (.A0(_0725_),
    .A1(_0726_),
    .S(_0790_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _2814_ (.A0(_0727_),
    .A1(_0728_),
    .S(_0790_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _2815_ (.A0(_0729_),
    .A1(_0730_),
    .S(_0790_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _2816_ (.A0(_0731_),
    .A1(_0732_),
    .S(_0790_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _2817_ (.A0(_0733_),
    .A1(_0734_),
    .S(_0790_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _2818_ (.A0(_0735_),
    .A1(_0736_),
    .S(_0790_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _2819_ (.A0(_0737_),
    .A1(_0738_),
    .S(_0790_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _2820_ (.A0(_0739_),
    .A1(_0740_),
    .S(_0790_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _2821_ (.A0(_0741_),
    .A1(_0742_),
    .S(_0790_),
    .X(_0271_));
 sky130_fd_sc_hd__buf_6 _2822_ (.A(_0789_),
    .X(_0791_));
 sky130_fd_sc_hd__mux2_1 _2823_ (.A0(_0744_),
    .A1(_0745_),
    .S(_0791_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _2824_ (.A0(_0746_),
    .A1(_0747_),
    .S(_0791_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _2825_ (.A0(_0748_),
    .A1(_0749_),
    .S(_0791_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _2826_ (.A0(_0750_),
    .A1(_0751_),
    .S(_0791_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _2827_ (.A0(_0752_),
    .A1(_0753_),
    .S(_0791_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _2828_ (.A0(_0754_),
    .A1(_0755_),
    .S(_0791_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _2829_ (.A0(_0756_),
    .A1(_0757_),
    .S(_0791_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _2830_ (.A0(_0758_),
    .A1(_0759_),
    .S(_0791_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _2831_ (.A0(_0760_),
    .A1(_0761_),
    .S(_0791_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _2832_ (.A0(_0762_),
    .A1(_0763_),
    .S(_0791_),
    .X(_0250_));
 sky130_fd_sc_hd__buf_6 _2833_ (.A(_0789_),
    .X(_0792_));
 sky130_fd_sc_hd__mux2_1 _2834_ (.A0(_0765_),
    .A1(_0766_),
    .S(_0792_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _2835_ (.A0(_0767_),
    .A1(_0768_),
    .S(_0792_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _2836_ (.A0(_0769_),
    .A1(_0770_),
    .S(_0792_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _2837_ (.A0(_0771_),
    .A1(_0772_),
    .S(_0792_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _2838_ (.A0(_0773_),
    .A1(_0774_),
    .S(_0792_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _2839_ (.A0(_0775_),
    .A1(_0776_),
    .S(_0792_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _2840_ (.A0(_0777_),
    .A1(_0778_),
    .S(_0792_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _2841_ (.A0(_0779_),
    .A1(_0780_),
    .S(_0792_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _2842_ (.A0(_0781_),
    .A1(_0782_),
    .S(_0792_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _2843_ (.A0(_0783_),
    .A1(_0784_),
    .S(_0792_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _2844_ (.A0(_0785_),
    .A1(_0786_),
    .S(_0789_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _2845_ (.A0(_0787_),
    .A1(_0788_),
    .S(_0789_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _2846_ (.A0(_0723_),
    .A1(_0724_),
    .S(_0642_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _2847_ (.A0(_0725_),
    .A1(_0726_),
    .S(_0642_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _2848_ (.A0(_0727_),
    .A1(_0728_),
    .S(_0642_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _2849_ (.A0(_0729_),
    .A1(_0730_),
    .S(_0642_),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _2850_ (.A0(_0731_),
    .A1(_0732_),
    .S(_0642_),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _2851_ (.A0(_0733_),
    .A1(_0734_),
    .S(_0642_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _2852_ (.A0(_0735_),
    .A1(_0736_),
    .S(_0642_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _2853_ (.A0(_0737_),
    .A1(_0738_),
    .S(_0642_),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _2854_ (.A0(_0739_),
    .A1(_0740_),
    .S(_0642_),
    .X(_0302_));
 sky130_fd_sc_hd__buf_6 _2855_ (.A(_0641_),
    .X(_0793_));
 sky130_fd_sc_hd__mux2_1 _2856_ (.A0(_0741_),
    .A1(_0742_),
    .S(_0793_),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _2857_ (.A0(_0744_),
    .A1(_0745_),
    .S(_0793_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _2858_ (.A0(_0746_),
    .A1(_0747_),
    .S(_0793_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _2859_ (.A0(_0748_),
    .A1(_0749_),
    .S(_0793_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _2860_ (.A0(_0750_),
    .A1(_0751_),
    .S(_0793_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _2861_ (.A0(_0752_),
    .A1(_0753_),
    .S(_0793_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _2862_ (.A0(_0754_),
    .A1(_0755_),
    .S(_0793_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _2863_ (.A0(_0756_),
    .A1(_0757_),
    .S(_0793_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _2864_ (.A0(_0758_),
    .A1(_0759_),
    .S(_0793_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _2865_ (.A0(_0760_),
    .A1(_0761_),
    .S(_0793_),
    .X(_0281_));
 sky130_fd_sc_hd__buf_4 _2866_ (.A(_0641_),
    .X(_0794_));
 sky130_fd_sc_hd__mux2_1 _2867_ (.A0(_0762_),
    .A1(_0763_),
    .S(_0794_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _2868_ (.A0(_0765_),
    .A1(_0766_),
    .S(_0794_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _2869_ (.A0(_0767_),
    .A1(_0768_),
    .S(_0794_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _2870_ (.A0(_0769_),
    .A1(_0770_),
    .S(_0794_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _2871_ (.A0(_0771_),
    .A1(_0772_),
    .S(_0794_),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _2872_ (.A0(_0773_),
    .A1(_0774_),
    .S(_0794_),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _2873_ (.A0(_0775_),
    .A1(_0776_),
    .S(_0794_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _2874_ (.A0(_0777_),
    .A1(_0778_),
    .S(_0794_),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _2875_ (.A0(_0779_),
    .A1(_0780_),
    .S(_0794_),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _2876_ (.A0(_0781_),
    .A1(_0782_),
    .S(_0794_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _2877_ (.A0(_0783_),
    .A1(_0784_),
    .S(_0641_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _2878_ (.A0(_0785_),
    .A1(_0786_),
    .S(_0641_),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _2879_ (.A0(_0787_),
    .A1(_0788_),
    .S(_0641_),
    .X(_0296_));
 sky130_fd_sc_hd__nor2_4 _2880_ (.A(_0704_),
    .B(_0646_),
    .Y(_0795_));
 sky130_fd_sc_hd__buf_6 _2881_ (.A(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__mux2_1 _2882_ (.A0(_0723_),
    .A1(_0724_),
    .S(_0796_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _2883_ (.A0(_0725_),
    .A1(_0726_),
    .S(_0796_),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _2884_ (.A0(_0727_),
    .A1(_0728_),
    .S(_0796_),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _2885_ (.A0(_0729_),
    .A1(_0730_),
    .S(_0796_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _2886_ (.A0(_0731_),
    .A1(_0732_),
    .S(_0796_),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _2887_ (.A0(_0733_),
    .A1(_0734_),
    .S(_0796_),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _2888_ (.A0(_0735_),
    .A1(_0736_),
    .S(_0796_),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _2889_ (.A0(_0737_),
    .A1(_0738_),
    .S(_0796_),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _2890_ (.A0(_0739_),
    .A1(_0740_),
    .S(_0796_),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _2891_ (.A0(_0741_),
    .A1(_0742_),
    .S(_0796_),
    .X(_0335_));
 sky130_fd_sc_hd__buf_6 _2892_ (.A(_0795_),
    .X(_0797_));
 sky130_fd_sc_hd__mux2_1 _2893_ (.A0(_0744_),
    .A1(_0745_),
    .S(_0797_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _2894_ (.A0(_0746_),
    .A1(_0747_),
    .S(_0797_),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _2895_ (.A0(_0748_),
    .A1(_0749_),
    .S(_0797_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _2896_ (.A0(_0750_),
    .A1(_0751_),
    .S(_0797_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _2897_ (.A0(_0752_),
    .A1(_0753_),
    .S(_0797_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _2898_ (.A0(_0754_),
    .A1(_0755_),
    .S(_0797_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _2899_ (.A0(_0756_),
    .A1(_0757_),
    .S(_0797_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _2900_ (.A0(_0758_),
    .A1(_0759_),
    .S(_0797_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _2901_ (.A0(_0760_),
    .A1(_0761_),
    .S(_0797_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _2902_ (.A0(_0762_),
    .A1(_0763_),
    .S(_0797_),
    .X(_0314_));
 sky130_fd_sc_hd__clkbuf_8 _2903_ (.A(_0795_),
    .X(_0798_));
 sky130_fd_sc_hd__mux2_1 _2904_ (.A0(_0765_),
    .A1(_0766_),
    .S(_0798_),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _2905_ (.A0(_0767_),
    .A1(_0768_),
    .S(_0798_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _2906_ (.A0(_0769_),
    .A1(_0770_),
    .S(_0798_),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _2907_ (.A0(_0771_),
    .A1(_0772_),
    .S(_0798_),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _2908_ (.A0(_0773_),
    .A1(_0774_),
    .S(_0798_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _2909_ (.A0(_0775_),
    .A1(_0776_),
    .S(_0798_),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _2910_ (.A0(_0777_),
    .A1(_0778_),
    .S(_0798_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _2911_ (.A0(_0779_),
    .A1(_0780_),
    .S(_0798_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _2912_ (.A0(_0781_),
    .A1(_0782_),
    .S(_0798_),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _2913_ (.A0(_0783_),
    .A1(_0784_),
    .S(_0798_),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _2914_ (.A0(_0785_),
    .A1(_0786_),
    .S(_0795_),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _2915_ (.A0(_0787_),
    .A1(_0788_),
    .S(_0795_),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _2916_ (.A0(_0723_),
    .A1(_0724_),
    .S(_0703_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _2917_ (.A0(_0725_),
    .A1(_0726_),
    .S(_0703_),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _2918_ (.A0(_0727_),
    .A1(_0728_),
    .S(_0703_),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _2919_ (.A0(_0729_),
    .A1(_0730_),
    .S(_0703_),
    .X(_0361_));
 sky130_fd_sc_hd__mux2_1 _2920_ (.A0(_0731_),
    .A1(_0732_),
    .S(_0703_),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_1 _2921_ (.A0(_0733_),
    .A1(_0734_),
    .S(_0703_),
    .X(_0363_));
 sky130_fd_sc_hd__mux2_1 _2922_ (.A0(_0735_),
    .A1(_0736_),
    .S(_0703_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _2923_ (.A0(_0737_),
    .A1(_0738_),
    .S(_0703_),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _2924_ (.A0(_0739_),
    .A1(_0740_),
    .S(_0703_),
    .X(_0366_));
 sky130_fd_sc_hd__buf_6 _2925_ (.A(_0702_),
    .X(_0799_));
 sky130_fd_sc_hd__mux2_1 _2926_ (.A0(_0741_),
    .A1(_0742_),
    .S(_0799_),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _2927_ (.A0(_0744_),
    .A1(_0745_),
    .S(_0799_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _2928_ (.A0(_0746_),
    .A1(_0747_),
    .S(_0799_),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _2929_ (.A0(_0748_),
    .A1(_0749_),
    .S(_0799_),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _2930_ (.A0(_0750_),
    .A1(_0751_),
    .S(_0799_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _2931_ (.A0(_0752_),
    .A1(_0753_),
    .S(_0799_),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _2932_ (.A0(_0754_),
    .A1(_0755_),
    .S(_0799_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _2933_ (.A0(_0756_),
    .A1(_0757_),
    .S(_0799_),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _2934_ (.A0(_0758_),
    .A1(_0759_),
    .S(_0799_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _2935_ (.A0(_0760_),
    .A1(_0761_),
    .S(_0799_),
    .X(_0345_));
 sky130_fd_sc_hd__clkbuf_8 _2936_ (.A(_0702_),
    .X(_0800_));
 sky130_fd_sc_hd__mux2_1 _2937_ (.A0(_0762_),
    .A1(_0763_),
    .S(_0800_),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _2938_ (.A0(_0765_),
    .A1(_0766_),
    .S(_0800_),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _2939_ (.A0(_0767_),
    .A1(_0768_),
    .S(_0800_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _2940_ (.A0(_0769_),
    .A1(_0770_),
    .S(_0800_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _2941_ (.A0(_0771_),
    .A1(_0772_),
    .S(_0800_),
    .X(_0351_));
 sky130_fd_sc_hd__mux2_1 _2942_ (.A0(_0773_),
    .A1(_0774_),
    .S(_0800_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _2943_ (.A0(_0775_),
    .A1(_0776_),
    .S(_0800_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _2944_ (.A0(_0777_),
    .A1(_0778_),
    .S(_0800_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _2945_ (.A0(_0779_),
    .A1(_0780_),
    .S(_0800_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _2946_ (.A0(_0781_),
    .A1(_0782_),
    .S(_0800_),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _2947_ (.A0(_0783_),
    .A1(_0784_),
    .S(_0702_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _2948_ (.A0(_0785_),
    .A1(_0786_),
    .S(_0702_),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _2949_ (.A0(_0787_),
    .A1(_0788_),
    .S(_0702_),
    .X(_0360_));
 sky130_fd_sc_hd__nor2_4 _2950_ (.A(_0646_),
    .B(_0700_),
    .Y(_0801_));
 sky130_fd_sc_hd__buf_6 _2951_ (.A(_0801_),
    .X(_0802_));
 sky130_fd_sc_hd__mux2_1 _2952_ (.A0(_0723_),
    .A1(_0724_),
    .S(_0802_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _2953_ (.A0(_0725_),
    .A1(_0726_),
    .S(_0802_),
    .X(_0379_));
 sky130_fd_sc_hd__mux2_1 _2954_ (.A0(_0727_),
    .A1(_0728_),
    .S(_0802_),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_1 _2955_ (.A0(_0729_),
    .A1(_0730_),
    .S(_0802_),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_1 _2956_ (.A0(_0731_),
    .A1(_0732_),
    .S(_0802_),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _2957_ (.A0(_0733_),
    .A1(_0734_),
    .S(_0802_),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _2958_ (.A0(_0735_),
    .A1(_0736_),
    .S(_0802_),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _2959_ (.A0(_0737_),
    .A1(_0738_),
    .S(_0802_),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _2960_ (.A0(_0739_),
    .A1(_0740_),
    .S(_0802_),
    .X(_0398_));
 sky130_fd_sc_hd__mux2_1 _2961_ (.A0(_0741_),
    .A1(_0742_),
    .S(_0802_),
    .X(_0399_));
 sky130_fd_sc_hd__buf_6 _2962_ (.A(_0801_),
    .X(_0803_));
 sky130_fd_sc_hd__mux2_1 _2963_ (.A0(_0744_),
    .A1(_0745_),
    .S(_0803_),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _2964_ (.A0(_0746_),
    .A1(_0747_),
    .S(_0803_),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _2965_ (.A0(_0748_),
    .A1(_0749_),
    .S(_0803_),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_1 _2966_ (.A0(_0750_),
    .A1(_0751_),
    .S(_0803_),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _2967_ (.A0(_0752_),
    .A1(_0753_),
    .S(_0803_),
    .X(_0373_));
 sky130_fd_sc_hd__mux2_1 _2968_ (.A0(_0754_),
    .A1(_0755_),
    .S(_0803_),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_1 _2969_ (.A0(_0756_),
    .A1(_0757_),
    .S(_0803_),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_1 _2970_ (.A0(_0758_),
    .A1(_0759_),
    .S(_0803_),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _2971_ (.A0(_0760_),
    .A1(_0761_),
    .S(_0803_),
    .X(_0377_));
 sky130_fd_sc_hd__mux2_1 _2972_ (.A0(_0762_),
    .A1(_0763_),
    .S(_0803_),
    .X(_0378_));
 sky130_fd_sc_hd__buf_6 _2973_ (.A(_0801_),
    .X(_0804_));
 sky130_fd_sc_hd__mux2_1 _2974_ (.A0(_0765_),
    .A1(_0766_),
    .S(_0804_),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_1 _2975_ (.A0(_0767_),
    .A1(_0768_),
    .S(_0804_),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _2976_ (.A0(_0769_),
    .A1(_0770_),
    .S(_0804_),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _2977_ (.A0(_0771_),
    .A1(_0772_),
    .S(_0804_),
    .X(_0383_));
 sky130_fd_sc_hd__mux2_1 _2978_ (.A0(_0773_),
    .A1(_0774_),
    .S(_0804_),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_1 _2979_ (.A0(_0775_),
    .A1(_0776_),
    .S(_0804_),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_1 _2980_ (.A0(_0777_),
    .A1(_0778_),
    .S(_0804_),
    .X(_0386_));
 sky130_fd_sc_hd__mux2_1 _2981_ (.A0(_0779_),
    .A1(_0780_),
    .S(_0804_),
    .X(_0387_));
 sky130_fd_sc_hd__mux2_1 _2982_ (.A0(_0781_),
    .A1(_0782_),
    .S(_0804_),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _2983_ (.A0(_0783_),
    .A1(_0784_),
    .S(_0804_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _2984_ (.A0(_0785_),
    .A1(_0786_),
    .S(_0801_),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_1 _2985_ (.A0(_0787_),
    .A1(_0788_),
    .S(_0801_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _2986_ (.A0(_0723_),
    .A1(_0724_),
    .S(_0699_),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_1 _2987_ (.A0(_0725_),
    .A1(_0726_),
    .S(_0699_),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _2988_ (.A0(_0727_),
    .A1(_0728_),
    .S(_0699_),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_1 _2989_ (.A0(_0729_),
    .A1(_0730_),
    .S(_0699_),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _2990_ (.A0(_0731_),
    .A1(_0732_),
    .S(_0699_),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _2991_ (.A0(_0733_),
    .A1(_0734_),
    .S(_0699_),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _2992_ (.A0(_0735_),
    .A1(_0736_),
    .S(_0699_),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_1 _2993_ (.A0(_0737_),
    .A1(_0738_),
    .S(_0699_),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _2994_ (.A0(_0739_),
    .A1(_0740_),
    .S(_0699_),
    .X(_0430_));
 sky130_fd_sc_hd__buf_6 _2995_ (.A(_0698_),
    .X(_0805_));
 sky130_fd_sc_hd__mux2_1 _2996_ (.A0(_0741_),
    .A1(_0742_),
    .S(_0805_),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _2997_ (.A0(_0744_),
    .A1(_0745_),
    .S(_0805_),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_1 _2998_ (.A0(_0746_),
    .A1(_0747_),
    .S(_0805_),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_1 _2999_ (.A0(_0748_),
    .A1(_0749_),
    .S(_0805_),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_1 _3000_ (.A0(_0750_),
    .A1(_0751_),
    .S(_0805_),
    .X(_0404_));
 sky130_fd_sc_hd__mux2_1 _3001_ (.A0(_0752_),
    .A1(_0753_),
    .S(_0805_),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _3002_ (.A0(_0754_),
    .A1(_0755_),
    .S(_0805_),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _3003_ (.A0(_0756_),
    .A1(_0757_),
    .S(_0805_),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _3004_ (.A0(_0758_),
    .A1(_0759_),
    .S(_0805_),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_1 _3005_ (.A0(_0760_),
    .A1(_0761_),
    .S(_0805_),
    .X(_0409_));
 sky130_fd_sc_hd__clkbuf_8 _3006_ (.A(_0698_),
    .X(_0806_));
 sky130_fd_sc_hd__mux2_1 _3007_ (.A0(_0762_),
    .A1(_0763_),
    .S(_0806_),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _3008_ (.A0(_0765_),
    .A1(_0766_),
    .S(_0806_),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _3009_ (.A0(_0767_),
    .A1(_0768_),
    .S(_0806_),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _3010_ (.A0(_0769_),
    .A1(_0770_),
    .S(_0806_),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _3011_ (.A0(_0771_),
    .A1(_0772_),
    .S(_0806_),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _3012_ (.A0(_0773_),
    .A1(_0774_),
    .S(_0806_),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _3013_ (.A0(_0775_),
    .A1(_0776_),
    .S(_0806_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _3014_ (.A0(_0777_),
    .A1(_0778_),
    .S(_0806_),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _3015_ (.A0(_0779_),
    .A1(_0780_),
    .S(_0806_),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_1 _3016_ (.A0(_0781_),
    .A1(_0782_),
    .S(_0806_),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _3017_ (.A0(_0783_),
    .A1(_0784_),
    .S(_0698_),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _3018_ (.A0(_0785_),
    .A1(_0786_),
    .S(_0698_),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _3019_ (.A0(_0787_),
    .A1(_0788_),
    .S(_0698_),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _3020_ (.A0(_0723_),
    .A1(_0724_),
    .S(_0689_),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_1 _3021_ (.A0(_0725_),
    .A1(_0726_),
    .S(_0689_),
    .X(_0443_));
 sky130_fd_sc_hd__mux2_1 _3022_ (.A0(_0727_),
    .A1(_0728_),
    .S(_0689_),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_1 _3023_ (.A0(_0729_),
    .A1(_0730_),
    .S(_0689_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _3024_ (.A0(_0731_),
    .A1(_0732_),
    .S(_0689_),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _3025_ (.A0(_0733_),
    .A1(_0734_),
    .S(_0689_),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _3026_ (.A0(_0735_),
    .A1(_0736_),
    .S(_0689_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _3027_ (.A0(_0737_),
    .A1(_0738_),
    .S(_0689_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _3028_ (.A0(_0739_),
    .A1(_0740_),
    .S(_0689_),
    .X(_0462_));
 sky130_fd_sc_hd__buf_6 _3029_ (.A(_0688_),
    .X(_0807_));
 sky130_fd_sc_hd__mux2_1 _3030_ (.A0(_0741_),
    .A1(_0742_),
    .S(_0807_),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _3031_ (.A0(_0744_),
    .A1(_0745_),
    .S(_0807_),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _3032_ (.A0(_0746_),
    .A1(_0747_),
    .S(_0807_),
    .X(_0434_));
 sky130_fd_sc_hd__mux2_1 _3033_ (.A0(_0748_),
    .A1(_0749_),
    .S(_0807_),
    .X(_0435_));
 sky130_fd_sc_hd__mux2_1 _3034_ (.A0(_0750_),
    .A1(_0751_),
    .S(_0807_),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_1 _3035_ (.A0(_0752_),
    .A1(_0753_),
    .S(_0807_),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _3036_ (.A0(_0754_),
    .A1(_0755_),
    .S(_0807_),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_1 _3037_ (.A0(_0756_),
    .A1(_0757_),
    .S(_0807_),
    .X(_0439_));
 sky130_fd_sc_hd__mux2_1 _3038_ (.A0(_0758_),
    .A1(_0759_),
    .S(_0807_),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _3039_ (.A0(_0760_),
    .A1(_0761_),
    .S(_0807_),
    .X(_0441_));
 sky130_fd_sc_hd__clkbuf_8 _3040_ (.A(_0688_),
    .X(_0808_));
 sky130_fd_sc_hd__mux2_1 _3041_ (.A0(_0762_),
    .A1(_0763_),
    .S(_0808_),
    .X(_0442_));
 sky130_fd_sc_hd__mux2_1 _3042_ (.A0(_0765_),
    .A1(_0766_),
    .S(_0808_),
    .X(_0444_));
 sky130_fd_sc_hd__mux2_1 _3043_ (.A0(_0767_),
    .A1(_0768_),
    .S(_0808_),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _3044_ (.A0(_0769_),
    .A1(_0770_),
    .S(_0808_),
    .X(_0446_));
 sky130_fd_sc_hd__mux2_1 _3045_ (.A0(_0771_),
    .A1(_0772_),
    .S(_0808_),
    .X(_0447_));
 sky130_fd_sc_hd__mux2_1 _3046_ (.A0(_0773_),
    .A1(_0774_),
    .S(_0808_),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _3047_ (.A0(_0775_),
    .A1(_0776_),
    .S(_0808_),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _3048_ (.A0(_0777_),
    .A1(_0778_),
    .S(_0808_),
    .X(_0450_));
 sky130_fd_sc_hd__mux2_1 _3049_ (.A0(_0779_),
    .A1(_0780_),
    .S(_0808_),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _3050_ (.A0(_0781_),
    .A1(_0782_),
    .S(_0808_),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _3051_ (.A0(_0783_),
    .A1(_0784_),
    .S(_0688_),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _3052_ (.A0(_0785_),
    .A1(_0786_),
    .S(_0688_),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _3053_ (.A0(_0787_),
    .A1(_0788_),
    .S(_0688_),
    .X(_0456_));
 sky130_fd_sc_hd__mux2_1 _3054_ (.A0(_0723_),
    .A1(_0724_),
    .S(_0707_),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _3055_ (.A0(_0725_),
    .A1(_0726_),
    .S(_0707_),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _3056_ (.A0(_0727_),
    .A1(_0728_),
    .S(_0707_),
    .X(_0486_));
 sky130_fd_sc_hd__mux2_1 _3057_ (.A0(_0729_),
    .A1(_0730_),
    .S(_0707_),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_1 _3058_ (.A0(_0731_),
    .A1(_0732_),
    .S(_0707_),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _3059_ (.A0(_0733_),
    .A1(_0734_),
    .S(_0707_),
    .X(_0491_));
 sky130_fd_sc_hd__mux2_1 _3060_ (.A0(_0735_),
    .A1(_0736_),
    .S(_0707_),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_1 _3061_ (.A0(_0737_),
    .A1(_0738_),
    .S(_0707_),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _3062_ (.A0(_0739_),
    .A1(_0740_),
    .S(_0707_),
    .X(_0494_));
 sky130_fd_sc_hd__buf_6 _3063_ (.A(_0706_),
    .X(_0809_));
 sky130_fd_sc_hd__mux2_1 _3064_ (.A0(_0741_),
    .A1(_0742_),
    .S(_0809_),
    .X(_0495_));
 sky130_fd_sc_hd__mux2_1 _3065_ (.A0(_0744_),
    .A1(_0745_),
    .S(_0809_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _3066_ (.A0(_0746_),
    .A1(_0747_),
    .S(_0809_),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_1 _3067_ (.A0(_0748_),
    .A1(_0749_),
    .S(_0809_),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _3068_ (.A0(_0750_),
    .A1(_0751_),
    .S(_0809_),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_1 _3069_ (.A0(_0752_),
    .A1(_0753_),
    .S(_0809_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _3070_ (.A0(_0754_),
    .A1(_0755_),
    .S(_0809_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _3071_ (.A0(_0756_),
    .A1(_0757_),
    .S(_0809_),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_1 _3072_ (.A0(_0758_),
    .A1(_0759_),
    .S(_0809_),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _3073_ (.A0(_0760_),
    .A1(_0761_),
    .S(_0809_),
    .X(_0473_));
 sky130_fd_sc_hd__buf_6 _3074_ (.A(_0706_),
    .X(_0810_));
 sky130_fd_sc_hd__mux2_1 _3075_ (.A0(_0762_),
    .A1(_0763_),
    .S(_0810_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _3076_ (.A0(_0765_),
    .A1(_0766_),
    .S(_0810_),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_1 _3077_ (.A0(_0767_),
    .A1(_0768_),
    .S(_0810_),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _3078_ (.A0(_0769_),
    .A1(_0770_),
    .S(_0810_),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _3079_ (.A0(_0771_),
    .A1(_0772_),
    .S(_0810_),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _3080_ (.A0(_0773_),
    .A1(_0774_),
    .S(_0810_),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_1 _3081_ (.A0(_0775_),
    .A1(_0776_),
    .S(_0810_),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _3082_ (.A0(_0777_),
    .A1(_0778_),
    .S(_0810_),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _3083_ (.A0(_0779_),
    .A1(_0780_),
    .S(_0810_),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_1 _3084_ (.A0(_0781_),
    .A1(_0782_),
    .S(_0810_),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_1 _3085_ (.A0(_0783_),
    .A1(_0784_),
    .S(_0706_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _3086_ (.A0(_0785_),
    .A1(_0786_),
    .S(_0706_),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _3087_ (.A0(_0787_),
    .A1(_0788_),
    .S(_0706_),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_1 _3088_ (.A0(_0723_),
    .A1(net28),
    .S(_0710_),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_1 _3089_ (.A0(_0725_),
    .A1(net29),
    .S(_0710_),
    .X(_0507_));
 sky130_fd_sc_hd__mux2_1 _3090_ (.A0(_0727_),
    .A1(net30),
    .S(_0710_),
    .X(_0518_));
 sky130_fd_sc_hd__mux2_1 _3091_ (.A0(_0729_),
    .A1(net31),
    .S(_0710_),
    .X(_0521_));
 sky130_fd_sc_hd__mux2_1 _3092_ (.A0(_0731_),
    .A1(net32),
    .S(_0710_),
    .X(_0522_));
 sky130_fd_sc_hd__mux2_1 _3093_ (.A0(_0733_),
    .A1(net33),
    .S(_0710_),
    .X(_0523_));
 sky130_fd_sc_hd__mux2_1 _3094_ (.A0(_0735_),
    .A1(net34),
    .S(_0710_),
    .X(_0524_));
 sky130_fd_sc_hd__mux2_1 _3095_ (.A0(_0737_),
    .A1(net35),
    .S(_0710_),
    .X(_0525_));
 sky130_fd_sc_hd__mux2_1 _3096_ (.A0(_0739_),
    .A1(net37),
    .S(_0710_),
    .X(_0526_));
 sky130_fd_sc_hd__buf_6 _3097_ (.A(_0709_),
    .X(_0811_));
 sky130_fd_sc_hd__mux2_1 _3098_ (.A0(_0741_),
    .A1(net38),
    .S(_0811_),
    .X(_0527_));
 sky130_fd_sc_hd__mux2_1 _3099_ (.A0(_0744_),
    .A1(net39),
    .S(_0811_),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _3100_ (.A0(_0746_),
    .A1(net40),
    .S(_0811_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _3101_ (.A0(_0748_),
    .A1(net41),
    .S(_0811_),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _3102_ (.A0(_0750_),
    .A1(net42),
    .S(_0811_),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_1 _3103_ (.A0(_0752_),
    .A1(net43),
    .S(_0811_),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _3104_ (.A0(_0754_),
    .A1(net44),
    .S(_0811_),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_1 _3105_ (.A0(_0756_),
    .A1(net45),
    .S(_0811_),
    .X(_0503_));
 sky130_fd_sc_hd__mux2_1 _3106_ (.A0(_0758_),
    .A1(net46),
    .S(_0811_),
    .X(_0504_));
 sky130_fd_sc_hd__mux2_1 _3107_ (.A0(_0760_),
    .A1(net48),
    .S(_0811_),
    .X(_0505_));
 sky130_fd_sc_hd__buf_8 _3108_ (.A(_0709_),
    .X(_0812_));
 sky130_fd_sc_hd__mux2_1 _3109_ (.A0(_0762_),
    .A1(net49),
    .S(_0812_),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_1 _3110_ (.A0(_0765_),
    .A1(net50),
    .S(_0812_),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _3111_ (.A0(_0767_),
    .A1(net51),
    .S(_0812_),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _3112_ (.A0(_0769_),
    .A1(net52),
    .S(_0812_),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _3113_ (.A0(_0771_),
    .A1(net53),
    .S(_0812_),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _3114_ (.A0(_0773_),
    .A1(net54),
    .S(_0812_),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _3115_ (.A0(_0775_),
    .A1(net55),
    .S(_0812_),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _3116_ (.A0(_0777_),
    .A1(net56),
    .S(_0812_),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_1 _3117_ (.A0(_0779_),
    .A1(net57),
    .S(_0812_),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _3118_ (.A0(_0781_),
    .A1(net59),
    .S(_0812_),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _3119_ (.A0(_0783_),
    .A1(net60),
    .S(_0709_),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_1 _3120_ (.A0(_0785_),
    .A1(net61),
    .S(_0709_),
    .X(_0519_));
 sky130_fd_sc_hd__mux2_1 _3121_ (.A0(_0787_),
    .A1(net62),
    .S(_0709_),
    .X(_0520_));
 sky130_fd_sc_hd__mux2_1 _3122_ (.A0(net3),
    .A1(net28),
    .S(_0685_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _3123_ (.A0(net14),
    .A1(net29),
    .S(_0685_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _3124_ (.A0(net25),
    .A1(net30),
    .S(_0685_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _3125_ (.A0(net36),
    .A1(net31),
    .S(_0685_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _3126_ (.A0(net47),
    .A1(net32),
    .S(_0685_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _3127_ (.A0(net58),
    .A1(net33),
    .S(_0685_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _3128_ (.A0(net63),
    .A1(net34),
    .S(_0685_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _3129_ (.A0(net64),
    .A1(net35),
    .S(_0685_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _3130_ (.A0(net65),
    .A1(net37),
    .S(_0685_),
    .X(_0078_));
 sky130_fd_sc_hd__buf_8 _3131_ (.A(_0684_),
    .X(_0813_));
 sky130_fd_sc_hd__mux2_1 _3132_ (.A0(net66),
    .A1(net38),
    .S(_0813_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _3133_ (.A0(net4),
    .A1(net39),
    .S(_0813_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _3134_ (.A0(net5),
    .A1(net40),
    .S(_0813_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _3135_ (.A0(net6),
    .A1(net41),
    .S(_0813_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _3136_ (.A0(net7),
    .A1(net42),
    .S(_0813_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _3137_ (.A0(net8),
    .A1(net43),
    .S(_0813_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _3138_ (.A0(net9),
    .A1(net44),
    .S(_0813_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _3139_ (.A0(net10),
    .A1(net45),
    .S(_0813_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _3140_ (.A0(net11),
    .A1(net46),
    .S(_0813_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _3141_ (.A0(net12),
    .A1(net48),
    .S(_0813_),
    .X(_0057_));
 sky130_fd_sc_hd__buf_6 _3142_ (.A(_0684_),
    .X(_0814_));
 sky130_fd_sc_hd__mux2_1 _3143_ (.A0(net13),
    .A1(net49),
    .S(_0814_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _3144_ (.A0(net15),
    .A1(net50),
    .S(_0814_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _3145_ (.A0(net16),
    .A1(net51),
    .S(_0814_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _3146_ (.A0(net17),
    .A1(net52),
    .S(_0814_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _3147_ (.A0(net18),
    .A1(net53),
    .S(_0814_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _3148_ (.A0(net19),
    .A1(net54),
    .S(_0814_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _3149_ (.A0(net20),
    .A1(net55),
    .S(_0814_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _3150_ (.A0(net21),
    .A1(net56),
    .S(_0814_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _3151_ (.A0(net22),
    .A1(net57),
    .S(_0814_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _3152_ (.A0(net23),
    .A1(net59),
    .S(_0814_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _3153_ (.A0(net24),
    .A1(net60),
    .S(_0684_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _3154_ (.A0(net26),
    .A1(net61),
    .S(_0684_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _3155_ (.A0(net27),
    .A1(net62),
    .S(_0684_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _3156_ (.A0(net3),
    .A1(net28),
    .S(_0692_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _3157_ (.A0(net14),
    .A1(net29),
    .S(_0692_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _3158_ (.A0(net25),
    .A1(net30),
    .S(_0692_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _3159_ (.A0(net36),
    .A1(net31),
    .S(_0692_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _3160_ (.A0(net47),
    .A1(net32),
    .S(_0692_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _3161_ (.A0(net58),
    .A1(net33),
    .S(_0692_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _3162_ (.A0(net63),
    .A1(net34),
    .S(_0692_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _3163_ (.A0(net64),
    .A1(net35),
    .S(_0692_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _3164_ (.A0(net65),
    .A1(net37),
    .S(_0692_),
    .X(_0110_));
 sky130_fd_sc_hd__buf_6 _3165_ (.A(_0691_),
    .X(_0815_));
 sky130_fd_sc_hd__mux2_1 _3166_ (.A0(net66),
    .A1(net38),
    .S(_0815_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _3167_ (.A0(net4),
    .A1(net39),
    .S(_0815_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _3168_ (.A0(net5),
    .A1(net40),
    .S(_0815_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _3169_ (.A0(net6),
    .A1(net41),
    .S(_0815_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _3170_ (.A0(net7),
    .A1(net42),
    .S(_0815_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _3171_ (.A0(net8),
    .A1(net43),
    .S(_0815_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _3172_ (.A0(net9),
    .A1(net44),
    .S(_0815_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _3173_ (.A0(net10),
    .A1(net45),
    .S(_0815_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _3174_ (.A0(net11),
    .A1(net46),
    .S(_0815_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _3175_ (.A0(net12),
    .A1(net48),
    .S(_0815_),
    .X(_0089_));
 sky130_fd_sc_hd__buf_6 _3176_ (.A(_0691_),
    .X(_0816_));
 sky130_fd_sc_hd__mux2_1 _3177_ (.A0(net13),
    .A1(net49),
    .S(_0816_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _3178_ (.A0(net15),
    .A1(net50),
    .S(_0816_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _3179_ (.A0(net16),
    .A1(net51),
    .S(_0816_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _3180_ (.A0(net17),
    .A1(net52),
    .S(_0816_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _3181_ (.A0(net18),
    .A1(net53),
    .S(_0816_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _3182_ (.A0(net19),
    .A1(net54),
    .S(_0816_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _3183_ (.A0(net20),
    .A1(net55),
    .S(_0816_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _3184_ (.A0(net21),
    .A1(net56),
    .S(_0816_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _3185_ (.A0(net22),
    .A1(net57),
    .S(_0816_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _3186_ (.A0(net23),
    .A1(net59),
    .S(_0816_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _3187_ (.A0(net24),
    .A1(net60),
    .S(_0691_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _3188_ (.A0(net26),
    .A1(net61),
    .S(_0691_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _3189_ (.A0(net27),
    .A1(net62),
    .S(_0691_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _3190_ (.A0(net3),
    .A1(net28),
    .S(_0681_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _3191_ (.A0(net14),
    .A1(net29),
    .S(_0681_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _3192_ (.A0(net25),
    .A1(net30),
    .S(_0681_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _3193_ (.A0(net36),
    .A1(net31),
    .S(_0681_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _3194_ (.A0(net47),
    .A1(net32),
    .S(_0681_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _3195_ (.A0(net58),
    .A1(net33),
    .S(_0681_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _3196_ (.A0(net63),
    .A1(net34),
    .S(_0681_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _3197_ (.A0(net64),
    .A1(net35),
    .S(_0681_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _3198_ (.A0(net65),
    .A1(net37),
    .S(_0681_),
    .X(_0142_));
 sky130_fd_sc_hd__buf_6 _3199_ (.A(_0680_),
    .X(_0817_));
 sky130_fd_sc_hd__mux2_1 _3200_ (.A0(net66),
    .A1(net38),
    .S(_0817_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _3201_ (.A0(net4),
    .A1(net39),
    .S(_0817_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _3202_ (.A0(net5),
    .A1(net40),
    .S(_0817_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _3203_ (.A0(net6),
    .A1(net41),
    .S(_0817_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _3204_ (.A0(net7),
    .A1(net42),
    .S(_0817_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _3205_ (.A0(net8),
    .A1(net43),
    .S(_0817_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _3206_ (.A0(net9),
    .A1(net44),
    .S(_0817_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _3207_ (.A0(net10),
    .A1(net45),
    .S(_0817_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _3208_ (.A0(net11),
    .A1(net46),
    .S(_0817_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _3209_ (.A0(net12),
    .A1(net48),
    .S(_0817_),
    .X(_0121_));
 sky130_fd_sc_hd__buf_8 _3210_ (.A(_0680_),
    .X(_0818_));
 sky130_fd_sc_hd__mux2_1 _3211_ (.A0(net13),
    .A1(net49),
    .S(_0818_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _3212_ (.A0(net15),
    .A1(net50),
    .S(_0818_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _3213_ (.A0(net16),
    .A1(net51),
    .S(_0818_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _3214_ (.A0(net17),
    .A1(net52),
    .S(_0818_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _3215_ (.A0(net18),
    .A1(net53),
    .S(_0818_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _3216_ (.A0(net19),
    .A1(net54),
    .S(_0818_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _3217_ (.A0(net20),
    .A1(net55),
    .S(_0818_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _3218_ (.A0(net21),
    .A1(net56),
    .S(_0818_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _3219_ (.A0(net22),
    .A1(net57),
    .S(_0818_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _3220_ (.A0(net23),
    .A1(net59),
    .S(_0818_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _3221_ (.A0(net24),
    .A1(net60),
    .S(_0680_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _3222_ (.A0(net26),
    .A1(net61),
    .S(_0680_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _3223_ (.A0(net27),
    .A1(net62),
    .S(_0680_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _3224_ (.A0(net3),
    .A1(net28),
    .S(_0677_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _3225_ (.A0(net14),
    .A1(net29),
    .S(_0677_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _3226_ (.A0(net25),
    .A1(net30),
    .S(_0677_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _3227_ (.A0(net36),
    .A1(net31),
    .S(_0677_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _3228_ (.A0(net47),
    .A1(net32),
    .S(_0677_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _3229_ (.A0(net58),
    .A1(net33),
    .S(_0677_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _3230_ (.A0(net63),
    .A1(net34),
    .S(_0677_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _3231_ (.A0(net64),
    .A1(net35),
    .S(_0677_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _3232_ (.A0(net65),
    .A1(net37),
    .S(_0677_),
    .X(_0174_));
 sky130_fd_sc_hd__buf_8 _3233_ (.A(_0676_),
    .X(_0819_));
 sky130_fd_sc_hd__mux2_1 _3234_ (.A0(net66),
    .A1(net38),
    .S(_0819_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _3235_ (.A0(net4),
    .A1(net39),
    .S(_0819_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _3236_ (.A0(net5),
    .A1(net40),
    .S(_0819_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _3237_ (.A0(net6),
    .A1(net41),
    .S(_0819_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _3238_ (.A0(net7),
    .A1(net42),
    .S(_0819_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _3239_ (.A0(net8),
    .A1(net43),
    .S(_0819_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _3240_ (.A0(net9),
    .A1(net44),
    .S(_0819_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _3241_ (.A0(net10),
    .A1(net45),
    .S(_0819_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _3242_ (.A0(net11),
    .A1(net46),
    .S(_0819_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _3243_ (.A0(net12),
    .A1(net48),
    .S(_0819_),
    .X(_0153_));
 sky130_fd_sc_hd__buf_8 _3244_ (.A(_0676_),
    .X(_0820_));
 sky130_fd_sc_hd__mux2_1 _3245_ (.A0(net13),
    .A1(net49),
    .S(_0820_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _3246_ (.A0(net15),
    .A1(net50),
    .S(_0820_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _3247_ (.A0(net16),
    .A1(net51),
    .S(_0820_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _3248_ (.A0(net17),
    .A1(net52),
    .S(_0820_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _3249_ (.A0(net18),
    .A1(net53),
    .S(_0820_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _3250_ (.A0(net19),
    .A1(net54),
    .S(_0820_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _3251_ (.A0(net20),
    .A1(net55),
    .S(_0820_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _3252_ (.A0(net21),
    .A1(net56),
    .S(_0820_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _3253_ (.A0(net22),
    .A1(net57),
    .S(_0820_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _3254_ (.A0(net23),
    .A1(net59),
    .S(_0820_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _3255_ (.A0(net24),
    .A1(net60),
    .S(_0676_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _3256_ (.A0(net26),
    .A1(net61),
    .S(_0676_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _3257_ (.A0(net27),
    .A1(net62),
    .S(_0676_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _3258_ (.A0(net3),
    .A1(net28),
    .S(_0671_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _3259_ (.A0(net14),
    .A1(net29),
    .S(_0671_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _3260_ (.A0(net25),
    .A1(net30),
    .S(_0671_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _3261_ (.A0(net36),
    .A1(net31),
    .S(_0671_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _3262_ (.A0(net47),
    .A1(net32),
    .S(_0671_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _3263_ (.A0(net58),
    .A1(net33),
    .S(_0671_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _3264_ (.A0(net63),
    .A1(net34),
    .S(_0671_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _3265_ (.A0(net64),
    .A1(net35),
    .S(_0671_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _3266_ (.A0(net65),
    .A1(net37),
    .S(_0671_),
    .X(_0206_));
 sky130_fd_sc_hd__buf_6 _3267_ (.A(_0670_),
    .X(_0821_));
 sky130_fd_sc_hd__mux2_1 _3268_ (.A0(net66),
    .A1(net38),
    .S(_0821_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _3269_ (.A0(net4),
    .A1(net39),
    .S(_0821_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _3270_ (.A0(net5),
    .A1(net40),
    .S(_0821_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _3271_ (.A0(net6),
    .A1(net41),
    .S(_0821_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _3272_ (.A0(net7),
    .A1(net42),
    .S(_0821_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _3273_ (.A0(net8),
    .A1(net43),
    .S(_0821_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _3274_ (.A0(net9),
    .A1(net44),
    .S(_0821_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _3275_ (.A0(net10),
    .A1(net45),
    .S(_0821_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _3276_ (.A0(net11),
    .A1(net46),
    .S(_0821_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _3277_ (.A0(net12),
    .A1(net48),
    .S(_0821_),
    .X(_0185_));
 sky130_fd_sc_hd__buf_8 _3278_ (.A(_0670_),
    .X(_0822_));
 sky130_fd_sc_hd__mux2_1 _3279_ (.A0(net13),
    .A1(net49),
    .S(_0822_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _3280_ (.A0(net15),
    .A1(net50),
    .S(_0822_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _3281_ (.A0(net16),
    .A1(net51),
    .S(_0822_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _3282_ (.A0(net17),
    .A1(net52),
    .S(_0822_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _3283_ (.A0(net18),
    .A1(net53),
    .S(_0822_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _3284_ (.A0(net19),
    .A1(net54),
    .S(_0822_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _3285_ (.A0(net20),
    .A1(net55),
    .S(_0822_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _3286_ (.A0(net21),
    .A1(net56),
    .S(_0822_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _3287_ (.A0(net22),
    .A1(net57),
    .S(_0822_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _3288_ (.A0(net23),
    .A1(net59),
    .S(_0822_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _3289_ (.A0(net24),
    .A1(net60),
    .S(_0670_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _3290_ (.A0(net26),
    .A1(net61),
    .S(_0670_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _3291_ (.A0(net27),
    .A1(net62),
    .S(_0670_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _3292_ (.A0(_0724_),
    .A1(net3),
    .S(_0663_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _3293_ (.A0(_0726_),
    .A1(net14),
    .S(_0663_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _3294_ (.A0(_0728_),
    .A1(net25),
    .S(_0663_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _3295_ (.A0(_0730_),
    .A1(net36),
    .S(_0663_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _3296_ (.A0(_0732_),
    .A1(net47),
    .S(_0663_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _3297_ (.A0(_0734_),
    .A1(net58),
    .S(_0663_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _3298_ (.A0(_0736_),
    .A1(net63),
    .S(_0663_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _3299_ (.A0(_0738_),
    .A1(net64),
    .S(_0663_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _3300_ (.A0(_0740_),
    .A1(net65),
    .S(_0663_),
    .X(_0238_));
 sky130_fd_sc_hd__buf_6 _3301_ (.A(_0662_),
    .X(_0823_));
 sky130_fd_sc_hd__mux2_1 _3302_ (.A0(_0742_),
    .A1(net66),
    .S(_0823_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _3303_ (.A0(_0745_),
    .A1(net4),
    .S(_0823_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _3304_ (.A0(_0747_),
    .A1(net5),
    .S(_0823_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _3305_ (.A0(_0749_),
    .A1(net6),
    .S(_0823_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _3306_ (.A0(_0751_),
    .A1(net7),
    .S(_0823_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _3307_ (.A0(_0753_),
    .A1(net8),
    .S(_0823_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _3308_ (.A0(_0755_),
    .A1(net9),
    .S(_0823_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _3309_ (.A0(_0757_),
    .A1(net10),
    .S(_0823_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _3310_ (.A0(_0759_),
    .A1(net11),
    .S(_0823_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _3311_ (.A0(_0761_),
    .A1(net12),
    .S(_0823_),
    .X(_0217_));
 sky130_fd_sc_hd__buf_6 _3312_ (.A(_0662_),
    .X(_0824_));
 sky130_fd_sc_hd__mux2_1 _3313_ (.A0(_0763_),
    .A1(net13),
    .S(_0824_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _3314_ (.A0(_0766_),
    .A1(net15),
    .S(_0824_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _3315_ (.A0(_0768_),
    .A1(net16),
    .S(_0824_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _3316_ (.A0(_0770_),
    .A1(net17),
    .S(_0824_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _3317_ (.A0(_0772_),
    .A1(net18),
    .S(_0824_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _3318_ (.A0(_0774_),
    .A1(net19),
    .S(_0824_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _3319_ (.A0(_0776_),
    .A1(net20),
    .S(_0824_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _3320_ (.A0(_0778_),
    .A1(net21),
    .S(_0824_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _3321_ (.A0(_0780_),
    .A1(net22),
    .S(_0824_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _3322_ (.A0(_0782_),
    .A1(net23),
    .S(_0824_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _3323_ (.A0(_0784_),
    .A1(net24),
    .S(_0662_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _3324_ (.A0(_0786_),
    .A1(net26),
    .S(_0662_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _3325_ (.A0(_0788_),
    .A1(net27),
    .S(_0662_),
    .X(_0232_));
 sky130_fd_sc_hd__inv_1 _3326_ (.A(_2539_),
    .Y(_2493_));
 sky130_fd_sc_hd__buf_8 _3327_ (.A(_0720_),
    .X(_2534_));
 sky130_fd_sc_hd__xor2_1 _3328_ (.A(_0609_),
    .B(_2523_),
    .X(_2540_));
 sky130_fd_sc_hd__inv_1 _3329_ (.A(_2544_),
    .Y(_2497_));
 sky130_fd_sc_hd__inv_1 _3330_ (.A(net73),
    .Y(_2546_));
 sky130_fd_sc_hd__inv_2 _3331_ (.A(net74),
    .Y(_2547_));
 sky130_fd_sc_hd__inv_1 _3332_ (.A(_2545_),
    .Y(_2567_));
 sky130_fd_sc_hd__nand3_1 _3333_ (.A(_0609_),
    .B(_0607_),
    .C(_2552_),
    .Y(_2511_));
 sky130_fd_sc_hd__xor2_1 _3334_ (.A(_0613_),
    .B(_2523_),
    .X(_2529_));
 sky130_fd_sc_hd__buf_4 _3335_ (.A(_0714_),
    .X(_0825_));
 sky130_fd_sc_hd__buf_6 _3336_ (.A(_0825_),
    .X(_2535_));
 sky130_fd_sc_hd__inv_2 _3337_ (.A(_2531_),
    .Y(_2494_));
 sky130_fd_sc_hd__a21o_1 _3338_ (.A1(_0609_),
    .A2(_2521_),
    .B1(_2541_),
    .X(_2554_));
 sky130_fd_sc_hd__buf_2 _3339_ (.A(\rd_ptr[2] ),
    .X(_0826_));
 sky130_fd_sc_hd__buf_6 _3340_ (.A(_0826_),
    .X(_0827_));
 sky130_fd_sc_hd__buf_4 _3341_ (.A(_0827_),
    .X(_0828_));
 sky130_fd_sc_hd__buf_6 _3342_ (.A(_0828_),
    .X(_0829_));
 sky130_fd_sc_hd__buf_8 _3343_ (.A(_0722_),
    .X(_0830_));
 sky130_fd_sc_hd__buf_8 _3344_ (.A(_0830_),
    .X(_0831_));
 sky130_fd_sc_hd__mux2i_1 _3345_ (.A0(\mem[5][0] ),
    .A1(\mem[7][0] ),
    .S(_0831_),
    .Y(_0832_));
 sky130_fd_sc_hd__buf_8 _3346_ (.A(_0722_),
    .X(_0833_));
 sky130_fd_sc_hd__mux2i_1 _3347_ (.A0(\mem[4][0] ),
    .A1(\mem[6][0] ),
    .S(_0833_),
    .Y(_0834_));
 sky130_fd_sc_hd__buf_6 _3348_ (.A(_0722_),
    .X(_0835_));
 sky130_fd_sc_hd__mux2i_2 _3349_ (.A0(\mem[13][0] ),
    .A1(\mem[15][0] ),
    .S(_0835_),
    .Y(_0836_));
 sky130_fd_sc_hd__buf_16 _3350_ (.A(_0830_),
    .X(_0837_));
 sky130_fd_sc_hd__mux2i_2 _3351_ (.A0(\mem[12][0] ),
    .A1(\mem[14][0] ),
    .S(_0837_),
    .Y(_0838_));
 sky130_fd_sc_hd__buf_6 _3352_ (.A(\rd_ptr[0] ),
    .X(_0839_));
 sky130_fd_sc_hd__inv_4 _3353_ (.A(_0839_),
    .Y(_0840_));
 sky130_fd_sc_hd__clkbuf_4 _3354_ (.A(\rd_ptr[3] ),
    .X(_0841_));
 sky130_fd_sc_hd__buf_6 _3355_ (.A(_0841_),
    .X(_0842_));
 sky130_fd_sc_hd__mux4_1 _3356_ (.A0(_0832_),
    .A1(_0834_),
    .A2(_0836_),
    .A3(_0838_),
    .S0(_0840_),
    .S1(_0842_),
    .X(_0843_));
 sky130_fd_sc_hd__buf_8 _3357_ (.A(_0841_),
    .X(_0844_));
 sky130_fd_sc_hd__buf_6 _3358_ (.A(_0840_),
    .X(_0845_));
 sky130_fd_sc_hd__buf_6 _3359_ (.A(_0833_),
    .X(_0846_));
 sky130_fd_sc_hd__mux2i_1 _3360_ (.A0(\mem[8][0] ),
    .A1(\mem[10][0] ),
    .S(_0846_),
    .Y(_0847_));
 sky130_fd_sc_hd__nand2_1 _3361_ (.A(_0845_),
    .B(_0847_),
    .Y(_0848_));
 sky130_fd_sc_hd__buf_6 _3362_ (.A(_0839_),
    .X(_0849_));
 sky130_fd_sc_hd__clkbuf_8 _3363_ (.A(_0849_),
    .X(_0850_));
 sky130_fd_sc_hd__buf_8 _3364_ (.A(_0837_),
    .X(_0851_));
 sky130_fd_sc_hd__mux2i_1 _3365_ (.A0(\mem[9][0] ),
    .A1(\mem[11][0] ),
    .S(_0851_),
    .Y(_0852_));
 sky130_fd_sc_hd__nand2_1 _3366_ (.A(_0850_),
    .B(_0852_),
    .Y(_0853_));
 sky130_fd_sc_hd__clkbuf_8 _3367_ (.A(_0839_),
    .X(_0854_));
 sky130_fd_sc_hd__buf_6 _3368_ (.A(_0835_),
    .X(_0855_));
 sky130_fd_sc_hd__mux2i_2 _3369_ (.A0(\mem[1][0] ),
    .A1(\mem[3][0] ),
    .S(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__mux2_1 _3370_ (.A0(\mem[0][0] ),
    .A1(\mem[2][0] ),
    .S(_0835_),
    .X(_0857_));
 sky130_fd_sc_hd__nor2_1 _3371_ (.A(_0849_),
    .B(_0857_),
    .Y(_0858_));
 sky130_fd_sc_hd__a211oi_1 _3372_ (.A1(_0854_),
    .A2(_0856_),
    .B1(_0858_),
    .C1(_0842_),
    .Y(_0859_));
 sky130_fd_sc_hd__buf_4 _3373_ (.A(_0826_),
    .X(_0860_));
 sky130_fd_sc_hd__buf_8 _3374_ (.A(_0860_),
    .X(_0861_));
 sky130_fd_sc_hd__a311oi_1 _3375_ (.A1(_0844_),
    .A2(_0848_),
    .A3(_0853_),
    .B1(_0859_),
    .C1(_0861_),
    .Y(_0862_));
 sky130_fd_sc_hd__a211oi_2 _3376_ (.A1(_0829_),
    .A2(_0843_),
    .B1(_0862_),
    .C1(_0825_),
    .Y(_0863_));
 sky130_fd_sc_hd__a21o_1 _3377_ (.A1(net78),
    .A2(_0825_),
    .B1(_0863_),
    .X(_0535_));
 sky130_fd_sc_hd__buf_6 _3378_ (.A(_0825_),
    .X(_0864_));
 sky130_fd_sc_hd__buf_6 _3379_ (.A(_0860_),
    .X(_0865_));
 sky130_fd_sc_hd__clkbuf_8 _3380_ (.A(_0865_),
    .X(_0866_));
 sky130_fd_sc_hd__buf_6 _3381_ (.A(_0844_),
    .X(_0867_));
 sky130_fd_sc_hd__buf_6 _3382_ (.A(_0854_),
    .X(_0868_));
 sky130_fd_sc_hd__buf_6 _3383_ (.A(_0833_),
    .X(_0869_));
 sky130_fd_sc_hd__mux2_1 _3384_ (.A0(\mem[4][10] ),
    .A1(\mem[6][10] ),
    .S(_0869_),
    .X(_0870_));
 sky130_fd_sc_hd__buf_6 _3385_ (.A(_0849_),
    .X(_0871_));
 sky130_fd_sc_hd__buf_8 _3386_ (.A(_0831_),
    .X(_0872_));
 sky130_fd_sc_hd__mux2i_1 _3387_ (.A0(\mem[5][10] ),
    .A1(\mem[7][10] ),
    .S(_0872_),
    .Y(_0873_));
 sky130_fd_sc_hd__nand2_1 _3388_ (.A(_0871_),
    .B(_0873_),
    .Y(_0874_));
 sky130_fd_sc_hd__o21ai_0 _3389_ (.A1(_0868_),
    .A2(_0870_),
    .B1(_0874_),
    .Y(_0875_));
 sky130_fd_sc_hd__buf_4 _3390_ (.A(_0854_),
    .X(_0876_));
 sky130_fd_sc_hd__mux2_1 _3391_ (.A0(\mem[12][10] ),
    .A1(\mem[14][10] ),
    .S(_0831_),
    .X(_0877_));
 sky130_fd_sc_hd__clkbuf_8 _3392_ (.A(_0854_),
    .X(_0878_));
 sky130_fd_sc_hd__buf_8 _3393_ (.A(_0855_),
    .X(_0879_));
 sky130_fd_sc_hd__mux2i_1 _3394_ (.A0(\mem[13][10] ),
    .A1(\mem[15][10] ),
    .S(_0879_),
    .Y(_0880_));
 sky130_fd_sc_hd__nand2_1 _3395_ (.A(_0878_),
    .B(_0880_),
    .Y(_0881_));
 sky130_fd_sc_hd__clkbuf_8 _3396_ (.A(_0842_),
    .X(_0882_));
 sky130_fd_sc_hd__o211ai_1 _3397_ (.A1(_0876_),
    .A2(_0877_),
    .B1(_0881_),
    .C1(_0882_),
    .Y(_0883_));
 sky130_fd_sc_hd__o21ai_0 _3398_ (.A1(_0867_),
    .A2(_0875_),
    .B1(_0883_),
    .Y(_0884_));
 sky130_fd_sc_hd__buf_8 _3399_ (.A(_0830_),
    .X(_0885_));
 sky130_fd_sc_hd__mux2i_2 _3400_ (.A0(\mem[0][10] ),
    .A1(\mem[2][10] ),
    .S(_0885_),
    .Y(_0886_));
 sky130_fd_sc_hd__buf_6 _3401_ (.A(_0835_),
    .X(_0887_));
 sky130_fd_sc_hd__mux2i_1 _3402_ (.A0(\mem[1][10] ),
    .A1(\mem[3][10] ),
    .S(_0887_),
    .Y(_0888_));
 sky130_fd_sc_hd__mux2i_1 _3403_ (.A0(\mem[8][10] ),
    .A1(\mem[10][10] ),
    .S(_0837_),
    .Y(_0889_));
 sky130_fd_sc_hd__buf_8 _3404_ (.A(_0835_),
    .X(_0890_));
 sky130_fd_sc_hd__mux2i_1 _3405_ (.A0(\mem[9][10] ),
    .A1(\mem[11][10] ),
    .S(_0890_),
    .Y(_0891_));
 sky130_fd_sc_hd__mux4_1 _3406_ (.A0(_0886_),
    .A1(_0888_),
    .A2(_0889_),
    .A3(_0891_),
    .S0(_0849_),
    .S1(_0844_),
    .X(_0892_));
 sky130_fd_sc_hd__nor2_1 _3407_ (.A(_0829_),
    .B(_0892_),
    .Y(_0893_));
 sky130_fd_sc_hd__a21oi_1 _3408_ (.A1(_0866_),
    .A2(_0884_),
    .B1(_0893_),
    .Y(_0894_));
 sky130_fd_sc_hd__nand2_1 _3409_ (.A(net79),
    .B(_2535_),
    .Y(_0895_));
 sky130_fd_sc_hd__o21ai_0 _3410_ (.A1(_0864_),
    .A2(_0894_),
    .B1(_0895_),
    .Y(_0536_));
 sky130_fd_sc_hd__inv_4 _3411_ (.A(_0826_),
    .Y(_0896_));
 sky130_fd_sc_hd__buf_4 _3412_ (.A(_0896_),
    .X(_0897_));
 sky130_fd_sc_hd__buf_4 _3413_ (.A(_0897_),
    .X(_0898_));
 sky130_fd_sc_hd__mux2_1 _3414_ (.A0(\mem[0][11] ),
    .A1(\mem[2][11] ),
    .S(_0722_),
    .X(_0899_));
 sky130_fd_sc_hd__mux2i_2 _3415_ (.A0(\mem[1][11] ),
    .A1(\mem[3][11] ),
    .S(_0872_),
    .Y(_0900_));
 sky130_fd_sc_hd__nand2_1 _3416_ (.A(_0871_),
    .B(_0900_),
    .Y(_0901_));
 sky130_fd_sc_hd__o21ai_0 _3417_ (.A1(_0868_),
    .A2(_0899_),
    .B1(_0901_),
    .Y(_0902_));
 sky130_fd_sc_hd__buf_4 _3418_ (.A(_0845_),
    .X(_0903_));
 sky130_fd_sc_hd__mux2i_1 _3419_ (.A0(\mem[8][11] ),
    .A1(\mem[10][11] ),
    .S(_0851_),
    .Y(_0904_));
 sky130_fd_sc_hd__nand2_1 _3420_ (.A(_0903_),
    .B(_0904_),
    .Y(_0905_));
 sky130_fd_sc_hd__buf_6 _3421_ (.A(_0854_),
    .X(_0906_));
 sky130_fd_sc_hd__buf_6 _3422_ (.A(_0855_),
    .X(_0907_));
 sky130_fd_sc_hd__mux2i_1 _3423_ (.A0(\mem[9][11] ),
    .A1(\mem[11][11] ),
    .S(_0907_),
    .Y(_0908_));
 sky130_fd_sc_hd__nand2_1 _3424_ (.A(_0906_),
    .B(_0908_),
    .Y(_0909_));
 sky130_fd_sc_hd__nand3_1 _3425_ (.A(_0882_),
    .B(_0905_),
    .C(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__o21ai_0 _3426_ (.A1(_0867_),
    .A2(_0902_),
    .B1(_0910_),
    .Y(_0911_));
 sky130_fd_sc_hd__mux2i_1 _3427_ (.A0(\mem[5][11] ),
    .A1(\mem[7][11] ),
    .S(_0890_),
    .Y(_0912_));
 sky130_fd_sc_hd__mux2i_2 _3428_ (.A0(\mem[4][11] ),
    .A1(\mem[6][11] ),
    .S(_0831_),
    .Y(_0913_));
 sky130_fd_sc_hd__buf_16 _3429_ (.A(_0830_),
    .X(_0914_));
 sky130_fd_sc_hd__mux2i_1 _3430_ (.A0(\mem[13][11] ),
    .A1(\mem[15][11] ),
    .S(_0914_),
    .Y(_0915_));
 sky130_fd_sc_hd__buf_8 _3431_ (.A(_0835_),
    .X(_0916_));
 sky130_fd_sc_hd__mux2i_1 _3432_ (.A0(\mem[12][11] ),
    .A1(\mem[14][11] ),
    .S(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__mux4_1 _3433_ (.A0(_0912_),
    .A1(_0913_),
    .A2(_0915_),
    .A3(_0917_),
    .S0(_0845_),
    .S1(_0844_),
    .X(_0918_));
 sky130_fd_sc_hd__nor2_1 _3434_ (.A(_0898_),
    .B(_0918_),
    .Y(_0919_));
 sky130_fd_sc_hd__a21oi_1 _3435_ (.A1(_0898_),
    .A2(_0911_),
    .B1(_0919_),
    .Y(_0920_));
 sky130_fd_sc_hd__nand2_1 _3436_ (.A(net80),
    .B(_2535_),
    .Y(_0921_));
 sky130_fd_sc_hd__o21ai_0 _3437_ (.A1(_0864_),
    .A2(_0920_),
    .B1(_0921_),
    .Y(_0537_));
 sky130_fd_sc_hd__mux2_1 _3438_ (.A0(\mem[4][12] ),
    .A1(\mem[6][12] ),
    .S(_0869_),
    .X(_0922_));
 sky130_fd_sc_hd__mux2i_1 _3439_ (.A0(\mem[5][12] ),
    .A1(\mem[7][12] ),
    .S(_0872_),
    .Y(_0923_));
 sky130_fd_sc_hd__nand2_1 _3440_ (.A(_0871_),
    .B(_0923_),
    .Y(_0924_));
 sky130_fd_sc_hd__o21ai_0 _3441_ (.A1(_0868_),
    .A2(_0922_),
    .B1(_0924_),
    .Y(_0925_));
 sky130_fd_sc_hd__buf_6 _3442_ (.A(_0722_),
    .X(_0926_));
 sky130_fd_sc_hd__mux2_1 _3443_ (.A0(\mem[12][12] ),
    .A1(\mem[14][12] ),
    .S(_0926_),
    .X(_0927_));
 sky130_fd_sc_hd__mux2i_1 _3444_ (.A0(\mem[13][12] ),
    .A1(\mem[15][12] ),
    .S(_0879_),
    .Y(_0928_));
 sky130_fd_sc_hd__nand2_1 _3445_ (.A(_0878_),
    .B(_0928_),
    .Y(_0929_));
 sky130_fd_sc_hd__clkbuf_8 _3446_ (.A(_0842_),
    .X(_0930_));
 sky130_fd_sc_hd__o211ai_1 _3447_ (.A1(_0876_),
    .A2(_0927_),
    .B1(_0929_),
    .C1(_0930_),
    .Y(_0931_));
 sky130_fd_sc_hd__o21ai_0 _3448_ (.A1(_0867_),
    .A2(_0925_),
    .B1(_0931_),
    .Y(_0932_));
 sky130_fd_sc_hd__mux2i_2 _3449_ (.A0(\mem[0][12] ),
    .A1(\mem[2][12] ),
    .S(_0885_),
    .Y(_0933_));
 sky130_fd_sc_hd__mux2i_1 _3450_ (.A0(\mem[1][12] ),
    .A1(\mem[3][12] ),
    .S(_0887_),
    .Y(_0934_));
 sky130_fd_sc_hd__mux2i_1 _3451_ (.A0(\mem[8][12] ),
    .A1(\mem[10][12] ),
    .S(_0837_),
    .Y(_0935_));
 sky130_fd_sc_hd__mux2i_1 _3452_ (.A0(\mem[9][12] ),
    .A1(\mem[11][12] ),
    .S(_0890_),
    .Y(_0936_));
 sky130_fd_sc_hd__mux4_1 _3453_ (.A0(_0933_),
    .A1(_0934_),
    .A2(_0935_),
    .A3(_0936_),
    .S0(_0849_),
    .S1(_0844_),
    .X(_0937_));
 sky130_fd_sc_hd__nor2_1 _3454_ (.A(_0829_),
    .B(_0937_),
    .Y(_0938_));
 sky130_fd_sc_hd__a21oi_1 _3455_ (.A1(_0866_),
    .A2(_0932_),
    .B1(_0938_),
    .Y(_0939_));
 sky130_fd_sc_hd__nand2_1 _3456_ (.A(net81),
    .B(_2535_),
    .Y(_0940_));
 sky130_fd_sc_hd__o21ai_0 _3457_ (.A1(_0864_),
    .A2(_0939_),
    .B1(_0940_),
    .Y(_0538_));
 sky130_fd_sc_hd__mux2_1 _3458_ (.A0(\mem[4][13] ),
    .A1(\mem[6][13] ),
    .S(_0869_),
    .X(_0941_));
 sky130_fd_sc_hd__mux2i_1 _3459_ (.A0(\mem[5][13] ),
    .A1(\mem[7][13] ),
    .S(_0872_),
    .Y(_0942_));
 sky130_fd_sc_hd__nand2_1 _3460_ (.A(_0871_),
    .B(_0942_),
    .Y(_0943_));
 sky130_fd_sc_hd__o21ai_0 _3461_ (.A1(_0868_),
    .A2(_0941_),
    .B1(_0943_),
    .Y(_0944_));
 sky130_fd_sc_hd__mux2_1 _3462_ (.A0(\mem[12][13] ),
    .A1(\mem[14][13] ),
    .S(_0926_),
    .X(_0945_));
 sky130_fd_sc_hd__mux2i_1 _3463_ (.A0(\mem[13][13] ),
    .A1(\mem[15][13] ),
    .S(_0879_),
    .Y(_0946_));
 sky130_fd_sc_hd__nand2_1 _3464_ (.A(_0878_),
    .B(_0946_),
    .Y(_0947_));
 sky130_fd_sc_hd__o211ai_1 _3465_ (.A1(_0876_),
    .A2(_0945_),
    .B1(_0947_),
    .C1(_0930_),
    .Y(_0948_));
 sky130_fd_sc_hd__o21ai_0 _3466_ (.A1(_0867_),
    .A2(_0944_),
    .B1(_0948_),
    .Y(_0949_));
 sky130_fd_sc_hd__mux2i_2 _3467_ (.A0(\mem[0][13] ),
    .A1(\mem[2][13] ),
    .S(_0885_),
    .Y(_0950_));
 sky130_fd_sc_hd__mux2i_1 _3468_ (.A0(\mem[1][13] ),
    .A1(\mem[3][13] ),
    .S(_0887_),
    .Y(_0951_));
 sky130_fd_sc_hd__clkbuf_16 _3469_ (.A(_0830_),
    .X(_0952_));
 sky130_fd_sc_hd__mux2i_1 _3470_ (.A0(\mem[8][13] ),
    .A1(\mem[10][13] ),
    .S(_0952_),
    .Y(_0953_));
 sky130_fd_sc_hd__clkbuf_16 _3471_ (.A(_0830_),
    .X(_0954_));
 sky130_fd_sc_hd__mux2i_1 _3472_ (.A0(\mem[9][13] ),
    .A1(\mem[11][13] ),
    .S(_0954_),
    .Y(_0955_));
 sky130_fd_sc_hd__mux4_1 _3473_ (.A0(_0950_),
    .A1(_0951_),
    .A2(_0953_),
    .A3(_0955_),
    .S0(_0849_),
    .S1(_0844_),
    .X(_0956_));
 sky130_fd_sc_hd__nor2_1 _3474_ (.A(_0829_),
    .B(_0956_),
    .Y(_0957_));
 sky130_fd_sc_hd__a21oi_1 _3475_ (.A1(_0866_),
    .A2(_0949_),
    .B1(_0957_),
    .Y(_0958_));
 sky130_fd_sc_hd__nand2_1 _3476_ (.A(net82),
    .B(_2535_),
    .Y(_0959_));
 sky130_fd_sc_hd__o21ai_0 _3477_ (.A1(_0864_),
    .A2(_0958_),
    .B1(_0959_),
    .Y(_0539_));
 sky130_fd_sc_hd__mux2_1 _3478_ (.A0(\mem[4][14] ),
    .A1(\mem[6][14] ),
    .S(_0869_),
    .X(_0960_));
 sky130_fd_sc_hd__mux2i_1 _3479_ (.A0(\mem[5][14] ),
    .A1(\mem[7][14] ),
    .S(_0872_),
    .Y(_0961_));
 sky130_fd_sc_hd__nand2_1 _3480_ (.A(_0871_),
    .B(_0961_),
    .Y(_0962_));
 sky130_fd_sc_hd__o21ai_0 _3481_ (.A1(_0868_),
    .A2(_0960_),
    .B1(_0962_),
    .Y(_0963_));
 sky130_fd_sc_hd__mux2_1 _3482_ (.A0(\mem[12][14] ),
    .A1(\mem[14][14] ),
    .S(_0926_),
    .X(_0964_));
 sky130_fd_sc_hd__mux2i_1 _3483_ (.A0(\mem[13][14] ),
    .A1(\mem[15][14] ),
    .S(_0879_),
    .Y(_0965_));
 sky130_fd_sc_hd__nand2_1 _3484_ (.A(_0878_),
    .B(_0965_),
    .Y(_0966_));
 sky130_fd_sc_hd__o211ai_1 _3485_ (.A1(_0876_),
    .A2(_0964_),
    .B1(_0966_),
    .C1(_0930_),
    .Y(_0967_));
 sky130_fd_sc_hd__o21ai_0 _3486_ (.A1(_0867_),
    .A2(_0963_),
    .B1(_0967_),
    .Y(_0968_));
 sky130_fd_sc_hd__mux2i_2 _3487_ (.A0(\mem[0][14] ),
    .A1(\mem[2][14] ),
    .S(_0885_),
    .Y(_0969_));
 sky130_fd_sc_hd__mux2i_1 _3488_ (.A0(\mem[1][14] ),
    .A1(\mem[3][14] ),
    .S(_0887_),
    .Y(_0970_));
 sky130_fd_sc_hd__mux2i_2 _3489_ (.A0(\mem[8][14] ),
    .A1(\mem[10][14] ),
    .S(_0952_),
    .Y(_0971_));
 sky130_fd_sc_hd__mux2i_2 _3490_ (.A0(\mem[9][14] ),
    .A1(\mem[11][14] ),
    .S(_0954_),
    .Y(_0972_));
 sky130_fd_sc_hd__mux4_1 _3491_ (.A0(_0969_),
    .A1(_0970_),
    .A2(_0971_),
    .A3(_0972_),
    .S0(_0849_),
    .S1(_0844_),
    .X(_0973_));
 sky130_fd_sc_hd__nor2_1 _3492_ (.A(_0829_),
    .B(_0973_),
    .Y(_0974_));
 sky130_fd_sc_hd__a21oi_1 _3493_ (.A1(_0866_),
    .A2(_0968_),
    .B1(_0974_),
    .Y(_0975_));
 sky130_fd_sc_hd__nand2_1 _3494_ (.A(net83),
    .B(_2535_),
    .Y(_0976_));
 sky130_fd_sc_hd__o21ai_0 _3495_ (.A1(_0864_),
    .A2(_0975_),
    .B1(_0976_),
    .Y(_0540_));
 sky130_fd_sc_hd__mux2_1 _3496_ (.A0(\mem[0][15] ),
    .A1(\mem[2][15] ),
    .S(_0833_),
    .X(_0977_));
 sky130_fd_sc_hd__clkbuf_8 _3497_ (.A(_0849_),
    .X(_0978_));
 sky130_fd_sc_hd__mux2i_1 _3498_ (.A0(\mem[1][15] ),
    .A1(\mem[3][15] ),
    .S(_0846_),
    .Y(_0979_));
 sky130_fd_sc_hd__nand2_1 _3499_ (.A(_0978_),
    .B(_0979_),
    .Y(_0980_));
 sky130_fd_sc_hd__o21ai_1 _3500_ (.A1(_0868_),
    .A2(_0977_),
    .B1(_0980_),
    .Y(_0981_));
 sky130_fd_sc_hd__mux2i_1 _3501_ (.A0(\mem[8][15] ),
    .A1(\mem[10][15] ),
    .S(_0907_),
    .Y(_0982_));
 sky130_fd_sc_hd__nand2_1 _3502_ (.A(_0903_),
    .B(_0982_),
    .Y(_0983_));
 sky130_fd_sc_hd__mux2i_1 _3503_ (.A0(\mem[9][15] ),
    .A1(\mem[11][15] ),
    .S(_0907_),
    .Y(_0984_));
 sky130_fd_sc_hd__nand2_1 _3504_ (.A(_0876_),
    .B(_0984_),
    .Y(_0985_));
 sky130_fd_sc_hd__nand3_1 _3505_ (.A(_0882_),
    .B(_0983_),
    .C(_0985_),
    .Y(_0986_));
 sky130_fd_sc_hd__o21ai_0 _3506_ (.A1(_0867_),
    .A2(_0981_),
    .B1(_0986_),
    .Y(_0987_));
 sky130_fd_sc_hd__mux2i_1 _3507_ (.A0(\mem[5][15] ),
    .A1(\mem[7][15] ),
    .S(_0890_),
    .Y(_0988_));
 sky130_fd_sc_hd__mux2i_1 _3508_ (.A0(\mem[4][15] ),
    .A1(\mem[6][15] ),
    .S(_0914_),
    .Y(_0989_));
 sky130_fd_sc_hd__mux2i_1 _3509_ (.A0(\mem[13][15] ),
    .A1(\mem[15][15] ),
    .S(_0952_),
    .Y(_0990_));
 sky130_fd_sc_hd__mux2i_1 _3510_ (.A0(\mem[12][15] ),
    .A1(\mem[14][15] ),
    .S(_0916_),
    .Y(_0991_));
 sky130_fd_sc_hd__buf_8 _3511_ (.A(_0841_),
    .X(_0992_));
 sky130_fd_sc_hd__mux4_1 _3512_ (.A0(_0988_),
    .A1(_0989_),
    .A2(_0990_),
    .A3(_0991_),
    .S0(_0845_),
    .S1(_0992_),
    .X(_0993_));
 sky130_fd_sc_hd__nor2_1 _3513_ (.A(_0898_),
    .B(_0993_),
    .Y(_0994_));
 sky130_fd_sc_hd__a21oi_1 _3514_ (.A1(_0898_),
    .A2(_0987_),
    .B1(_0994_),
    .Y(_0995_));
 sky130_fd_sc_hd__nand2_1 _3515_ (.A(net84),
    .B(_2535_),
    .Y(_0996_));
 sky130_fd_sc_hd__o21ai_0 _3516_ (.A1(_0864_),
    .A2(_0995_),
    .B1(_0996_),
    .Y(_0541_));
 sky130_fd_sc_hd__buf_6 _3517_ (.A(_0839_),
    .X(_0997_));
 sky130_fd_sc_hd__mux2_1 _3518_ (.A0(\mem[4][16] ),
    .A1(\mem[6][16] ),
    .S(_0869_),
    .X(_0998_));
 sky130_fd_sc_hd__mux2i_1 _3519_ (.A0(\mem[5][16] ),
    .A1(\mem[7][16] ),
    .S(_0872_),
    .Y(_0999_));
 sky130_fd_sc_hd__nand2_1 _3520_ (.A(_0978_),
    .B(_0999_),
    .Y(_1000_));
 sky130_fd_sc_hd__o21ai_0 _3521_ (.A1(_0997_),
    .A2(_0998_),
    .B1(_1000_),
    .Y(_1001_));
 sky130_fd_sc_hd__buf_4 _3522_ (.A(_0854_),
    .X(_1002_));
 sky130_fd_sc_hd__mux2_1 _3523_ (.A0(\mem[12][16] ),
    .A1(\mem[14][16] ),
    .S(_0926_),
    .X(_1003_));
 sky130_fd_sc_hd__mux2i_1 _3524_ (.A0(\mem[13][16] ),
    .A1(\mem[15][16] ),
    .S(_0879_),
    .Y(_1004_));
 sky130_fd_sc_hd__nand2_1 _3525_ (.A(_0878_),
    .B(_1004_),
    .Y(_1005_));
 sky130_fd_sc_hd__o211ai_1 _3526_ (.A1(_1002_),
    .A2(_1003_),
    .B1(_1005_),
    .C1(_0930_),
    .Y(_1006_));
 sky130_fd_sc_hd__o21ai_0 _3527_ (.A1(_0867_),
    .A2(_1001_),
    .B1(_1006_),
    .Y(_1007_));
 sky130_fd_sc_hd__mux2i_1 _3528_ (.A0(\mem[0][16] ),
    .A1(\mem[2][16] ),
    .S(_0885_),
    .Y(_1008_));
 sky130_fd_sc_hd__mux2i_1 _3529_ (.A0(\mem[1][16] ),
    .A1(\mem[3][16] ),
    .S(_0887_),
    .Y(_1009_));
 sky130_fd_sc_hd__mux2i_2 _3530_ (.A0(\mem[8][16] ),
    .A1(\mem[10][16] ),
    .S(_0952_),
    .Y(_1010_));
 sky130_fd_sc_hd__mux2i_4 _3531_ (.A0(\mem[9][16] ),
    .A1(\mem[11][16] ),
    .S(_0954_),
    .Y(_1011_));
 sky130_fd_sc_hd__buf_6 _3532_ (.A(_0839_),
    .X(_1012_));
 sky130_fd_sc_hd__mux4_1 _3533_ (.A0(_1008_),
    .A1(_1009_),
    .A2(_1010_),
    .A3(_1011_),
    .S0(_1012_),
    .S1(_0992_),
    .X(_1013_));
 sky130_fd_sc_hd__nor2_1 _3534_ (.A(_0829_),
    .B(_1013_),
    .Y(_1014_));
 sky130_fd_sc_hd__a21oi_1 _3535_ (.A1(_0866_),
    .A2(_1007_),
    .B1(_1014_),
    .Y(_1015_));
 sky130_fd_sc_hd__nand2_1 _3536_ (.A(net85),
    .B(_2535_),
    .Y(_1016_));
 sky130_fd_sc_hd__o21ai_0 _3537_ (.A1(_0864_),
    .A2(_1015_),
    .B1(_1016_),
    .Y(_0542_));
 sky130_fd_sc_hd__mux2_1 _3538_ (.A0(\mem[4][17] ),
    .A1(\mem[6][17] ),
    .S(_0869_),
    .X(_1017_));
 sky130_fd_sc_hd__mux2i_1 _3539_ (.A0(\mem[5][17] ),
    .A1(\mem[7][17] ),
    .S(_0872_),
    .Y(_1018_));
 sky130_fd_sc_hd__nand2_1 _3540_ (.A(_0978_),
    .B(_1018_),
    .Y(_1019_));
 sky130_fd_sc_hd__o21ai_0 _3541_ (.A1(_0997_),
    .A2(_1017_),
    .B1(_1019_),
    .Y(_1020_));
 sky130_fd_sc_hd__mux2_1 _3542_ (.A0(\mem[12][17] ),
    .A1(\mem[14][17] ),
    .S(_0926_),
    .X(_1021_));
 sky130_fd_sc_hd__mux2i_1 _3543_ (.A0(\mem[13][17] ),
    .A1(\mem[15][17] ),
    .S(_0879_),
    .Y(_1022_));
 sky130_fd_sc_hd__nand2_1 _3544_ (.A(_0878_),
    .B(_1022_),
    .Y(_1023_));
 sky130_fd_sc_hd__o211ai_1 _3545_ (.A1(_1002_),
    .A2(_1021_),
    .B1(_1023_),
    .C1(_0930_),
    .Y(_1024_));
 sky130_fd_sc_hd__o21ai_0 _3546_ (.A1(_0867_),
    .A2(_1020_),
    .B1(_1024_),
    .Y(_1025_));
 sky130_fd_sc_hd__buf_4 _3547_ (.A(_0828_),
    .X(_1026_));
 sky130_fd_sc_hd__mux2i_2 _3548_ (.A0(\mem[0][17] ),
    .A1(\mem[2][17] ),
    .S(_0885_),
    .Y(_1027_));
 sky130_fd_sc_hd__mux2i_1 _3549_ (.A0(\mem[1][17] ),
    .A1(\mem[3][17] ),
    .S(_0887_),
    .Y(_1028_));
 sky130_fd_sc_hd__mux2i_2 _3550_ (.A0(\mem[8][17] ),
    .A1(\mem[10][17] ),
    .S(_0952_),
    .Y(_1029_));
 sky130_fd_sc_hd__mux2i_2 _3551_ (.A0(\mem[9][17] ),
    .A1(\mem[11][17] ),
    .S(_0954_),
    .Y(_1030_));
 sky130_fd_sc_hd__mux4_1 _3552_ (.A0(_1027_),
    .A1(_1028_),
    .A2(_1029_),
    .A3(_1030_),
    .S0(_1012_),
    .S1(_0992_),
    .X(_1031_));
 sky130_fd_sc_hd__nor2_1 _3553_ (.A(_1026_),
    .B(_1031_),
    .Y(_1032_));
 sky130_fd_sc_hd__a21oi_1 _3554_ (.A1(_0866_),
    .A2(_1025_),
    .B1(_1032_),
    .Y(_1033_));
 sky130_fd_sc_hd__nand2_1 _3555_ (.A(net86),
    .B(_2535_),
    .Y(_1034_));
 sky130_fd_sc_hd__o21ai_0 _3556_ (.A1(_0864_),
    .A2(_1033_),
    .B1(_1034_),
    .Y(_0543_));
 sky130_fd_sc_hd__buf_6 _3557_ (.A(net221),
    .X(_1035_));
 sky130_fd_sc_hd__mux2_1 _3558_ (.A0(\mem[4][18] ),
    .A1(\mem[6][18] ),
    .S(_0869_),
    .X(_1036_));
 sky130_fd_sc_hd__mux2i_1 _3559_ (.A0(\mem[5][18] ),
    .A1(\mem[7][18] ),
    .S(_0872_),
    .Y(_1037_));
 sky130_fd_sc_hd__nand2_1 _3560_ (.A(_0978_),
    .B(_1037_),
    .Y(_1038_));
 sky130_fd_sc_hd__o21ai_0 _3561_ (.A1(_0997_),
    .A2(_1036_),
    .B1(_1038_),
    .Y(_1039_));
 sky130_fd_sc_hd__mux2_1 _3562_ (.A0(\mem[12][18] ),
    .A1(\mem[14][18] ),
    .S(_0926_),
    .X(_1040_));
 sky130_fd_sc_hd__buf_8 _3563_ (.A(_0855_),
    .X(_1041_));
 sky130_fd_sc_hd__mux2i_1 _3564_ (.A0(\mem[13][18] ),
    .A1(\mem[15][18] ),
    .S(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__nand2_1 _3565_ (.A(_0878_),
    .B(_1042_),
    .Y(_1043_));
 sky130_fd_sc_hd__o211ai_1 _3566_ (.A1(_1002_),
    .A2(_1040_),
    .B1(_1043_),
    .C1(_0930_),
    .Y(_1044_));
 sky130_fd_sc_hd__o21ai_0 _3567_ (.A1(_0867_),
    .A2(_1039_),
    .B1(_1044_),
    .Y(_1045_));
 sky130_fd_sc_hd__mux2i_2 _3568_ (.A0(\mem[0][18] ),
    .A1(\mem[2][18] ),
    .S(_0885_),
    .Y(_1046_));
 sky130_fd_sc_hd__mux2i_1 _3569_ (.A0(\mem[1][18] ),
    .A1(\mem[3][18] ),
    .S(_0887_),
    .Y(_1047_));
 sky130_fd_sc_hd__mux2i_1 _3570_ (.A0(\mem[8][18] ),
    .A1(\mem[10][18] ),
    .S(_0952_),
    .Y(_1048_));
 sky130_fd_sc_hd__mux2i_2 _3571_ (.A0(\mem[9][18] ),
    .A1(\mem[11][18] ),
    .S(_0954_),
    .Y(_1049_));
 sky130_fd_sc_hd__mux4_1 _3572_ (.A0(_1046_),
    .A1(_1047_),
    .A2(_1048_),
    .A3(_1049_),
    .S0(_1012_),
    .S1(_0992_),
    .X(_1050_));
 sky130_fd_sc_hd__nor2_1 _3573_ (.A(_1026_),
    .B(_1050_),
    .Y(_1051_));
 sky130_fd_sc_hd__a21oi_1 _3574_ (.A1(_0866_),
    .A2(_1045_),
    .B1(_1051_),
    .Y(_1052_));
 sky130_fd_sc_hd__nand2_1 _3575_ (.A(net87),
    .B(_2535_),
    .Y(_1053_));
 sky130_fd_sc_hd__o21ai_0 _3576_ (.A1(_1035_),
    .A2(_1052_),
    .B1(_1053_),
    .Y(_0544_));
 sky130_fd_sc_hd__buf_6 _3577_ (.A(_0841_),
    .X(_1054_));
 sky130_fd_sc_hd__mux2_1 _3578_ (.A0(\mem[4][19] ),
    .A1(\mem[6][19] ),
    .S(_0869_),
    .X(_1055_));
 sky130_fd_sc_hd__mux2i_1 _3579_ (.A0(\mem[5][19] ),
    .A1(\mem[7][19] ),
    .S(_0872_),
    .Y(_1056_));
 sky130_fd_sc_hd__nand2_1 _3580_ (.A(_0978_),
    .B(_1056_),
    .Y(_1057_));
 sky130_fd_sc_hd__o21ai_0 _3581_ (.A1(_0997_),
    .A2(_1055_),
    .B1(_1057_),
    .Y(_1058_));
 sky130_fd_sc_hd__mux2_1 _3582_ (.A0(\mem[12][19] ),
    .A1(\mem[14][19] ),
    .S(_0926_),
    .X(_1059_));
 sky130_fd_sc_hd__mux2i_1 _3583_ (.A0(\mem[13][19] ),
    .A1(\mem[15][19] ),
    .S(_1041_),
    .Y(_1060_));
 sky130_fd_sc_hd__nand2_1 _3584_ (.A(_0878_),
    .B(_1060_),
    .Y(_1061_));
 sky130_fd_sc_hd__o211ai_1 _3585_ (.A1(_1002_),
    .A2(_1059_),
    .B1(_1061_),
    .C1(_0930_),
    .Y(_1062_));
 sky130_fd_sc_hd__o21ai_0 _3586_ (.A1(_1054_),
    .A2(_1058_),
    .B1(_1062_),
    .Y(_1063_));
 sky130_fd_sc_hd__mux2i_2 _3587_ (.A0(\mem[0][19] ),
    .A1(\mem[2][19] ),
    .S(_0885_),
    .Y(_1064_));
 sky130_fd_sc_hd__mux2i_1 _3588_ (.A0(\mem[1][19] ),
    .A1(\mem[3][19] ),
    .S(_0887_),
    .Y(_1065_));
 sky130_fd_sc_hd__mux2i_1 _3589_ (.A0(\mem[8][19] ),
    .A1(\mem[10][19] ),
    .S(_0952_),
    .Y(_1066_));
 sky130_fd_sc_hd__mux2i_2 _3590_ (.A0(\mem[9][19] ),
    .A1(\mem[11][19] ),
    .S(_0954_),
    .Y(_1067_));
 sky130_fd_sc_hd__mux4_1 _3591_ (.A0(_1064_),
    .A1(_1065_),
    .A2(_1066_),
    .A3(_1067_),
    .S0(_1012_),
    .S1(_0992_),
    .X(_1068_));
 sky130_fd_sc_hd__nor2_1 _3592_ (.A(_1026_),
    .B(_1068_),
    .Y(_1069_));
 sky130_fd_sc_hd__a21oi_1 _3593_ (.A1(_0866_),
    .A2(_1063_),
    .B1(_1069_),
    .Y(_1070_));
 sky130_fd_sc_hd__buf_8 _3594_ (.A(_0825_),
    .X(_1071_));
 sky130_fd_sc_hd__nand2_1 _3595_ (.A(net88),
    .B(_1071_),
    .Y(_1072_));
 sky130_fd_sc_hd__o21ai_0 _3596_ (.A1(_1035_),
    .A2(_1070_),
    .B1(_1072_),
    .Y(_0545_));
 sky130_fd_sc_hd__mux2_1 _3597_ (.A0(\mem[0][1] ),
    .A1(\mem[2][1] ),
    .S(_0833_),
    .X(_1073_));
 sky130_fd_sc_hd__mux2i_1 _3598_ (.A0(\mem[1][1] ),
    .A1(\mem[3][1] ),
    .S(_0846_),
    .Y(_1074_));
 sky130_fd_sc_hd__nand2_1 _3599_ (.A(_0978_),
    .B(_1074_),
    .Y(_1075_));
 sky130_fd_sc_hd__o21ai_0 _3600_ (.A1(_0997_),
    .A2(_1073_),
    .B1(_1075_),
    .Y(_1076_));
 sky130_fd_sc_hd__mux2i_1 _3601_ (.A0(\mem[8][1] ),
    .A1(\mem[10][1] ),
    .S(_0907_),
    .Y(_1077_));
 sky130_fd_sc_hd__nand2_1 _3602_ (.A(_0903_),
    .B(_1077_),
    .Y(_1078_));
 sky130_fd_sc_hd__mux2i_1 _3603_ (.A0(\mem[9][1] ),
    .A1(\mem[11][1] ),
    .S(_0907_),
    .Y(_1079_));
 sky130_fd_sc_hd__nand2_1 _3604_ (.A(_0876_),
    .B(_1079_),
    .Y(_1080_));
 sky130_fd_sc_hd__nand3_1 _3605_ (.A(_0882_),
    .B(_1078_),
    .C(_1080_),
    .Y(_1081_));
 sky130_fd_sc_hd__o21ai_0 _3606_ (.A1(_1054_),
    .A2(_1076_),
    .B1(_1081_),
    .Y(_1082_));
 sky130_fd_sc_hd__mux2i_1 _3607_ (.A0(\mem[5][1] ),
    .A1(\mem[7][1] ),
    .S(_0890_),
    .Y(_1083_));
 sky130_fd_sc_hd__mux2i_2 _3608_ (.A0(\mem[4][1] ),
    .A1(\mem[6][1] ),
    .S(_0831_),
    .Y(_1084_));
 sky130_fd_sc_hd__mux2i_1 _3609_ (.A0(\mem[13][1] ),
    .A1(\mem[15][1] ),
    .S(_0952_),
    .Y(_1085_));
 sky130_fd_sc_hd__mux2i_1 _3610_ (.A0(\mem[12][1] ),
    .A1(\mem[14][1] ),
    .S(_0916_),
    .Y(_1086_));
 sky130_fd_sc_hd__mux4_1 _3611_ (.A0(_1083_),
    .A1(_1084_),
    .A2(_1085_),
    .A3(_1086_),
    .S0(_0845_),
    .S1(_0992_),
    .X(_1087_));
 sky130_fd_sc_hd__nor2_1 _3612_ (.A(_0897_),
    .B(_1087_),
    .Y(_1088_));
 sky130_fd_sc_hd__a21oi_2 _3613_ (.A1(_0898_),
    .A2(_1082_),
    .B1(_1088_),
    .Y(_1089_));
 sky130_fd_sc_hd__nand2_1 _3614_ (.A(net89),
    .B(_1071_),
    .Y(_1090_));
 sky130_fd_sc_hd__o21ai_0 _3615_ (.A1(_1035_),
    .A2(_1089_),
    .B1(_1090_),
    .Y(_0546_));
 sky130_fd_sc_hd__buf_4 _3616_ (.A(_0835_),
    .X(_1091_));
 sky130_fd_sc_hd__mux2_1 _3617_ (.A0(\mem[4][20] ),
    .A1(\mem[6][20] ),
    .S(_1091_),
    .X(_1092_));
 sky130_fd_sc_hd__mux2i_1 _3618_ (.A0(\mem[5][20] ),
    .A1(\mem[7][20] ),
    .S(_0872_),
    .Y(_1093_));
 sky130_fd_sc_hd__nand2_1 _3619_ (.A(_0978_),
    .B(_1093_),
    .Y(_1094_));
 sky130_fd_sc_hd__o21ai_0 _3620_ (.A1(_0997_),
    .A2(_1092_),
    .B1(_1094_),
    .Y(_1095_));
 sky130_fd_sc_hd__mux2_1 _3621_ (.A0(\mem[12][20] ),
    .A1(\mem[14][20] ),
    .S(_0926_),
    .X(_1096_));
 sky130_fd_sc_hd__mux2i_1 _3622_ (.A0(\mem[13][20] ),
    .A1(\mem[15][20] ),
    .S(_1041_),
    .Y(_1097_));
 sky130_fd_sc_hd__nand2_1 _3623_ (.A(_0878_),
    .B(_1097_),
    .Y(_1098_));
 sky130_fd_sc_hd__o211ai_1 _3624_ (.A1(_1002_),
    .A2(_1096_),
    .B1(_1098_),
    .C1(_0930_),
    .Y(_1099_));
 sky130_fd_sc_hd__o21ai_0 _3625_ (.A1(_1054_),
    .A2(_1095_),
    .B1(_1099_),
    .Y(_1100_));
 sky130_fd_sc_hd__buf_8 _3626_ (.A(_0830_),
    .X(_1101_));
 sky130_fd_sc_hd__mux2i_2 _3627_ (.A0(\mem[0][20] ),
    .A1(\mem[2][20] ),
    .S(_1101_),
    .Y(_1102_));
 sky130_fd_sc_hd__mux2i_2 _3628_ (.A0(\mem[1][20] ),
    .A1(\mem[3][20] ),
    .S(_0887_),
    .Y(_1103_));
 sky130_fd_sc_hd__mux2i_1 _3629_ (.A0(\mem[8][20] ),
    .A1(\mem[10][20] ),
    .S(_0952_),
    .Y(_1104_));
 sky130_fd_sc_hd__mux2i_2 _3630_ (.A0(\mem[9][20] ),
    .A1(\mem[11][20] ),
    .S(_0954_),
    .Y(_1105_));
 sky130_fd_sc_hd__mux4_1 _3631_ (.A0(_1102_),
    .A1(_1103_),
    .A2(_1104_),
    .A3(_1105_),
    .S0(_1012_),
    .S1(_0992_),
    .X(_1106_));
 sky130_fd_sc_hd__nor2_1 _3632_ (.A(_1026_),
    .B(_1106_),
    .Y(_1107_));
 sky130_fd_sc_hd__a21oi_1 _3633_ (.A1(_0866_),
    .A2(_1100_),
    .B1(_1107_),
    .Y(_1108_));
 sky130_fd_sc_hd__nand2_1 _3634_ (.A(net90),
    .B(_1071_),
    .Y(_1109_));
 sky130_fd_sc_hd__o21ai_0 _3635_ (.A1(_1035_),
    .A2(_1108_),
    .B1(_1109_),
    .Y(_0547_));
 sky130_fd_sc_hd__mux2_1 _3636_ (.A0(\mem[4][21] ),
    .A1(\mem[6][21] ),
    .S(_1091_),
    .X(_1110_));
 sky130_fd_sc_hd__buf_6 _3637_ (.A(_0831_),
    .X(_1111_));
 sky130_fd_sc_hd__mux2i_1 _3638_ (.A0(\mem[5][21] ),
    .A1(\mem[7][21] ),
    .S(_1111_),
    .Y(_1112_));
 sky130_fd_sc_hd__nand2_1 _3639_ (.A(_0978_),
    .B(_1112_),
    .Y(_1113_));
 sky130_fd_sc_hd__o21ai_0 _3640_ (.A1(_0997_),
    .A2(_1110_),
    .B1(_1113_),
    .Y(_1114_));
 sky130_fd_sc_hd__mux2_1 _3641_ (.A0(\mem[12][21] ),
    .A1(\mem[14][21] ),
    .S(_0926_),
    .X(_1115_));
 sky130_fd_sc_hd__mux2i_1 _3642_ (.A0(\mem[13][21] ),
    .A1(\mem[15][21] ),
    .S(_1041_),
    .Y(_1116_));
 sky130_fd_sc_hd__nand2_1 _3643_ (.A(_0878_),
    .B(_1116_),
    .Y(_1117_));
 sky130_fd_sc_hd__o211ai_1 _3644_ (.A1(_1002_),
    .A2(_1115_),
    .B1(_1117_),
    .C1(_0930_),
    .Y(_1118_));
 sky130_fd_sc_hd__o21ai_0 _3645_ (.A1(_1054_),
    .A2(_1114_),
    .B1(_1118_),
    .Y(_1119_));
 sky130_fd_sc_hd__mux2i_2 _3646_ (.A0(\mem[0][21] ),
    .A1(\mem[2][21] ),
    .S(_1101_),
    .Y(_1120_));
 sky130_fd_sc_hd__mux2i_1 _3647_ (.A0(\mem[1][21] ),
    .A1(\mem[3][21] ),
    .S(_0887_),
    .Y(_1121_));
 sky130_fd_sc_hd__mux2i_1 _3648_ (.A0(\mem[8][21] ),
    .A1(\mem[10][21] ),
    .S(_0952_),
    .Y(_1122_));
 sky130_fd_sc_hd__mux2i_2 _3649_ (.A0(\mem[9][21] ),
    .A1(\mem[11][21] ),
    .S(_0954_),
    .Y(_1123_));
 sky130_fd_sc_hd__mux4_1 _3650_ (.A0(_1120_),
    .A1(_1121_),
    .A2(_1122_),
    .A3(_1123_),
    .S0(_1012_),
    .S1(_0992_),
    .X(_1124_));
 sky130_fd_sc_hd__nor2_1 _3651_ (.A(_1026_),
    .B(_1124_),
    .Y(_1125_));
 sky130_fd_sc_hd__a21oi_2 _3652_ (.A1(_0866_),
    .A2(_1119_),
    .B1(_1125_),
    .Y(_1126_));
 sky130_fd_sc_hd__nand2_1 _3653_ (.A(net91),
    .B(_1071_),
    .Y(_1127_));
 sky130_fd_sc_hd__o21ai_0 _3654_ (.A1(_1035_),
    .A2(_1126_),
    .B1(_1127_),
    .Y(_0548_));
 sky130_fd_sc_hd__buf_4 _3655_ (.A(_0861_),
    .X(_1128_));
 sky130_fd_sc_hd__mux2_1 _3656_ (.A0(\mem[4][22] ),
    .A1(\mem[6][22] ),
    .S(_1091_),
    .X(_1129_));
 sky130_fd_sc_hd__mux2i_1 _3657_ (.A0(\mem[5][22] ),
    .A1(\mem[7][22] ),
    .S(_1111_),
    .Y(_1130_));
 sky130_fd_sc_hd__nand2_1 _3658_ (.A(_0978_),
    .B(_1130_),
    .Y(_1131_));
 sky130_fd_sc_hd__o21ai_0 _3659_ (.A1(_0997_),
    .A2(_1129_),
    .B1(_1131_),
    .Y(_1132_));
 sky130_fd_sc_hd__mux2_1 _3660_ (.A0(\mem[12][22] ),
    .A1(\mem[14][22] ),
    .S(_0926_),
    .X(_1133_));
 sky130_fd_sc_hd__buf_4 _3661_ (.A(_0854_),
    .X(_1134_));
 sky130_fd_sc_hd__mux2i_1 _3662_ (.A0(\mem[13][22] ),
    .A1(\mem[15][22] ),
    .S(_1041_),
    .Y(_1135_));
 sky130_fd_sc_hd__nand2_1 _3663_ (.A(_1134_),
    .B(_1135_),
    .Y(_1136_));
 sky130_fd_sc_hd__o211ai_1 _3664_ (.A1(_1002_),
    .A2(_1133_),
    .B1(_1136_),
    .C1(_0930_),
    .Y(_1137_));
 sky130_fd_sc_hd__o21ai_0 _3665_ (.A1(_1054_),
    .A2(_1132_),
    .B1(_1137_),
    .Y(_1138_));
 sky130_fd_sc_hd__mux2i_2 _3666_ (.A0(\mem[0][22] ),
    .A1(\mem[2][22] ),
    .S(_1101_),
    .Y(_1139_));
 sky130_fd_sc_hd__buf_6 _3667_ (.A(_0835_),
    .X(_1140_));
 sky130_fd_sc_hd__mux2i_1 _3668_ (.A0(\mem[1][22] ),
    .A1(\mem[3][22] ),
    .S(_1140_),
    .Y(_1141_));
 sky130_fd_sc_hd__buf_8 _3669_ (.A(_0830_),
    .X(_1142_));
 sky130_fd_sc_hd__mux2i_2 _3670_ (.A0(\mem[8][22] ),
    .A1(\mem[10][22] ),
    .S(_1142_),
    .Y(_1143_));
 sky130_fd_sc_hd__mux2i_2 _3671_ (.A0(\mem[9][22] ),
    .A1(\mem[11][22] ),
    .S(_0954_),
    .Y(_1144_));
 sky130_fd_sc_hd__mux4_1 _3672_ (.A0(_1139_),
    .A1(_1141_),
    .A2(_1143_),
    .A3(_1144_),
    .S0(_1012_),
    .S1(_0992_),
    .X(_1145_));
 sky130_fd_sc_hd__nor2_1 _3673_ (.A(_1026_),
    .B(_1145_),
    .Y(_1146_));
 sky130_fd_sc_hd__a21oi_2 _3674_ (.A1(_1128_),
    .A2(_1138_),
    .B1(_1146_),
    .Y(_1147_));
 sky130_fd_sc_hd__nand2_1 _3675_ (.A(net92),
    .B(_1071_),
    .Y(_1148_));
 sky130_fd_sc_hd__o21ai_0 _3676_ (.A1(_1035_),
    .A2(_1147_),
    .B1(_1148_),
    .Y(_0549_));
 sky130_fd_sc_hd__mux2_1 _3677_ (.A0(\mem[4][23] ),
    .A1(\mem[6][23] ),
    .S(_1091_),
    .X(_1149_));
 sky130_fd_sc_hd__mux2i_1 _3678_ (.A0(\mem[5][23] ),
    .A1(\mem[7][23] ),
    .S(_1111_),
    .Y(_1150_));
 sky130_fd_sc_hd__nand2_1 _3679_ (.A(_0978_),
    .B(_1150_),
    .Y(_1151_));
 sky130_fd_sc_hd__o21ai_1 _3680_ (.A1(_0997_),
    .A2(_1149_),
    .B1(_1151_),
    .Y(_1152_));
 sky130_fd_sc_hd__buf_6 _3681_ (.A(_0722_),
    .X(_1153_));
 sky130_fd_sc_hd__mux2_1 _3682_ (.A0(\mem[12][23] ),
    .A1(\mem[14][23] ),
    .S(_1153_),
    .X(_1154_));
 sky130_fd_sc_hd__mux2i_1 _3683_ (.A0(\mem[13][23] ),
    .A1(\mem[15][23] ),
    .S(_1041_),
    .Y(_1155_));
 sky130_fd_sc_hd__nand2_1 _3684_ (.A(_1134_),
    .B(_1155_),
    .Y(_1156_));
 sky130_fd_sc_hd__buf_4 _3685_ (.A(_0841_),
    .X(_1157_));
 sky130_fd_sc_hd__o211ai_1 _3686_ (.A1(_1002_),
    .A2(_1154_),
    .B1(_1156_),
    .C1(_1157_),
    .Y(_1158_));
 sky130_fd_sc_hd__o21ai_0 _3687_ (.A1(_1054_),
    .A2(_1152_),
    .B1(_1158_),
    .Y(_1159_));
 sky130_fd_sc_hd__mux2i_2 _3688_ (.A0(\mem[0][23] ),
    .A1(\mem[2][23] ),
    .S(_1101_),
    .Y(_1160_));
 sky130_fd_sc_hd__mux2i_1 _3689_ (.A0(\mem[1][23] ),
    .A1(\mem[3][23] ),
    .S(_1140_),
    .Y(_1161_));
 sky130_fd_sc_hd__mux2i_2 _3690_ (.A0(\mem[8][23] ),
    .A1(\mem[10][23] ),
    .S(_1142_),
    .Y(_1162_));
 sky130_fd_sc_hd__mux2i_2 _3691_ (.A0(\mem[9][23] ),
    .A1(\mem[11][23] ),
    .S(_0954_),
    .Y(_1163_));
 sky130_fd_sc_hd__mux4_1 _3692_ (.A0(_1160_),
    .A1(_1161_),
    .A2(_1162_),
    .A3(_1163_),
    .S0(_1012_),
    .S1(_0992_),
    .X(_1164_));
 sky130_fd_sc_hd__nor2_1 _3693_ (.A(_1026_),
    .B(_1164_),
    .Y(_1165_));
 sky130_fd_sc_hd__a21oi_1 _3694_ (.A1(_1128_),
    .A2(_1159_),
    .B1(_1165_),
    .Y(_1166_));
 sky130_fd_sc_hd__nand2_1 _3695_ (.A(net93),
    .B(_1071_),
    .Y(_1167_));
 sky130_fd_sc_hd__o21ai_0 _3696_ (.A1(_1035_),
    .A2(_1166_),
    .B1(_1167_),
    .Y(_0550_));
 sky130_fd_sc_hd__mux2_1 _3697_ (.A0(\mem[0][24] ),
    .A1(\mem[2][24] ),
    .S(_0833_),
    .X(_1168_));
 sky130_fd_sc_hd__buf_6 _3698_ (.A(_0849_),
    .X(_1169_));
 sky130_fd_sc_hd__mux2i_1 _3699_ (.A0(\mem[1][24] ),
    .A1(\mem[3][24] ),
    .S(_0846_),
    .Y(_1170_));
 sky130_fd_sc_hd__nand2_1 _3700_ (.A(_1169_),
    .B(_1170_),
    .Y(_1171_));
 sky130_fd_sc_hd__o21ai_0 _3701_ (.A1(_0997_),
    .A2(_1168_),
    .B1(_1171_),
    .Y(_1172_));
 sky130_fd_sc_hd__mux2i_2 _3702_ (.A0(\mem[8][24] ),
    .A1(\mem[10][24] ),
    .S(_0879_),
    .Y(_1173_));
 sky130_fd_sc_hd__nand2_1 _3703_ (.A(_0903_),
    .B(_1173_),
    .Y(_1174_));
 sky130_fd_sc_hd__mux2i_1 _3704_ (.A0(\mem[9][24] ),
    .A1(\mem[11][24] ),
    .S(_0907_),
    .Y(_1175_));
 sky130_fd_sc_hd__nand2_1 _3705_ (.A(_0876_),
    .B(_1175_),
    .Y(_1176_));
 sky130_fd_sc_hd__nand3_1 _3706_ (.A(_0882_),
    .B(_1174_),
    .C(_1176_),
    .Y(_1177_));
 sky130_fd_sc_hd__o21ai_0 _3707_ (.A1(_1054_),
    .A2(_1172_),
    .B1(_1177_),
    .Y(_1178_));
 sky130_fd_sc_hd__mux2i_2 _3708_ (.A0(\mem[5][24] ),
    .A1(\mem[7][24] ),
    .S(_0890_),
    .Y(_1179_));
 sky130_fd_sc_hd__mux2i_2 _3709_ (.A0(\mem[4][24] ),
    .A1(\mem[6][24] ),
    .S(_0831_),
    .Y(_1180_));
 sky130_fd_sc_hd__mux2i_1 _3710_ (.A0(\mem[13][24] ),
    .A1(\mem[15][24] ),
    .S(_1142_),
    .Y(_1181_));
 sky130_fd_sc_hd__mux2i_1 _3711_ (.A0(\mem[12][24] ),
    .A1(\mem[14][24] ),
    .S(_0916_),
    .Y(_1182_));
 sky130_fd_sc_hd__clkbuf_8 _3712_ (.A(_0841_),
    .X(_1183_));
 sky130_fd_sc_hd__mux4_1 _3713_ (.A0(_1179_),
    .A1(_1180_),
    .A2(_1181_),
    .A3(_1182_),
    .S0(_0845_),
    .S1(_1183_),
    .X(_1184_));
 sky130_fd_sc_hd__nor2_1 _3714_ (.A(_0897_),
    .B(_1184_),
    .Y(_1185_));
 sky130_fd_sc_hd__a21oi_2 _3715_ (.A1(_0898_),
    .A2(_1178_),
    .B1(_1185_),
    .Y(_1186_));
 sky130_fd_sc_hd__nand2_1 _3716_ (.A(net94),
    .B(_1071_),
    .Y(_1187_));
 sky130_fd_sc_hd__o21ai_0 _3717_ (.A1(_1035_),
    .A2(_1186_),
    .B1(_1187_),
    .Y(_0551_));
 sky130_fd_sc_hd__buf_6 _3718_ (.A(_0839_),
    .X(_1188_));
 sky130_fd_sc_hd__mux2_1 _3719_ (.A0(\mem[4][25] ),
    .A1(\mem[6][25] ),
    .S(_1091_),
    .X(_1189_));
 sky130_fd_sc_hd__mux2i_2 _3720_ (.A0(\mem[5][25] ),
    .A1(\mem[7][25] ),
    .S(_1111_),
    .Y(_1190_));
 sky130_fd_sc_hd__nand2_1 _3721_ (.A(_1169_),
    .B(_1190_),
    .Y(_1191_));
 sky130_fd_sc_hd__o21ai_1 _3722_ (.A1(_1188_),
    .A2(_1189_),
    .B1(_1191_),
    .Y(_1192_));
 sky130_fd_sc_hd__mux2_1 _3723_ (.A0(\mem[12][25] ),
    .A1(\mem[14][25] ),
    .S(_1153_),
    .X(_1193_));
 sky130_fd_sc_hd__mux2i_1 _3724_ (.A0(\mem[13][25] ),
    .A1(\mem[15][25] ),
    .S(_1041_),
    .Y(_1194_));
 sky130_fd_sc_hd__nand2_1 _3725_ (.A(_1134_),
    .B(_1194_),
    .Y(_1195_));
 sky130_fd_sc_hd__o211ai_1 _3726_ (.A1(_1002_),
    .A2(_1193_),
    .B1(_1195_),
    .C1(_1157_),
    .Y(_1196_));
 sky130_fd_sc_hd__o21ai_0 _3727_ (.A1(_1054_),
    .A2(_1192_),
    .B1(_1196_),
    .Y(_1197_));
 sky130_fd_sc_hd__mux2i_2 _3728_ (.A0(\mem[0][25] ),
    .A1(\mem[2][25] ),
    .S(_1101_),
    .Y(_1198_));
 sky130_fd_sc_hd__mux2i_1 _3729_ (.A0(\mem[1][25] ),
    .A1(\mem[3][25] ),
    .S(_1140_),
    .Y(_1199_));
 sky130_fd_sc_hd__mux2i_2 _3730_ (.A0(\mem[8][25] ),
    .A1(\mem[10][25] ),
    .S(_1142_),
    .Y(_1200_));
 sky130_fd_sc_hd__buf_8 _3731_ (.A(_0830_),
    .X(_1201_));
 sky130_fd_sc_hd__mux2i_2 _3732_ (.A0(\mem[9][25] ),
    .A1(\mem[11][25] ),
    .S(_1201_),
    .Y(_1202_));
 sky130_fd_sc_hd__mux4_1 _3733_ (.A0(_1198_),
    .A1(_1199_),
    .A2(_1200_),
    .A3(_1202_),
    .S0(_1012_),
    .S1(_1183_),
    .X(_1203_));
 sky130_fd_sc_hd__nor2_1 _3734_ (.A(_1026_),
    .B(_1203_),
    .Y(_1204_));
 sky130_fd_sc_hd__a21oi_1 _3735_ (.A1(_1128_),
    .A2(_1197_),
    .B1(_1204_),
    .Y(_1205_));
 sky130_fd_sc_hd__nand2_1 _3736_ (.A(net95),
    .B(_1071_),
    .Y(_1206_));
 sky130_fd_sc_hd__o21ai_0 _3737_ (.A1(_1035_),
    .A2(_1205_),
    .B1(_1206_),
    .Y(_0552_));
 sky130_fd_sc_hd__mux2_1 _3738_ (.A0(\mem[4][26] ),
    .A1(\mem[6][26] ),
    .S(_1091_),
    .X(_1207_));
 sky130_fd_sc_hd__mux2i_1 _3739_ (.A0(\mem[5][26] ),
    .A1(\mem[7][26] ),
    .S(_1111_),
    .Y(_1208_));
 sky130_fd_sc_hd__nand2_1 _3740_ (.A(_1169_),
    .B(_1208_),
    .Y(_1209_));
 sky130_fd_sc_hd__o21ai_1 _3741_ (.A1(_1188_),
    .A2(_1207_),
    .B1(_1209_),
    .Y(_1210_));
 sky130_fd_sc_hd__mux2_1 _3742_ (.A0(\mem[12][26] ),
    .A1(\mem[14][26] ),
    .S(_1153_),
    .X(_1211_));
 sky130_fd_sc_hd__mux2i_1 _3743_ (.A0(\mem[13][26] ),
    .A1(\mem[15][26] ),
    .S(_1041_),
    .Y(_1212_));
 sky130_fd_sc_hd__nand2_1 _3744_ (.A(_1134_),
    .B(_1212_),
    .Y(_1213_));
 sky130_fd_sc_hd__o211ai_1 _3745_ (.A1(_1002_),
    .A2(_1211_),
    .B1(_1213_),
    .C1(_1157_),
    .Y(_1214_));
 sky130_fd_sc_hd__o21ai_0 _3746_ (.A1(_1054_),
    .A2(_1210_),
    .B1(_1214_),
    .Y(_1215_));
 sky130_fd_sc_hd__mux2i_2 _3747_ (.A0(\mem[0][26] ),
    .A1(\mem[2][26] ),
    .S(_1101_),
    .Y(_1216_));
 sky130_fd_sc_hd__mux2i_1 _3748_ (.A0(\mem[1][26] ),
    .A1(\mem[3][26] ),
    .S(_1140_),
    .Y(_1217_));
 sky130_fd_sc_hd__mux2i_1 _3749_ (.A0(\mem[8][26] ),
    .A1(\mem[10][26] ),
    .S(_1142_),
    .Y(_1218_));
 sky130_fd_sc_hd__mux2i_2 _3750_ (.A0(\mem[9][26] ),
    .A1(\mem[11][26] ),
    .S(_1201_),
    .Y(_1219_));
 sky130_fd_sc_hd__mux4_1 _3751_ (.A0(_1216_),
    .A1(_1217_),
    .A2(_1218_),
    .A3(_1219_),
    .S0(_1012_),
    .S1(_1183_),
    .X(_1220_));
 sky130_fd_sc_hd__nor2_1 _3752_ (.A(_1026_),
    .B(_1220_),
    .Y(_1221_));
 sky130_fd_sc_hd__a21oi_1 _3753_ (.A1(_1128_),
    .A2(_1215_),
    .B1(_1221_),
    .Y(_1222_));
 sky130_fd_sc_hd__nand2_1 _3754_ (.A(net96),
    .B(_1071_),
    .Y(_1223_));
 sky130_fd_sc_hd__o21ai_0 _3755_ (.A1(_1035_),
    .A2(_1222_),
    .B1(_1223_),
    .Y(_0553_));
 sky130_fd_sc_hd__clkbuf_8 _3756_ (.A(_0714_),
    .X(_1224_));
 sky130_fd_sc_hd__mux2_1 _3757_ (.A0(\mem[4][27] ),
    .A1(\mem[6][27] ),
    .S(_1091_),
    .X(_1225_));
 sky130_fd_sc_hd__mux2i_1 _3758_ (.A0(\mem[5][27] ),
    .A1(\mem[7][27] ),
    .S(_1111_),
    .Y(_1226_));
 sky130_fd_sc_hd__nand2_1 _3759_ (.A(_1169_),
    .B(_1226_),
    .Y(_1227_));
 sky130_fd_sc_hd__o21ai_1 _3760_ (.A1(_1188_),
    .A2(_1225_),
    .B1(_1227_),
    .Y(_1228_));
 sky130_fd_sc_hd__buf_6 _3761_ (.A(_0854_),
    .X(_1229_));
 sky130_fd_sc_hd__mux2_1 _3762_ (.A0(\mem[12][27] ),
    .A1(\mem[14][27] ),
    .S(_1153_),
    .X(_1230_));
 sky130_fd_sc_hd__mux2i_1 _3763_ (.A0(\mem[13][27] ),
    .A1(\mem[15][27] ),
    .S(_1041_),
    .Y(_1231_));
 sky130_fd_sc_hd__nand2_1 _3764_ (.A(_1134_),
    .B(_1231_),
    .Y(_1232_));
 sky130_fd_sc_hd__o211ai_1 _3765_ (.A1(_1229_),
    .A2(_1230_),
    .B1(_1232_),
    .C1(_1157_),
    .Y(_1233_));
 sky130_fd_sc_hd__o21ai_0 _3766_ (.A1(_1054_),
    .A2(_1228_),
    .B1(_1233_),
    .Y(_1234_));
 sky130_fd_sc_hd__mux2i_2 _3767_ (.A0(\mem[0][27] ),
    .A1(\mem[2][27] ),
    .S(_1101_),
    .Y(_1235_));
 sky130_fd_sc_hd__mux2i_1 _3768_ (.A0(\mem[1][27] ),
    .A1(\mem[3][27] ),
    .S(_1140_),
    .Y(_1236_));
 sky130_fd_sc_hd__mux2i_1 _3769_ (.A0(\mem[8][27] ),
    .A1(\mem[10][27] ),
    .S(_1142_),
    .Y(_1237_));
 sky130_fd_sc_hd__mux2i_2 _3770_ (.A0(\mem[9][27] ),
    .A1(\mem[11][27] ),
    .S(_1201_),
    .Y(_1238_));
 sky130_fd_sc_hd__buf_8 _3771_ (.A(_0839_),
    .X(_1239_));
 sky130_fd_sc_hd__mux4_1 _3772_ (.A0(_1235_),
    .A1(_1236_),
    .A2(_1237_),
    .A3(_1238_),
    .S0(_1239_),
    .S1(_1183_),
    .X(_1240_));
 sky130_fd_sc_hd__nor2_1 _3773_ (.A(_1026_),
    .B(_1240_),
    .Y(_1241_));
 sky130_fd_sc_hd__a21oi_1 _3774_ (.A1(_1128_),
    .A2(_1234_),
    .B1(_1241_),
    .Y(_1242_));
 sky130_fd_sc_hd__nand2_1 _3775_ (.A(net97),
    .B(_1071_),
    .Y(_1243_));
 sky130_fd_sc_hd__o21ai_0 _3776_ (.A1(_1224_),
    .A2(_1242_),
    .B1(_1243_),
    .Y(_0554_));
 sky130_fd_sc_hd__clkbuf_8 _3777_ (.A(_0841_),
    .X(_1244_));
 sky130_fd_sc_hd__mux2_1 _3778_ (.A0(\mem[4][28] ),
    .A1(\mem[6][28] ),
    .S(_1091_),
    .X(_1245_));
 sky130_fd_sc_hd__mux2i_1 _3779_ (.A0(\mem[5][28] ),
    .A1(\mem[7][28] ),
    .S(_1111_),
    .Y(_1246_));
 sky130_fd_sc_hd__nand2_1 _3780_ (.A(_1169_),
    .B(_1246_),
    .Y(_1247_));
 sky130_fd_sc_hd__o21ai_1 _3781_ (.A1(_1188_),
    .A2(_1245_),
    .B1(_1247_),
    .Y(_1248_));
 sky130_fd_sc_hd__mux2_1 _3782_ (.A0(\mem[12][28] ),
    .A1(\mem[14][28] ),
    .S(_1153_),
    .X(_1249_));
 sky130_fd_sc_hd__mux2i_1 _3783_ (.A0(\mem[13][28] ),
    .A1(\mem[15][28] ),
    .S(_1041_),
    .Y(_1250_));
 sky130_fd_sc_hd__nand2_1 _3784_ (.A(_1134_),
    .B(_1250_),
    .Y(_1251_));
 sky130_fd_sc_hd__o211ai_1 _3785_ (.A1(_1229_),
    .A2(_1249_),
    .B1(_1251_),
    .C1(_1157_),
    .Y(_1252_));
 sky130_fd_sc_hd__o21ai_0 _3786_ (.A1(_1244_),
    .A2(_1248_),
    .B1(_1252_),
    .Y(_1253_));
 sky130_fd_sc_hd__mux2i_2 _3787_ (.A0(\mem[0][28] ),
    .A1(\mem[2][28] ),
    .S(_1101_),
    .Y(_1254_));
 sky130_fd_sc_hd__mux2i_1 _3788_ (.A0(\mem[1][28] ),
    .A1(\mem[3][28] ),
    .S(_1140_),
    .Y(_1255_));
 sky130_fd_sc_hd__mux2i_1 _3789_ (.A0(\mem[8][28] ),
    .A1(\mem[10][28] ),
    .S(_1142_),
    .Y(_1256_));
 sky130_fd_sc_hd__mux2i_1 _3790_ (.A0(\mem[9][28] ),
    .A1(\mem[11][28] ),
    .S(_1201_),
    .Y(_1257_));
 sky130_fd_sc_hd__mux4_1 _3791_ (.A0(_1254_),
    .A1(_1255_),
    .A2(_1256_),
    .A3(_1257_),
    .S0(_1239_),
    .S1(_1183_),
    .X(_1258_));
 sky130_fd_sc_hd__nor2_1 _3792_ (.A(_0865_),
    .B(_1258_),
    .Y(_1259_));
 sky130_fd_sc_hd__a21oi_1 _3793_ (.A1(_1128_),
    .A2(_1253_),
    .B1(_1259_),
    .Y(_1260_));
 sky130_fd_sc_hd__buf_4 _3794_ (.A(_0825_),
    .X(_1261_));
 sky130_fd_sc_hd__nand2_1 _3795_ (.A(net98),
    .B(_1261_),
    .Y(_1262_));
 sky130_fd_sc_hd__o21ai_0 _3796_ (.A1(_1224_),
    .A2(_1260_),
    .B1(_1262_),
    .Y(_0555_));
 sky130_fd_sc_hd__mux2_1 _3797_ (.A0(\mem[0][29] ),
    .A1(\mem[2][29] ),
    .S(_0833_),
    .X(_1263_));
 sky130_fd_sc_hd__mux2i_1 _3798_ (.A0(\mem[1][29] ),
    .A1(\mem[3][29] ),
    .S(_0846_),
    .Y(_1264_));
 sky130_fd_sc_hd__nand2_1 _3799_ (.A(_1169_),
    .B(_1264_),
    .Y(_1265_));
 sky130_fd_sc_hd__o21ai_0 _3800_ (.A1(_1188_),
    .A2(_1263_),
    .B1(_1265_),
    .Y(_1266_));
 sky130_fd_sc_hd__mux2i_1 _3801_ (.A0(\mem[8][29] ),
    .A1(\mem[10][29] ),
    .S(_0879_),
    .Y(_1267_));
 sky130_fd_sc_hd__nand2_1 _3802_ (.A(_0903_),
    .B(_1267_),
    .Y(_1268_));
 sky130_fd_sc_hd__mux2i_1 _3803_ (.A0(\mem[9][29] ),
    .A1(\mem[11][29] ),
    .S(_0907_),
    .Y(_1269_));
 sky130_fd_sc_hd__nand2_1 _3804_ (.A(_0876_),
    .B(_1269_),
    .Y(_1270_));
 sky130_fd_sc_hd__nand3_1 _3805_ (.A(_0882_),
    .B(_1268_),
    .C(_1270_),
    .Y(_1271_));
 sky130_fd_sc_hd__o21ai_0 _3806_ (.A1(_1244_),
    .A2(_1266_),
    .B1(_1271_),
    .Y(_1272_));
 sky130_fd_sc_hd__mux2i_2 _3807_ (.A0(\mem[5][29] ),
    .A1(\mem[7][29] ),
    .S(_0890_),
    .Y(_1273_));
 sky130_fd_sc_hd__mux2i_1 _3808_ (.A0(\mem[4][29] ),
    .A1(\mem[6][29] ),
    .S(_0831_),
    .Y(_1274_));
 sky130_fd_sc_hd__mux2i_2 _3809_ (.A0(\mem[13][29] ),
    .A1(\mem[15][29] ),
    .S(_1142_),
    .Y(_1275_));
 sky130_fd_sc_hd__mux2i_2 _3810_ (.A0(\mem[12][29] ),
    .A1(\mem[14][29] ),
    .S(_0916_),
    .Y(_1276_));
 sky130_fd_sc_hd__mux4_1 _3811_ (.A0(_1273_),
    .A1(_1274_),
    .A2(_1275_),
    .A3(_1276_),
    .S0(_0840_),
    .S1(_1183_),
    .X(_1277_));
 sky130_fd_sc_hd__nor2_1 _3812_ (.A(_0897_),
    .B(_1277_),
    .Y(_1278_));
 sky130_fd_sc_hd__a21oi_2 _3813_ (.A1(_0898_),
    .A2(_1272_),
    .B1(_1278_),
    .Y(_1279_));
 sky130_fd_sc_hd__nand2_1 _3814_ (.A(net99),
    .B(_1261_),
    .Y(_1280_));
 sky130_fd_sc_hd__o21ai_0 _3815_ (.A1(_1224_),
    .A2(_1279_),
    .B1(_1280_),
    .Y(_0556_));
 sky130_fd_sc_hd__mux2_1 _3816_ (.A0(\mem[4][2] ),
    .A1(\mem[6][2] ),
    .S(_1091_),
    .X(_1281_));
 sky130_fd_sc_hd__mux2i_1 _3817_ (.A0(\mem[5][2] ),
    .A1(\mem[7][2] ),
    .S(_1111_),
    .Y(_1282_));
 sky130_fd_sc_hd__nand2_1 _3818_ (.A(_1169_),
    .B(_1282_),
    .Y(_1283_));
 sky130_fd_sc_hd__o21ai_1 _3819_ (.A1(_1188_),
    .A2(_1281_),
    .B1(_1283_),
    .Y(_1284_));
 sky130_fd_sc_hd__mux2_1 _3820_ (.A0(\mem[12][2] ),
    .A1(\mem[14][2] ),
    .S(_1153_),
    .X(_1285_));
 sky130_fd_sc_hd__mux2i_1 _3821_ (.A0(\mem[13][2] ),
    .A1(\mem[15][2] ),
    .S(_0851_),
    .Y(_1286_));
 sky130_fd_sc_hd__nand2_1 _3822_ (.A(_1134_),
    .B(_1286_),
    .Y(_1287_));
 sky130_fd_sc_hd__o211ai_1 _3823_ (.A1(_1229_),
    .A2(_1285_),
    .B1(_1287_),
    .C1(_1157_),
    .Y(_1288_));
 sky130_fd_sc_hd__o21ai_0 _3824_ (.A1(_1244_),
    .A2(_1284_),
    .B1(_1288_),
    .Y(_1289_));
 sky130_fd_sc_hd__mux2i_4 _3825_ (.A0(\mem[0][2] ),
    .A1(\mem[2][2] ),
    .S(_1101_),
    .Y(_1290_));
 sky130_fd_sc_hd__mux2i_2 _3826_ (.A0(\mem[1][2] ),
    .A1(\mem[3][2] ),
    .S(_1140_),
    .Y(_1291_));
 sky130_fd_sc_hd__mux2i_1 _3827_ (.A0(\mem[8][2] ),
    .A1(\mem[10][2] ),
    .S(_1142_),
    .Y(_1292_));
 sky130_fd_sc_hd__mux2i_1 _3828_ (.A0(\mem[9][2] ),
    .A1(\mem[11][2] ),
    .S(_1201_),
    .Y(_1293_));
 sky130_fd_sc_hd__mux4_1 _3829_ (.A0(_1290_),
    .A1(_1291_),
    .A2(_1292_),
    .A3(_1293_),
    .S0(_1239_),
    .S1(_1183_),
    .X(_1294_));
 sky130_fd_sc_hd__nor2_1 _3830_ (.A(_0865_),
    .B(_1294_),
    .Y(_1295_));
 sky130_fd_sc_hd__a21oi_1 _3831_ (.A1(_1128_),
    .A2(_1289_),
    .B1(_1295_),
    .Y(_1296_));
 sky130_fd_sc_hd__nand2_1 _3832_ (.A(net100),
    .B(_1261_),
    .Y(_1297_));
 sky130_fd_sc_hd__o21ai_0 _3833_ (.A1(_1224_),
    .A2(_1296_),
    .B1(_1297_),
    .Y(_0557_));
 sky130_fd_sc_hd__mux2_1 _3834_ (.A0(\mem[4][30] ),
    .A1(\mem[6][30] ),
    .S(_1091_),
    .X(_1298_));
 sky130_fd_sc_hd__mux2i_1 _3835_ (.A0(\mem[5][30] ),
    .A1(\mem[7][30] ),
    .S(_1111_),
    .Y(_1299_));
 sky130_fd_sc_hd__nand2_1 _3836_ (.A(_1169_),
    .B(_1299_),
    .Y(_1300_));
 sky130_fd_sc_hd__o21ai_1 _3837_ (.A1(_1188_),
    .A2(_1298_),
    .B1(_1300_),
    .Y(_1301_));
 sky130_fd_sc_hd__mux2_1 _3838_ (.A0(\mem[12][30] ),
    .A1(\mem[14][30] ),
    .S(_1153_),
    .X(_1302_));
 sky130_fd_sc_hd__mux2i_1 _3839_ (.A0(\mem[13][30] ),
    .A1(\mem[15][30] ),
    .S(_0851_),
    .Y(_1303_));
 sky130_fd_sc_hd__nand2_1 _3840_ (.A(_1134_),
    .B(_1303_),
    .Y(_1304_));
 sky130_fd_sc_hd__o211ai_1 _3841_ (.A1(_1229_),
    .A2(_1302_),
    .B1(_1304_),
    .C1(_1157_),
    .Y(_1305_));
 sky130_fd_sc_hd__o21ai_0 _3842_ (.A1(_1244_),
    .A2(_1301_),
    .B1(_1305_),
    .Y(_1306_));
 sky130_fd_sc_hd__mux2i_2 _3843_ (.A0(\mem[0][30] ),
    .A1(\mem[2][30] ),
    .S(_1101_),
    .Y(_1307_));
 sky130_fd_sc_hd__mux2i_1 _3844_ (.A0(\mem[1][30] ),
    .A1(\mem[3][30] ),
    .S(_1140_),
    .Y(_1308_));
 sky130_fd_sc_hd__mux2i_1 _3845_ (.A0(\mem[8][30] ),
    .A1(\mem[10][30] ),
    .S(_1142_),
    .Y(_1309_));
 sky130_fd_sc_hd__mux2i_1 _3846_ (.A0(\mem[9][30] ),
    .A1(\mem[11][30] ),
    .S(_1201_),
    .Y(_1310_));
 sky130_fd_sc_hd__mux4_1 _3847_ (.A0(_1307_),
    .A1(_1308_),
    .A2(_1309_),
    .A3(_1310_),
    .S0(_1239_),
    .S1(_1183_),
    .X(_1311_));
 sky130_fd_sc_hd__nor2_1 _3848_ (.A(_0865_),
    .B(_1311_),
    .Y(_1312_));
 sky130_fd_sc_hd__a21oi_1 _3849_ (.A1(_1128_),
    .A2(_1306_),
    .B1(_1312_),
    .Y(_1313_));
 sky130_fd_sc_hd__nand2_1 _3850_ (.A(net101),
    .B(_1261_),
    .Y(_1314_));
 sky130_fd_sc_hd__o21ai_0 _3851_ (.A1(_1224_),
    .A2(_1313_),
    .B1(_1314_),
    .Y(_0558_));
 sky130_fd_sc_hd__mux2_1 _3852_ (.A0(\mem[4][31] ),
    .A1(\mem[6][31] ),
    .S(_0855_),
    .X(_1315_));
 sky130_fd_sc_hd__mux2i_1 _3853_ (.A0(\mem[5][31] ),
    .A1(\mem[7][31] ),
    .S(_1111_),
    .Y(_1316_));
 sky130_fd_sc_hd__nand2_1 _3854_ (.A(_1169_),
    .B(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hd__o21ai_1 _3855_ (.A1(_1188_),
    .A2(_1315_),
    .B1(_1317_),
    .Y(_1318_));
 sky130_fd_sc_hd__mux2_1 _3856_ (.A0(\mem[12][31] ),
    .A1(\mem[14][31] ),
    .S(_1153_),
    .X(_1319_));
 sky130_fd_sc_hd__mux2i_1 _3857_ (.A0(\mem[13][31] ),
    .A1(\mem[15][31] ),
    .S(_0851_),
    .Y(_1320_));
 sky130_fd_sc_hd__nand2_1 _3858_ (.A(_1134_),
    .B(_1320_),
    .Y(_1321_));
 sky130_fd_sc_hd__o211ai_1 _3859_ (.A1(_1229_),
    .A2(_1319_),
    .B1(_1321_),
    .C1(_1157_),
    .Y(_1322_));
 sky130_fd_sc_hd__o21ai_0 _3860_ (.A1(_1244_),
    .A2(_1318_),
    .B1(_1322_),
    .Y(_1323_));
 sky130_fd_sc_hd__mux2i_2 _3861_ (.A0(\mem[0][31] ),
    .A1(\mem[2][31] ),
    .S(_0837_),
    .Y(_1324_));
 sky130_fd_sc_hd__mux2i_1 _3862_ (.A0(\mem[1][31] ),
    .A1(\mem[3][31] ),
    .S(_1140_),
    .Y(_1325_));
 sky130_fd_sc_hd__mux2i_1 _3863_ (.A0(\mem[8][31] ),
    .A1(\mem[10][31] ),
    .S(_0914_),
    .Y(_1326_));
 sky130_fd_sc_hd__mux2i_2 _3864_ (.A0(\mem[9][31] ),
    .A1(\mem[11][31] ),
    .S(_1201_),
    .Y(_1327_));
 sky130_fd_sc_hd__mux4_1 _3865_ (.A0(_1324_),
    .A1(_1325_),
    .A2(_1326_),
    .A3(_1327_),
    .S0(_1239_),
    .S1(_1183_),
    .X(_1328_));
 sky130_fd_sc_hd__nor2_1 _3866_ (.A(_0865_),
    .B(_1328_),
    .Y(_1329_));
 sky130_fd_sc_hd__a21oi_1 _3867_ (.A1(_1128_),
    .A2(_1323_),
    .B1(_1329_),
    .Y(_1330_));
 sky130_fd_sc_hd__nand2_1 _3868_ (.A(net102),
    .B(_1261_),
    .Y(_1331_));
 sky130_fd_sc_hd__o21ai_0 _3869_ (.A1(_1224_),
    .A2(_1330_),
    .B1(_1331_),
    .Y(_0559_));
 sky130_fd_sc_hd__mux2_1 _3870_ (.A0(\mem[4][3] ),
    .A1(\mem[6][3] ),
    .S(_0855_),
    .X(_1332_));
 sky130_fd_sc_hd__mux2i_1 _3871_ (.A0(\mem[5][3] ),
    .A1(\mem[7][3] ),
    .S(_0846_),
    .Y(_1333_));
 sky130_fd_sc_hd__nand2_1 _3872_ (.A(_1169_),
    .B(_1333_),
    .Y(_1334_));
 sky130_fd_sc_hd__o21ai_0 _3873_ (.A1(_1188_),
    .A2(_1332_),
    .B1(_1334_),
    .Y(_1335_));
 sky130_fd_sc_hd__mux2_1 _3874_ (.A0(\mem[12][3] ),
    .A1(\mem[14][3] ),
    .S(_1153_),
    .X(_1336_));
 sky130_fd_sc_hd__mux2i_1 _3875_ (.A0(\mem[13][3] ),
    .A1(\mem[15][3] ),
    .S(_0851_),
    .Y(_1337_));
 sky130_fd_sc_hd__nand2_1 _3876_ (.A(_1134_),
    .B(_1337_),
    .Y(_1338_));
 sky130_fd_sc_hd__o211ai_1 _3877_ (.A1(_1229_),
    .A2(_1336_),
    .B1(_1338_),
    .C1(_1157_),
    .Y(_1339_));
 sky130_fd_sc_hd__o21ai_0 _3878_ (.A1(_1244_),
    .A2(_1335_),
    .B1(_1339_),
    .Y(_1340_));
 sky130_fd_sc_hd__mux2i_2 _3879_ (.A0(\mem[0][3] ),
    .A1(\mem[2][3] ),
    .S(_0837_),
    .Y(_1341_));
 sky130_fd_sc_hd__mux2i_1 _3880_ (.A0(\mem[1][3] ),
    .A1(\mem[3][3] ),
    .S(_1140_),
    .Y(_1342_));
 sky130_fd_sc_hd__mux2i_2 _3881_ (.A0(\mem[8][3] ),
    .A1(\mem[10][3] ),
    .S(_0914_),
    .Y(_1343_));
 sky130_fd_sc_hd__mux2i_1 _3882_ (.A0(\mem[9][3] ),
    .A1(\mem[11][3] ),
    .S(_1201_),
    .Y(_1344_));
 sky130_fd_sc_hd__mux4_1 _3883_ (.A0(_1341_),
    .A1(_1342_),
    .A2(_1343_),
    .A3(_1344_),
    .S0(_1239_),
    .S1(_1183_),
    .X(_1345_));
 sky130_fd_sc_hd__nor2_1 _3884_ (.A(_0865_),
    .B(_1345_),
    .Y(_1346_));
 sky130_fd_sc_hd__a21oi_2 _3885_ (.A1(_1128_),
    .A2(_1340_),
    .B1(_1346_),
    .Y(_1347_));
 sky130_fd_sc_hd__nand2_1 _3886_ (.A(net111),
    .B(_1261_),
    .Y(_1348_));
 sky130_fd_sc_hd__o21ai_0 _3887_ (.A1(_1224_),
    .A2(_1347_),
    .B1(_1348_),
    .Y(_0560_));
 sky130_fd_sc_hd__mux2_1 _3888_ (.A0(\mem[0][4] ),
    .A1(\mem[2][4] ),
    .S(_0835_),
    .X(_1349_));
 sky130_fd_sc_hd__mux2i_1 _3889_ (.A0(\mem[1][4] ),
    .A1(\mem[3][4] ),
    .S(_0869_),
    .Y(_1350_));
 sky130_fd_sc_hd__nand2_1 _3890_ (.A(_0850_),
    .B(_1350_),
    .Y(_1351_));
 sky130_fd_sc_hd__o21ai_0 _3891_ (.A1(_1188_),
    .A2(_1349_),
    .B1(_1351_),
    .Y(_1352_));
 sky130_fd_sc_hd__mux2i_1 _3892_ (.A0(\mem[8][4] ),
    .A1(\mem[10][4] ),
    .S(_0879_),
    .Y(_1353_));
 sky130_fd_sc_hd__nand2_1 _3893_ (.A(_0845_),
    .B(_1353_),
    .Y(_1354_));
 sky130_fd_sc_hd__mux2i_1 _3894_ (.A0(\mem[9][4] ),
    .A1(\mem[11][4] ),
    .S(_0907_),
    .Y(_1355_));
 sky130_fd_sc_hd__nand2_1 _3895_ (.A(_0876_),
    .B(_1355_),
    .Y(_1356_));
 sky130_fd_sc_hd__nand3_1 _3896_ (.A(_0882_),
    .B(_1354_),
    .C(_1356_),
    .Y(_1357_));
 sky130_fd_sc_hd__o21ai_0 _3897_ (.A1(_1244_),
    .A2(_1352_),
    .B1(_1357_),
    .Y(_1358_));
 sky130_fd_sc_hd__mux2i_1 _3898_ (.A0(\mem[5][4] ),
    .A1(\mem[7][4] ),
    .S(_0890_),
    .Y(_1359_));
 sky130_fd_sc_hd__mux2i_2 _3899_ (.A0(\mem[4][4] ),
    .A1(\mem[6][4] ),
    .S(_0831_),
    .Y(_1360_));
 sky130_fd_sc_hd__mux2i_1 _3900_ (.A0(\mem[13][4] ),
    .A1(\mem[15][4] ),
    .S(_0914_),
    .Y(_1361_));
 sky130_fd_sc_hd__mux2i_1 _3901_ (.A0(\mem[12][4] ),
    .A1(\mem[14][4] ),
    .S(_0916_),
    .Y(_1362_));
 sky130_fd_sc_hd__mux4_1 _3902_ (.A0(_1359_),
    .A1(_1360_),
    .A2(_1361_),
    .A3(_1362_),
    .S0(_0840_),
    .S1(_0842_),
    .X(_1363_));
 sky130_fd_sc_hd__nor2_1 _3903_ (.A(_0897_),
    .B(_1363_),
    .Y(_1364_));
 sky130_fd_sc_hd__a21oi_2 _3904_ (.A1(_0898_),
    .A2(_1358_),
    .B1(_1364_),
    .Y(_1365_));
 sky130_fd_sc_hd__nand2_1 _3905_ (.A(net122),
    .B(_1261_),
    .Y(_1366_));
 sky130_fd_sc_hd__o21ai_0 _3906_ (.A1(_1224_),
    .A2(_1365_),
    .B1(_1366_),
    .Y(_0561_));
 sky130_fd_sc_hd__mux2_1 _3907_ (.A0(\mem[4][5] ),
    .A1(\mem[6][5] ),
    .S(_0855_),
    .X(_1367_));
 sky130_fd_sc_hd__mux2i_1 _3908_ (.A0(\mem[5][5] ),
    .A1(\mem[7][5] ),
    .S(_0846_),
    .Y(_1368_));
 sky130_fd_sc_hd__nand2_1 _3909_ (.A(_0850_),
    .B(_1368_),
    .Y(_1369_));
 sky130_fd_sc_hd__o21ai_0 _3910_ (.A1(_0871_),
    .A2(_1367_),
    .B1(_1369_),
    .Y(_1370_));
 sky130_fd_sc_hd__mux2_1 _3911_ (.A0(\mem[12][5] ),
    .A1(\mem[14][5] ),
    .S(_1153_),
    .X(_1371_));
 sky130_fd_sc_hd__mux2i_1 _3912_ (.A0(\mem[13][5] ),
    .A1(\mem[15][5] ),
    .S(_0851_),
    .Y(_1372_));
 sky130_fd_sc_hd__nand2_1 _3913_ (.A(_0868_),
    .B(_1372_),
    .Y(_1373_));
 sky130_fd_sc_hd__o211ai_1 _3914_ (.A1(_1229_),
    .A2(_1371_),
    .B1(_1373_),
    .C1(_1157_),
    .Y(_1374_));
 sky130_fd_sc_hd__o21ai_0 _3915_ (.A1(_1244_),
    .A2(_1370_),
    .B1(_1374_),
    .Y(_1375_));
 sky130_fd_sc_hd__mux2i_2 _3916_ (.A0(\mem[0][5] ),
    .A1(\mem[2][5] ),
    .S(_0837_),
    .Y(_1376_));
 sky130_fd_sc_hd__mux2i_2 _3917_ (.A0(\mem[1][5] ),
    .A1(\mem[3][5] ),
    .S(_0916_),
    .Y(_1377_));
 sky130_fd_sc_hd__mux2i_2 _3918_ (.A0(\mem[8][5] ),
    .A1(\mem[10][5] ),
    .S(_0914_),
    .Y(_1378_));
 sky130_fd_sc_hd__mux2i_2 _3919_ (.A0(\mem[9][5] ),
    .A1(\mem[11][5] ),
    .S(_1201_),
    .Y(_1379_));
 sky130_fd_sc_hd__mux4_1 _3920_ (.A0(_1376_),
    .A1(_1377_),
    .A2(_1378_),
    .A3(_1379_),
    .S0(_1239_),
    .S1(_0842_),
    .X(_1380_));
 sky130_fd_sc_hd__nor2_1 _3921_ (.A(_0865_),
    .B(_1380_),
    .Y(_1381_));
 sky130_fd_sc_hd__a21oi_1 _3922_ (.A1(_0829_),
    .A2(_1375_),
    .B1(_1381_),
    .Y(_1382_));
 sky130_fd_sc_hd__nand2_1 _3923_ (.A(net133),
    .B(_1261_),
    .Y(_1383_));
 sky130_fd_sc_hd__o21ai_0 _3924_ (.A1(_1224_),
    .A2(_1382_),
    .B1(_1383_),
    .Y(_0562_));
 sky130_fd_sc_hd__mux2_1 _3925_ (.A0(\mem[4][6] ),
    .A1(\mem[6][6] ),
    .S(_0855_),
    .X(_1384_));
 sky130_fd_sc_hd__mux2i_1 _3926_ (.A0(\mem[5][6] ),
    .A1(\mem[7][6] ),
    .S(_0846_),
    .Y(_1385_));
 sky130_fd_sc_hd__nand2_1 _3927_ (.A(_0850_),
    .B(_1385_),
    .Y(_1386_));
 sky130_fd_sc_hd__o21ai_0 _3928_ (.A1(_0871_),
    .A2(_1384_),
    .B1(_1386_),
    .Y(_1387_));
 sky130_fd_sc_hd__mux2_1 _3929_ (.A0(\mem[12][6] ),
    .A1(\mem[14][6] ),
    .S(_0833_),
    .X(_1388_));
 sky130_fd_sc_hd__mux2i_1 _3930_ (.A0(\mem[13][6] ),
    .A1(\mem[15][6] ),
    .S(_0851_),
    .Y(_1389_));
 sky130_fd_sc_hd__nand2_1 _3931_ (.A(_0868_),
    .B(_1389_),
    .Y(_1390_));
 sky130_fd_sc_hd__o211ai_1 _3932_ (.A1(_1229_),
    .A2(_1388_),
    .B1(_1390_),
    .C1(_0844_),
    .Y(_1391_));
 sky130_fd_sc_hd__o21ai_0 _3933_ (.A1(_1244_),
    .A2(_1387_),
    .B1(_1391_),
    .Y(_1392_));
 sky130_fd_sc_hd__mux2i_2 _3934_ (.A0(\mem[0][6] ),
    .A1(\mem[2][6] ),
    .S(_0837_),
    .Y(_1393_));
 sky130_fd_sc_hd__mux2i_1 _3935_ (.A0(\mem[1][6] ),
    .A1(\mem[3][6] ),
    .S(_0916_),
    .Y(_1394_));
 sky130_fd_sc_hd__mux2i_1 _3936_ (.A0(\mem[8][6] ),
    .A1(\mem[10][6] ),
    .S(_0914_),
    .Y(_1395_));
 sky130_fd_sc_hd__mux2i_1 _3937_ (.A0(\mem[9][6] ),
    .A1(\mem[11][6] ),
    .S(_1201_),
    .Y(_1396_));
 sky130_fd_sc_hd__mux4_1 _3938_ (.A0(_1393_),
    .A1(_1394_),
    .A2(_1395_),
    .A3(_1396_),
    .S0(_1239_),
    .S1(_0842_),
    .X(_1397_));
 sky130_fd_sc_hd__nor2_1 _3939_ (.A(_0865_),
    .B(_1397_),
    .Y(_1398_));
 sky130_fd_sc_hd__a21oi_1 _3940_ (.A1(_0829_),
    .A2(_1392_),
    .B1(_1398_),
    .Y(_1399_));
 sky130_fd_sc_hd__nand2_1 _3941_ (.A(net138),
    .B(_1261_),
    .Y(_1400_));
 sky130_fd_sc_hd__o21ai_0 _3942_ (.A1(_1224_),
    .A2(_1399_),
    .B1(_1400_),
    .Y(_0563_));
 sky130_fd_sc_hd__mux2_1 _3943_ (.A0(\mem[4][7] ),
    .A1(\mem[6][7] ),
    .S(_0855_),
    .X(_1401_));
 sky130_fd_sc_hd__mux2i_1 _3944_ (.A0(\mem[5][7] ),
    .A1(\mem[7][7] ),
    .S(_0846_),
    .Y(_1402_));
 sky130_fd_sc_hd__nand2_1 _3945_ (.A(_0850_),
    .B(_1402_),
    .Y(_1403_));
 sky130_fd_sc_hd__o21ai_0 _3946_ (.A1(_0871_),
    .A2(_1401_),
    .B1(_1403_),
    .Y(_1404_));
 sky130_fd_sc_hd__mux2_1 _3947_ (.A0(\mem[12][7] ),
    .A1(\mem[14][7] ),
    .S(_0833_),
    .X(_1405_));
 sky130_fd_sc_hd__mux2i_1 _3948_ (.A0(\mem[13][7] ),
    .A1(\mem[15][7] ),
    .S(_0851_),
    .Y(_1406_));
 sky130_fd_sc_hd__nand2_1 _3949_ (.A(_0868_),
    .B(_1406_),
    .Y(_1407_));
 sky130_fd_sc_hd__o211ai_1 _3950_ (.A1(_1229_),
    .A2(_1405_),
    .B1(_1407_),
    .C1(_0844_),
    .Y(_1408_));
 sky130_fd_sc_hd__o21ai_0 _3951_ (.A1(_1244_),
    .A2(_1404_),
    .B1(_1408_),
    .Y(_1409_));
 sky130_fd_sc_hd__mux2i_2 _3952_ (.A0(\mem[0][7] ),
    .A1(\mem[2][7] ),
    .S(_0837_),
    .Y(_1410_));
 sky130_fd_sc_hd__mux2i_1 _3953_ (.A0(\mem[1][7] ),
    .A1(\mem[3][7] ),
    .S(_0916_),
    .Y(_1411_));
 sky130_fd_sc_hd__mux2i_1 _3954_ (.A0(\mem[8][7] ),
    .A1(\mem[10][7] ),
    .S(_0914_),
    .Y(_1412_));
 sky130_fd_sc_hd__mux2i_1 _3955_ (.A0(\mem[9][7] ),
    .A1(\mem[11][7] ),
    .S(_0885_),
    .Y(_1413_));
 sky130_fd_sc_hd__mux4_1 _3956_ (.A0(_1410_),
    .A1(_1411_),
    .A2(_1412_),
    .A3(_1413_),
    .S0(_1239_),
    .S1(_0842_),
    .X(_1414_));
 sky130_fd_sc_hd__nor2_1 _3957_ (.A(_0865_),
    .B(_1414_),
    .Y(_1415_));
 sky130_fd_sc_hd__a21oi_1 _3958_ (.A1(_0829_),
    .A2(_1409_),
    .B1(_1415_),
    .Y(_1416_));
 sky130_fd_sc_hd__nand2_1 _3959_ (.A(net139),
    .B(_1261_),
    .Y(_1417_));
 sky130_fd_sc_hd__o21ai_0 _3960_ (.A1(_0825_),
    .A2(_1416_),
    .B1(_1417_),
    .Y(_0564_));
 sky130_fd_sc_hd__mux2_1 _3961_ (.A0(\mem[4][8] ),
    .A1(\mem[6][8] ),
    .S(_0855_),
    .X(_1418_));
 sky130_fd_sc_hd__mux2i_1 _3962_ (.A0(\mem[5][8] ),
    .A1(\mem[7][8] ),
    .S(_0846_),
    .Y(_1419_));
 sky130_fd_sc_hd__nand2_1 _3963_ (.A(_0850_),
    .B(_1419_),
    .Y(_1420_));
 sky130_fd_sc_hd__o21ai_0 _3964_ (.A1(_0871_),
    .A2(_1418_),
    .B1(_1420_),
    .Y(_1421_));
 sky130_fd_sc_hd__mux2_1 _3965_ (.A0(\mem[12][8] ),
    .A1(\mem[14][8] ),
    .S(_0833_),
    .X(_1422_));
 sky130_fd_sc_hd__mux2i_1 _3966_ (.A0(\mem[13][8] ),
    .A1(\mem[15][8] ),
    .S(_0851_),
    .Y(_1423_));
 sky130_fd_sc_hd__nand2_1 _3967_ (.A(_0868_),
    .B(_1423_),
    .Y(_1424_));
 sky130_fd_sc_hd__o211ai_1 _3968_ (.A1(_1229_),
    .A2(_1422_),
    .B1(_1424_),
    .C1(_0844_),
    .Y(_1425_));
 sky130_fd_sc_hd__o21ai_0 _3969_ (.A1(_0882_),
    .A2(_1421_),
    .B1(_1425_),
    .Y(_1426_));
 sky130_fd_sc_hd__mux2i_2 _3970_ (.A0(\mem[0][8] ),
    .A1(\mem[2][8] ),
    .S(_0837_),
    .Y(_1427_));
 sky130_fd_sc_hd__mux2i_1 _3971_ (.A0(\mem[1][8] ),
    .A1(\mem[3][8] ),
    .S(_0916_),
    .Y(_1428_));
 sky130_fd_sc_hd__mux2i_1 _3972_ (.A0(\mem[8][8] ),
    .A1(\mem[10][8] ),
    .S(_0914_),
    .Y(_1429_));
 sky130_fd_sc_hd__mux2i_1 _3973_ (.A0(\mem[9][8] ),
    .A1(\mem[11][8] ),
    .S(_0885_),
    .Y(_1430_));
 sky130_fd_sc_hd__mux4_1 _3974_ (.A0(_1427_),
    .A1(_1428_),
    .A2(_1429_),
    .A3(_1430_),
    .S0(_1239_),
    .S1(_0842_),
    .X(_1431_));
 sky130_fd_sc_hd__nor2_1 _3975_ (.A(_0865_),
    .B(_1431_),
    .Y(_1432_));
 sky130_fd_sc_hd__a21oi_1 _3976_ (.A1(_0829_),
    .A2(_1426_),
    .B1(_1432_),
    .Y(_1433_));
 sky130_fd_sc_hd__nand2_1 _3977_ (.A(net140),
    .B(_0864_),
    .Y(_1434_));
 sky130_fd_sc_hd__o21ai_0 _3978_ (.A1(_0825_),
    .A2(_1433_),
    .B1(_1434_),
    .Y(_0565_));
 sky130_fd_sc_hd__mux2_1 _3979_ (.A0(\mem[0][9] ),
    .A1(\mem[2][9] ),
    .S(_0835_),
    .X(_1435_));
 sky130_fd_sc_hd__mux2i_1 _3980_ (.A0(\mem[1][9] ),
    .A1(\mem[3][9] ),
    .S(_0869_),
    .Y(_1436_));
 sky130_fd_sc_hd__nand2_1 _3981_ (.A(_0850_),
    .B(_1436_),
    .Y(_1437_));
 sky130_fd_sc_hd__o21ai_0 _3982_ (.A1(_0871_),
    .A2(_1435_),
    .B1(_1437_),
    .Y(_1438_));
 sky130_fd_sc_hd__mux2i_1 _3983_ (.A0(\mem[8][9] ),
    .A1(\mem[10][9] ),
    .S(_0879_),
    .Y(_1439_));
 sky130_fd_sc_hd__nand2_1 _3984_ (.A(_0845_),
    .B(_1439_),
    .Y(_1440_));
 sky130_fd_sc_hd__mux2i_1 _3985_ (.A0(\mem[9][9] ),
    .A1(\mem[11][9] ),
    .S(_0907_),
    .Y(_1441_));
 sky130_fd_sc_hd__nand2_1 _3986_ (.A(_0876_),
    .B(_1441_),
    .Y(_1442_));
 sky130_fd_sc_hd__nand3_1 _3987_ (.A(_0882_),
    .B(_1440_),
    .C(_1442_),
    .Y(_1443_));
 sky130_fd_sc_hd__o21ai_0 _3988_ (.A1(_0882_),
    .A2(_1438_),
    .B1(_1443_),
    .Y(_1444_));
 sky130_fd_sc_hd__mux2i_1 _3989_ (.A0(\mem[5][9] ),
    .A1(\mem[7][9] ),
    .S(_0890_),
    .Y(_1445_));
 sky130_fd_sc_hd__mux2i_1 _3990_ (.A0(\mem[4][9] ),
    .A1(\mem[6][9] ),
    .S(_0831_),
    .Y(_1446_));
 sky130_fd_sc_hd__mux2i_1 _3991_ (.A0(\mem[13][9] ),
    .A1(\mem[15][9] ),
    .S(_0914_),
    .Y(_1447_));
 sky130_fd_sc_hd__mux2i_2 _3992_ (.A0(\mem[12][9] ),
    .A1(\mem[14][9] ),
    .S(_0890_),
    .Y(_1448_));
 sky130_fd_sc_hd__mux4_1 _3993_ (.A0(_1445_),
    .A1(_1446_),
    .A2(_1447_),
    .A3(_1448_),
    .S0(_0840_),
    .S1(_0842_),
    .X(_1449_));
 sky130_fd_sc_hd__nor2_1 _3994_ (.A(_0897_),
    .B(_1449_),
    .Y(_1450_));
 sky130_fd_sc_hd__a21oi_2 _3995_ (.A1(_0898_),
    .A2(_1444_),
    .B1(_1450_),
    .Y(_1451_));
 sky130_fd_sc_hd__nand2_1 _3996_ (.A(net141),
    .B(_0864_),
    .Y(_1452_));
 sky130_fd_sc_hd__o21ai_0 _3997_ (.A1(_0825_),
    .A2(_1451_),
    .B1(_1452_),
    .Y(_0566_));
 sky130_fd_sc_hd__inv_2 _3998_ (.A(_0711_),
    .Y(_1453_));
 sky130_fd_sc_hd__nor4b_4 _3999_ (.A(_0609_),
    .B(_0607_),
    .C(net73),
    .D_N(_2557_),
    .Y(_1454_));
 sky130_fd_sc_hd__o21ai_4 _4000_ (.A1(_1453_),
    .A2(_1454_),
    .B1(_2492_),
    .Y(_1455_));
 sky130_fd_sc_hd__buf_6 _4001_ (.A(_1455_),
    .X(_1456_));
 sky130_fd_sc_hd__buf_6 _4002_ (.A(_2518_),
    .X(_1457_));
 sky130_fd_sc_hd__or3_1 _4003_ (.A(_1453_),
    .B(_1457_),
    .C(_1454_),
    .X(_1458_));
 sky130_fd_sc_hd__clkbuf_2 _4004_ (.A(_1458_),
    .X(_1459_));
 sky130_fd_sc_hd__buf_6 _4005_ (.A(_1459_),
    .X(_1460_));
 sky130_fd_sc_hd__o22ai_1 _4006_ (.A1(\mem[9][0] ),
    .A2(_1456_),
    .B1(_1460_),
    .B2(\mem[8][0] ),
    .Y(_1461_));
 sky130_fd_sc_hd__nand3_4 _4007_ (.A(_0711_),
    .B(_1457_),
    .C(net219),
    .Y(_1462_));
 sky130_fd_sc_hd__buf_6 _4008_ (.A(_1462_),
    .X(_1463_));
 sky130_fd_sc_hd__o21ai_4 _4009_ (.A1(_1453_),
    .A2(_1454_),
    .B1(_0830_),
    .Y(_1464_));
 sky130_fd_sc_hd__buf_6 _4010_ (.A(_1464_),
    .X(_1465_));
 sky130_fd_sc_hd__o22ai_1 _4011_ (.A1(\mem[10][0] ),
    .A2(_1463_),
    .B1(_1465_),
    .B2(\mem[11][0] ),
    .Y(_1466_));
 sky130_fd_sc_hd__buf_4 _4012_ (.A(_2517_),
    .X(_1467_));
 sky130_fd_sc_hd__inv_2 _4013_ (.A(_1467_),
    .Y(_1468_));
 sky130_fd_sc_hd__nor2_2 _4014_ (.A(_0826_),
    .B(_1468_),
    .Y(_1469_));
 sky130_fd_sc_hd__a31oi_2 _4015_ (.A1(_0711_),
    .A2(_1467_),
    .A3(net166),
    .B1(_0896_),
    .Y(_1470_));
 sky130_fd_sc_hd__a211o_4 _4016_ (.A1(_0715_),
    .A2(_1469_),
    .B1(_1470_),
    .C1(_0840_),
    .X(_1471_));
 sky130_fd_sc_hd__clkbuf_8 _4017_ (.A(_1471_),
    .X(_1472_));
 sky130_fd_sc_hd__nor3_1 _4018_ (.A(_1461_),
    .B(_1466_),
    .C(_1472_),
    .Y(_1473_));
 sky130_fd_sc_hd__and3_1 _4019_ (.A(_0840_),
    .B(\rd_ptr[3] ),
    .C(_0721_),
    .X(_1474_));
 sky130_fd_sc_hd__buf_4 _4020_ (.A(_1474_),
    .X(_1475_));
 sky130_fd_sc_hd__buf_6 _4021_ (.A(_1475_),
    .X(_1476_));
 sky130_fd_sc_hd__xnor2_1 _4022_ (.A(_0826_),
    .B(_1467_),
    .Y(_1477_));
 sky130_fd_sc_hd__buf_4 _4023_ (.A(_1477_),
    .X(_1478_));
 sky130_fd_sc_hd__buf_4 _4024_ (.A(_1478_),
    .X(_1479_));
 sky130_fd_sc_hd__buf_8 _4025_ (.A(_1457_),
    .X(_1480_));
 sky130_fd_sc_hd__buf_8 _4026_ (.A(_1480_),
    .X(_1481_));
 sky130_fd_sc_hd__mux2i_1 _4027_ (.A0(\mem[13][0] ),
    .A1(\mem[15][0] ),
    .S(_1481_),
    .Y(_1482_));
 sky130_fd_sc_hd__buf_6 _4028_ (.A(_1457_),
    .X(_1483_));
 sky130_fd_sc_hd__mux2_1 _4029_ (.A0(\mem[9][0] ),
    .A1(\mem[11][0] ),
    .S(_1483_),
    .X(_1484_));
 sky130_fd_sc_hd__nand3_1 _4030_ (.A(_0897_),
    .B(_1468_),
    .C(_1484_),
    .Y(_1485_));
 sky130_fd_sc_hd__o21ai_0 _4031_ (.A1(_1479_),
    .A2(_1482_),
    .B1(_1485_),
    .Y(_1486_));
 sky130_fd_sc_hd__nand2_1 _4032_ (.A(net222),
    .B(_1486_),
    .Y(_1487_));
 sky130_fd_sc_hd__buf_6 _4033_ (.A(_0827_),
    .X(_1488_));
 sky130_fd_sc_hd__clkbuf_4 _4034_ (.A(_0715_),
    .X(_1489_));
 sky130_fd_sc_hd__buf_6 _4035_ (.A(_0711_),
    .X(_1490_));
 sky130_fd_sc_hd__buf_6 _4036_ (.A(net220),
    .X(_1491_));
 sky130_fd_sc_hd__nand4_1 _4037_ (.A(_1490_),
    .B(_1467_),
    .C(_1491_),
    .D(_1484_),
    .Y(_1492_));
 sky130_fd_sc_hd__o21ai_0 _4038_ (.A1(_1489_),
    .A2(_0838_),
    .B1(_1492_),
    .Y(_1493_));
 sky130_fd_sc_hd__o21ai_4 _4039_ (.A1(_1453_),
    .A2(_1454_),
    .B1(_0896_),
    .Y(_1494_));
 sky130_fd_sc_hd__buf_6 _4040_ (.A(_1494_),
    .X(_1495_));
 sky130_fd_sc_hd__nor2_1 _4041_ (.A(_0847_),
    .B(_1495_),
    .Y(_1496_));
 sky130_fd_sc_hd__a21oi_1 _4042_ (.A1(_1488_),
    .A2(_1493_),
    .B1(_1496_),
    .Y(_1497_));
 sky130_fd_sc_hd__nand4_1 _4043_ (.A(_0711_),
    .B(_0839_),
    .C(_0826_),
    .D(_0722_),
    .Y(_1498_));
 sky130_fd_sc_hd__o21ai_2 _4044_ (.A1(_1454_),
    .A2(_1498_),
    .B1(_0841_),
    .Y(_1499_));
 sky130_fd_sc_hd__or3_2 _4045_ (.A(_0841_),
    .B(_1454_),
    .C(_1498_),
    .X(_1500_));
 sky130_fd_sc_hd__a211oi_4 _4046_ (.A1(_1499_),
    .A2(_1500_),
    .B1(_0840_),
    .C1(net164),
    .Y(_1501_));
 sky130_fd_sc_hd__nor2_1 _4047_ (.A(_0896_),
    .B(_1467_),
    .Y(_1502_));
 sky130_fd_sc_hd__mux2_1 _4048_ (.A0(\mem[12][0] ),
    .A1(\mem[14][0] ),
    .S(_1480_),
    .X(_1503_));
 sky130_fd_sc_hd__o211ai_1 _4049_ (.A1(_1502_),
    .A2(_1469_),
    .B1(_1503_),
    .C1(_1489_),
    .Y(_1504_));
 sky130_fd_sc_hd__or3_1 _4050_ (.A(_0896_),
    .B(_0715_),
    .C(_0836_),
    .X(_1505_));
 sky130_fd_sc_hd__and3_1 _4051_ (.A(_1501_),
    .B(_1504_),
    .C(_1505_),
    .X(_1506_));
 sky130_fd_sc_hd__a31oi_1 _4052_ (.A1(_1476_),
    .A2(_1487_),
    .A3(_1497_),
    .B1(_1506_),
    .Y(_1507_));
 sky130_fd_sc_hd__nand2_2 _4053_ (.A(_1499_),
    .B(_1500_),
    .Y(_1508_));
 sky130_fd_sc_hd__nor3_4 _4054_ (.A(_0845_),
    .B(_2534_),
    .C(_1508_),
    .Y(_1509_));
 sky130_fd_sc_hd__buf_8 _4055_ (.A(_1483_),
    .X(_1510_));
 sky130_fd_sc_hd__mux4_1 _4056_ (.A0(\mem[4][0] ),
    .A1(\mem[6][0] ),
    .A2(\mem[0][0] ),
    .A3(\mem[2][0] ),
    .S0(_1510_),
    .S1(_1478_),
    .X(_1511_));
 sky130_fd_sc_hd__nand2_1 _4057_ (.A(_0529_),
    .B(_1511_),
    .Y(_1512_));
 sky130_fd_sc_hd__nand2_1 _4058_ (.A(_0897_),
    .B(_0856_),
    .Y(_1513_));
 sky130_fd_sc_hd__buf_8 _4059_ (.A(_0827_),
    .X(_1514_));
 sky130_fd_sc_hd__nand2_1 _4060_ (.A(_1514_),
    .B(_0832_),
    .Y(_1515_));
 sky130_fd_sc_hd__nand3_1 _4061_ (.A(_0825_),
    .B(_1513_),
    .C(_1515_),
    .Y(_1516_));
 sky130_fd_sc_hd__mux4_1 _4062_ (.A0(\mem[5][0] ),
    .A1(\mem[7][0] ),
    .A2(\mem[1][0] ),
    .A3(\mem[3][0] ),
    .S0(_1480_),
    .S1(_1478_),
    .X(_1517_));
 sky130_fd_sc_hd__nor2_1 _4063_ (.A(_0827_),
    .B(_0857_),
    .Y(_1518_));
 sky130_fd_sc_hd__buf_4 _4064_ (.A(_0715_),
    .X(_1519_));
 sky130_fd_sc_hd__a211oi_1 _4065_ (.A1(_0828_),
    .A2(_0834_),
    .B1(_1518_),
    .C1(_1519_),
    .Y(_1520_));
 sky130_fd_sc_hd__or3_1 _4066_ (.A(_0839_),
    .B(_0841_),
    .C(net164),
    .X(_1521_));
 sky130_fd_sc_hd__clkbuf_4 _4067_ (.A(_1521_),
    .X(_1522_));
 sky130_fd_sc_hd__a211oi_1 _4068_ (.A1(_0529_),
    .A2(_1517_),
    .B1(_1520_),
    .C1(_1522_),
    .Y(_1523_));
 sky130_fd_sc_hd__a31oi_1 _4069_ (.A1(_1509_),
    .A2(_1512_),
    .A3(_1516_),
    .B1(_1523_),
    .Y(_1524_));
 sky130_fd_sc_hd__o221a_1 _4070_ (.A1(net103),
    .A2(_2537_),
    .B1(_1473_),
    .B2(_1507_),
    .C1(_1524_),
    .X(_0567_));
 sky130_fd_sc_hd__buf_6 _4071_ (.A(_0850_),
    .X(_1525_));
 sky130_fd_sc_hd__nor2_4 _4072_ (.A(_0896_),
    .B(_0715_),
    .Y(_1526_));
 sky130_fd_sc_hd__buf_4 _4073_ (.A(_1526_),
    .X(_1527_));
 sky130_fd_sc_hd__or3_1 _4074_ (.A(_1453_),
    .B(_1454_),
    .C(_1477_),
    .X(_1528_));
 sky130_fd_sc_hd__clkbuf_4 _4075_ (.A(_1528_),
    .X(_1529_));
 sky130_fd_sc_hd__buf_4 _4076_ (.A(_1529_),
    .X(_1530_));
 sky130_fd_sc_hd__buf_6 _4077_ (.A(_1530_),
    .X(_1531_));
 sky130_fd_sc_hd__buf_6 _4078_ (.A(_1483_),
    .X(_1532_));
 sky130_fd_sc_hd__buf_6 _4079_ (.A(_1532_),
    .X(_1533_));
 sky130_fd_sc_hd__mux2i_1 _4080_ (.A0(\mem[5][10] ),
    .A1(\mem[7][10] ),
    .S(_1533_),
    .Y(_1534_));
 sky130_fd_sc_hd__nor2_1 _4081_ (.A(_1531_),
    .B(_1534_),
    .Y(_1535_));
 sky130_fd_sc_hd__a21oi_1 _4082_ (.A1(_0870_),
    .A2(_1527_),
    .B1(_1535_),
    .Y(_1536_));
 sky130_fd_sc_hd__buf_4 _4083_ (.A(_0849_),
    .X(_1537_));
 sky130_fd_sc_hd__buf_6 _4084_ (.A(_0827_),
    .X(_1538_));
 sky130_fd_sc_hd__buf_6 _4085_ (.A(_0715_),
    .X(_1539_));
 sky130_fd_sc_hd__buf_4 _4086_ (.A(_0711_),
    .X(_1540_));
 sky130_fd_sc_hd__buf_4 _4087_ (.A(_1540_),
    .X(_1541_));
 sky130_fd_sc_hd__buf_4 _4088_ (.A(net220),
    .X(_1542_));
 sky130_fd_sc_hd__buf_4 _4089_ (.A(_1542_),
    .X(_1543_));
 sky130_fd_sc_hd__mux2_1 _4090_ (.A0(\mem[1][10] ),
    .A1(\mem[3][10] ),
    .S(_1510_),
    .X(_1544_));
 sky130_fd_sc_hd__nand4_1 _4091_ (.A(_1541_),
    .B(_1543_),
    .C(_1479_),
    .D(_1544_),
    .Y(_1545_));
 sky130_fd_sc_hd__o31ai_1 _4092_ (.A1(_1538_),
    .A2(_1539_),
    .A3(_0886_),
    .B1(_1545_),
    .Y(_1546_));
 sky130_fd_sc_hd__o21ai_1 _4093_ (.A1(_1453_),
    .A2(_1454_),
    .B1(_0826_),
    .Y(_1547_));
 sky130_fd_sc_hd__buf_6 _4094_ (.A(_1547_),
    .X(_1548_));
 sky130_fd_sc_hd__buf_4 _4095_ (.A(_1529_),
    .X(_1549_));
 sky130_fd_sc_hd__buf_16 _4096_ (.A(_1510_),
    .X(_1550_));
 sky130_fd_sc_hd__mux2i_1 _4097_ (.A0(\mem[4][10] ),
    .A1(\mem[6][10] ),
    .S(_1550_),
    .Y(_1551_));
 sky130_fd_sc_hd__buf_6 _4098_ (.A(_0854_),
    .X(_1552_));
 sky130_fd_sc_hd__o221ai_1 _4099_ (.A1(_0873_),
    .A2(_1548_),
    .B1(_1549_),
    .B2(_1551_),
    .C1(_1552_),
    .Y(_1553_));
 sky130_fd_sc_hd__o21ai_0 _4100_ (.A1(_1537_),
    .A2(_1546_),
    .B1(_1553_),
    .Y(_1554_));
 sky130_fd_sc_hd__buf_6 _4101_ (.A(_1455_),
    .X(_1555_));
 sky130_fd_sc_hd__buf_6 _4102_ (.A(_1459_),
    .X(_1556_));
 sky130_fd_sc_hd__o22ai_1 _4103_ (.A1(\mem[1][10] ),
    .A2(_1555_),
    .B1(_1556_),
    .B2(\mem[0][10] ),
    .Y(_1557_));
 sky130_fd_sc_hd__o22ai_1 _4104_ (.A1(\mem[2][10] ),
    .A2(_1463_),
    .B1(_1465_),
    .B2(\mem[3][10] ),
    .Y(_1558_));
 sky130_fd_sc_hd__or3_1 _4105_ (.A(_1472_),
    .B(_1557_),
    .C(_1558_),
    .X(_1559_));
 sky130_fd_sc_hd__nor2_4 _4106_ (.A(_2534_),
    .B(_1508_),
    .Y(_1560_));
 sky130_fd_sc_hd__buf_4 _4107_ (.A(_1560_),
    .X(_1561_));
 sky130_fd_sc_hd__o2111ai_1 _4108_ (.A1(_1525_),
    .A2(_1536_),
    .B1(_1554_),
    .C1(_1559_),
    .D1(_1561_),
    .Y(_1562_));
 sky130_fd_sc_hd__buf_6 _4109_ (.A(_1530_),
    .X(_1563_));
 sky130_fd_sc_hd__buf_4 _4110_ (.A(_1563_),
    .X(_1564_));
 sky130_fd_sc_hd__clkbuf_16 _4111_ (.A(_1550_),
    .X(_1565_));
 sky130_fd_sc_hd__mux2i_1 _4112_ (.A0(\mem[12][10] ),
    .A1(\mem[14][10] ),
    .S(_1565_),
    .Y(_1566_));
 sky130_fd_sc_hd__buf_4 _4113_ (.A(_0715_),
    .X(_1567_));
 sky130_fd_sc_hd__buf_6 _4114_ (.A(_1540_),
    .X(_1568_));
 sky130_fd_sc_hd__buf_6 _4115_ (.A(_1542_),
    .X(_1569_));
 sky130_fd_sc_hd__mux2_1 _4116_ (.A0(\mem[8][10] ),
    .A1(\mem[10][10] ),
    .S(_1480_),
    .X(_1570_));
 sky130_fd_sc_hd__nand3_1 _4117_ (.A(_1568_),
    .B(_1569_),
    .C(_1570_),
    .Y(_1571_));
 sky130_fd_sc_hd__buf_6 _4118_ (.A(_1467_),
    .X(_1572_));
 sky130_fd_sc_hd__o22ai_1 _4119_ (.A1(_1567_),
    .A2(_0891_),
    .B1(_1571_),
    .B2(_1572_),
    .Y(_1573_));
 sky130_fd_sc_hd__buf_6 _4120_ (.A(_1468_),
    .X(_1574_));
 sky130_fd_sc_hd__nor2_1 _4121_ (.A(_1574_),
    .B(_1571_),
    .Y(_1575_));
 sky130_fd_sc_hd__o21ai_0 _4122_ (.A1(net222),
    .A2(_0880_),
    .B1(_1488_),
    .Y(_1576_));
 sky130_fd_sc_hd__o22ai_1 _4123_ (.A1(_0861_),
    .A2(_1573_),
    .B1(_1575_),
    .B2(_1576_),
    .Y(_1577_));
 sky130_fd_sc_hd__buf_6 _4124_ (.A(_1501_),
    .X(_1578_));
 sky130_fd_sc_hd__o211ai_1 _4125_ (.A1(_1564_),
    .A2(_1566_),
    .B1(_1577_),
    .C1(_1578_),
    .Y(_1579_));
 sky130_fd_sc_hd__buf_6 _4126_ (.A(_1529_),
    .X(_1580_));
 sky130_fd_sc_hd__buf_8 _4127_ (.A(_1510_),
    .X(_1581_));
 sky130_fd_sc_hd__mux2i_1 _4128_ (.A0(\mem[13][10] ),
    .A1(\mem[15][10] ),
    .S(_1581_),
    .Y(_1582_));
 sky130_fd_sc_hd__clkbuf_8 _4129_ (.A(net221),
    .X(_1583_));
 sky130_fd_sc_hd__nand3_1 _4130_ (.A(_0828_),
    .B(_1583_),
    .C(_0877_),
    .Y(_1584_));
 sky130_fd_sc_hd__o221ai_1 _4131_ (.A1(_0889_),
    .A2(_1495_),
    .B1(_1580_),
    .B2(_1582_),
    .C1(_1584_),
    .Y(_1585_));
 sky130_fd_sc_hd__mux2i_1 _4132_ (.A0(\mem[9][10] ),
    .A1(\mem[11][10] ),
    .S(_1581_),
    .Y(_1586_));
 sky130_fd_sc_hd__nand3_1 _4133_ (.A(_0711_),
    .B(net166),
    .C(_1478_),
    .Y(_1587_));
 sky130_fd_sc_hd__buf_6 _4134_ (.A(_1587_),
    .X(_1588_));
 sky130_fd_sc_hd__clkbuf_8 _4135_ (.A(_1588_),
    .X(_1589_));
 sky130_fd_sc_hd__o21ai_0 _4136_ (.A1(_1586_),
    .A2(_1589_),
    .B1(_1476_),
    .Y(_1590_));
 sky130_fd_sc_hd__o22a_1 _4137_ (.A1(net114),
    .A2(_2537_),
    .B1(_1585_),
    .B2(_1590_),
    .X(_1591_));
 sky130_fd_sc_hd__and3_1 _4138_ (.A(_1562_),
    .B(_1579_),
    .C(_1591_),
    .X(_0568_));
 sky130_fd_sc_hd__and2_0 _4139_ (.A(_1499_),
    .B(_1500_),
    .X(_1592_));
 sky130_fd_sc_hd__clkbuf_4 _4140_ (.A(_1592_),
    .X(_1593_));
 sky130_fd_sc_hd__nor2_1 _4141_ (.A(net163),
    .B(_1593_),
    .Y(_1594_));
 sky130_fd_sc_hd__buf_4 _4142_ (.A(_0845_),
    .X(_1595_));
 sky130_fd_sc_hd__buf_4 _4143_ (.A(_1547_),
    .X(_1596_));
 sky130_fd_sc_hd__buf_4 _4144_ (.A(_1596_),
    .X(_1597_));
 sky130_fd_sc_hd__buf_4 _4145_ (.A(_1530_),
    .X(_1598_));
 sky130_fd_sc_hd__buf_6 _4146_ (.A(_1532_),
    .X(_1599_));
 sky130_fd_sc_hd__mux2i_1 _4147_ (.A0(\mem[13][11] ),
    .A1(\mem[15][11] ),
    .S(_1599_),
    .Y(_1600_));
 sky130_fd_sc_hd__o22ai_1 _4148_ (.A1(_0917_),
    .A2(_1597_),
    .B1(_1598_),
    .B2(_1600_),
    .Y(_1601_));
 sky130_fd_sc_hd__nand2_1 _4149_ (.A(_1595_),
    .B(_1601_),
    .Y(_1602_));
 sky130_fd_sc_hd__o22ai_1 _4150_ (.A1(\mem[9][11] ),
    .A2(_1555_),
    .B1(_1556_),
    .B2(\mem[8][11] ),
    .Y(_1603_));
 sky130_fd_sc_hd__o22ai_1 _4151_ (.A1(\mem[10][11] ),
    .A2(_1463_),
    .B1(_1465_),
    .B2(\mem[11][11] ),
    .Y(_1604_));
 sky130_fd_sc_hd__or3_1 _4152_ (.A(_1472_),
    .B(_1603_),
    .C(_1604_),
    .X(_1605_));
 sky130_fd_sc_hd__mux2i_1 _4153_ (.A0(\mem[12][11] ),
    .A1(\mem[14][11] ),
    .S(_1533_),
    .Y(_1606_));
 sky130_fd_sc_hd__o22ai_1 _4154_ (.A1(_0915_),
    .A2(_1548_),
    .B1(_1563_),
    .B2(_1606_),
    .Y(_1607_));
 sky130_fd_sc_hd__buf_8 _4155_ (.A(_1532_),
    .X(_1608_));
 sky130_fd_sc_hd__mux2i_1 _4156_ (.A0(\mem[9][11] ),
    .A1(\mem[11][11] ),
    .S(_1608_),
    .Y(_1609_));
 sky130_fd_sc_hd__o221ai_1 _4157_ (.A1(_0904_),
    .A2(_1495_),
    .B1(_1589_),
    .B2(_1609_),
    .C1(_0903_),
    .Y(_1610_));
 sky130_fd_sc_hd__o21ai_0 _4158_ (.A1(_0903_),
    .A2(_1607_),
    .B1(_1610_),
    .Y(_1611_));
 sky130_fd_sc_hd__nand4_1 _4159_ (.A(_1594_),
    .B(_1602_),
    .C(_1605_),
    .D(_1611_),
    .Y(_1612_));
 sky130_fd_sc_hd__mux2i_1 _4160_ (.A0(\mem[4][11] ),
    .A1(\mem[6][11] ),
    .S(_1565_),
    .Y(_1613_));
 sky130_fd_sc_hd__mux2_1 _4161_ (.A0(\mem[0][11] ),
    .A1(\mem[2][11] ),
    .S(_1480_),
    .X(_1614_));
 sky130_fd_sc_hd__nand3_1 _4162_ (.A(_1568_),
    .B(_1569_),
    .C(_1614_),
    .Y(_1615_));
 sky130_fd_sc_hd__o22ai_1 _4163_ (.A1(_1567_),
    .A2(_0900_),
    .B1(_1615_),
    .B2(_1572_),
    .Y(_1616_));
 sky130_fd_sc_hd__nor2_1 _4164_ (.A(_1574_),
    .B(_1615_),
    .Y(_1617_));
 sky130_fd_sc_hd__o21ai_0 _4165_ (.A1(net222),
    .A2(_0912_),
    .B1(_1488_),
    .Y(_1618_));
 sky130_fd_sc_hd__o22ai_1 _4166_ (.A1(_0861_),
    .A2(_1616_),
    .B1(_1617_),
    .B2(_1618_),
    .Y(_1619_));
 sky130_fd_sc_hd__o211ai_1 _4167_ (.A1(_1564_),
    .A2(_1613_),
    .B1(_1619_),
    .C1(_1509_),
    .Y(_1620_));
 sky130_fd_sc_hd__mux2i_1 _4168_ (.A0(\mem[1][11] ),
    .A1(\mem[3][11] ),
    .S(_1481_),
    .Y(_1621_));
 sky130_fd_sc_hd__nor2_1 _4169_ (.A(_1588_),
    .B(_1621_),
    .Y(_1622_));
 sky130_fd_sc_hd__mux2_1 _4170_ (.A0(\mem[5][11] ),
    .A1(\mem[7][11] ),
    .S(_1480_),
    .X(_1623_));
 sky130_fd_sc_hd__o211ai_1 _4171_ (.A1(_1502_),
    .A2(_1469_),
    .B1(_1623_),
    .C1(_1489_),
    .Y(_1624_));
 sky130_fd_sc_hd__and2_0 _4172_ (.A(_0896_),
    .B(_0899_),
    .X(_1625_));
 sky130_fd_sc_hd__nor2_1 _4173_ (.A(_0896_),
    .B(_0913_),
    .Y(_1626_));
 sky130_fd_sc_hd__clkbuf_8 _4174_ (.A(net221),
    .X(_1627_));
 sky130_fd_sc_hd__o21ai_0 _4175_ (.A1(_1625_),
    .A2(_1626_),
    .B1(_1627_),
    .Y(_1628_));
 sky130_fd_sc_hd__nand2_1 _4176_ (.A(_1624_),
    .B(_1628_),
    .Y(_1629_));
 sky130_fd_sc_hd__o32a_1 _4177_ (.A1(_1522_),
    .A2(_1622_),
    .A3(_1629_),
    .B1(_2537_),
    .B2(net115),
    .X(_1630_));
 sky130_fd_sc_hd__and3_1 _4178_ (.A(_1612_),
    .B(_1620_),
    .C(_1630_),
    .X(_0569_));
 sky130_fd_sc_hd__mux2i_1 _4179_ (.A0(\mem[5][12] ),
    .A1(\mem[7][12] ),
    .S(_1533_),
    .Y(_1631_));
 sky130_fd_sc_hd__nor2_1 _4180_ (.A(_1531_),
    .B(_1631_),
    .Y(_1632_));
 sky130_fd_sc_hd__a21oi_1 _4181_ (.A1(_0922_),
    .A2(_1527_),
    .B1(_1632_),
    .Y(_1633_));
 sky130_fd_sc_hd__mux2_1 _4182_ (.A0(\mem[1][12] ),
    .A1(\mem[3][12] ),
    .S(_1510_),
    .X(_1634_));
 sky130_fd_sc_hd__nand4_1 _4183_ (.A(_1541_),
    .B(_1543_),
    .C(_1479_),
    .D(_1634_),
    .Y(_1635_));
 sky130_fd_sc_hd__o31ai_1 _4184_ (.A1(_1538_),
    .A2(_1539_),
    .A3(_0933_),
    .B1(_1635_),
    .Y(_1636_));
 sky130_fd_sc_hd__mux2i_1 _4185_ (.A0(\mem[4][12] ),
    .A1(\mem[6][12] ),
    .S(_1550_),
    .Y(_1637_));
 sky130_fd_sc_hd__o221ai_1 _4186_ (.A1(_0923_),
    .A2(_1548_),
    .B1(_1549_),
    .B2(_1637_),
    .C1(_1552_),
    .Y(_1638_));
 sky130_fd_sc_hd__o21ai_0 _4187_ (.A1(_1537_),
    .A2(_1636_),
    .B1(_1638_),
    .Y(_1639_));
 sky130_fd_sc_hd__o22ai_1 _4188_ (.A1(\mem[1][12] ),
    .A2(_1555_),
    .B1(_1556_),
    .B2(\mem[0][12] ),
    .Y(_1640_));
 sky130_fd_sc_hd__o22ai_1 _4189_ (.A1(\mem[2][12] ),
    .A2(_1463_),
    .B1(_1465_),
    .B2(\mem[3][12] ),
    .Y(_1641_));
 sky130_fd_sc_hd__or3_1 _4190_ (.A(_1472_),
    .B(_1640_),
    .C(_1641_),
    .X(_1642_));
 sky130_fd_sc_hd__o2111ai_1 _4191_ (.A1(_1525_),
    .A2(_1633_),
    .B1(_1639_),
    .C1(_1642_),
    .D1(_1561_),
    .Y(_1643_));
 sky130_fd_sc_hd__mux2i_1 _4192_ (.A0(\mem[12][12] ),
    .A1(\mem[14][12] ),
    .S(_1565_),
    .Y(_1644_));
 sky130_fd_sc_hd__mux2_1 _4193_ (.A0(\mem[8][12] ),
    .A1(\mem[10][12] ),
    .S(_1480_),
    .X(_1645_));
 sky130_fd_sc_hd__nand3_1 _4194_ (.A(_1568_),
    .B(_1569_),
    .C(_1645_),
    .Y(_1646_));
 sky130_fd_sc_hd__o22ai_1 _4195_ (.A1(_1567_),
    .A2(_0936_),
    .B1(_1646_),
    .B2(_1572_),
    .Y(_1647_));
 sky130_fd_sc_hd__nor2_1 _4196_ (.A(_1574_),
    .B(_1646_),
    .Y(_1648_));
 sky130_fd_sc_hd__o21ai_0 _4197_ (.A1(net222),
    .A2(_0928_),
    .B1(_1488_),
    .Y(_1649_));
 sky130_fd_sc_hd__o22ai_1 _4198_ (.A1(_0861_),
    .A2(_1647_),
    .B1(_1648_),
    .B2(_1649_),
    .Y(_1650_));
 sky130_fd_sc_hd__o211ai_1 _4199_ (.A1(_1564_),
    .A2(_1644_),
    .B1(_1650_),
    .C1(_1578_),
    .Y(_1651_));
 sky130_fd_sc_hd__buf_6 _4200_ (.A(_0721_),
    .X(_1652_));
 sky130_fd_sc_hd__mux2i_1 _4201_ (.A0(\mem[13][12] ),
    .A1(\mem[15][12] ),
    .S(_1581_),
    .Y(_1653_));
 sky130_fd_sc_hd__buf_4 _4202_ (.A(_0827_),
    .X(_1654_));
 sky130_fd_sc_hd__nand3_1 _4203_ (.A(_1654_),
    .B(_1583_),
    .C(_0927_),
    .Y(_1655_));
 sky130_fd_sc_hd__o221ai_1 _4204_ (.A1(_0935_),
    .A2(_1495_),
    .B1(_1580_),
    .B2(_1653_),
    .C1(_1655_),
    .Y(_1656_));
 sky130_fd_sc_hd__mux2i_1 _4205_ (.A0(\mem[9][12] ),
    .A1(\mem[11][12] ),
    .S(_1608_),
    .Y(_1657_));
 sky130_fd_sc_hd__o21ai_0 _4206_ (.A1(_1589_),
    .A2(_1657_),
    .B1(_1476_),
    .Y(_1658_));
 sky130_fd_sc_hd__o22a_1 _4207_ (.A1(net116),
    .A2(_1652_),
    .B1(_1656_),
    .B2(_1658_),
    .X(_1659_));
 sky130_fd_sc_hd__and3_1 _4208_ (.A(_1643_),
    .B(_1651_),
    .C(_1659_),
    .X(_0570_));
 sky130_fd_sc_hd__mux2i_1 _4209_ (.A0(\mem[5][13] ),
    .A1(\mem[7][13] ),
    .S(_1533_),
    .Y(_1660_));
 sky130_fd_sc_hd__nor2_1 _4210_ (.A(_1531_),
    .B(_1660_),
    .Y(_1661_));
 sky130_fd_sc_hd__a21oi_1 _4211_ (.A1(_0941_),
    .A2(_1527_),
    .B1(_1661_),
    .Y(_1662_));
 sky130_fd_sc_hd__buf_4 _4212_ (.A(_1457_),
    .X(_1663_));
 sky130_fd_sc_hd__mux2_1 _4213_ (.A0(\mem[1][13] ),
    .A1(\mem[3][13] ),
    .S(_1663_),
    .X(_1664_));
 sky130_fd_sc_hd__nand4_1 _4214_ (.A(_1541_),
    .B(_1543_),
    .C(_1479_),
    .D(_1664_),
    .Y(_1665_));
 sky130_fd_sc_hd__o31ai_1 _4215_ (.A1(_1538_),
    .A2(_1539_),
    .A3(_0950_),
    .B1(_1665_),
    .Y(_1666_));
 sky130_fd_sc_hd__mux2i_1 _4216_ (.A0(\mem[4][13] ),
    .A1(\mem[6][13] ),
    .S(_1550_),
    .Y(_1667_));
 sky130_fd_sc_hd__o221ai_1 _4217_ (.A1(_0942_),
    .A2(_1548_),
    .B1(_1549_),
    .B2(_1667_),
    .C1(_1552_),
    .Y(_1668_));
 sky130_fd_sc_hd__o21ai_0 _4218_ (.A1(_1537_),
    .A2(_1666_),
    .B1(_1668_),
    .Y(_1669_));
 sky130_fd_sc_hd__clkbuf_4 _4219_ (.A(_1471_),
    .X(_1670_));
 sky130_fd_sc_hd__o22ai_1 _4220_ (.A1(\mem[1][13] ),
    .A2(_1555_),
    .B1(_1556_),
    .B2(\mem[0][13] ),
    .Y(_1671_));
 sky130_fd_sc_hd__buf_4 _4221_ (.A(_1462_),
    .X(_1672_));
 sky130_fd_sc_hd__buf_4 _4222_ (.A(_1464_),
    .X(_1673_));
 sky130_fd_sc_hd__o22ai_1 _4223_ (.A1(\mem[2][13] ),
    .A2(_1672_),
    .B1(_1673_),
    .B2(\mem[3][13] ),
    .Y(_1674_));
 sky130_fd_sc_hd__or3_1 _4224_ (.A(_1670_),
    .B(_1671_),
    .C(_1674_),
    .X(_1675_));
 sky130_fd_sc_hd__o2111ai_2 _4225_ (.A1(_1525_),
    .A2(_1662_),
    .B1(_1669_),
    .C1(_1675_),
    .D1(_1561_),
    .Y(_1676_));
 sky130_fd_sc_hd__mux2i_1 _4226_ (.A0(\mem[12][13] ),
    .A1(\mem[14][13] ),
    .S(_1565_),
    .Y(_1677_));
 sky130_fd_sc_hd__mux2_1 _4227_ (.A0(\mem[8][13] ),
    .A1(\mem[10][13] ),
    .S(_1480_),
    .X(_1678_));
 sky130_fd_sc_hd__nand3_1 _4228_ (.A(_1568_),
    .B(_1569_),
    .C(_1678_),
    .Y(_1679_));
 sky130_fd_sc_hd__o22ai_1 _4229_ (.A1(_1567_),
    .A2(_0955_),
    .B1(_1679_),
    .B2(_1572_),
    .Y(_1680_));
 sky130_fd_sc_hd__nor2_1 _4230_ (.A(_1574_),
    .B(_1679_),
    .Y(_1681_));
 sky130_fd_sc_hd__o21ai_0 _4231_ (.A1(net222),
    .A2(_0946_),
    .B1(_1488_),
    .Y(_1682_));
 sky130_fd_sc_hd__o22ai_1 _4232_ (.A1(_0861_),
    .A2(_1680_),
    .B1(_1681_),
    .B2(_1682_),
    .Y(_1683_));
 sky130_fd_sc_hd__o211ai_1 _4233_ (.A1(_1564_),
    .A2(_1677_),
    .B1(_1683_),
    .C1(_1578_),
    .Y(_1684_));
 sky130_fd_sc_hd__buf_4 _4234_ (.A(_1494_),
    .X(_1685_));
 sky130_fd_sc_hd__mux2i_1 _4235_ (.A0(\mem[13][13] ),
    .A1(\mem[15][13] ),
    .S(_1581_),
    .Y(_1686_));
 sky130_fd_sc_hd__nand3_1 _4236_ (.A(_1654_),
    .B(_1583_),
    .C(_0945_),
    .Y(_1687_));
 sky130_fd_sc_hd__o221ai_1 _4237_ (.A1(_0953_),
    .A2(_1685_),
    .B1(_1580_),
    .B2(_1686_),
    .C1(_1687_),
    .Y(_1688_));
 sky130_fd_sc_hd__mux2i_1 _4238_ (.A0(\mem[9][13] ),
    .A1(\mem[11][13] ),
    .S(_1608_),
    .Y(_1689_));
 sky130_fd_sc_hd__o21ai_0 _4239_ (.A1(_1589_),
    .A2(_1689_),
    .B1(_1476_),
    .Y(_1690_));
 sky130_fd_sc_hd__o22a_1 _4240_ (.A1(net117),
    .A2(_1652_),
    .B1(_1688_),
    .B2(_1690_),
    .X(_1691_));
 sky130_fd_sc_hd__and3_1 _4241_ (.A(_1676_),
    .B(_1684_),
    .C(_1691_),
    .X(_0571_));
 sky130_fd_sc_hd__buf_6 _4242_ (.A(_1532_),
    .X(_1692_));
 sky130_fd_sc_hd__mux2i_1 _4243_ (.A0(\mem[5][14] ),
    .A1(\mem[7][14] ),
    .S(_1692_),
    .Y(_1693_));
 sky130_fd_sc_hd__nor2_1 _4244_ (.A(_1531_),
    .B(_1693_),
    .Y(_1694_));
 sky130_fd_sc_hd__a21oi_1 _4245_ (.A1(_0960_),
    .A2(_1527_),
    .B1(_1694_),
    .Y(_1695_));
 sky130_fd_sc_hd__mux2_1 _4246_ (.A0(\mem[1][14] ),
    .A1(\mem[3][14] ),
    .S(_1663_),
    .X(_1696_));
 sky130_fd_sc_hd__nand4_1 _4247_ (.A(_1541_),
    .B(_1543_),
    .C(_1479_),
    .D(_1696_),
    .Y(_1697_));
 sky130_fd_sc_hd__o31ai_1 _4248_ (.A1(_1538_),
    .A2(_1539_),
    .A3(_0969_),
    .B1(_1697_),
    .Y(_1698_));
 sky130_fd_sc_hd__buf_6 _4249_ (.A(_1510_),
    .X(_1699_));
 sky130_fd_sc_hd__mux2i_1 _4250_ (.A0(\mem[4][14] ),
    .A1(\mem[6][14] ),
    .S(_1699_),
    .Y(_1700_));
 sky130_fd_sc_hd__o221ai_1 _4251_ (.A1(_0961_),
    .A2(_1548_),
    .B1(_1549_),
    .B2(_1700_),
    .C1(_1552_),
    .Y(_1701_));
 sky130_fd_sc_hd__o21ai_0 _4252_ (.A1(_1537_),
    .A2(_1698_),
    .B1(_1701_),
    .Y(_1702_));
 sky130_fd_sc_hd__o22ai_1 _4253_ (.A1(\mem[1][14] ),
    .A2(_1555_),
    .B1(_1556_),
    .B2(\mem[0][14] ),
    .Y(_1703_));
 sky130_fd_sc_hd__o22ai_1 _4254_ (.A1(\mem[2][14] ),
    .A2(_1672_),
    .B1(_1673_),
    .B2(\mem[3][14] ),
    .Y(_1704_));
 sky130_fd_sc_hd__or3_1 _4255_ (.A(_1670_),
    .B(_1703_),
    .C(_1704_),
    .X(_1705_));
 sky130_fd_sc_hd__o2111ai_2 _4256_ (.A1(_1525_),
    .A2(_1695_),
    .B1(_1702_),
    .C1(_1705_),
    .D1(_1561_),
    .Y(_1706_));
 sky130_fd_sc_hd__mux2i_1 _4257_ (.A0(\mem[12][14] ),
    .A1(\mem[14][14] ),
    .S(_1565_),
    .Y(_1707_));
 sky130_fd_sc_hd__buf_6 _4258_ (.A(_0715_),
    .X(_1708_));
 sky130_fd_sc_hd__clkbuf_8 _4259_ (.A(_1457_),
    .X(_1709_));
 sky130_fd_sc_hd__mux2_1 _4260_ (.A0(\mem[8][14] ),
    .A1(\mem[10][14] ),
    .S(_1709_),
    .X(_1710_));
 sky130_fd_sc_hd__nand3_1 _4261_ (.A(_1568_),
    .B(_1569_),
    .C(_1710_),
    .Y(_1711_));
 sky130_fd_sc_hd__o22ai_1 _4262_ (.A1(_1708_),
    .A2(_0972_),
    .B1(_1711_),
    .B2(_1572_),
    .Y(_1712_));
 sky130_fd_sc_hd__nor2_1 _4263_ (.A(_1574_),
    .B(_1711_),
    .Y(_1713_));
 sky130_fd_sc_hd__o21ai_0 _4264_ (.A1(net222),
    .A2(_0965_),
    .B1(_1488_),
    .Y(_1714_));
 sky130_fd_sc_hd__o22ai_1 _4265_ (.A1(_0861_),
    .A2(_1712_),
    .B1(_1713_),
    .B2(_1714_),
    .Y(_1715_));
 sky130_fd_sc_hd__o211ai_1 _4266_ (.A1(_1564_),
    .A2(_1707_),
    .B1(_1715_),
    .C1(_1578_),
    .Y(_1716_));
 sky130_fd_sc_hd__mux2i_1 _4267_ (.A0(\mem[13][14] ),
    .A1(\mem[15][14] ),
    .S(_1581_),
    .Y(_1717_));
 sky130_fd_sc_hd__nand3_1 _4268_ (.A(_1654_),
    .B(_1583_),
    .C(_0964_),
    .Y(_1718_));
 sky130_fd_sc_hd__o221ai_1 _4269_ (.A1(_0971_),
    .A2(_1685_),
    .B1(_1580_),
    .B2(_1717_),
    .C1(_1718_),
    .Y(_1719_));
 sky130_fd_sc_hd__mux2i_1 _4270_ (.A0(\mem[9][14] ),
    .A1(\mem[11][14] ),
    .S(_1608_),
    .Y(_1720_));
 sky130_fd_sc_hd__o21ai_0 _4271_ (.A1(_1589_),
    .A2(_1720_),
    .B1(_1476_),
    .Y(_1721_));
 sky130_fd_sc_hd__o22a_1 _4272_ (.A1(net118),
    .A2(_1652_),
    .B1(_1719_),
    .B2(_1721_),
    .X(_1722_));
 sky130_fd_sc_hd__and3_1 _4273_ (.A(_1706_),
    .B(_1716_),
    .C(_1722_),
    .X(_0572_));
 sky130_fd_sc_hd__mux2i_1 _4274_ (.A0(\mem[13][15] ),
    .A1(\mem[15][15] ),
    .S(_1599_),
    .Y(_1723_));
 sky130_fd_sc_hd__o22ai_1 _4275_ (.A1(_0991_),
    .A2(_1597_),
    .B1(_1598_),
    .B2(_1723_),
    .Y(_1724_));
 sky130_fd_sc_hd__a211oi_1 _4276_ (.A1(_1595_),
    .A2(_1724_),
    .B1(_1593_),
    .C1(_2534_),
    .Y(_1725_));
 sky130_fd_sc_hd__buf_4 _4277_ (.A(_1588_),
    .X(_1726_));
 sky130_fd_sc_hd__buf_6 _4278_ (.A(_1481_),
    .X(_1727_));
 sky130_fd_sc_hd__mux2i_1 _4279_ (.A0(\mem[9][15] ),
    .A1(\mem[11][15] ),
    .S(_1727_),
    .Y(_1728_));
 sky130_fd_sc_hd__o221ai_1 _4280_ (.A1(_0982_),
    .A2(_1495_),
    .B1(_1726_),
    .B2(_1728_),
    .C1(_1595_),
    .Y(_1729_));
 sky130_fd_sc_hd__mux2i_1 _4281_ (.A0(\mem[12][15] ),
    .A1(\mem[14][15] ),
    .S(_1533_),
    .Y(_1730_));
 sky130_fd_sc_hd__buf_6 _4282_ (.A(_0850_),
    .X(_1731_));
 sky130_fd_sc_hd__o221ai_1 _4283_ (.A1(_0990_),
    .A2(_1597_),
    .B1(_1598_),
    .B2(_1730_),
    .C1(_1731_),
    .Y(_1732_));
 sky130_fd_sc_hd__o22ai_1 _4284_ (.A1(\mem[10][15] ),
    .A2(_1463_),
    .B1(_1465_),
    .B2(\mem[11][15] ),
    .Y(_1733_));
 sky130_fd_sc_hd__o22ai_1 _4285_ (.A1(\mem[9][15] ),
    .A2(_1456_),
    .B1(_1460_),
    .B2(\mem[8][15] ),
    .Y(_1734_));
 sky130_fd_sc_hd__nor3_1 _4286_ (.A(_1472_),
    .B(_1733_),
    .C(_1734_),
    .Y(_1735_));
 sky130_fd_sc_hd__a21oi_1 _4287_ (.A1(_1729_),
    .A2(_1732_),
    .B1(_1735_),
    .Y(_1736_));
 sky130_fd_sc_hd__buf_6 _4288_ (.A(_1580_),
    .X(_1737_));
 sky130_fd_sc_hd__clkbuf_16 _4289_ (.A(_1581_),
    .X(_1738_));
 sky130_fd_sc_hd__mux2i_1 _4290_ (.A0(\mem[4][15] ),
    .A1(\mem[6][15] ),
    .S(_1738_),
    .Y(_1739_));
 sky130_fd_sc_hd__buf_4 _4291_ (.A(_0715_),
    .X(_1740_));
 sky130_fd_sc_hd__mux2_1 _4292_ (.A0(\mem[0][15] ),
    .A1(\mem[2][15] ),
    .S(_1483_),
    .X(_1741_));
 sky130_fd_sc_hd__nand3_1 _4293_ (.A(_1540_),
    .B(_1542_),
    .C(_1741_),
    .Y(_1742_));
 sky130_fd_sc_hd__buf_6 _4294_ (.A(_1467_),
    .X(_1743_));
 sky130_fd_sc_hd__o22ai_1 _4295_ (.A1(_1740_),
    .A2(_0979_),
    .B1(_1742_),
    .B2(_1743_),
    .Y(_1744_));
 sky130_fd_sc_hd__buf_6 _4296_ (.A(_1468_),
    .X(_1745_));
 sky130_fd_sc_hd__nor2_1 _4297_ (.A(_1745_),
    .B(_1742_),
    .Y(_1746_));
 sky130_fd_sc_hd__o21ai_0 _4298_ (.A1(_1567_),
    .A2(_0988_),
    .B1(_0828_),
    .Y(_1747_));
 sky130_fd_sc_hd__o22ai_1 _4299_ (.A1(_1514_),
    .A2(_1744_),
    .B1(_1746_),
    .B2(_1747_),
    .Y(_1748_));
 sky130_fd_sc_hd__o211a_1 _4300_ (.A1(_1737_),
    .A2(_1739_),
    .B1(_1748_),
    .C1(_1509_),
    .X(_1749_));
 sky130_fd_sc_hd__mux2i_1 _4301_ (.A0(\mem[5][15] ),
    .A1(\mem[7][15] ),
    .S(_1532_),
    .Y(_1750_));
 sky130_fd_sc_hd__nor2_1 _4302_ (.A(_1530_),
    .B(_1750_),
    .Y(_1751_));
 sky130_fd_sc_hd__clkbuf_4 _4303_ (.A(_0896_),
    .X(_1752_));
 sky130_fd_sc_hd__nor3_1 _4304_ (.A(_1752_),
    .B(_1489_),
    .C(_0989_),
    .Y(_1753_));
 sky130_fd_sc_hd__a311o_1 _4305_ (.A1(_0897_),
    .A2(_1627_),
    .A3(_0977_),
    .B1(_1751_),
    .C1(_1753_),
    .X(_1754_));
 sky130_fd_sc_hd__mux2i_1 _4306_ (.A0(\mem[1][15] ),
    .A1(\mem[3][15] ),
    .S(_1727_),
    .Y(_1755_));
 sky130_fd_sc_hd__nor2_1 _4307_ (.A(_1726_),
    .B(_1755_),
    .Y(_1756_));
 sky130_fd_sc_hd__o32ai_1 _4308_ (.A1(_1522_),
    .A2(_1754_),
    .A3(_1756_),
    .B1(_2537_),
    .B2(net119),
    .Y(_1757_));
 sky130_fd_sc_hd__a211oi_1 _4309_ (.A1(_1725_),
    .A2(_1736_),
    .B1(_1749_),
    .C1(_1757_),
    .Y(_0573_));
 sky130_fd_sc_hd__mux2i_1 _4310_ (.A0(\mem[5][16] ),
    .A1(\mem[7][16] ),
    .S(_1692_),
    .Y(_1758_));
 sky130_fd_sc_hd__nor2_1 _4311_ (.A(_1531_),
    .B(_1758_),
    .Y(_1759_));
 sky130_fd_sc_hd__a21oi_1 _4312_ (.A1(_0998_),
    .A2(_1527_),
    .B1(_1759_),
    .Y(_1760_));
 sky130_fd_sc_hd__mux2_1 _4313_ (.A0(\mem[1][16] ),
    .A1(\mem[3][16] ),
    .S(_1663_),
    .X(_1761_));
 sky130_fd_sc_hd__nand4_1 _4314_ (.A(_1541_),
    .B(_1543_),
    .C(_1479_),
    .D(_1761_),
    .Y(_1762_));
 sky130_fd_sc_hd__o31ai_1 _4315_ (.A1(_1538_),
    .A2(_1539_),
    .A3(_1008_),
    .B1(_1762_),
    .Y(_1763_));
 sky130_fd_sc_hd__mux2i_1 _4316_ (.A0(\mem[4][16] ),
    .A1(\mem[6][16] ),
    .S(_1699_),
    .Y(_1764_));
 sky130_fd_sc_hd__o221ai_1 _4317_ (.A1(_0999_),
    .A2(_1548_),
    .B1(_1549_),
    .B2(_1764_),
    .C1(_1552_),
    .Y(_1765_));
 sky130_fd_sc_hd__o21ai_0 _4318_ (.A1(_1537_),
    .A2(_1763_),
    .B1(_1765_),
    .Y(_1766_));
 sky130_fd_sc_hd__buf_6 _4319_ (.A(_1462_),
    .X(_1767_));
 sky130_fd_sc_hd__buf_6 _4320_ (.A(_1464_),
    .X(_1768_));
 sky130_fd_sc_hd__o22ai_1 _4321_ (.A1(\mem[2][16] ),
    .A2(_1767_),
    .B1(_1768_),
    .B2(\mem[3][16] ),
    .Y(_1769_));
 sky130_fd_sc_hd__o22ai_1 _4322_ (.A1(\mem[1][16] ),
    .A2(_1456_),
    .B1(_1460_),
    .B2(\mem[0][16] ),
    .Y(_1770_));
 sky130_fd_sc_hd__or3_1 _4323_ (.A(_1670_),
    .B(_1769_),
    .C(_1770_),
    .X(_1771_));
 sky130_fd_sc_hd__o2111ai_1 _4324_ (.A1(_1525_),
    .A2(_1760_),
    .B1(_1766_),
    .C1(_1771_),
    .D1(_1561_),
    .Y(_1772_));
 sky130_fd_sc_hd__mux2i_1 _4325_ (.A0(\mem[12][16] ),
    .A1(\mem[14][16] ),
    .S(_1565_),
    .Y(_1773_));
 sky130_fd_sc_hd__mux2_1 _4326_ (.A0(\mem[8][16] ),
    .A1(\mem[10][16] ),
    .S(_1709_),
    .X(_1774_));
 sky130_fd_sc_hd__nand3_1 _4327_ (.A(_1568_),
    .B(_1569_),
    .C(_1774_),
    .Y(_1775_));
 sky130_fd_sc_hd__o22ai_1 _4328_ (.A1(_1708_),
    .A2(_1011_),
    .B1(_1775_),
    .B2(_1572_),
    .Y(_1776_));
 sky130_fd_sc_hd__nor2_1 _4329_ (.A(_1574_),
    .B(_1775_),
    .Y(_1777_));
 sky130_fd_sc_hd__buf_4 _4330_ (.A(_0827_),
    .X(_1778_));
 sky130_fd_sc_hd__o21ai_0 _4331_ (.A1(net222),
    .A2(_1004_),
    .B1(_1778_),
    .Y(_1779_));
 sky130_fd_sc_hd__o22ai_1 _4332_ (.A1(_0861_),
    .A2(_1776_),
    .B1(_1777_),
    .B2(_1779_),
    .Y(_1780_));
 sky130_fd_sc_hd__o211ai_1 _4333_ (.A1(_1564_),
    .A2(_1773_),
    .B1(_1780_),
    .C1(_1578_),
    .Y(_1781_));
 sky130_fd_sc_hd__clkbuf_8 _4334_ (.A(_1529_),
    .X(_1782_));
 sky130_fd_sc_hd__mux2i_1 _4335_ (.A0(\mem[13][16] ),
    .A1(\mem[15][16] ),
    .S(_1581_),
    .Y(_1783_));
 sky130_fd_sc_hd__nand3_1 _4336_ (.A(_1654_),
    .B(_1583_),
    .C(_1003_),
    .Y(_1784_));
 sky130_fd_sc_hd__o221ai_1 _4337_ (.A1(_1010_),
    .A2(_1685_),
    .B1(_1782_),
    .B2(_1783_),
    .C1(_1784_),
    .Y(_1785_));
 sky130_fd_sc_hd__mux2i_1 _4338_ (.A0(\mem[9][16] ),
    .A1(\mem[11][16] ),
    .S(_1608_),
    .Y(_1786_));
 sky130_fd_sc_hd__o21ai_0 _4339_ (.A1(_1589_),
    .A2(_1786_),
    .B1(_1476_),
    .Y(_1787_));
 sky130_fd_sc_hd__o22a_1 _4340_ (.A1(net120),
    .A2(_1652_),
    .B1(_1785_),
    .B2(_1787_),
    .X(_1788_));
 sky130_fd_sc_hd__and3_1 _4341_ (.A(_1772_),
    .B(_1781_),
    .C(_1788_),
    .X(_0574_));
 sky130_fd_sc_hd__mux2i_1 _4342_ (.A0(\mem[5][17] ),
    .A1(\mem[7][17] ),
    .S(_1692_),
    .Y(_1789_));
 sky130_fd_sc_hd__nor2_1 _4343_ (.A(_1531_),
    .B(_1789_),
    .Y(_1790_));
 sky130_fd_sc_hd__a21oi_1 _4344_ (.A1(_1017_),
    .A2(_1527_),
    .B1(_1790_),
    .Y(_1791_));
 sky130_fd_sc_hd__mux2_1 _4345_ (.A0(\mem[1][17] ),
    .A1(\mem[3][17] ),
    .S(_1663_),
    .X(_1792_));
 sky130_fd_sc_hd__nand4_1 _4346_ (.A(_1541_),
    .B(_1543_),
    .C(_1479_),
    .D(_1792_),
    .Y(_1793_));
 sky130_fd_sc_hd__o31ai_1 _4347_ (.A1(_1538_),
    .A2(_1539_),
    .A3(_1027_),
    .B1(_1793_),
    .Y(_1794_));
 sky130_fd_sc_hd__mux2i_1 _4348_ (.A0(\mem[4][17] ),
    .A1(\mem[6][17] ),
    .S(_1699_),
    .Y(_1795_));
 sky130_fd_sc_hd__buf_4 _4349_ (.A(_0854_),
    .X(_1796_));
 sky130_fd_sc_hd__o221ai_1 _4350_ (.A1(_1018_),
    .A2(_1548_),
    .B1(_1549_),
    .B2(_1795_),
    .C1(_1796_),
    .Y(_1797_));
 sky130_fd_sc_hd__o21ai_0 _4351_ (.A1(_1537_),
    .A2(_1794_),
    .B1(_1797_),
    .Y(_1798_));
 sky130_fd_sc_hd__o22ai_1 _4352_ (.A1(\mem[1][17] ),
    .A2(_1555_),
    .B1(_1556_),
    .B2(\mem[0][17] ),
    .Y(_1799_));
 sky130_fd_sc_hd__o22ai_1 _4353_ (.A1(\mem[2][17] ),
    .A2(_1672_),
    .B1(_1673_),
    .B2(\mem[3][17] ),
    .Y(_1800_));
 sky130_fd_sc_hd__or3_1 _4354_ (.A(_1670_),
    .B(_1799_),
    .C(_1800_),
    .X(_1801_));
 sky130_fd_sc_hd__o2111ai_1 _4355_ (.A1(_1525_),
    .A2(_1791_),
    .B1(_1798_),
    .C1(_1801_),
    .D1(_1561_),
    .Y(_1802_));
 sky130_fd_sc_hd__mux2i_1 _4356_ (.A0(\mem[12][17] ),
    .A1(\mem[14][17] ),
    .S(_1565_),
    .Y(_1803_));
 sky130_fd_sc_hd__buf_4 _4357_ (.A(_1540_),
    .X(_1804_));
 sky130_fd_sc_hd__clkbuf_8 _4358_ (.A(_1542_),
    .X(_1805_));
 sky130_fd_sc_hd__mux2_1 _4359_ (.A0(\mem[8][17] ),
    .A1(\mem[10][17] ),
    .S(_1709_),
    .X(_1806_));
 sky130_fd_sc_hd__nand3_1 _4360_ (.A(_1804_),
    .B(_1805_),
    .C(_1806_),
    .Y(_1807_));
 sky130_fd_sc_hd__o22ai_1 _4361_ (.A1(_1708_),
    .A2(_1030_),
    .B1(_1807_),
    .B2(_1572_),
    .Y(_1808_));
 sky130_fd_sc_hd__nor2_1 _4362_ (.A(_1574_),
    .B(_1807_),
    .Y(_1809_));
 sky130_fd_sc_hd__buf_6 _4363_ (.A(_0715_),
    .X(_1810_));
 sky130_fd_sc_hd__o21ai_0 _4364_ (.A1(_1810_),
    .A2(_1022_),
    .B1(_1778_),
    .Y(_1811_));
 sky130_fd_sc_hd__o22ai_1 _4365_ (.A1(_0861_),
    .A2(_1808_),
    .B1(_1809_),
    .B2(_1811_),
    .Y(_1812_));
 sky130_fd_sc_hd__o211ai_1 _4366_ (.A1(_1564_),
    .A2(_1803_),
    .B1(_1812_),
    .C1(_1578_),
    .Y(_1813_));
 sky130_fd_sc_hd__mux2i_1 _4367_ (.A0(\mem[13][17] ),
    .A1(\mem[15][17] ),
    .S(_1581_),
    .Y(_1814_));
 sky130_fd_sc_hd__nand3_1 _4368_ (.A(_1654_),
    .B(_1583_),
    .C(_1021_),
    .Y(_1815_));
 sky130_fd_sc_hd__o221ai_1 _4369_ (.A1(_1029_),
    .A2(_1685_),
    .B1(_1782_),
    .B2(_1814_),
    .C1(_1815_),
    .Y(_1816_));
 sky130_fd_sc_hd__mux2i_1 _4370_ (.A0(\mem[9][17] ),
    .A1(\mem[11][17] ),
    .S(_1608_),
    .Y(_1817_));
 sky130_fd_sc_hd__o21ai_0 _4371_ (.A1(_1589_),
    .A2(_1817_),
    .B1(_1476_),
    .Y(_1818_));
 sky130_fd_sc_hd__o22a_1 _4372_ (.A1(net121),
    .A2(_1652_),
    .B1(_1816_),
    .B2(_1818_),
    .X(_1819_));
 sky130_fd_sc_hd__and3_1 _4373_ (.A(_1802_),
    .B(_1813_),
    .C(_1819_),
    .X(_0575_));
 sky130_fd_sc_hd__buf_4 _4374_ (.A(_1530_),
    .X(_1820_));
 sky130_fd_sc_hd__mux2i_1 _4375_ (.A0(\mem[5][18] ),
    .A1(\mem[7][18] ),
    .S(_1692_),
    .Y(_1821_));
 sky130_fd_sc_hd__nor2_1 _4376_ (.A(_1820_),
    .B(_1821_),
    .Y(_1822_));
 sky130_fd_sc_hd__a21oi_1 _4377_ (.A1(_1036_),
    .A2(_1527_),
    .B1(_1822_),
    .Y(_1823_));
 sky130_fd_sc_hd__mux2_1 _4378_ (.A0(\mem[1][18] ),
    .A1(\mem[3][18] ),
    .S(_1663_),
    .X(_1824_));
 sky130_fd_sc_hd__nand4_1 _4379_ (.A(_1541_),
    .B(_1543_),
    .C(_1479_),
    .D(_1824_),
    .Y(_1825_));
 sky130_fd_sc_hd__o31ai_1 _4380_ (.A1(_1538_),
    .A2(_1539_),
    .A3(_1046_),
    .B1(_1825_),
    .Y(_1826_));
 sky130_fd_sc_hd__buf_4 _4381_ (.A(_1596_),
    .X(_1827_));
 sky130_fd_sc_hd__mux2i_1 _4382_ (.A0(\mem[4][18] ),
    .A1(\mem[6][18] ),
    .S(_1699_),
    .Y(_1828_));
 sky130_fd_sc_hd__o221ai_1 _4383_ (.A1(_1037_),
    .A2(_1827_),
    .B1(_1549_),
    .B2(_1828_),
    .C1(_1796_),
    .Y(_1829_));
 sky130_fd_sc_hd__o21ai_0 _4384_ (.A1(_1537_),
    .A2(_1826_),
    .B1(_1829_),
    .Y(_1830_));
 sky130_fd_sc_hd__o22ai_1 _4385_ (.A1(\mem[1][18] ),
    .A2(_1555_),
    .B1(_1556_),
    .B2(\mem[0][18] ),
    .Y(_1831_));
 sky130_fd_sc_hd__o22ai_1 _4386_ (.A1(\mem[2][18] ),
    .A2(_1672_),
    .B1(_1673_),
    .B2(\mem[3][18] ),
    .Y(_1832_));
 sky130_fd_sc_hd__or3_1 _4387_ (.A(_1670_),
    .B(_1831_),
    .C(_1832_),
    .X(_1833_));
 sky130_fd_sc_hd__o2111ai_1 _4388_ (.A1(_1525_),
    .A2(_1823_),
    .B1(_1830_),
    .C1(_1833_),
    .D1(_1561_),
    .Y(_1834_));
 sky130_fd_sc_hd__mux2i_1 _4389_ (.A0(\mem[12][18] ),
    .A1(\mem[14][18] ),
    .S(_1565_),
    .Y(_1835_));
 sky130_fd_sc_hd__mux2_1 _4390_ (.A0(\mem[8][18] ),
    .A1(\mem[10][18] ),
    .S(_1709_),
    .X(_1836_));
 sky130_fd_sc_hd__nand3_1 _4391_ (.A(_1804_),
    .B(_1805_),
    .C(_1836_),
    .Y(_1837_));
 sky130_fd_sc_hd__o22ai_1 _4392_ (.A1(_1708_),
    .A2(_1049_),
    .B1(_1837_),
    .B2(_1572_),
    .Y(_1838_));
 sky130_fd_sc_hd__nor2_1 _4393_ (.A(_1574_),
    .B(_1837_),
    .Y(_1839_));
 sky130_fd_sc_hd__o21ai_0 _4394_ (.A1(_1810_),
    .A2(_1042_),
    .B1(_1778_),
    .Y(_1840_));
 sky130_fd_sc_hd__o22ai_1 _4395_ (.A1(_0861_),
    .A2(_1838_),
    .B1(_1839_),
    .B2(_1840_),
    .Y(_1841_));
 sky130_fd_sc_hd__o211ai_1 _4396_ (.A1(_1564_),
    .A2(_1835_),
    .B1(_1841_),
    .C1(_1578_),
    .Y(_1842_));
 sky130_fd_sc_hd__mux2i_1 _4397_ (.A0(\mem[13][18] ),
    .A1(\mem[15][18] ),
    .S(_1581_),
    .Y(_1843_));
 sky130_fd_sc_hd__nand3_1 _4398_ (.A(_1654_),
    .B(_1583_),
    .C(_1040_),
    .Y(_1844_));
 sky130_fd_sc_hd__o221ai_1 _4399_ (.A1(_1048_),
    .A2(_1685_),
    .B1(_1782_),
    .B2(_1843_),
    .C1(_1844_),
    .Y(_1845_));
 sky130_fd_sc_hd__mux2i_1 _4400_ (.A0(\mem[9][18] ),
    .A1(\mem[11][18] ),
    .S(_1608_),
    .Y(_1846_));
 sky130_fd_sc_hd__o21ai_0 _4401_ (.A1(_1589_),
    .A2(_1846_),
    .B1(_1476_),
    .Y(_1847_));
 sky130_fd_sc_hd__o22a_1 _4402_ (.A1(net123),
    .A2(_1652_),
    .B1(_1845_),
    .B2(_1847_),
    .X(_1848_));
 sky130_fd_sc_hd__and3_1 _4403_ (.A(_1834_),
    .B(_1842_),
    .C(_1848_),
    .X(_0576_));
 sky130_fd_sc_hd__mux2i_1 _4404_ (.A0(\mem[5][19] ),
    .A1(\mem[7][19] ),
    .S(_1692_),
    .Y(_1849_));
 sky130_fd_sc_hd__nor2_1 _4405_ (.A(_1820_),
    .B(_1849_),
    .Y(_1850_));
 sky130_fd_sc_hd__a21oi_1 _4406_ (.A1(_1055_),
    .A2(_1527_),
    .B1(_1850_),
    .Y(_1851_));
 sky130_fd_sc_hd__buf_4 _4407_ (.A(_0827_),
    .X(_1852_));
 sky130_fd_sc_hd__mux2_1 _4408_ (.A0(\mem[1][19] ),
    .A1(\mem[3][19] ),
    .S(_1663_),
    .X(_1853_));
 sky130_fd_sc_hd__nand4_1 _4409_ (.A(_1541_),
    .B(_1543_),
    .C(_1479_),
    .D(_1853_),
    .Y(_1854_));
 sky130_fd_sc_hd__o31ai_1 _4410_ (.A1(_1852_),
    .A2(_1539_),
    .A3(_1064_),
    .B1(_1854_),
    .Y(_1855_));
 sky130_fd_sc_hd__mux2i_1 _4411_ (.A0(\mem[4][19] ),
    .A1(\mem[6][19] ),
    .S(_1699_),
    .Y(_1856_));
 sky130_fd_sc_hd__o221ai_1 _4412_ (.A1(_1056_),
    .A2(_1827_),
    .B1(_1549_),
    .B2(_1856_),
    .C1(_1796_),
    .Y(_1857_));
 sky130_fd_sc_hd__o21ai_0 _4413_ (.A1(_1537_),
    .A2(_1855_),
    .B1(_1857_),
    .Y(_1858_));
 sky130_fd_sc_hd__o22ai_1 _4414_ (.A1(\mem[1][19] ),
    .A2(_1555_),
    .B1(_1556_),
    .B2(\mem[0][19] ),
    .Y(_1859_));
 sky130_fd_sc_hd__o22ai_1 _4415_ (.A1(\mem[2][19] ),
    .A2(_1672_),
    .B1(_1673_),
    .B2(\mem[3][19] ),
    .Y(_1860_));
 sky130_fd_sc_hd__or3_1 _4416_ (.A(_1670_),
    .B(_1859_),
    .C(_1860_),
    .X(_1861_));
 sky130_fd_sc_hd__o2111ai_1 _4417_ (.A1(_1525_),
    .A2(_1851_),
    .B1(_1858_),
    .C1(_1861_),
    .D1(_1561_),
    .Y(_1862_));
 sky130_fd_sc_hd__mux2i_1 _4418_ (.A0(\mem[12][19] ),
    .A1(\mem[14][19] ),
    .S(_1565_),
    .Y(_1863_));
 sky130_fd_sc_hd__buf_6 _4419_ (.A(_0860_),
    .X(_1864_));
 sky130_fd_sc_hd__mux2_1 _4420_ (.A0(\mem[8][19] ),
    .A1(\mem[10][19] ),
    .S(_1709_),
    .X(_1865_));
 sky130_fd_sc_hd__nand3_1 _4421_ (.A(_1804_),
    .B(_1805_),
    .C(_1865_),
    .Y(_1866_));
 sky130_fd_sc_hd__o22ai_1 _4422_ (.A1(_1708_),
    .A2(_1067_),
    .B1(_1866_),
    .B2(_1572_),
    .Y(_1867_));
 sky130_fd_sc_hd__nor2_1 _4423_ (.A(_1574_),
    .B(_1866_),
    .Y(_1868_));
 sky130_fd_sc_hd__o21ai_0 _4424_ (.A1(_1810_),
    .A2(_1060_),
    .B1(_1778_),
    .Y(_1869_));
 sky130_fd_sc_hd__o22ai_1 _4425_ (.A1(_1864_),
    .A2(_1867_),
    .B1(_1868_),
    .B2(_1869_),
    .Y(_1870_));
 sky130_fd_sc_hd__o211ai_1 _4426_ (.A1(_1564_),
    .A2(_1863_),
    .B1(_1870_),
    .C1(_1578_),
    .Y(_1871_));
 sky130_fd_sc_hd__buf_8 _4427_ (.A(_1510_),
    .X(_1872_));
 sky130_fd_sc_hd__mux2i_1 _4428_ (.A0(\mem[13][19] ),
    .A1(\mem[15][19] ),
    .S(_1872_),
    .Y(_1873_));
 sky130_fd_sc_hd__nand3_1 _4429_ (.A(_1654_),
    .B(_1583_),
    .C(_1059_),
    .Y(_1874_));
 sky130_fd_sc_hd__o221ai_1 _4430_ (.A1(_1066_),
    .A2(_1685_),
    .B1(_1782_),
    .B2(_1873_),
    .C1(_1874_),
    .Y(_1875_));
 sky130_fd_sc_hd__buf_6 _4431_ (.A(_1587_),
    .X(_1876_));
 sky130_fd_sc_hd__mux2i_1 _4432_ (.A0(\mem[9][19] ),
    .A1(\mem[11][19] ),
    .S(_1608_),
    .Y(_1877_));
 sky130_fd_sc_hd__o21ai_0 _4433_ (.A1(_1876_),
    .A2(_1877_),
    .B1(_1476_),
    .Y(_1878_));
 sky130_fd_sc_hd__o22a_1 _4434_ (.A1(net124),
    .A2(_1652_),
    .B1(_1875_),
    .B2(_1878_),
    .X(_1879_));
 sky130_fd_sc_hd__and3_1 _4435_ (.A(_1862_),
    .B(_1871_),
    .C(_1879_),
    .X(_0577_));
 sky130_fd_sc_hd__mux2i_1 _4436_ (.A0(\mem[13][1] ),
    .A1(\mem[15][1] ),
    .S(_1599_),
    .Y(_1880_));
 sky130_fd_sc_hd__o22ai_1 _4437_ (.A1(_1086_),
    .A2(_1597_),
    .B1(_1598_),
    .B2(_1880_),
    .Y(_1881_));
 sky130_fd_sc_hd__a211oi_1 _4438_ (.A1(_1595_),
    .A2(_1881_),
    .B1(_1593_),
    .C1(net163),
    .Y(_1882_));
 sky130_fd_sc_hd__mux2i_1 _4439_ (.A0(\mem[9][1] ),
    .A1(\mem[11][1] ),
    .S(_1727_),
    .Y(_1883_));
 sky130_fd_sc_hd__o221ai_1 _4440_ (.A1(_1077_),
    .A2(_1495_),
    .B1(_1726_),
    .B2(_1883_),
    .C1(_1595_),
    .Y(_1884_));
 sky130_fd_sc_hd__mux2i_1 _4441_ (.A0(\mem[12][1] ),
    .A1(\mem[14][1] ),
    .S(_1533_),
    .Y(_1885_));
 sky130_fd_sc_hd__o221ai_1 _4442_ (.A1(_1085_),
    .A2(_1597_),
    .B1(_1598_),
    .B2(_1885_),
    .C1(_1731_),
    .Y(_1886_));
 sky130_fd_sc_hd__o22ai_1 _4443_ (.A1(\mem[10][1] ),
    .A2(_1463_),
    .B1(_1465_),
    .B2(\mem[11][1] ),
    .Y(_1887_));
 sky130_fd_sc_hd__o22ai_1 _4444_ (.A1(\mem[9][1] ),
    .A2(_1456_),
    .B1(_1460_),
    .B2(\mem[8][1] ),
    .Y(_1888_));
 sky130_fd_sc_hd__nor3_1 _4445_ (.A(_1472_),
    .B(_1887_),
    .C(_1888_),
    .Y(_1889_));
 sky130_fd_sc_hd__a21oi_1 _4446_ (.A1(_1884_),
    .A2(_1886_),
    .B1(_1889_),
    .Y(_1890_));
 sky130_fd_sc_hd__mux2i_1 _4447_ (.A0(\mem[4][1] ),
    .A1(\mem[6][1] ),
    .S(_1738_),
    .Y(_1891_));
 sky130_fd_sc_hd__mux2_1 _4448_ (.A0(\mem[0][1] ),
    .A1(\mem[2][1] ),
    .S(_1483_),
    .X(_1892_));
 sky130_fd_sc_hd__nand3_1 _4449_ (.A(_1540_),
    .B(_1542_),
    .C(_1892_),
    .Y(_1893_));
 sky130_fd_sc_hd__o22ai_1 _4450_ (.A1(_1740_),
    .A2(_1074_),
    .B1(_1893_),
    .B2(_1743_),
    .Y(_1894_));
 sky130_fd_sc_hd__nor2_1 _4451_ (.A(_1745_),
    .B(_1893_),
    .Y(_1895_));
 sky130_fd_sc_hd__o21ai_0 _4452_ (.A1(_1567_),
    .A2(_1083_),
    .B1(_0828_),
    .Y(_1896_));
 sky130_fd_sc_hd__o22ai_1 _4453_ (.A1(_1514_),
    .A2(_1894_),
    .B1(_1895_),
    .B2(_1896_),
    .Y(_1897_));
 sky130_fd_sc_hd__o211a_1 _4454_ (.A1(_1737_),
    .A2(_1891_),
    .B1(_1897_),
    .C1(_1509_),
    .X(_1898_));
 sky130_fd_sc_hd__mux2i_1 _4455_ (.A0(\mem[5][1] ),
    .A1(\mem[7][1] ),
    .S(_1532_),
    .Y(_1899_));
 sky130_fd_sc_hd__nor2_1 _4456_ (.A(_1530_),
    .B(_1899_),
    .Y(_1900_));
 sky130_fd_sc_hd__nor3_1 _4457_ (.A(_1752_),
    .B(_1489_),
    .C(_1084_),
    .Y(_1901_));
 sky130_fd_sc_hd__a311o_1 _4458_ (.A1(_1752_),
    .A2(_1627_),
    .A3(_1073_),
    .B1(_1900_),
    .C1(_1901_),
    .X(_1902_));
 sky130_fd_sc_hd__mux2i_1 _4459_ (.A0(\mem[1][1] ),
    .A1(\mem[3][1] ),
    .S(_1727_),
    .Y(_1903_));
 sky130_fd_sc_hd__nor2_1 _4460_ (.A(_1726_),
    .B(_1903_),
    .Y(_1904_));
 sky130_fd_sc_hd__o32ai_1 _4461_ (.A1(_1522_),
    .A2(_1902_),
    .A3(_1904_),
    .B1(_2537_),
    .B2(net104),
    .Y(_1905_));
 sky130_fd_sc_hd__a211oi_1 _4462_ (.A1(_1882_),
    .A2(_1890_),
    .B1(_1898_),
    .C1(_1905_),
    .Y(_0578_));
 sky130_fd_sc_hd__mux2i_1 _4463_ (.A0(\mem[5][20] ),
    .A1(\mem[7][20] ),
    .S(_1692_),
    .Y(_1906_));
 sky130_fd_sc_hd__nor2_1 _4464_ (.A(_1820_),
    .B(_1906_),
    .Y(_1907_));
 sky130_fd_sc_hd__a21oi_1 _4465_ (.A1(_1092_),
    .A2(_1527_),
    .B1(_1907_),
    .Y(_1908_));
 sky130_fd_sc_hd__mux2_1 _4466_ (.A0(\mem[1][20] ),
    .A1(\mem[3][20] ),
    .S(_1663_),
    .X(_1909_));
 sky130_fd_sc_hd__nand4_1 _4467_ (.A(_1541_),
    .B(_1543_),
    .C(_1479_),
    .D(_1909_),
    .Y(_1910_));
 sky130_fd_sc_hd__o31ai_1 _4468_ (.A1(_1852_),
    .A2(_1539_),
    .A3(_1102_),
    .B1(_1910_),
    .Y(_1911_));
 sky130_fd_sc_hd__mux2i_1 _4469_ (.A0(\mem[4][20] ),
    .A1(\mem[6][20] ),
    .S(_1699_),
    .Y(_1912_));
 sky130_fd_sc_hd__o221ai_1 _4470_ (.A1(_1093_),
    .A2(_1827_),
    .B1(_1549_),
    .B2(_1912_),
    .C1(_1796_),
    .Y(_1913_));
 sky130_fd_sc_hd__o21ai_0 _4471_ (.A1(_1537_),
    .A2(_1911_),
    .B1(_1913_),
    .Y(_1914_));
 sky130_fd_sc_hd__o22ai_1 _4472_ (.A1(\mem[2][20] ),
    .A2(_1767_),
    .B1(_1768_),
    .B2(\mem[3][20] ),
    .Y(_1915_));
 sky130_fd_sc_hd__o22ai_1 _4473_ (.A1(\mem[1][20] ),
    .A2(_1456_),
    .B1(_1460_),
    .B2(\mem[0][20] ),
    .Y(_1916_));
 sky130_fd_sc_hd__or3_1 _4474_ (.A(_1670_),
    .B(_1915_),
    .C(_1916_),
    .X(_1917_));
 sky130_fd_sc_hd__o2111ai_1 _4475_ (.A1(_1525_),
    .A2(_1908_),
    .B1(_1914_),
    .C1(_1917_),
    .D1(_1561_),
    .Y(_1918_));
 sky130_fd_sc_hd__mux2i_1 _4476_ (.A0(\mem[12][20] ),
    .A1(\mem[14][20] ),
    .S(_1565_),
    .Y(_1919_));
 sky130_fd_sc_hd__mux2_1 _4477_ (.A0(\mem[8][20] ),
    .A1(\mem[10][20] ),
    .S(_1709_),
    .X(_1920_));
 sky130_fd_sc_hd__nand3_1 _4478_ (.A(_1804_),
    .B(_1805_),
    .C(_1920_),
    .Y(_1921_));
 sky130_fd_sc_hd__o22ai_1 _4479_ (.A1(_1708_),
    .A2(_1105_),
    .B1(_1921_),
    .B2(_1572_),
    .Y(_1922_));
 sky130_fd_sc_hd__nor2_1 _4480_ (.A(_1574_),
    .B(_1921_),
    .Y(_1923_));
 sky130_fd_sc_hd__o21ai_0 _4481_ (.A1(_1810_),
    .A2(_1097_),
    .B1(_1778_),
    .Y(_1924_));
 sky130_fd_sc_hd__o22ai_1 _4482_ (.A1(_1864_),
    .A2(_1922_),
    .B1(_1923_),
    .B2(_1924_),
    .Y(_1925_));
 sky130_fd_sc_hd__o211ai_1 _4483_ (.A1(_1564_),
    .A2(_1919_),
    .B1(_1925_),
    .C1(_1578_),
    .Y(_1926_));
 sky130_fd_sc_hd__mux2i_1 _4484_ (.A0(\mem[13][20] ),
    .A1(\mem[15][20] ),
    .S(_1872_),
    .Y(_1927_));
 sky130_fd_sc_hd__nand3_1 _4485_ (.A(_1654_),
    .B(_1583_),
    .C(_1096_),
    .Y(_1928_));
 sky130_fd_sc_hd__o221ai_1 _4486_ (.A1(_1104_),
    .A2(_1685_),
    .B1(_1782_),
    .B2(_1927_),
    .C1(_1928_),
    .Y(_1929_));
 sky130_fd_sc_hd__mux2i_1 _4487_ (.A0(\mem[9][20] ),
    .A1(\mem[11][20] ),
    .S(_1608_),
    .Y(_1930_));
 sky130_fd_sc_hd__o21ai_0 _4488_ (.A1(_1876_),
    .A2(_1930_),
    .B1(_1476_),
    .Y(_1931_));
 sky130_fd_sc_hd__o22a_1 _4489_ (.A1(net125),
    .A2(_1652_),
    .B1(_1929_),
    .B2(_1931_),
    .X(_1932_));
 sky130_fd_sc_hd__and3_1 _4490_ (.A(_1918_),
    .B(_1926_),
    .C(_1932_),
    .X(_0579_));
 sky130_fd_sc_hd__buf_6 _4491_ (.A(_0850_),
    .X(_1933_));
 sky130_fd_sc_hd__mux2i_1 _4492_ (.A0(\mem[5][21] ),
    .A1(\mem[7][21] ),
    .S(_1692_),
    .Y(_1934_));
 sky130_fd_sc_hd__nor2_1 _4493_ (.A(_1820_),
    .B(_1934_),
    .Y(_1935_));
 sky130_fd_sc_hd__a21oi_1 _4494_ (.A1(_1110_),
    .A2(_1527_),
    .B1(_1935_),
    .Y(_1936_));
 sky130_fd_sc_hd__buf_4 _4495_ (.A(_0839_),
    .X(_1937_));
 sky130_fd_sc_hd__buf_4 _4496_ (.A(_0715_),
    .X(_1938_));
 sky130_fd_sc_hd__clkbuf_4 _4497_ (.A(_1478_),
    .X(_1939_));
 sky130_fd_sc_hd__mux2_1 _4498_ (.A0(\mem[1][21] ),
    .A1(\mem[3][21] ),
    .S(_1663_),
    .X(_1940_));
 sky130_fd_sc_hd__nand4_1 _4499_ (.A(_1541_),
    .B(_1543_),
    .C(_1939_),
    .D(_1940_),
    .Y(_1941_));
 sky130_fd_sc_hd__o31ai_1 _4500_ (.A1(_1852_),
    .A2(_1938_),
    .A3(_1120_),
    .B1(_1941_),
    .Y(_1942_));
 sky130_fd_sc_hd__buf_4 _4501_ (.A(_1529_),
    .X(_1943_));
 sky130_fd_sc_hd__mux2i_1 _4502_ (.A0(\mem[4][21] ),
    .A1(\mem[6][21] ),
    .S(_1699_),
    .Y(_1944_));
 sky130_fd_sc_hd__o221ai_1 _4503_ (.A1(_1112_),
    .A2(_1827_),
    .B1(_1943_),
    .B2(_1944_),
    .C1(_1796_),
    .Y(_1945_));
 sky130_fd_sc_hd__o21ai_0 _4504_ (.A1(_1937_),
    .A2(_1942_),
    .B1(_1945_),
    .Y(_1946_));
 sky130_fd_sc_hd__buf_4 _4505_ (.A(_1455_),
    .X(_1947_));
 sky130_fd_sc_hd__buf_4 _4506_ (.A(_1459_),
    .X(_1948_));
 sky130_fd_sc_hd__o22ai_1 _4507_ (.A1(\mem[1][21] ),
    .A2(_1947_),
    .B1(_1948_),
    .B2(\mem[0][21] ),
    .Y(_1949_));
 sky130_fd_sc_hd__o22ai_1 _4508_ (.A1(\mem[2][21] ),
    .A2(_1672_),
    .B1(_1673_),
    .B2(\mem[3][21] ),
    .Y(_1950_));
 sky130_fd_sc_hd__or3_1 _4509_ (.A(_1670_),
    .B(_1949_),
    .C(_1950_),
    .X(_1951_));
 sky130_fd_sc_hd__o2111ai_2 _4510_ (.A1(_1933_),
    .A2(_1936_),
    .B1(_1946_),
    .C1(_1951_),
    .D1(_1561_),
    .Y(_1952_));
 sky130_fd_sc_hd__clkbuf_8 _4511_ (.A(_1549_),
    .X(_1953_));
 sky130_fd_sc_hd__buf_8 _4512_ (.A(_1550_),
    .X(_1954_));
 sky130_fd_sc_hd__mux2i_1 _4513_ (.A0(\mem[12][21] ),
    .A1(\mem[14][21] ),
    .S(_1954_),
    .Y(_1955_));
 sky130_fd_sc_hd__mux2_1 _4514_ (.A0(\mem[8][21] ),
    .A1(\mem[10][21] ),
    .S(_1709_),
    .X(_1956_));
 sky130_fd_sc_hd__nand3_1 _4515_ (.A(_1804_),
    .B(_1805_),
    .C(_1956_),
    .Y(_1957_));
 sky130_fd_sc_hd__clkbuf_8 _4516_ (.A(_1467_),
    .X(_1958_));
 sky130_fd_sc_hd__o22ai_1 _4517_ (.A1(_1708_),
    .A2(_1123_),
    .B1(_1957_),
    .B2(_1958_),
    .Y(_1959_));
 sky130_fd_sc_hd__clkbuf_8 _4518_ (.A(_1468_),
    .X(_1960_));
 sky130_fd_sc_hd__nor2_1 _4519_ (.A(_1960_),
    .B(_1957_),
    .Y(_1961_));
 sky130_fd_sc_hd__o21ai_0 _4520_ (.A1(_1810_),
    .A2(_1116_),
    .B1(_1778_),
    .Y(_1962_));
 sky130_fd_sc_hd__o22ai_1 _4521_ (.A1(_1864_),
    .A2(_1959_),
    .B1(_1961_),
    .B2(_1962_),
    .Y(_1963_));
 sky130_fd_sc_hd__o211ai_1 _4522_ (.A1(_1953_),
    .A2(_1955_),
    .B1(_1963_),
    .C1(_1578_),
    .Y(_1964_));
 sky130_fd_sc_hd__mux2i_1 _4523_ (.A0(\mem[13][21] ),
    .A1(\mem[15][21] ),
    .S(_1872_),
    .Y(_1965_));
 sky130_fd_sc_hd__nand3_1 _4524_ (.A(_1654_),
    .B(_1583_),
    .C(_1115_),
    .Y(_1966_));
 sky130_fd_sc_hd__o221ai_1 _4525_ (.A1(_1122_),
    .A2(_1685_),
    .B1(_1782_),
    .B2(_1965_),
    .C1(_1966_),
    .Y(_1967_));
 sky130_fd_sc_hd__buf_6 _4526_ (.A(_1532_),
    .X(_1968_));
 sky130_fd_sc_hd__mux2i_1 _4527_ (.A0(\mem[9][21] ),
    .A1(\mem[11][21] ),
    .S(_1968_),
    .Y(_1969_));
 sky130_fd_sc_hd__buf_4 _4528_ (.A(_1475_),
    .X(_1970_));
 sky130_fd_sc_hd__o21ai_0 _4529_ (.A1(_1876_),
    .A2(_1969_),
    .B1(_1970_),
    .Y(_1971_));
 sky130_fd_sc_hd__o22a_1 _4530_ (.A1(net126),
    .A2(_1652_),
    .B1(_1967_),
    .B2(_1971_),
    .X(_1972_));
 sky130_fd_sc_hd__and3_1 _4531_ (.A(_1952_),
    .B(_1964_),
    .C(_1972_),
    .X(_0580_));
 sky130_fd_sc_hd__buf_4 _4532_ (.A(_1526_),
    .X(_1973_));
 sky130_fd_sc_hd__mux2i_1 _4533_ (.A0(\mem[5][22] ),
    .A1(\mem[7][22] ),
    .S(_1692_),
    .Y(_1974_));
 sky130_fd_sc_hd__nor2_1 _4534_ (.A(_1820_),
    .B(_1974_),
    .Y(_1975_));
 sky130_fd_sc_hd__a21oi_1 _4535_ (.A1(_1129_),
    .A2(_1973_),
    .B1(_1975_),
    .Y(_1976_));
 sky130_fd_sc_hd__buf_4 _4536_ (.A(_1540_),
    .X(_1977_));
 sky130_fd_sc_hd__buf_4 _4537_ (.A(_1542_),
    .X(_1978_));
 sky130_fd_sc_hd__mux2_1 _4538_ (.A0(\mem[1][22] ),
    .A1(\mem[3][22] ),
    .S(_1663_),
    .X(_1979_));
 sky130_fd_sc_hd__nand4_1 _4539_ (.A(_1977_),
    .B(_1978_),
    .C(_1939_),
    .D(_1979_),
    .Y(_1980_));
 sky130_fd_sc_hd__o31ai_1 _4540_ (.A1(_1852_),
    .A2(_1938_),
    .A3(_1139_),
    .B1(_1980_),
    .Y(_1981_));
 sky130_fd_sc_hd__mux2i_1 _4541_ (.A0(\mem[4][22] ),
    .A1(\mem[6][22] ),
    .S(_1699_),
    .Y(_1982_));
 sky130_fd_sc_hd__o221ai_1 _4542_ (.A1(_1130_),
    .A2(_1827_),
    .B1(_1943_),
    .B2(_1982_),
    .C1(_1796_),
    .Y(_1983_));
 sky130_fd_sc_hd__o21ai_0 _4543_ (.A1(_1937_),
    .A2(_1981_),
    .B1(_1983_),
    .Y(_1984_));
 sky130_fd_sc_hd__o22ai_1 _4544_ (.A1(\mem[1][22] ),
    .A2(_1947_),
    .B1(_1948_),
    .B2(\mem[0][22] ),
    .Y(_1985_));
 sky130_fd_sc_hd__o22ai_1 _4545_ (.A1(\mem[2][22] ),
    .A2(_1672_),
    .B1(_1673_),
    .B2(\mem[3][22] ),
    .Y(_1986_));
 sky130_fd_sc_hd__or3_1 _4546_ (.A(_1670_),
    .B(_1985_),
    .C(_1986_),
    .X(_1987_));
 sky130_fd_sc_hd__buf_6 _4547_ (.A(_1560_),
    .X(_1988_));
 sky130_fd_sc_hd__o2111ai_2 _4548_ (.A1(_1933_),
    .A2(_1976_),
    .B1(_1984_),
    .C1(_1987_),
    .D1(_1988_),
    .Y(_1989_));
 sky130_fd_sc_hd__mux2i_1 _4549_ (.A0(\mem[12][22] ),
    .A1(\mem[14][22] ),
    .S(_1954_),
    .Y(_1990_));
 sky130_fd_sc_hd__mux2_1 _4550_ (.A0(\mem[8][22] ),
    .A1(\mem[10][22] ),
    .S(_1709_),
    .X(_1991_));
 sky130_fd_sc_hd__nand3_1 _4551_ (.A(_1804_),
    .B(_1805_),
    .C(_1991_),
    .Y(_1992_));
 sky130_fd_sc_hd__o22ai_1 _4552_ (.A1(_1708_),
    .A2(_1144_),
    .B1(_1992_),
    .B2(_1958_),
    .Y(_1993_));
 sky130_fd_sc_hd__nor2_1 _4553_ (.A(_1960_),
    .B(_1992_),
    .Y(_1994_));
 sky130_fd_sc_hd__o21ai_0 _4554_ (.A1(_1810_),
    .A2(_1135_),
    .B1(_1778_),
    .Y(_1995_));
 sky130_fd_sc_hd__o22ai_1 _4555_ (.A1(_1864_),
    .A2(_1993_),
    .B1(_1994_),
    .B2(_1995_),
    .Y(_1996_));
 sky130_fd_sc_hd__buf_4 _4556_ (.A(_1501_),
    .X(_1997_));
 sky130_fd_sc_hd__o211ai_1 _4557_ (.A1(_1953_),
    .A2(_1990_),
    .B1(_1996_),
    .C1(_1997_),
    .Y(_1998_));
 sky130_fd_sc_hd__mux2i_1 _4558_ (.A0(\mem[13][22] ),
    .A1(\mem[15][22] ),
    .S(_1872_),
    .Y(_1999_));
 sky130_fd_sc_hd__clkbuf_8 _4559_ (.A(_0714_),
    .X(_2000_));
 sky130_fd_sc_hd__nand3_1 _4560_ (.A(_1654_),
    .B(_2000_),
    .C(_1133_),
    .Y(_2001_));
 sky130_fd_sc_hd__o221ai_1 _4561_ (.A1(_1143_),
    .A2(_1685_),
    .B1(_1782_),
    .B2(_1999_),
    .C1(_2001_),
    .Y(_2002_));
 sky130_fd_sc_hd__mux2i_1 _4562_ (.A0(\mem[9][22] ),
    .A1(\mem[11][22] ),
    .S(_1968_),
    .Y(_2003_));
 sky130_fd_sc_hd__o21ai_0 _4563_ (.A1(_1876_),
    .A2(_2003_),
    .B1(_1970_),
    .Y(_2004_));
 sky130_fd_sc_hd__o22a_1 _4564_ (.A1(net127),
    .A2(_1652_),
    .B1(_2002_),
    .B2(_2004_),
    .X(_2005_));
 sky130_fd_sc_hd__and3_1 _4565_ (.A(_1989_),
    .B(_1998_),
    .C(_2005_),
    .X(_0581_));
 sky130_fd_sc_hd__mux2i_1 _4566_ (.A0(\mem[5][23] ),
    .A1(\mem[7][23] ),
    .S(_1692_),
    .Y(_2006_));
 sky130_fd_sc_hd__nor2_1 _4567_ (.A(_1820_),
    .B(_2006_),
    .Y(_2007_));
 sky130_fd_sc_hd__a21oi_1 _4568_ (.A1(_1149_),
    .A2(_1973_),
    .B1(_2007_),
    .Y(_2008_));
 sky130_fd_sc_hd__mux2_1 _4569_ (.A0(\mem[1][23] ),
    .A1(\mem[3][23] ),
    .S(_1663_),
    .X(_2009_));
 sky130_fd_sc_hd__nand4_1 _4570_ (.A(_1977_),
    .B(_1978_),
    .C(_1939_),
    .D(_2009_),
    .Y(_2010_));
 sky130_fd_sc_hd__o31ai_1 _4571_ (.A1(_1852_),
    .A2(_1938_),
    .A3(_1160_),
    .B1(_2010_),
    .Y(_2011_));
 sky130_fd_sc_hd__mux2i_1 _4572_ (.A0(\mem[4][23] ),
    .A1(\mem[6][23] ),
    .S(_1699_),
    .Y(_2012_));
 sky130_fd_sc_hd__o221ai_1 _4573_ (.A1(_1150_),
    .A2(_1827_),
    .B1(_1943_),
    .B2(_2012_),
    .C1(_1796_),
    .Y(_2013_));
 sky130_fd_sc_hd__o21ai_0 _4574_ (.A1(_1937_),
    .A2(_2011_),
    .B1(_2013_),
    .Y(_2014_));
 sky130_fd_sc_hd__o22ai_1 _4575_ (.A1(\mem[1][23] ),
    .A2(_1947_),
    .B1(_1948_),
    .B2(\mem[0][23] ),
    .Y(_2015_));
 sky130_fd_sc_hd__o22ai_1 _4576_ (.A1(\mem[2][23] ),
    .A2(_1672_),
    .B1(_1673_),
    .B2(\mem[3][23] ),
    .Y(_2016_));
 sky130_fd_sc_hd__or3_1 _4577_ (.A(_1670_),
    .B(_2015_),
    .C(_2016_),
    .X(_2017_));
 sky130_fd_sc_hd__o2111ai_2 _4578_ (.A1(_1933_),
    .A2(_2008_),
    .B1(_2014_),
    .C1(_2017_),
    .D1(_1988_),
    .Y(_2018_));
 sky130_fd_sc_hd__mux2i_1 _4579_ (.A0(\mem[12][23] ),
    .A1(\mem[14][23] ),
    .S(_1954_),
    .Y(_2019_));
 sky130_fd_sc_hd__mux2_1 _4580_ (.A0(\mem[8][23] ),
    .A1(\mem[10][23] ),
    .S(_1709_),
    .X(_2020_));
 sky130_fd_sc_hd__nand3_1 _4581_ (.A(_1804_),
    .B(_1805_),
    .C(_2020_),
    .Y(_2021_));
 sky130_fd_sc_hd__o22ai_1 _4582_ (.A1(_1708_),
    .A2(_1163_),
    .B1(_2021_),
    .B2(_1958_),
    .Y(_2022_));
 sky130_fd_sc_hd__nor2_1 _4583_ (.A(_1960_),
    .B(_2021_),
    .Y(_2023_));
 sky130_fd_sc_hd__o21ai_0 _4584_ (.A1(_1810_),
    .A2(_1155_),
    .B1(_1778_),
    .Y(_2024_));
 sky130_fd_sc_hd__o22ai_1 _4585_ (.A1(_1864_),
    .A2(_2022_),
    .B1(_2023_),
    .B2(_2024_),
    .Y(_2025_));
 sky130_fd_sc_hd__o211ai_1 _4586_ (.A1(_1953_),
    .A2(_2019_),
    .B1(_2025_),
    .C1(_1997_),
    .Y(_2026_));
 sky130_fd_sc_hd__buf_4 _4587_ (.A(_0721_),
    .X(_2027_));
 sky130_fd_sc_hd__mux2i_1 _4588_ (.A0(\mem[13][23] ),
    .A1(\mem[15][23] ),
    .S(_1872_),
    .Y(_2028_));
 sky130_fd_sc_hd__clkbuf_8 _4589_ (.A(_0827_),
    .X(_2029_));
 sky130_fd_sc_hd__nand3_1 _4590_ (.A(_2029_),
    .B(_2000_),
    .C(_1154_),
    .Y(_2030_));
 sky130_fd_sc_hd__o221ai_1 _4591_ (.A1(_1162_),
    .A2(_1685_),
    .B1(_1782_),
    .B2(_2028_),
    .C1(_2030_),
    .Y(_2031_));
 sky130_fd_sc_hd__mux2i_1 _4592_ (.A0(\mem[9][23] ),
    .A1(\mem[11][23] ),
    .S(_1968_),
    .Y(_2032_));
 sky130_fd_sc_hd__o21ai_0 _4593_ (.A1(_1876_),
    .A2(_2032_),
    .B1(_1970_),
    .Y(_2033_));
 sky130_fd_sc_hd__o22a_1 _4594_ (.A1(net128),
    .A2(_2027_),
    .B1(_2031_),
    .B2(_2033_),
    .X(_2034_));
 sky130_fd_sc_hd__and3_1 _4595_ (.A(_2018_),
    .B(_2026_),
    .C(_2034_),
    .X(_0582_));
 sky130_fd_sc_hd__mux2i_1 _4596_ (.A0(\mem[13][24] ),
    .A1(\mem[15][24] ),
    .S(_1599_),
    .Y(_2035_));
 sky130_fd_sc_hd__o22ai_1 _4597_ (.A1(_1182_),
    .A2(_1597_),
    .B1(_1598_),
    .B2(_2035_),
    .Y(_2036_));
 sky130_fd_sc_hd__a211oi_1 _4598_ (.A1(_1595_),
    .A2(_2036_),
    .B1(_1593_),
    .C1(net163),
    .Y(_2037_));
 sky130_fd_sc_hd__mux2i_1 _4599_ (.A0(\mem[9][24] ),
    .A1(\mem[11][24] ),
    .S(_1727_),
    .Y(_2038_));
 sky130_fd_sc_hd__o221ai_1 _4600_ (.A1(_1173_),
    .A2(_1495_),
    .B1(_1726_),
    .B2(_2038_),
    .C1(_1595_),
    .Y(_2039_));
 sky130_fd_sc_hd__mux2i_1 _4601_ (.A0(\mem[12][24] ),
    .A1(\mem[14][24] ),
    .S(_1533_),
    .Y(_2040_));
 sky130_fd_sc_hd__o221ai_1 _4602_ (.A1(_1181_),
    .A2(_1597_),
    .B1(_1531_),
    .B2(_2040_),
    .C1(_1731_),
    .Y(_2041_));
 sky130_fd_sc_hd__o22ai_1 _4603_ (.A1(\mem[10][24] ),
    .A2(_1463_),
    .B1(_1465_),
    .B2(\mem[11][24] ),
    .Y(_2042_));
 sky130_fd_sc_hd__o22ai_1 _4604_ (.A1(\mem[9][24] ),
    .A2(_1456_),
    .B1(_1460_),
    .B2(\mem[8][24] ),
    .Y(_2043_));
 sky130_fd_sc_hd__nor3_1 _4605_ (.A(_1472_),
    .B(_2042_),
    .C(_2043_),
    .Y(_2044_));
 sky130_fd_sc_hd__a21oi_1 _4606_ (.A1(_2039_),
    .A2(_2041_),
    .B1(_2044_),
    .Y(_2045_));
 sky130_fd_sc_hd__mux2i_2 _4607_ (.A0(\mem[4][24] ),
    .A1(\mem[6][24] ),
    .S(_1738_),
    .Y(_2046_));
 sky130_fd_sc_hd__mux2_1 _4608_ (.A0(\mem[0][24] ),
    .A1(\mem[2][24] ),
    .S(_1483_),
    .X(_2047_));
 sky130_fd_sc_hd__nand3_1 _4609_ (.A(_1540_),
    .B(_1542_),
    .C(_2047_),
    .Y(_2048_));
 sky130_fd_sc_hd__o22ai_1 _4610_ (.A1(_1740_),
    .A2(_1170_),
    .B1(_2048_),
    .B2(_1743_),
    .Y(_2049_));
 sky130_fd_sc_hd__nor2_1 _4611_ (.A(_1745_),
    .B(_2048_),
    .Y(_2050_));
 sky130_fd_sc_hd__o21ai_0 _4612_ (.A1(_1567_),
    .A2(_1179_),
    .B1(_0828_),
    .Y(_2051_));
 sky130_fd_sc_hd__o22ai_1 _4613_ (.A1(_1488_),
    .A2(_2049_),
    .B1(_2050_),
    .B2(_2051_),
    .Y(_2052_));
 sky130_fd_sc_hd__o211a_1 _4614_ (.A1(_1737_),
    .A2(_2046_),
    .B1(_2052_),
    .C1(_1509_),
    .X(_2053_));
 sky130_fd_sc_hd__mux2i_1 _4615_ (.A0(\mem[5][24] ),
    .A1(\mem[7][24] ),
    .S(_1532_),
    .Y(_2054_));
 sky130_fd_sc_hd__nor2_1 _4616_ (.A(_1530_),
    .B(_2054_),
    .Y(_2055_));
 sky130_fd_sc_hd__nor3_1 _4617_ (.A(_1752_),
    .B(_1489_),
    .C(_1180_),
    .Y(_2056_));
 sky130_fd_sc_hd__a311o_1 _4618_ (.A1(_1752_),
    .A2(_1627_),
    .A3(_1168_),
    .B1(_2055_),
    .C1(_2056_),
    .X(_2057_));
 sky130_fd_sc_hd__mux2i_1 _4619_ (.A0(\mem[1][24] ),
    .A1(\mem[3][24] ),
    .S(_1727_),
    .Y(_2058_));
 sky130_fd_sc_hd__nor2_1 _4620_ (.A(_1726_),
    .B(_2058_),
    .Y(_2059_));
 sky130_fd_sc_hd__o32ai_1 _4621_ (.A1(_1522_),
    .A2(_2057_),
    .A3(_2059_),
    .B1(_2537_),
    .B2(net129),
    .Y(_2060_));
 sky130_fd_sc_hd__a211oi_1 _4622_ (.A1(_2037_),
    .A2(_2045_),
    .B1(_2053_),
    .C1(_2060_),
    .Y(_0583_));
 sky130_fd_sc_hd__mux2i_1 _4623_ (.A0(\mem[5][25] ),
    .A1(\mem[7][25] ),
    .S(_1692_),
    .Y(_2061_));
 sky130_fd_sc_hd__nor2_1 _4624_ (.A(_1820_),
    .B(_2061_),
    .Y(_2062_));
 sky130_fd_sc_hd__a21oi_1 _4625_ (.A1(_1189_),
    .A2(_1973_),
    .B1(_2062_),
    .Y(_2063_));
 sky130_fd_sc_hd__buf_6 _4626_ (.A(_1457_),
    .X(_2064_));
 sky130_fd_sc_hd__mux2_1 _4627_ (.A0(\mem[1][25] ),
    .A1(\mem[3][25] ),
    .S(_2064_),
    .X(_2065_));
 sky130_fd_sc_hd__nand4_1 _4628_ (.A(_1977_),
    .B(_1978_),
    .C(_1939_),
    .D(_2065_),
    .Y(_2066_));
 sky130_fd_sc_hd__o31ai_1 _4629_ (.A1(_1852_),
    .A2(_1938_),
    .A3(_1198_),
    .B1(_2066_),
    .Y(_2067_));
 sky130_fd_sc_hd__mux2i_1 _4630_ (.A0(\mem[4][25] ),
    .A1(\mem[6][25] ),
    .S(_1699_),
    .Y(_2068_));
 sky130_fd_sc_hd__o221ai_1 _4631_ (.A1(_1190_),
    .A2(_1827_),
    .B1(_1943_),
    .B2(_2068_),
    .C1(_1796_),
    .Y(_2069_));
 sky130_fd_sc_hd__o21ai_0 _4632_ (.A1(_1937_),
    .A2(_2067_),
    .B1(_2069_),
    .Y(_2070_));
 sky130_fd_sc_hd__buf_4 _4633_ (.A(_1471_),
    .X(_2071_));
 sky130_fd_sc_hd__o22ai_1 _4634_ (.A1(\mem[2][25] ),
    .A2(_1767_),
    .B1(_1768_),
    .B2(\mem[3][25] ),
    .Y(_2072_));
 sky130_fd_sc_hd__o22ai_1 _4635_ (.A1(\mem[1][25] ),
    .A2(_1456_),
    .B1(_1460_),
    .B2(\mem[0][25] ),
    .Y(_2073_));
 sky130_fd_sc_hd__or3_1 _4636_ (.A(_2071_),
    .B(_2072_),
    .C(_2073_),
    .X(_2074_));
 sky130_fd_sc_hd__o2111ai_2 _4637_ (.A1(_1933_),
    .A2(_2063_),
    .B1(_2070_),
    .C1(_2074_),
    .D1(_1988_),
    .Y(_2075_));
 sky130_fd_sc_hd__mux2i_1 _4638_ (.A0(\mem[12][25] ),
    .A1(\mem[14][25] ),
    .S(_1954_),
    .Y(_2076_));
 sky130_fd_sc_hd__mux2_1 _4639_ (.A0(\mem[8][25] ),
    .A1(\mem[10][25] ),
    .S(_1709_),
    .X(_2077_));
 sky130_fd_sc_hd__nand3_1 _4640_ (.A(_1804_),
    .B(_1805_),
    .C(_2077_),
    .Y(_2078_));
 sky130_fd_sc_hd__o22ai_1 _4641_ (.A1(_1708_),
    .A2(_1202_),
    .B1(_2078_),
    .B2(_1958_),
    .Y(_2079_));
 sky130_fd_sc_hd__nor2_1 _4642_ (.A(_1960_),
    .B(_2078_),
    .Y(_2080_));
 sky130_fd_sc_hd__o21ai_0 _4643_ (.A1(_1810_),
    .A2(_1194_),
    .B1(_1778_),
    .Y(_2081_));
 sky130_fd_sc_hd__o22ai_1 _4644_ (.A1(_1864_),
    .A2(_2079_),
    .B1(_2080_),
    .B2(_2081_),
    .Y(_2082_));
 sky130_fd_sc_hd__o211ai_1 _4645_ (.A1(_1953_),
    .A2(_2076_),
    .B1(_2082_),
    .C1(_1997_),
    .Y(_2083_));
 sky130_fd_sc_hd__buf_6 _4646_ (.A(_1494_),
    .X(_2084_));
 sky130_fd_sc_hd__mux2i_1 _4647_ (.A0(\mem[13][25] ),
    .A1(\mem[15][25] ),
    .S(_1872_),
    .Y(_2085_));
 sky130_fd_sc_hd__nand3_1 _4648_ (.A(_2029_),
    .B(_2000_),
    .C(_1193_),
    .Y(_2086_));
 sky130_fd_sc_hd__o221ai_1 _4649_ (.A1(_1200_),
    .A2(_2084_),
    .B1(_1782_),
    .B2(_2085_),
    .C1(_2086_),
    .Y(_2087_));
 sky130_fd_sc_hd__mux2i_1 _4650_ (.A0(\mem[9][25] ),
    .A1(\mem[11][25] ),
    .S(_1968_),
    .Y(_2088_));
 sky130_fd_sc_hd__o21ai_0 _4651_ (.A1(_1876_),
    .A2(_2088_),
    .B1(_1970_),
    .Y(_2089_));
 sky130_fd_sc_hd__o22a_1 _4652_ (.A1(net130),
    .A2(_2027_),
    .B1(_2087_),
    .B2(_2089_),
    .X(_2090_));
 sky130_fd_sc_hd__and3_1 _4653_ (.A(_2075_),
    .B(_2083_),
    .C(_2090_),
    .X(_0584_));
 sky130_fd_sc_hd__buf_6 _4654_ (.A(_1532_),
    .X(_2091_));
 sky130_fd_sc_hd__mux2i_1 _4655_ (.A0(\mem[5][26] ),
    .A1(\mem[7][26] ),
    .S(_2091_),
    .Y(_2092_));
 sky130_fd_sc_hd__nor2_1 _4656_ (.A(_1820_),
    .B(_2092_),
    .Y(_2093_));
 sky130_fd_sc_hd__a21oi_1 _4657_ (.A1(_1207_),
    .A2(_1973_),
    .B1(_2093_),
    .Y(_2094_));
 sky130_fd_sc_hd__mux2_1 _4658_ (.A0(\mem[1][26] ),
    .A1(\mem[3][26] ),
    .S(_2064_),
    .X(_2095_));
 sky130_fd_sc_hd__nand4_1 _4659_ (.A(_1977_),
    .B(_1978_),
    .C(_1939_),
    .D(_2095_),
    .Y(_2096_));
 sky130_fd_sc_hd__o31ai_1 _4660_ (.A1(_1852_),
    .A2(_1938_),
    .A3(_1216_),
    .B1(_2096_),
    .Y(_2097_));
 sky130_fd_sc_hd__buf_6 _4661_ (.A(_1510_),
    .X(_2098_));
 sky130_fd_sc_hd__mux2i_1 _4662_ (.A0(\mem[4][26] ),
    .A1(\mem[6][26] ),
    .S(_2098_),
    .Y(_2099_));
 sky130_fd_sc_hd__o221ai_1 _4663_ (.A1(_1208_),
    .A2(_1827_),
    .B1(_1943_),
    .B2(_2099_),
    .C1(_1796_),
    .Y(_2100_));
 sky130_fd_sc_hd__o21ai_0 _4664_ (.A1(_1937_),
    .A2(_2097_),
    .B1(_2100_),
    .Y(_2101_));
 sky130_fd_sc_hd__o22ai_1 _4665_ (.A1(\mem[1][26] ),
    .A2(_1947_),
    .B1(_1948_),
    .B2(\mem[0][26] ),
    .Y(_2102_));
 sky130_fd_sc_hd__o22ai_1 _4666_ (.A1(\mem[2][26] ),
    .A2(_1672_),
    .B1(_1673_),
    .B2(\mem[3][26] ),
    .Y(_2103_));
 sky130_fd_sc_hd__or3_1 _4667_ (.A(_2071_),
    .B(_2102_),
    .C(_2103_),
    .X(_2104_));
 sky130_fd_sc_hd__o2111ai_2 _4668_ (.A1(_1933_),
    .A2(_2094_),
    .B1(_2101_),
    .C1(_2104_),
    .D1(_1988_),
    .Y(_2105_));
 sky130_fd_sc_hd__mux2i_1 _4669_ (.A0(\mem[12][26] ),
    .A1(\mem[14][26] ),
    .S(_1954_),
    .Y(_2106_));
 sky130_fd_sc_hd__buf_6 _4670_ (.A(_0715_),
    .X(_2107_));
 sky130_fd_sc_hd__buf_6 _4671_ (.A(_1457_),
    .X(_2108_));
 sky130_fd_sc_hd__mux2_1 _4672_ (.A0(\mem[8][26] ),
    .A1(\mem[10][26] ),
    .S(_2108_),
    .X(_2109_));
 sky130_fd_sc_hd__nand3_1 _4673_ (.A(_1804_),
    .B(_1805_),
    .C(_2109_),
    .Y(_2110_));
 sky130_fd_sc_hd__o22ai_1 _4674_ (.A1(_2107_),
    .A2(_1219_),
    .B1(_2110_),
    .B2(_1958_),
    .Y(_2111_));
 sky130_fd_sc_hd__nor2_1 _4675_ (.A(_1960_),
    .B(_2110_),
    .Y(_2112_));
 sky130_fd_sc_hd__o21ai_0 _4676_ (.A1(_1810_),
    .A2(_1212_),
    .B1(_1778_),
    .Y(_2113_));
 sky130_fd_sc_hd__o22ai_1 _4677_ (.A1(_1864_),
    .A2(_2111_),
    .B1(_2112_),
    .B2(_2113_),
    .Y(_2114_));
 sky130_fd_sc_hd__o211ai_1 _4678_ (.A1(_1953_),
    .A2(_2106_),
    .B1(_2114_),
    .C1(_1997_),
    .Y(_2115_));
 sky130_fd_sc_hd__mux2i_1 _4679_ (.A0(\mem[13][26] ),
    .A1(\mem[15][26] ),
    .S(_1872_),
    .Y(_2116_));
 sky130_fd_sc_hd__nand3_1 _4680_ (.A(_2029_),
    .B(_2000_),
    .C(_1211_),
    .Y(_2117_));
 sky130_fd_sc_hd__o221ai_1 _4681_ (.A1(_1218_),
    .A2(_2084_),
    .B1(_1782_),
    .B2(_2116_),
    .C1(_2117_),
    .Y(_2118_));
 sky130_fd_sc_hd__mux2i_1 _4682_ (.A0(\mem[9][26] ),
    .A1(\mem[11][26] ),
    .S(_1968_),
    .Y(_2119_));
 sky130_fd_sc_hd__o21ai_0 _4683_ (.A1(_1876_),
    .A2(_2119_),
    .B1(_1970_),
    .Y(_2120_));
 sky130_fd_sc_hd__o22a_1 _4684_ (.A1(net131),
    .A2(_2027_),
    .B1(_2118_),
    .B2(_2120_),
    .X(_2121_));
 sky130_fd_sc_hd__and3_1 _4685_ (.A(_2105_),
    .B(_2115_),
    .C(_2121_),
    .X(_0585_));
 sky130_fd_sc_hd__mux2i_1 _4686_ (.A0(\mem[5][27] ),
    .A1(\mem[7][27] ),
    .S(_2091_),
    .Y(_2122_));
 sky130_fd_sc_hd__nor2_1 _4687_ (.A(_1820_),
    .B(_2122_),
    .Y(_2123_));
 sky130_fd_sc_hd__a21oi_1 _4688_ (.A1(_1225_),
    .A2(_1973_),
    .B1(_2123_),
    .Y(_2124_));
 sky130_fd_sc_hd__mux2_1 _4689_ (.A0(\mem[1][27] ),
    .A1(\mem[3][27] ),
    .S(_2064_),
    .X(_2125_));
 sky130_fd_sc_hd__nand4_1 _4690_ (.A(_1977_),
    .B(_1978_),
    .C(_1939_),
    .D(_2125_),
    .Y(_2126_));
 sky130_fd_sc_hd__o31ai_1 _4691_ (.A1(_1852_),
    .A2(_1938_),
    .A3(_1235_),
    .B1(_2126_),
    .Y(_2127_));
 sky130_fd_sc_hd__mux2i_1 _4692_ (.A0(\mem[4][27] ),
    .A1(\mem[6][27] ),
    .S(_2098_),
    .Y(_2128_));
 sky130_fd_sc_hd__o221ai_1 _4693_ (.A1(_1226_),
    .A2(_1827_),
    .B1(_1943_),
    .B2(_2128_),
    .C1(_1796_),
    .Y(_2129_));
 sky130_fd_sc_hd__o21ai_0 _4694_ (.A1(_1937_),
    .A2(_2127_),
    .B1(_2129_),
    .Y(_2130_));
 sky130_fd_sc_hd__o22ai_1 _4695_ (.A1(\mem[1][27] ),
    .A2(_1947_),
    .B1(_1948_),
    .B2(\mem[0][27] ),
    .Y(_2131_));
 sky130_fd_sc_hd__o22ai_1 _4696_ (.A1(\mem[2][27] ),
    .A2(_1672_),
    .B1(_1673_),
    .B2(\mem[3][27] ),
    .Y(_2132_));
 sky130_fd_sc_hd__or3_1 _4697_ (.A(_2071_),
    .B(_2131_),
    .C(_2132_),
    .X(_2133_));
 sky130_fd_sc_hd__o2111ai_2 _4698_ (.A1(_1933_),
    .A2(_2124_),
    .B1(_2130_),
    .C1(_2133_),
    .D1(_1988_),
    .Y(_2134_));
 sky130_fd_sc_hd__mux2i_1 _4699_ (.A0(\mem[12][27] ),
    .A1(\mem[14][27] ),
    .S(_1954_),
    .Y(_2135_));
 sky130_fd_sc_hd__mux2_1 _4700_ (.A0(\mem[8][27] ),
    .A1(\mem[10][27] ),
    .S(_2108_),
    .X(_2136_));
 sky130_fd_sc_hd__nand3_1 _4701_ (.A(_1804_),
    .B(_1805_),
    .C(_2136_),
    .Y(_2137_));
 sky130_fd_sc_hd__o22ai_1 _4702_ (.A1(_2107_),
    .A2(_1238_),
    .B1(_2137_),
    .B2(_1958_),
    .Y(_2138_));
 sky130_fd_sc_hd__nor2_1 _4703_ (.A(_1960_),
    .B(_2137_),
    .Y(_2139_));
 sky130_fd_sc_hd__buf_4 _4704_ (.A(_0827_),
    .X(_2140_));
 sky130_fd_sc_hd__o21ai_0 _4705_ (.A1(_1810_),
    .A2(_1231_),
    .B1(_2140_),
    .Y(_2141_));
 sky130_fd_sc_hd__o22ai_1 _4706_ (.A1(_1864_),
    .A2(_2138_),
    .B1(_2139_),
    .B2(_2141_),
    .Y(_2142_));
 sky130_fd_sc_hd__o211ai_1 _4707_ (.A1(_1953_),
    .A2(_2135_),
    .B1(_2142_),
    .C1(_1997_),
    .Y(_2143_));
 sky130_fd_sc_hd__buf_6 _4708_ (.A(_1529_),
    .X(_2144_));
 sky130_fd_sc_hd__mux2i_1 _4709_ (.A0(\mem[13][27] ),
    .A1(\mem[15][27] ),
    .S(_1872_),
    .Y(_2145_));
 sky130_fd_sc_hd__nand3_1 _4710_ (.A(_2029_),
    .B(_2000_),
    .C(_1230_),
    .Y(_2146_));
 sky130_fd_sc_hd__o221ai_1 _4711_ (.A1(_1237_),
    .A2(_2084_),
    .B1(_2144_),
    .B2(_2145_),
    .C1(_2146_),
    .Y(_2147_));
 sky130_fd_sc_hd__mux2i_1 _4712_ (.A0(\mem[9][27] ),
    .A1(\mem[11][27] ),
    .S(_1968_),
    .Y(_2148_));
 sky130_fd_sc_hd__o21ai_0 _4713_ (.A1(_1876_),
    .A2(_2148_),
    .B1(_1970_),
    .Y(_2149_));
 sky130_fd_sc_hd__o22a_1 _4714_ (.A1(net132),
    .A2(_2027_),
    .B1(_2147_),
    .B2(_2149_),
    .X(_2150_));
 sky130_fd_sc_hd__and3_1 _4715_ (.A(_2134_),
    .B(_2143_),
    .C(_2150_),
    .X(_0586_));
 sky130_fd_sc_hd__mux2i_1 _4716_ (.A0(\mem[5][28] ),
    .A1(\mem[7][28] ),
    .S(_2091_),
    .Y(_2151_));
 sky130_fd_sc_hd__nor2_1 _4717_ (.A(_1820_),
    .B(_2151_),
    .Y(_2152_));
 sky130_fd_sc_hd__a21oi_1 _4718_ (.A1(_1245_),
    .A2(_1973_),
    .B1(_2152_),
    .Y(_2153_));
 sky130_fd_sc_hd__mux2_1 _4719_ (.A0(\mem[1][28] ),
    .A1(\mem[3][28] ),
    .S(_2064_),
    .X(_2154_));
 sky130_fd_sc_hd__nand4_1 _4720_ (.A(_1977_),
    .B(_1978_),
    .C(_1939_),
    .D(_2154_),
    .Y(_2155_));
 sky130_fd_sc_hd__o31ai_1 _4721_ (.A1(_1852_),
    .A2(_1938_),
    .A3(_1254_),
    .B1(_2155_),
    .Y(_2156_));
 sky130_fd_sc_hd__mux2i_1 _4722_ (.A0(\mem[4][28] ),
    .A1(\mem[6][28] ),
    .S(_2098_),
    .Y(_2157_));
 sky130_fd_sc_hd__o221ai_1 _4723_ (.A1(_1246_),
    .A2(_1827_),
    .B1(_1943_),
    .B2(_2157_),
    .C1(_0906_),
    .Y(_2158_));
 sky130_fd_sc_hd__o21ai_0 _4724_ (.A1(_1937_),
    .A2(_2156_),
    .B1(_2158_),
    .Y(_2159_));
 sky130_fd_sc_hd__o22ai_1 _4725_ (.A1(\mem[1][28] ),
    .A2(_1947_),
    .B1(_1948_),
    .B2(\mem[0][28] ),
    .Y(_2160_));
 sky130_fd_sc_hd__o22ai_1 _4726_ (.A1(\mem[2][28] ),
    .A2(_1767_),
    .B1(_1768_),
    .B2(\mem[3][28] ),
    .Y(_2161_));
 sky130_fd_sc_hd__or3_1 _4727_ (.A(_2071_),
    .B(_2160_),
    .C(_2161_),
    .X(_2162_));
 sky130_fd_sc_hd__o2111ai_2 _4728_ (.A1(_1933_),
    .A2(_2153_),
    .B1(_2159_),
    .C1(_2162_),
    .D1(_1988_),
    .Y(_2163_));
 sky130_fd_sc_hd__mux2i_1 _4729_ (.A0(\mem[12][28] ),
    .A1(\mem[14][28] ),
    .S(_1954_),
    .Y(_2164_));
 sky130_fd_sc_hd__mux2_1 _4730_ (.A0(\mem[8][28] ),
    .A1(\mem[10][28] ),
    .S(_2108_),
    .X(_2165_));
 sky130_fd_sc_hd__nand3_1 _4731_ (.A(_1490_),
    .B(_1491_),
    .C(_2165_),
    .Y(_2166_));
 sky130_fd_sc_hd__o22ai_1 _4732_ (.A1(_2107_),
    .A2(_1257_),
    .B1(_2166_),
    .B2(_1958_),
    .Y(_2167_));
 sky130_fd_sc_hd__nor2_1 _4733_ (.A(_1960_),
    .B(_2166_),
    .Y(_2168_));
 sky130_fd_sc_hd__o21ai_0 _4734_ (.A1(_1519_),
    .A2(_1250_),
    .B1(_2140_),
    .Y(_2169_));
 sky130_fd_sc_hd__o22ai_1 _4735_ (.A1(_1864_),
    .A2(_2167_),
    .B1(_2168_),
    .B2(_2169_),
    .Y(_2170_));
 sky130_fd_sc_hd__o211ai_1 _4736_ (.A1(_1953_),
    .A2(_2164_),
    .B1(_2170_),
    .C1(_1997_),
    .Y(_2171_));
 sky130_fd_sc_hd__mux2i_1 _4737_ (.A0(\mem[13][28] ),
    .A1(\mem[15][28] ),
    .S(_1872_),
    .Y(_2172_));
 sky130_fd_sc_hd__nand3_1 _4738_ (.A(_2029_),
    .B(_2000_),
    .C(_1249_),
    .Y(_2173_));
 sky130_fd_sc_hd__o221ai_1 _4739_ (.A1(_1256_),
    .A2(_2084_),
    .B1(_2144_),
    .B2(_2172_),
    .C1(_2173_),
    .Y(_2174_));
 sky130_fd_sc_hd__mux2i_1 _4740_ (.A0(\mem[9][28] ),
    .A1(\mem[11][28] ),
    .S(_1968_),
    .Y(_2175_));
 sky130_fd_sc_hd__o21ai_0 _4741_ (.A1(_1876_),
    .A2(_2175_),
    .B1(_1970_),
    .Y(_2176_));
 sky130_fd_sc_hd__o22a_1 _4742_ (.A1(net134),
    .A2(_2027_),
    .B1(_2174_),
    .B2(_2176_),
    .X(_2177_));
 sky130_fd_sc_hd__and3_1 _4743_ (.A(_2163_),
    .B(_2171_),
    .C(_2177_),
    .X(_0587_));
 sky130_fd_sc_hd__mux2i_1 _4744_ (.A0(\mem[13][29] ),
    .A1(\mem[15][29] ),
    .S(_1599_),
    .Y(_2178_));
 sky130_fd_sc_hd__o22ai_1 _4745_ (.A1(_1276_),
    .A2(_1597_),
    .B1(_1598_),
    .B2(_2178_),
    .Y(_2179_));
 sky130_fd_sc_hd__a211oi_1 _4746_ (.A1(_1595_),
    .A2(_2179_),
    .B1(_1593_),
    .C1(net163),
    .Y(_2180_));
 sky130_fd_sc_hd__mux2i_1 _4747_ (.A0(\mem[9][29] ),
    .A1(\mem[11][29] ),
    .S(_1599_),
    .Y(_2181_));
 sky130_fd_sc_hd__o221ai_1 _4748_ (.A1(_1267_),
    .A2(_1495_),
    .B1(_1726_),
    .B2(_2181_),
    .C1(_0903_),
    .Y(_2182_));
 sky130_fd_sc_hd__mux2i_1 _4749_ (.A0(\mem[12][29] ),
    .A1(\mem[14][29] ),
    .S(_1533_),
    .Y(_2183_));
 sky130_fd_sc_hd__o221ai_1 _4750_ (.A1(_1275_),
    .A2(_1548_),
    .B1(_1531_),
    .B2(_2183_),
    .C1(_1731_),
    .Y(_2184_));
 sky130_fd_sc_hd__o22ai_1 _4751_ (.A1(\mem[10][29] ),
    .A2(_1463_),
    .B1(_1465_),
    .B2(\mem[11][29] ),
    .Y(_2185_));
 sky130_fd_sc_hd__o22ai_1 _4752_ (.A1(\mem[9][29] ),
    .A2(_1456_),
    .B1(_1460_),
    .B2(\mem[8][29] ),
    .Y(_2186_));
 sky130_fd_sc_hd__nor3_1 _4753_ (.A(_1472_),
    .B(_2185_),
    .C(_2186_),
    .Y(_2187_));
 sky130_fd_sc_hd__a21oi_1 _4754_ (.A1(_2182_),
    .A2(_2184_),
    .B1(_2187_),
    .Y(_2188_));
 sky130_fd_sc_hd__mux2i_1 _4755_ (.A0(\mem[4][29] ),
    .A1(\mem[6][29] ),
    .S(_1738_),
    .Y(_2189_));
 sky130_fd_sc_hd__mux2_1 _4756_ (.A0(\mem[0][29] ),
    .A1(\mem[2][29] ),
    .S(_1483_),
    .X(_2190_));
 sky130_fd_sc_hd__nand3_1 _4757_ (.A(_1540_),
    .B(_1542_),
    .C(_2190_),
    .Y(_2191_));
 sky130_fd_sc_hd__o22ai_1 _4758_ (.A1(_1740_),
    .A2(_1264_),
    .B1(_2191_),
    .B2(_1743_),
    .Y(_2192_));
 sky130_fd_sc_hd__nor2_1 _4759_ (.A(_1745_),
    .B(_2191_),
    .Y(_2193_));
 sky130_fd_sc_hd__o21ai_0 _4760_ (.A1(_1567_),
    .A2(_1273_),
    .B1(_0828_),
    .Y(_2194_));
 sky130_fd_sc_hd__o22ai_1 _4761_ (.A1(_1488_),
    .A2(_2192_),
    .B1(_2193_),
    .B2(_2194_),
    .Y(_2195_));
 sky130_fd_sc_hd__o211a_1 _4762_ (.A1(_1737_),
    .A2(_2189_),
    .B1(_2195_),
    .C1(_1509_),
    .X(_2196_));
 sky130_fd_sc_hd__mux2i_1 _4763_ (.A0(\mem[5][29] ),
    .A1(\mem[7][29] ),
    .S(_1532_),
    .Y(_2197_));
 sky130_fd_sc_hd__nor2_1 _4764_ (.A(_1530_),
    .B(_2197_),
    .Y(_2198_));
 sky130_fd_sc_hd__nor3_1 _4765_ (.A(_1752_),
    .B(_1489_),
    .C(_1274_),
    .Y(_2199_));
 sky130_fd_sc_hd__a311o_1 _4766_ (.A1(_1752_),
    .A2(_1627_),
    .A3(_1263_),
    .B1(_2198_),
    .C1(_2199_),
    .X(_2200_));
 sky130_fd_sc_hd__mux2i_1 _4767_ (.A0(\mem[1][29] ),
    .A1(\mem[3][29] ),
    .S(_1727_),
    .Y(_2201_));
 sky130_fd_sc_hd__nor2_1 _4768_ (.A(_1726_),
    .B(_2201_),
    .Y(_2202_));
 sky130_fd_sc_hd__o32ai_1 _4769_ (.A1(_1522_),
    .A2(_2200_),
    .A3(_2202_),
    .B1(_2537_),
    .B2(net135),
    .Y(_2203_));
 sky130_fd_sc_hd__a211oi_1 _4770_ (.A1(_2180_),
    .A2(_2188_),
    .B1(_2196_),
    .C1(_2203_),
    .Y(_0588_));
 sky130_fd_sc_hd__mux2i_1 _4771_ (.A0(\mem[5][2] ),
    .A1(\mem[7][2] ),
    .S(_2091_),
    .Y(_2204_));
 sky130_fd_sc_hd__nor2_1 _4772_ (.A(_1563_),
    .B(_2204_),
    .Y(_2205_));
 sky130_fd_sc_hd__a21oi_1 _4773_ (.A1(_1281_),
    .A2(_1973_),
    .B1(_2205_),
    .Y(_2206_));
 sky130_fd_sc_hd__mux2_1 _4774_ (.A0(\mem[1][2] ),
    .A1(\mem[3][2] ),
    .S(_2064_),
    .X(_2207_));
 sky130_fd_sc_hd__nand4_1 _4775_ (.A(_1977_),
    .B(_1978_),
    .C(_1939_),
    .D(_2207_),
    .Y(_2208_));
 sky130_fd_sc_hd__o31ai_1 _4776_ (.A1(_1852_),
    .A2(_1938_),
    .A3(_1290_),
    .B1(_2208_),
    .Y(_2209_));
 sky130_fd_sc_hd__mux2i_1 _4777_ (.A0(\mem[4][2] ),
    .A1(\mem[6][2] ),
    .S(_2098_),
    .Y(_2210_));
 sky130_fd_sc_hd__o221ai_1 _4778_ (.A1(_1282_),
    .A2(_1596_),
    .B1(_1943_),
    .B2(_2210_),
    .C1(_0906_),
    .Y(_2211_));
 sky130_fd_sc_hd__o21ai_1 _4779_ (.A1(_1937_),
    .A2(_2209_),
    .B1(_2211_),
    .Y(_2212_));
 sky130_fd_sc_hd__o22ai_1 _4780_ (.A1(\mem[2][2] ),
    .A2(_1462_),
    .B1(_1464_),
    .B2(\mem[3][2] ),
    .Y(_2213_));
 sky130_fd_sc_hd__o22ai_1 _4781_ (.A1(\mem[1][2] ),
    .A2(_1555_),
    .B1(_1556_),
    .B2(\mem[0][2] ),
    .Y(_2214_));
 sky130_fd_sc_hd__or3_1 _4782_ (.A(_2071_),
    .B(_2213_),
    .C(_2214_),
    .X(_2215_));
 sky130_fd_sc_hd__o2111ai_4 _4783_ (.A1(_1933_),
    .A2(_2206_),
    .B1(_2212_),
    .C1(_2215_),
    .D1(_1988_),
    .Y(_2216_));
 sky130_fd_sc_hd__mux2i_1 _4784_ (.A0(\mem[12][2] ),
    .A1(\mem[14][2] ),
    .S(_1954_),
    .Y(_2217_));
 sky130_fd_sc_hd__mux2_1 _4785_ (.A0(\mem[8][2] ),
    .A1(\mem[10][2] ),
    .S(_2108_),
    .X(_2218_));
 sky130_fd_sc_hd__nand3_1 _4786_ (.A(_1490_),
    .B(_1491_),
    .C(_2218_),
    .Y(_2219_));
 sky130_fd_sc_hd__o22ai_1 _4787_ (.A1(_2107_),
    .A2(_1293_),
    .B1(_2219_),
    .B2(_1958_),
    .Y(_2220_));
 sky130_fd_sc_hd__nor2_1 _4788_ (.A(_1960_),
    .B(_2219_),
    .Y(_2221_));
 sky130_fd_sc_hd__o21ai_0 _4789_ (.A1(_1519_),
    .A2(_1286_),
    .B1(_2140_),
    .Y(_2222_));
 sky130_fd_sc_hd__o22ai_1 _4790_ (.A1(_1864_),
    .A2(_2220_),
    .B1(_2221_),
    .B2(_2222_),
    .Y(_2223_));
 sky130_fd_sc_hd__o211ai_1 _4791_ (.A1(_1953_),
    .A2(_2217_),
    .B1(_2223_),
    .C1(_1997_),
    .Y(_2224_));
 sky130_fd_sc_hd__mux2i_1 _4792_ (.A0(\mem[13][2] ),
    .A1(\mem[15][2] ),
    .S(_1872_),
    .Y(_2225_));
 sky130_fd_sc_hd__nand3_1 _4793_ (.A(_2029_),
    .B(_2000_),
    .C(_1285_),
    .Y(_2226_));
 sky130_fd_sc_hd__o221ai_1 _4794_ (.A1(_1292_),
    .A2(_2084_),
    .B1(_2144_),
    .B2(_2225_),
    .C1(_2226_),
    .Y(_2227_));
 sky130_fd_sc_hd__mux2i_1 _4795_ (.A0(\mem[9][2] ),
    .A1(\mem[11][2] ),
    .S(_1968_),
    .Y(_2228_));
 sky130_fd_sc_hd__o21ai_0 _4796_ (.A1(_1876_),
    .A2(_2228_),
    .B1(_1970_),
    .Y(_2229_));
 sky130_fd_sc_hd__o22a_1 _4797_ (.A1(net105),
    .A2(_2027_),
    .B1(_2227_),
    .B2(_2229_),
    .X(_2230_));
 sky130_fd_sc_hd__and3_1 _4798_ (.A(_2216_),
    .B(_2224_),
    .C(_2230_),
    .X(_0589_));
 sky130_fd_sc_hd__mux2i_1 _4799_ (.A0(\mem[5][30] ),
    .A1(\mem[7][30] ),
    .S(_2091_),
    .Y(_2231_));
 sky130_fd_sc_hd__nor2_1 _4800_ (.A(_1563_),
    .B(_2231_),
    .Y(_2232_));
 sky130_fd_sc_hd__a21oi_1 _4801_ (.A1(_1298_),
    .A2(_1973_),
    .B1(_2232_),
    .Y(_2233_));
 sky130_fd_sc_hd__mux2_1 _4802_ (.A0(\mem[1][30] ),
    .A1(\mem[3][30] ),
    .S(_2064_),
    .X(_2234_));
 sky130_fd_sc_hd__nand4_1 _4803_ (.A(_1977_),
    .B(_1978_),
    .C(_1939_),
    .D(_2234_),
    .Y(_2235_));
 sky130_fd_sc_hd__o31ai_1 _4804_ (.A1(_0860_),
    .A2(_1938_),
    .A3(_1307_),
    .B1(_2235_),
    .Y(_2236_));
 sky130_fd_sc_hd__mux2i_1 _4805_ (.A0(\mem[4][30] ),
    .A1(\mem[6][30] ),
    .S(_2098_),
    .Y(_2237_));
 sky130_fd_sc_hd__o221ai_1 _4806_ (.A1(_1299_),
    .A2(_1596_),
    .B1(_1943_),
    .B2(_2237_),
    .C1(_0906_),
    .Y(_2238_));
 sky130_fd_sc_hd__o21ai_0 _4807_ (.A1(_1937_),
    .A2(_2236_),
    .B1(_2238_),
    .Y(_2239_));
 sky130_fd_sc_hd__o22ai_1 _4808_ (.A1(\mem[1][30] ),
    .A2(_1947_),
    .B1(_1948_),
    .B2(\mem[0][30] ),
    .Y(_2240_));
 sky130_fd_sc_hd__o22ai_1 _4809_ (.A1(\mem[2][30] ),
    .A2(_1767_),
    .B1(_1768_),
    .B2(\mem[3][30] ),
    .Y(_2241_));
 sky130_fd_sc_hd__or3_1 _4810_ (.A(_2071_),
    .B(_2240_),
    .C(_2241_),
    .X(_2242_));
 sky130_fd_sc_hd__o2111ai_2 _4811_ (.A1(_1933_),
    .A2(_2233_),
    .B1(_2239_),
    .C1(_2242_),
    .D1(_1988_),
    .Y(_2243_));
 sky130_fd_sc_hd__mux2i_1 _4812_ (.A0(\mem[12][30] ),
    .A1(\mem[14][30] ),
    .S(_1954_),
    .Y(_2244_));
 sky130_fd_sc_hd__mux2_1 _4813_ (.A0(\mem[8][30] ),
    .A1(\mem[10][30] ),
    .S(_2108_),
    .X(_2245_));
 sky130_fd_sc_hd__nand3_1 _4814_ (.A(_1490_),
    .B(_1491_),
    .C(_2245_),
    .Y(_2246_));
 sky130_fd_sc_hd__o22ai_1 _4815_ (.A1(_2107_),
    .A2(_1310_),
    .B1(_2246_),
    .B2(_1958_),
    .Y(_2247_));
 sky130_fd_sc_hd__nor2_1 _4816_ (.A(_1960_),
    .B(_2246_),
    .Y(_2248_));
 sky130_fd_sc_hd__o21ai_0 _4817_ (.A1(_1519_),
    .A2(_1303_),
    .B1(_2140_),
    .Y(_2249_));
 sky130_fd_sc_hd__o22ai_1 _4818_ (.A1(_1514_),
    .A2(_2247_),
    .B1(_2248_),
    .B2(_2249_),
    .Y(_2250_));
 sky130_fd_sc_hd__o211ai_1 _4819_ (.A1(_1953_),
    .A2(_2244_),
    .B1(_2250_),
    .C1(_1997_),
    .Y(_2251_));
 sky130_fd_sc_hd__mux2i_1 _4820_ (.A0(\mem[13][30] ),
    .A1(\mem[15][30] ),
    .S(_1481_),
    .Y(_2252_));
 sky130_fd_sc_hd__nand3_1 _4821_ (.A(_2029_),
    .B(_2000_),
    .C(_1302_),
    .Y(_2253_));
 sky130_fd_sc_hd__o221ai_1 _4822_ (.A1(_1309_),
    .A2(_2084_),
    .B1(_2144_),
    .B2(_2252_),
    .C1(_2253_),
    .Y(_2254_));
 sky130_fd_sc_hd__mux2i_1 _4823_ (.A0(\mem[9][30] ),
    .A1(\mem[11][30] ),
    .S(_1968_),
    .Y(_2255_));
 sky130_fd_sc_hd__o21ai_0 _4824_ (.A1(_1588_),
    .A2(_2255_),
    .B1(_1970_),
    .Y(_2256_));
 sky130_fd_sc_hd__o22a_1 _4825_ (.A1(net136),
    .A2(_2027_),
    .B1(_2254_),
    .B2(_2256_),
    .X(_2257_));
 sky130_fd_sc_hd__and3_1 _4826_ (.A(_2243_),
    .B(_2251_),
    .C(_2257_),
    .X(_0590_));
 sky130_fd_sc_hd__mux2i_1 _4827_ (.A0(\mem[5][31] ),
    .A1(\mem[7][31] ),
    .S(_2091_),
    .Y(_2258_));
 sky130_fd_sc_hd__nor2_1 _4828_ (.A(_1563_),
    .B(_2258_),
    .Y(_2259_));
 sky130_fd_sc_hd__a21oi_1 _4829_ (.A1(_1315_),
    .A2(_1973_),
    .B1(_2259_),
    .Y(_2260_));
 sky130_fd_sc_hd__mux2_1 _4830_ (.A0(\mem[1][31] ),
    .A1(\mem[3][31] ),
    .S(_2064_),
    .X(_2261_));
 sky130_fd_sc_hd__nand4_1 _4831_ (.A(_1977_),
    .B(_1978_),
    .C(_1939_),
    .D(_2261_),
    .Y(_2262_));
 sky130_fd_sc_hd__o31ai_1 _4832_ (.A1(_0860_),
    .A2(_1938_),
    .A3(_1324_),
    .B1(_2262_),
    .Y(_2263_));
 sky130_fd_sc_hd__mux2i_1 _4833_ (.A0(\mem[4][31] ),
    .A1(\mem[6][31] ),
    .S(_2098_),
    .Y(_2264_));
 sky130_fd_sc_hd__o221ai_1 _4834_ (.A1(_1316_),
    .A2(_1596_),
    .B1(_1943_),
    .B2(_2264_),
    .C1(_0906_),
    .Y(_2265_));
 sky130_fd_sc_hd__o21ai_0 _4835_ (.A1(_1937_),
    .A2(_2263_),
    .B1(_2265_),
    .Y(_2266_));
 sky130_fd_sc_hd__o22ai_1 _4836_ (.A1(\mem[1][31] ),
    .A2(_1947_),
    .B1(_1948_),
    .B2(\mem[0][31] ),
    .Y(_2267_));
 sky130_fd_sc_hd__o22ai_1 _4837_ (.A1(\mem[2][31] ),
    .A2(_1767_),
    .B1(_1768_),
    .B2(\mem[3][31] ),
    .Y(_2268_));
 sky130_fd_sc_hd__or3_1 _4838_ (.A(_2071_),
    .B(_2267_),
    .C(_2268_),
    .X(_2269_));
 sky130_fd_sc_hd__o2111ai_2 _4839_ (.A1(_1933_),
    .A2(_2260_),
    .B1(_2266_),
    .C1(_2269_),
    .D1(_1988_),
    .Y(_2270_));
 sky130_fd_sc_hd__mux2i_1 _4840_ (.A0(\mem[12][31] ),
    .A1(\mem[14][31] ),
    .S(_1954_),
    .Y(_2271_));
 sky130_fd_sc_hd__mux2_1 _4841_ (.A0(\mem[8][31] ),
    .A1(\mem[10][31] ),
    .S(_2108_),
    .X(_2272_));
 sky130_fd_sc_hd__nand3_1 _4842_ (.A(_1490_),
    .B(_1491_),
    .C(_2272_),
    .Y(_2273_));
 sky130_fd_sc_hd__o22ai_1 _4843_ (.A1(_2107_),
    .A2(_1327_),
    .B1(_2273_),
    .B2(_1958_),
    .Y(_2274_));
 sky130_fd_sc_hd__nor2_1 _4844_ (.A(_1960_),
    .B(_2273_),
    .Y(_2275_));
 sky130_fd_sc_hd__o21ai_0 _4845_ (.A1(_1519_),
    .A2(_1320_),
    .B1(_2140_),
    .Y(_2276_));
 sky130_fd_sc_hd__o22ai_1 _4846_ (.A1(_1514_),
    .A2(_2274_),
    .B1(_2275_),
    .B2(_2276_),
    .Y(_2277_));
 sky130_fd_sc_hd__o211ai_1 _4847_ (.A1(_1953_),
    .A2(_2271_),
    .B1(_2277_),
    .C1(_1997_),
    .Y(_2278_));
 sky130_fd_sc_hd__mux2i_1 _4848_ (.A0(\mem[13][31] ),
    .A1(\mem[15][31] ),
    .S(_1481_),
    .Y(_2279_));
 sky130_fd_sc_hd__nand3_1 _4849_ (.A(_2029_),
    .B(_2000_),
    .C(_1319_),
    .Y(_2280_));
 sky130_fd_sc_hd__o221ai_1 _4850_ (.A1(_1326_),
    .A2(_2084_),
    .B1(_2144_),
    .B2(_2279_),
    .C1(_2280_),
    .Y(_2281_));
 sky130_fd_sc_hd__mux2i_1 _4851_ (.A0(\mem[9][31] ),
    .A1(\mem[11][31] ),
    .S(_1968_),
    .Y(_2282_));
 sky130_fd_sc_hd__o21ai_0 _4852_ (.A1(_1588_),
    .A2(_2282_),
    .B1(_1970_),
    .Y(_2283_));
 sky130_fd_sc_hd__o22a_1 _4853_ (.A1(net137),
    .A2(_2027_),
    .B1(_2281_),
    .B2(_2283_),
    .X(_2284_));
 sky130_fd_sc_hd__and3_1 _4854_ (.A(_2270_),
    .B(_2278_),
    .C(_2284_),
    .X(_0591_));
 sky130_fd_sc_hd__mux2i_1 _4855_ (.A0(\mem[5][3] ),
    .A1(\mem[7][3] ),
    .S(_2091_),
    .Y(_2285_));
 sky130_fd_sc_hd__nor2_1 _4856_ (.A(_1563_),
    .B(_2285_),
    .Y(_2286_));
 sky130_fd_sc_hd__a21oi_1 _4857_ (.A1(_1332_),
    .A2(_1973_),
    .B1(_2286_),
    .Y(_2287_));
 sky130_fd_sc_hd__mux2_1 _4858_ (.A0(\mem[1][3] ),
    .A1(\mem[3][3] ),
    .S(_2064_),
    .X(_2288_));
 sky130_fd_sc_hd__nand4_1 _4859_ (.A(_1977_),
    .B(_1978_),
    .C(_1478_),
    .D(_2288_),
    .Y(_2289_));
 sky130_fd_sc_hd__o31ai_1 _4860_ (.A1(_0860_),
    .A2(_1740_),
    .A3(_1341_),
    .B1(_2289_),
    .Y(_2290_));
 sky130_fd_sc_hd__mux2i_1 _4861_ (.A0(\mem[4][3] ),
    .A1(\mem[6][3] ),
    .S(_2098_),
    .Y(_2291_));
 sky130_fd_sc_hd__o221ai_1 _4862_ (.A1(_1333_),
    .A2(_1596_),
    .B1(_1580_),
    .B2(_2291_),
    .C1(_0906_),
    .Y(_2292_));
 sky130_fd_sc_hd__o21ai_0 _4863_ (.A1(_1552_),
    .A2(_2290_),
    .B1(_2292_),
    .Y(_2293_));
 sky130_fd_sc_hd__o22ai_1 _4864_ (.A1(\mem[1][3] ),
    .A2(_1947_),
    .B1(_1948_),
    .B2(\mem[0][3] ),
    .Y(_2294_));
 sky130_fd_sc_hd__o22ai_1 _4865_ (.A1(\mem[2][3] ),
    .A2(_1767_),
    .B1(_1768_),
    .B2(\mem[3][3] ),
    .Y(_2295_));
 sky130_fd_sc_hd__or3_1 _4866_ (.A(_2071_),
    .B(_2294_),
    .C(_2295_),
    .X(_2296_));
 sky130_fd_sc_hd__o2111ai_2 _4867_ (.A1(_1731_),
    .A2(_2287_),
    .B1(_2293_),
    .C1(_2296_),
    .D1(_1988_),
    .Y(_2297_));
 sky130_fd_sc_hd__mux2i_1 _4868_ (.A0(\mem[12][3] ),
    .A1(\mem[14][3] ),
    .S(_1738_),
    .Y(_2298_));
 sky130_fd_sc_hd__mux2_1 _4869_ (.A0(\mem[8][3] ),
    .A1(\mem[10][3] ),
    .S(_2108_),
    .X(_2299_));
 sky130_fd_sc_hd__nand3_1 _4870_ (.A(_1490_),
    .B(_1491_),
    .C(_2299_),
    .Y(_2300_));
 sky130_fd_sc_hd__o22ai_1 _4871_ (.A1(_2107_),
    .A2(_1344_),
    .B1(_2300_),
    .B2(_1743_),
    .Y(_2301_));
 sky130_fd_sc_hd__nor2_1 _4872_ (.A(_1745_),
    .B(_2300_),
    .Y(_2302_));
 sky130_fd_sc_hd__o21ai_0 _4873_ (.A1(_1519_),
    .A2(_1337_),
    .B1(_2140_),
    .Y(_2303_));
 sky130_fd_sc_hd__o22ai_1 _4874_ (.A1(_1514_),
    .A2(_2301_),
    .B1(_2302_),
    .B2(_2303_),
    .Y(_2304_));
 sky130_fd_sc_hd__o211ai_1 _4875_ (.A1(_1737_),
    .A2(_2298_),
    .B1(_2304_),
    .C1(_1997_),
    .Y(_2305_));
 sky130_fd_sc_hd__mux2i_1 _4876_ (.A0(\mem[13][3] ),
    .A1(\mem[15][3] ),
    .S(_1481_),
    .Y(_2306_));
 sky130_fd_sc_hd__nand3_1 _4877_ (.A(_2029_),
    .B(_2000_),
    .C(_1336_),
    .Y(_2307_));
 sky130_fd_sc_hd__o221ai_1 _4878_ (.A1(_1343_),
    .A2(_2084_),
    .B1(_2144_),
    .B2(_2306_),
    .C1(_2307_),
    .Y(_2308_));
 sky130_fd_sc_hd__mux2i_1 _4879_ (.A0(\mem[9][3] ),
    .A1(\mem[11][3] ),
    .S(_1550_),
    .Y(_2309_));
 sky130_fd_sc_hd__o21ai_0 _4880_ (.A1(_1588_),
    .A2(_2309_),
    .B1(_1475_),
    .Y(_2310_));
 sky130_fd_sc_hd__o22a_1 _4881_ (.A1(net106),
    .A2(_2027_),
    .B1(_2308_),
    .B2(_2310_),
    .X(_2311_));
 sky130_fd_sc_hd__and3_1 _4882_ (.A(_2297_),
    .B(_2305_),
    .C(_2311_),
    .X(_0592_));
 sky130_fd_sc_hd__mux2i_1 _4883_ (.A0(\mem[13][4] ),
    .A1(\mem[15][4] ),
    .S(_1599_),
    .Y(_2312_));
 sky130_fd_sc_hd__o22ai_1 _4884_ (.A1(_1362_),
    .A2(_1597_),
    .B1(_1598_),
    .B2(_2312_),
    .Y(_2313_));
 sky130_fd_sc_hd__a211oi_1 _4885_ (.A1(_1595_),
    .A2(_2313_),
    .B1(_1593_),
    .C1(net163),
    .Y(_2314_));
 sky130_fd_sc_hd__mux2i_1 _4886_ (.A0(\mem[9][4] ),
    .A1(\mem[11][4] ),
    .S(_1599_),
    .Y(_2315_));
 sky130_fd_sc_hd__o221ai_1 _4887_ (.A1(_1353_),
    .A2(_1495_),
    .B1(_1589_),
    .B2(_2315_),
    .C1(_0903_),
    .Y(_2316_));
 sky130_fd_sc_hd__mux2i_1 _4888_ (.A0(\mem[12][4] ),
    .A1(\mem[14][4] ),
    .S(_1533_),
    .Y(_2317_));
 sky130_fd_sc_hd__o221ai_1 _4889_ (.A1(_1361_),
    .A2(_1548_),
    .B1(_1531_),
    .B2(_2317_),
    .C1(_1731_),
    .Y(_2318_));
 sky130_fd_sc_hd__o22ai_1 _4890_ (.A1(\mem[10][4] ),
    .A2(_1463_),
    .B1(_1465_),
    .B2(\mem[11][4] ),
    .Y(_2319_));
 sky130_fd_sc_hd__o22ai_1 _4891_ (.A1(\mem[9][4] ),
    .A2(_1456_),
    .B1(_1460_),
    .B2(\mem[8][4] ),
    .Y(_2320_));
 sky130_fd_sc_hd__nor3_1 _4892_ (.A(_1472_),
    .B(_2319_),
    .C(_2320_),
    .Y(_2321_));
 sky130_fd_sc_hd__a21oi_1 _4893_ (.A1(_2316_),
    .A2(_2318_),
    .B1(_2321_),
    .Y(_2322_));
 sky130_fd_sc_hd__mux2i_1 _4894_ (.A0(\mem[4][4] ),
    .A1(\mem[6][4] ),
    .S(_1738_),
    .Y(_2323_));
 sky130_fd_sc_hd__mux2_1 _4895_ (.A0(\mem[0][4] ),
    .A1(\mem[2][4] ),
    .S(_1483_),
    .X(_2324_));
 sky130_fd_sc_hd__nand3_1 _4896_ (.A(_1540_),
    .B(_1542_),
    .C(_2324_),
    .Y(_2325_));
 sky130_fd_sc_hd__o22ai_1 _4897_ (.A1(_1740_),
    .A2(_1350_),
    .B1(_2325_),
    .B2(_1743_),
    .Y(_2326_));
 sky130_fd_sc_hd__nor2_1 _4898_ (.A(_1745_),
    .B(_2325_),
    .Y(_2327_));
 sky130_fd_sc_hd__o21ai_0 _4899_ (.A1(_1567_),
    .A2(_1359_),
    .B1(_0828_),
    .Y(_2328_));
 sky130_fd_sc_hd__o22ai_1 _4900_ (.A1(_1488_),
    .A2(_2326_),
    .B1(_2327_),
    .B2(_2328_),
    .Y(_2329_));
 sky130_fd_sc_hd__o211a_1 _4901_ (.A1(_1737_),
    .A2(_2323_),
    .B1(_2329_),
    .C1(_1509_),
    .X(_2330_));
 sky130_fd_sc_hd__mux2i_1 _4902_ (.A0(\mem[5][4] ),
    .A1(\mem[7][4] ),
    .S(_1510_),
    .Y(_2331_));
 sky130_fd_sc_hd__nor2_1 _4903_ (.A(_1530_),
    .B(_2331_),
    .Y(_2332_));
 sky130_fd_sc_hd__nor3_1 _4904_ (.A(_1752_),
    .B(_1489_),
    .C(_1360_),
    .Y(_2333_));
 sky130_fd_sc_hd__a311o_1 _4905_ (.A1(_1752_),
    .A2(_1627_),
    .A3(_1349_),
    .B1(_2332_),
    .C1(_2333_),
    .X(_2334_));
 sky130_fd_sc_hd__mux2i_1 _4906_ (.A0(\mem[1][4] ),
    .A1(\mem[3][4] ),
    .S(_1727_),
    .Y(_2335_));
 sky130_fd_sc_hd__nor2_1 _4907_ (.A(_1726_),
    .B(_2335_),
    .Y(_2336_));
 sky130_fd_sc_hd__o32ai_1 _4908_ (.A1(_1522_),
    .A2(_2334_),
    .A3(_2336_),
    .B1(_2537_),
    .B2(net107),
    .Y(_2337_));
 sky130_fd_sc_hd__a211oi_1 _4909_ (.A1(_2314_),
    .A2(_2322_),
    .B1(_2330_),
    .C1(_2337_),
    .Y(_0593_));
 sky130_fd_sc_hd__mux2i_1 _4910_ (.A0(\mem[5][5] ),
    .A1(\mem[7][5] ),
    .S(_2091_),
    .Y(_2338_));
 sky130_fd_sc_hd__nor2_1 _4911_ (.A(_1563_),
    .B(_2338_),
    .Y(_2339_));
 sky130_fd_sc_hd__a21oi_1 _4912_ (.A1(_1367_),
    .A2(_1526_),
    .B1(_2339_),
    .Y(_2340_));
 sky130_fd_sc_hd__mux2_1 _4913_ (.A0(\mem[1][5] ),
    .A1(\mem[3][5] ),
    .S(_2064_),
    .X(_2341_));
 sky130_fd_sc_hd__nand4_1 _4914_ (.A(_1568_),
    .B(_1569_),
    .C(_1478_),
    .D(_2341_),
    .Y(_2342_));
 sky130_fd_sc_hd__o31ai_1 _4915_ (.A1(_0860_),
    .A2(_1740_),
    .A3(_1376_),
    .B1(_2342_),
    .Y(_2343_));
 sky130_fd_sc_hd__mux2i_1 _4916_ (.A0(\mem[4][5] ),
    .A1(\mem[6][5] ),
    .S(_2098_),
    .Y(_2344_));
 sky130_fd_sc_hd__o221ai_1 _4917_ (.A1(_1368_),
    .A2(_1596_),
    .B1(_1580_),
    .B2(_2344_),
    .C1(_0906_),
    .Y(_2345_));
 sky130_fd_sc_hd__o21ai_0 _4918_ (.A1(_1552_),
    .A2(_2343_),
    .B1(_2345_),
    .Y(_2346_));
 sky130_fd_sc_hd__o22ai_1 _4919_ (.A1(\mem[2][5] ),
    .A2(_1462_),
    .B1(_1464_),
    .B2(\mem[3][5] ),
    .Y(_2347_));
 sky130_fd_sc_hd__o22ai_1 _4920_ (.A1(\mem[1][5] ),
    .A2(_1555_),
    .B1(_1556_),
    .B2(\mem[0][5] ),
    .Y(_2348_));
 sky130_fd_sc_hd__or3_1 _4921_ (.A(_2071_),
    .B(_2347_),
    .C(_2348_),
    .X(_2349_));
 sky130_fd_sc_hd__o2111ai_2 _4922_ (.A1(_1731_),
    .A2(_2340_),
    .B1(_2346_),
    .C1(_2349_),
    .D1(_1560_),
    .Y(_2350_));
 sky130_fd_sc_hd__mux2i_1 _4923_ (.A0(\mem[12][5] ),
    .A1(\mem[14][5] ),
    .S(_1738_),
    .Y(_2351_));
 sky130_fd_sc_hd__mux2_1 _4924_ (.A0(\mem[8][5] ),
    .A1(\mem[10][5] ),
    .S(_2108_),
    .X(_2352_));
 sky130_fd_sc_hd__nand3_1 _4925_ (.A(_1490_),
    .B(_1491_),
    .C(_2352_),
    .Y(_2353_));
 sky130_fd_sc_hd__o22ai_1 _4926_ (.A1(_2107_),
    .A2(_1379_),
    .B1(_2353_),
    .B2(_1743_),
    .Y(_2354_));
 sky130_fd_sc_hd__nor2_1 _4927_ (.A(_1745_),
    .B(_2353_),
    .Y(_2355_));
 sky130_fd_sc_hd__o21ai_0 _4928_ (.A1(_1519_),
    .A2(_1372_),
    .B1(_2140_),
    .Y(_2356_));
 sky130_fd_sc_hd__o22ai_1 _4929_ (.A1(_1514_),
    .A2(_2354_),
    .B1(_2355_),
    .B2(_2356_),
    .Y(_2357_));
 sky130_fd_sc_hd__o211ai_1 _4930_ (.A1(_1737_),
    .A2(_2351_),
    .B1(_2357_),
    .C1(_1501_),
    .Y(_2358_));
 sky130_fd_sc_hd__mux2i_1 _4931_ (.A0(\mem[13][5] ),
    .A1(\mem[15][5] ),
    .S(_1481_),
    .Y(_2359_));
 sky130_fd_sc_hd__nand3_1 _4932_ (.A(_2029_),
    .B(_1627_),
    .C(_1371_),
    .Y(_2360_));
 sky130_fd_sc_hd__o221ai_1 _4933_ (.A1(_1378_),
    .A2(_2084_),
    .B1(_2144_),
    .B2(_2359_),
    .C1(_2360_),
    .Y(_2361_));
 sky130_fd_sc_hd__mux2i_1 _4934_ (.A0(\mem[9][5] ),
    .A1(\mem[11][5] ),
    .S(_1550_),
    .Y(_2362_));
 sky130_fd_sc_hd__o21ai_0 _4935_ (.A1(_1588_),
    .A2(_2362_),
    .B1(_1475_),
    .Y(_2363_));
 sky130_fd_sc_hd__o22a_1 _4936_ (.A1(net108),
    .A2(_2027_),
    .B1(_2361_),
    .B2(_2363_),
    .X(_2364_));
 sky130_fd_sc_hd__and3_1 _4937_ (.A(_2350_),
    .B(_2358_),
    .C(_2364_),
    .X(_0594_));
 sky130_fd_sc_hd__mux2i_1 _4938_ (.A0(\mem[5][6] ),
    .A1(\mem[7][6] ),
    .S(_2091_),
    .Y(_2365_));
 sky130_fd_sc_hd__nor2_1 _4939_ (.A(_1563_),
    .B(_2365_),
    .Y(_2366_));
 sky130_fd_sc_hd__a21oi_1 _4940_ (.A1(_1384_),
    .A2(_1526_),
    .B1(_2366_),
    .Y(_2367_));
 sky130_fd_sc_hd__mux2_1 _4941_ (.A0(\mem[1][6] ),
    .A1(\mem[3][6] ),
    .S(_2064_),
    .X(_2368_));
 sky130_fd_sc_hd__nand4_1 _4942_ (.A(_1568_),
    .B(_1569_),
    .C(_1478_),
    .D(_2368_),
    .Y(_2369_));
 sky130_fd_sc_hd__o31ai_1 _4943_ (.A1(_0860_),
    .A2(_1740_),
    .A3(_1393_),
    .B1(_2369_),
    .Y(_2370_));
 sky130_fd_sc_hd__mux2i_1 _4944_ (.A0(\mem[4][6] ),
    .A1(\mem[6][6] ),
    .S(_2098_),
    .Y(_2371_));
 sky130_fd_sc_hd__o221ai_1 _4945_ (.A1(_1385_),
    .A2(_1596_),
    .B1(_1580_),
    .B2(_2371_),
    .C1(_0906_),
    .Y(_2372_));
 sky130_fd_sc_hd__o21ai_0 _4946_ (.A1(_1552_),
    .A2(_2370_),
    .B1(_2372_),
    .Y(_2373_));
 sky130_fd_sc_hd__o22ai_1 _4947_ (.A1(\mem[1][6] ),
    .A2(_1947_),
    .B1(_1948_),
    .B2(\mem[0][6] ),
    .Y(_2374_));
 sky130_fd_sc_hd__o22ai_1 _4948_ (.A1(\mem[2][6] ),
    .A2(_1767_),
    .B1(_1768_),
    .B2(\mem[3][6] ),
    .Y(_2375_));
 sky130_fd_sc_hd__or3_1 _4949_ (.A(_2071_),
    .B(_2374_),
    .C(_2375_),
    .X(_2376_));
 sky130_fd_sc_hd__o2111ai_1 _4950_ (.A1(_1731_),
    .A2(_2367_),
    .B1(_2373_),
    .C1(_2376_),
    .D1(_1560_),
    .Y(_2377_));
 sky130_fd_sc_hd__mux2i_1 _4951_ (.A0(\mem[12][6] ),
    .A1(\mem[14][6] ),
    .S(_1738_),
    .Y(_2378_));
 sky130_fd_sc_hd__mux2_1 _4952_ (.A0(\mem[8][6] ),
    .A1(\mem[10][6] ),
    .S(_2108_),
    .X(_2379_));
 sky130_fd_sc_hd__nand3_1 _4953_ (.A(_1490_),
    .B(_1491_),
    .C(_2379_),
    .Y(_2380_));
 sky130_fd_sc_hd__o22ai_1 _4954_ (.A1(_2107_),
    .A2(_1396_),
    .B1(_2380_),
    .B2(_1743_),
    .Y(_2381_));
 sky130_fd_sc_hd__nor2_1 _4955_ (.A(_1745_),
    .B(_2380_),
    .Y(_2382_));
 sky130_fd_sc_hd__o21ai_0 _4956_ (.A1(_1519_),
    .A2(_1389_),
    .B1(_2140_),
    .Y(_2383_));
 sky130_fd_sc_hd__o22ai_1 _4957_ (.A1(_1514_),
    .A2(_2381_),
    .B1(_2382_),
    .B2(_2383_),
    .Y(_2384_));
 sky130_fd_sc_hd__o211ai_1 _4958_ (.A1(_1737_),
    .A2(_2378_),
    .B1(_2384_),
    .C1(_1501_),
    .Y(_2385_));
 sky130_fd_sc_hd__mux2i_1 _4959_ (.A0(\mem[13][6] ),
    .A1(\mem[15][6] ),
    .S(_1481_),
    .Y(_2386_));
 sky130_fd_sc_hd__nand3_1 _4960_ (.A(_1538_),
    .B(_1627_),
    .C(_1388_),
    .Y(_2387_));
 sky130_fd_sc_hd__o221ai_1 _4961_ (.A1(_1395_),
    .A2(_2084_),
    .B1(_2144_),
    .B2(_2386_),
    .C1(_2387_),
    .Y(_2388_));
 sky130_fd_sc_hd__mux2i_1 _4962_ (.A0(\mem[9][6] ),
    .A1(\mem[11][6] ),
    .S(_1550_),
    .Y(_2389_));
 sky130_fd_sc_hd__o21ai_0 _4963_ (.A1(_1588_),
    .A2(_2389_),
    .B1(_1475_),
    .Y(_2390_));
 sky130_fd_sc_hd__o22a_1 _4964_ (.A1(net109),
    .A2(_0721_),
    .B1(_2388_),
    .B2(_2390_),
    .X(_2391_));
 sky130_fd_sc_hd__and3_1 _4965_ (.A(_2377_),
    .B(_2385_),
    .C(_2391_),
    .X(_0595_));
 sky130_fd_sc_hd__mux2i_1 _4966_ (.A0(\mem[5][7] ),
    .A1(\mem[7][7] ),
    .S(_2091_),
    .Y(_2392_));
 sky130_fd_sc_hd__nor2_1 _4967_ (.A(_1563_),
    .B(_2392_),
    .Y(_2393_));
 sky130_fd_sc_hd__a21oi_1 _4968_ (.A1(_1401_),
    .A2(_1526_),
    .B1(_2393_),
    .Y(_2394_));
 sky130_fd_sc_hd__mux2_1 _4969_ (.A0(\mem[1][7] ),
    .A1(\mem[3][7] ),
    .S(_1480_),
    .X(_2395_));
 sky130_fd_sc_hd__nand4_1 _4970_ (.A(_1568_),
    .B(_1569_),
    .C(_1478_),
    .D(_2395_),
    .Y(_2396_));
 sky130_fd_sc_hd__o31ai_1 _4971_ (.A1(_0860_),
    .A2(_1740_),
    .A3(_1410_),
    .B1(_2396_),
    .Y(_2397_));
 sky130_fd_sc_hd__mux2i_1 _4972_ (.A0(\mem[4][7] ),
    .A1(\mem[6][7] ),
    .S(_2098_),
    .Y(_2398_));
 sky130_fd_sc_hd__o221ai_1 _4973_ (.A1(_1402_),
    .A2(_1596_),
    .B1(_1580_),
    .B2(_2398_),
    .C1(_0906_),
    .Y(_2399_));
 sky130_fd_sc_hd__o21ai_0 _4974_ (.A1(_1552_),
    .A2(_2397_),
    .B1(_2399_),
    .Y(_2400_));
 sky130_fd_sc_hd__o22ai_1 _4975_ (.A1(\mem[1][7] ),
    .A2(_1455_),
    .B1(_1459_),
    .B2(\mem[0][7] ),
    .Y(_2401_));
 sky130_fd_sc_hd__o22ai_1 _4976_ (.A1(\mem[2][7] ),
    .A2(_1767_),
    .B1(_1768_),
    .B2(\mem[3][7] ),
    .Y(_2402_));
 sky130_fd_sc_hd__or3_1 _4977_ (.A(_1471_),
    .B(_2401_),
    .C(_2402_),
    .X(_2403_));
 sky130_fd_sc_hd__o2111ai_1 _4978_ (.A1(_1731_),
    .A2(_2394_),
    .B1(_2400_),
    .C1(_2403_),
    .D1(_1560_),
    .Y(_2404_));
 sky130_fd_sc_hd__mux2i_1 _4979_ (.A0(\mem[12][7] ),
    .A1(\mem[14][7] ),
    .S(_1738_),
    .Y(_2405_));
 sky130_fd_sc_hd__mux2_1 _4980_ (.A0(\mem[8][7] ),
    .A1(\mem[10][7] ),
    .S(_2108_),
    .X(_2406_));
 sky130_fd_sc_hd__nand3_1 _4981_ (.A(_1490_),
    .B(_1491_),
    .C(_2406_),
    .Y(_2407_));
 sky130_fd_sc_hd__o22ai_1 _4982_ (.A1(_2107_),
    .A2(_1413_),
    .B1(_2407_),
    .B2(_1743_),
    .Y(_2408_));
 sky130_fd_sc_hd__nor2_1 _4983_ (.A(_1745_),
    .B(_2407_),
    .Y(_2409_));
 sky130_fd_sc_hd__o21ai_0 _4984_ (.A1(_1519_),
    .A2(_1406_),
    .B1(_2140_),
    .Y(_2410_));
 sky130_fd_sc_hd__o22ai_1 _4985_ (.A1(_1514_),
    .A2(_2408_),
    .B1(_2409_),
    .B2(_2410_),
    .Y(_2411_));
 sky130_fd_sc_hd__o211ai_1 _4986_ (.A1(_1737_),
    .A2(_2405_),
    .B1(_2411_),
    .C1(_1501_),
    .Y(_2412_));
 sky130_fd_sc_hd__mux2i_1 _4987_ (.A0(\mem[13][7] ),
    .A1(\mem[15][7] ),
    .S(_1481_),
    .Y(_2413_));
 sky130_fd_sc_hd__nand3_1 _4988_ (.A(_1538_),
    .B(_1627_),
    .C(_1405_),
    .Y(_2414_));
 sky130_fd_sc_hd__o221ai_1 _4989_ (.A1(_1412_),
    .A2(_1494_),
    .B1(_2144_),
    .B2(_2413_),
    .C1(_2414_),
    .Y(_2415_));
 sky130_fd_sc_hd__mux2i_1 _4990_ (.A0(\mem[9][7] ),
    .A1(\mem[11][7] ),
    .S(_1550_),
    .Y(_2416_));
 sky130_fd_sc_hd__o21ai_0 _4991_ (.A1(_1588_),
    .A2(_2416_),
    .B1(_1475_),
    .Y(_2417_));
 sky130_fd_sc_hd__o22a_1 _4992_ (.A1(net110),
    .A2(_0721_),
    .B1(_2415_),
    .B2(_2417_),
    .X(_2418_));
 sky130_fd_sc_hd__and3_1 _4993_ (.A(_2404_),
    .B(_2412_),
    .C(_2418_),
    .X(_0596_));
 sky130_fd_sc_hd__mux2i_1 _4994_ (.A0(\mem[5][8] ),
    .A1(\mem[7][8] ),
    .S(_1608_),
    .Y(_2419_));
 sky130_fd_sc_hd__nor2_1 _4995_ (.A(_1563_),
    .B(_2419_),
    .Y(_2420_));
 sky130_fd_sc_hd__a21oi_1 _4996_ (.A1(_1418_),
    .A2(_1526_),
    .B1(_2420_),
    .Y(_2421_));
 sky130_fd_sc_hd__mux2_1 _4997_ (.A0(\mem[1][8] ),
    .A1(\mem[3][8] ),
    .S(_1480_),
    .X(_2422_));
 sky130_fd_sc_hd__nand4_1 _4998_ (.A(_1568_),
    .B(_1569_),
    .C(_1478_),
    .D(_2422_),
    .Y(_2423_));
 sky130_fd_sc_hd__o31ai_1 _4999_ (.A1(_0860_),
    .A2(_1740_),
    .A3(_1427_),
    .B1(_2423_),
    .Y(_2424_));
 sky130_fd_sc_hd__mux2i_1 _5000_ (.A0(\mem[4][8] ),
    .A1(\mem[6][8] ),
    .S(_1581_),
    .Y(_2425_));
 sky130_fd_sc_hd__o221ai_1 _5001_ (.A1(_1419_),
    .A2(_1596_),
    .B1(_1580_),
    .B2(_2425_),
    .C1(_0906_),
    .Y(_2426_));
 sky130_fd_sc_hd__o21ai_0 _5002_ (.A1(_1552_),
    .A2(_2424_),
    .B1(_2426_),
    .Y(_2427_));
 sky130_fd_sc_hd__o22ai_1 _5003_ (.A1(\mem[1][8] ),
    .A2(_1455_),
    .B1(_1459_),
    .B2(\mem[0][8] ),
    .Y(_2428_));
 sky130_fd_sc_hd__o22ai_1 _5004_ (.A1(\mem[2][8] ),
    .A2(_1767_),
    .B1(_1768_),
    .B2(\mem[3][8] ),
    .Y(_2429_));
 sky130_fd_sc_hd__or3_1 _5005_ (.A(_1471_),
    .B(_2428_),
    .C(_2429_),
    .X(_2430_));
 sky130_fd_sc_hd__o2111ai_1 _5006_ (.A1(_1731_),
    .A2(_2421_),
    .B1(_2427_),
    .C1(_2430_),
    .D1(_1560_),
    .Y(_2431_));
 sky130_fd_sc_hd__mux2i_1 _5007_ (.A0(\mem[12][8] ),
    .A1(\mem[14][8] ),
    .S(_1738_),
    .Y(_2432_));
 sky130_fd_sc_hd__mux2_1 _5008_ (.A0(\mem[8][8] ),
    .A1(\mem[10][8] ),
    .S(_1483_),
    .X(_2433_));
 sky130_fd_sc_hd__nand3_1 _5009_ (.A(_1490_),
    .B(_1491_),
    .C(_2433_),
    .Y(_2434_));
 sky130_fd_sc_hd__o22ai_1 _5010_ (.A1(_1539_),
    .A2(_1430_),
    .B1(_2434_),
    .B2(_1743_),
    .Y(_2435_));
 sky130_fd_sc_hd__nor2_1 _5011_ (.A(_1745_),
    .B(_2434_),
    .Y(_2436_));
 sky130_fd_sc_hd__o21ai_0 _5012_ (.A1(_1519_),
    .A2(_1423_),
    .B1(_2140_),
    .Y(_2437_));
 sky130_fd_sc_hd__o22ai_1 _5013_ (.A1(_1514_),
    .A2(_2435_),
    .B1(_2436_),
    .B2(_2437_),
    .Y(_2438_));
 sky130_fd_sc_hd__o211ai_1 _5014_ (.A1(_1737_),
    .A2(_2432_),
    .B1(_2438_),
    .C1(_1501_),
    .Y(_2439_));
 sky130_fd_sc_hd__mux2i_1 _5015_ (.A0(\mem[13][8] ),
    .A1(\mem[15][8] ),
    .S(_1481_),
    .Y(_2440_));
 sky130_fd_sc_hd__nand3_1 _5016_ (.A(_1538_),
    .B(_1627_),
    .C(_1422_),
    .Y(_2441_));
 sky130_fd_sc_hd__o221ai_1 _5017_ (.A1(_1429_),
    .A2(_1494_),
    .B1(_2144_),
    .B2(_2440_),
    .C1(_2441_),
    .Y(_2442_));
 sky130_fd_sc_hd__mux2i_1 _5018_ (.A0(\mem[9][8] ),
    .A1(\mem[11][8] ),
    .S(_1550_),
    .Y(_2443_));
 sky130_fd_sc_hd__o21ai_0 _5019_ (.A1(_1588_),
    .A2(_2443_),
    .B1(_1475_),
    .Y(_2444_));
 sky130_fd_sc_hd__o22a_1 _5020_ (.A1(net112),
    .A2(_0721_),
    .B1(_2442_),
    .B2(_2444_),
    .X(_2445_));
 sky130_fd_sc_hd__and3_1 _5021_ (.A(_2431_),
    .B(_2439_),
    .C(_2445_),
    .X(_0597_));
 sky130_fd_sc_hd__mux2i_1 _5022_ (.A0(\mem[13][9] ),
    .A1(\mem[15][9] ),
    .S(_1599_),
    .Y(_2446_));
 sky130_fd_sc_hd__o22ai_1 _5023_ (.A1(_1448_),
    .A2(_1597_),
    .B1(_1598_),
    .B2(_2446_),
    .Y(_2447_));
 sky130_fd_sc_hd__a211oi_1 _5024_ (.A1(_1595_),
    .A2(_2447_),
    .B1(_1593_),
    .C1(_2534_),
    .Y(_2448_));
 sky130_fd_sc_hd__mux2i_1 _5025_ (.A0(\mem[9][9] ),
    .A1(\mem[11][9] ),
    .S(_1599_),
    .Y(_2449_));
 sky130_fd_sc_hd__o221ai_1 _5026_ (.A1(_1439_),
    .A2(_1495_),
    .B1(_1589_),
    .B2(_2449_),
    .C1(_0903_),
    .Y(_2450_));
 sky130_fd_sc_hd__mux2i_1 _5027_ (.A0(\mem[12][9] ),
    .A1(\mem[14][9] ),
    .S(_1533_),
    .Y(_2451_));
 sky130_fd_sc_hd__o221ai_1 _5028_ (.A1(_1447_),
    .A2(_1548_),
    .B1(_1531_),
    .B2(_2451_),
    .C1(_1537_),
    .Y(_2452_));
 sky130_fd_sc_hd__o22ai_1 _5029_ (.A1(\mem[10][9] ),
    .A2(_1463_),
    .B1(_1465_),
    .B2(\mem[11][9] ),
    .Y(_2453_));
 sky130_fd_sc_hd__o22ai_1 _5030_ (.A1(\mem[9][9] ),
    .A2(_1456_),
    .B1(_1460_),
    .B2(\mem[8][9] ),
    .Y(_2454_));
 sky130_fd_sc_hd__nor3_1 _5031_ (.A(_1472_),
    .B(_2453_),
    .C(_2454_),
    .Y(_2455_));
 sky130_fd_sc_hd__a21oi_1 _5032_ (.A1(_2450_),
    .A2(_2452_),
    .B1(_2455_),
    .Y(_2456_));
 sky130_fd_sc_hd__mux2i_1 _5033_ (.A0(\mem[4][9] ),
    .A1(\mem[6][9] ),
    .S(_1727_),
    .Y(_2457_));
 sky130_fd_sc_hd__mux2_1 _5034_ (.A0(\mem[0][9] ),
    .A1(\mem[2][9] ),
    .S(_1483_),
    .X(_2458_));
 sky130_fd_sc_hd__nand3_1 _5035_ (.A(_1540_),
    .B(_1542_),
    .C(_2458_),
    .Y(_2459_));
 sky130_fd_sc_hd__o22ai_1 _5036_ (.A1(_1489_),
    .A2(_1436_),
    .B1(_2459_),
    .B2(_1467_),
    .Y(_2460_));
 sky130_fd_sc_hd__nor2_1 _5037_ (.A(_1468_),
    .B(_2459_),
    .Y(_2461_));
 sky130_fd_sc_hd__o21ai_0 _5038_ (.A1(_1567_),
    .A2(_1445_),
    .B1(_0828_),
    .Y(_2462_));
 sky130_fd_sc_hd__o22ai_1 _5039_ (.A1(_1488_),
    .A2(_2460_),
    .B1(_2461_),
    .B2(_2462_),
    .Y(_2463_));
 sky130_fd_sc_hd__o211a_1 _5040_ (.A1(_1598_),
    .A2(_2457_),
    .B1(_2463_),
    .C1(_1509_),
    .X(_2464_));
 sky130_fd_sc_hd__mux2i_1 _5041_ (.A0(\mem[5][9] ),
    .A1(\mem[7][9] ),
    .S(_1510_),
    .Y(_2465_));
 sky130_fd_sc_hd__nor2_1 _5042_ (.A(_1530_),
    .B(_2465_),
    .Y(_2466_));
 sky130_fd_sc_hd__nor3_1 _5043_ (.A(_0896_),
    .B(_1489_),
    .C(_1446_),
    .Y(_2467_));
 sky130_fd_sc_hd__a311o_1 _5044_ (.A1(_1752_),
    .A2(_0714_),
    .A3(_1435_),
    .B1(_2466_),
    .C1(_2467_),
    .X(_2468_));
 sky130_fd_sc_hd__mux2i_1 _5045_ (.A0(\mem[1][9] ),
    .A1(\mem[3][9] ),
    .S(_1727_),
    .Y(_2469_));
 sky130_fd_sc_hd__nor2_1 _5046_ (.A(_1726_),
    .B(_2469_),
    .Y(_2470_));
 sky130_fd_sc_hd__o32ai_1 _5047_ (.A1(_1522_),
    .A2(_2468_),
    .A3(_2470_),
    .B1(_2537_),
    .B2(net113),
    .Y(_2471_));
 sky130_fd_sc_hd__a211oi_1 _5048_ (.A1(_2448_),
    .A2(_2456_),
    .B1(_2464_),
    .C1(_2471_),
    .Y(_0598_));
 sky130_fd_sc_hd__mux2_1 _5049_ (.A0(_0533_),
    .A1(_1525_),
    .S(_0528_),
    .X(_0599_));
 sky130_fd_sc_hd__mux2_1 _5050_ (.A0(_0534_),
    .A1(_0907_),
    .S(_0528_),
    .X(_0600_));
 sky130_fd_sc_hd__nor2_1 _5051_ (.A(_2495_),
    .B(_0528_),
    .Y(_2472_));
 sky130_fd_sc_hd__xnor2_1 _5052_ (.A(_0898_),
    .B(_2472_),
    .Y(_0601_));
 sky130_fd_sc_hd__a21oi_1 _5053_ (.A1(_2539_),
    .A2(_2533_),
    .B1(_2532_),
    .Y(_2473_));
 sky130_fd_sc_hd__nor3_1 _5054_ (.A(_0897_),
    .B(_0528_),
    .C(_2473_),
    .Y(_2474_));
 sky130_fd_sc_hd__xor2_1 _5055_ (.A(_0867_),
    .B(_2474_),
    .X(_0602_));
 sky130_fd_sc_hd__mux2_1 _5056_ (.A0(_0531_),
    .A1(\wr_ptr[0] ),
    .S(_0530_),
    .X(_0603_));
 sky130_fd_sc_hd__mux2_1 _5057_ (.A0(_0532_),
    .A1(_0613_),
    .S(_0530_),
    .X(_0604_));
 sky130_fd_sc_hd__a21oi_1 _5058_ (.A1(_0613_),
    .A2(_2521_),
    .B1(_2530_),
    .Y(_2475_));
 sky130_fd_sc_hd__nor2_1 _5059_ (.A(_0530_),
    .B(_2475_),
    .Y(_2476_));
 sky130_fd_sc_hd__xor2_1 _5060_ (.A(_0622_),
    .B(_2476_),
    .X(_0605_));
 sky130_fd_sc_hd__nand2_1 _5061_ (.A(_2523_),
    .B(_2528_),
    .Y(_2477_));
 sky130_fd_sc_hd__nor2b_1 _5062_ (.A(_2523_),
    .B_N(_2528_),
    .Y(_2478_));
 sky130_fd_sc_hd__o21ai_0 _5063_ (.A1(_2521_),
    .A2(_2478_),
    .B1(_0613_),
    .Y(_2479_));
 sky130_fd_sc_hd__o21ai_0 _5064_ (.A1(_0613_),
    .A2(_2477_),
    .B1(_2479_),
    .Y(_2480_));
 sky130_fd_sc_hd__nand3b_1 _5065_ (.A_N(_0530_),
    .B(_2480_),
    .C(_0622_),
    .Y(_2481_));
 sky130_fd_sc_hd__xnor2_1 _5066_ (.A(_0621_),
    .B(_2481_),
    .Y(_0606_));
 sky130_fd_sc_hd__a32oi_1 _5067_ (.A1(_0609_),
    .A2(_2510_),
    .A3(_2548_),
    .B1(_2557_),
    .B2(_2546_),
    .Y(_2482_));
 sky130_fd_sc_hd__a21oi_1 _5068_ (.A1(_0609_),
    .A2(_0607_),
    .B1(_2482_),
    .Y(net69));
 sky130_fd_sc_hd__nand2_1 _5069_ (.A(_0607_),
    .B(net73),
    .Y(_2483_));
 sky130_fd_sc_hd__o22ai_1 _5070_ (.A1(_0607_),
    .A2(_0616_),
    .B1(_2483_),
    .B2(_2557_),
    .Y(_2484_));
 sky130_fd_sc_hd__nand2_1 _5071_ (.A(_0609_),
    .B(_2484_),
    .Y(_2485_));
 sky130_fd_sc_hd__o21ai_0 _5072_ (.A1(_2563_),
    .A2(_2557_),
    .B1(_2485_),
    .Y(net70));
 sky130_fd_sc_hd__nor4b_1 _5073_ (.A(_0609_),
    .B(_0607_),
    .C(net223),
    .D_N(_2548_),
    .Y(net76));
 sky130_fd_sc_hd__xor2_1 _5074_ (.A(_2556_),
    .B(_2499_),
    .X(\next_count[2] ));
 sky130_fd_sc_hd__a21o_1 _5075_ (.A1(_2496_),
    .A2(_2543_),
    .B1(_2542_),
    .X(_2486_));
 sky130_fd_sc_hd__a21oi_1 _5076_ (.A1(_2556_),
    .A2(_2486_),
    .B1(_2555_),
    .Y(_2487_));
 sky130_fd_sc_hd__xor2_1 _5077_ (.A(_2549_),
    .B(_2487_),
    .X(\next_count[3] ));
 sky130_fd_sc_hd__a21oi_1 _5078_ (.A1(_2556_),
    .A2(_2499_),
    .B1(_2555_),
    .Y(_2488_));
 sky130_fd_sc_hd__nor2_1 _5079_ (.A(_2549_),
    .B(_2488_),
    .Y(_2489_));
 sky130_fd_sc_hd__nor2_1 _5080_ (.A(_2550_),
    .B(_2489_),
    .Y(_2490_));
 sky130_fd_sc_hd__xor2_1 _5081_ (.A(_2490_),
    .B(_2558_),
    .X(\next_count[4] ));
 sky130_fd_sc_hd__nor2_1 _5082_ (.A(net77),
    .B(_0611_),
    .Y(net144));
 sky130_fd_sc_hd__nor2_1 _5083_ (.A(_0618_),
    .B(_0617_),
    .Y(_2491_));
 sky130_fd_sc_hd__nor3_1 _5084_ (.A(_2513_),
    .B(net77),
    .C(_2491_),
    .Y(net145));
 sky130_fd_sc_hd__fa_1 _5085_ (.A(_2492_),
    .B(_2493_),
    .CIN(_2494_),
    .COUT(_2495_),
    .SUM(_0534_));
 sky130_fd_sc_hd__fa_2 _5086_ (.A(_2496_),
    .B(_2497_),
    .CIN(_2498_),
    .COUT(_2499_),
    .SUM(\next_count[1] ));
 sky130_fd_sc_hd__ha_1 _5087_ (.A(_2500_),
    .B(_2501_),
    .COUT(_2502_),
    .SUM(_2503_));
 sky130_fd_sc_hd__ha_1 _5088_ (.A(_2500_),
    .B(\wr_ptr[1] ),
    .COUT(_2504_),
    .SUM(_2505_));
 sky130_fd_sc_hd__ha_1 _5089_ (.A(\wr_ptr[0] ),
    .B(_2501_),
    .COUT(_2506_),
    .SUM(_2507_));
 sky130_fd_sc_hd__ha_1 _5090_ (.A(\wr_ptr[0] ),
    .B(\wr_ptr[1] ),
    .COUT(_2508_),
    .SUM(_2509_));
 sky130_fd_sc_hd__ha_1 _5091_ (.A(_2510_),
    .B(_2511_),
    .COUT(_2512_),
    .SUM(_2513_));
 sky130_fd_sc_hd__ha_1 _5092_ (.A(_2514_),
    .B(_0529_),
    .COUT(_2515_),
    .SUM(_2516_));
 sky130_fd_sc_hd__ha_1 _5093_ (.A(\rd_ptr[0] ),
    .B(\rd_ptr[1] ),
    .COUT(_2517_),
    .SUM(_2518_));
 sky130_fd_sc_hd__ha_1 _5094_ (.A(_2519_),
    .B(_2520_),
    .COUT(_2521_),
    .SUM(_2522_));
 sky130_fd_sc_hd__ha_1 _5095_ (.A(_2519_),
    .B(_2520_),
    .COUT(_2523_),
    .SUM(_2524_));
 sky130_fd_sc_hd__ha_1 _5096_ (.A(_2525_),
    .B(_2526_),
    .COUT(_0530_),
    .SUM(_2527_));
 sky130_fd_sc_hd__ha_1 _5097_ (.A(_2528_),
    .B(_2529_),
    .COUT(_2530_),
    .SUM(_0532_));
 sky130_fd_sc_hd__ha_1 _5098_ (.A(\wr_ptr[0] ),
    .B(_2522_),
    .COUT(_2528_),
    .SUM(_0531_));
 sky130_fd_sc_hd__ha_1 _5099_ (.A(\rd_ptr[1] ),
    .B(_2531_),
    .COUT(_2532_),
    .SUM(_2533_));
 sky130_fd_sc_hd__ha_4 _5100_ (.A(_2534_),
    .B(_2535_),
    .COUT(_0528_),
    .SUM(_2536_));
 sky130_fd_sc_hd__ha_1 _5101_ (.A(_2537_),
    .B(_0529_),
    .COUT(_2531_),
    .SUM(_2538_));
 sky130_fd_sc_hd__ha_1 _5102_ (.A(\rd_ptr[0] ),
    .B(_2536_),
    .COUT(_2539_),
    .SUM(_0533_));
 sky130_fd_sc_hd__ha_1 _5103_ (.A(_2540_),
    .B(_2494_),
    .COUT(_2541_),
    .SUM(_2498_));
 sky130_fd_sc_hd__ha_1 _5104_ (.A(_2497_),
    .B(_2498_),
    .COUT(_2542_),
    .SUM(_2543_));
 sky130_fd_sc_hd__ha_1 _5105_ (.A(_2514_),
    .B(_2536_),
    .COUT(_2544_),
    .SUM(_2545_));
 sky130_fd_sc_hd__ha_1 _5106_ (.A(_2546_),
    .B(_2547_),
    .COUT(_2548_),
    .SUM(_2549_));
 sky130_fd_sc_hd__ha_1 _5107_ (.A(net73),
    .B(_2547_),
    .COUT(_2550_),
    .SUM(_2551_));
 sky130_fd_sc_hd__ha_1 _5108_ (.A(net73),
    .B(net169),
    .COUT(_2552_),
    .SUM(_2553_));
 sky130_fd_sc_hd__ha_1 _5109_ (.A(_2546_),
    .B(_2554_),
    .COUT(_2555_),
    .SUM(_2556_));
 sky130_fd_sc_hd__ha_4 _5110_ (.A(_2510_),
    .B(_2547_),
    .COUT(_2557_),
    .SUM(_2558_));
 sky130_fd_sc_hd__ha_1 _5111_ (.A(net167),
    .B(_2510_),
    .COUT(_2559_),
    .SUM(_2560_));
 sky130_fd_sc_hd__ha_1 _5112_ (.A(net167),
    .B(net168),
    .COUT(_2561_),
    .SUM(_2562_));
 sky130_fd_sc_hd__ha_1 _5113_ (.A(net169),
    .B(_2510_),
    .COUT(_2563_),
    .SUM(_2564_));
 sky130_fd_sc_hd__ha_1 _5114_ (.A(net170),
    .B(net168),
    .COUT(_2565_),
    .SUM(_2566_));
 sky130_fd_sc_hd__ha_1 _5115_ (.A(_2567_),
    .B(_2522_),
    .COUT(_2496_),
    .SUM(\next_count[0] ));
 sky130_fd_sc_hd__dfrtp_1 \fifo_count[0]$_DFF_PN0_  (.D(\next_count[0] ),
    .Q(net71),
    .RESET_B(net1),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_1 \fifo_count[1]$_DFF_PN0_  (.D(\next_count[1] ),
    .Q(net72),
    .RESET_B(net1),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_4 \fifo_count[2]$_DFF_PN0_  (.D(\next_count[2] ),
    .Q(net73),
    .RESET_B(net1),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_1 \fifo_count[3]$_DFF_PN0_  (.D(\next_count[3] ),
    .Q(net74),
    .RESET_B(net1),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_2 \fifo_count[4]$_DFF_PN0_  (.D(\next_count[4] ),
    .Q(net75),
    .RESET_B(net1),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][0]$_DFFE_PP_  (.D(_0016_),
    .DE(net217),
    .Q(\mem[0][0] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][10]$_DFFE_PP_  (.D(_0017_),
    .DE(net217),
    .Q(\mem[0][10] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][11]$_DFFE_PP_  (.D(_0018_),
    .DE(net217),
    .Q(\mem[0][11] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][12]$_DFFE_PP_  (.D(_0019_),
    .DE(net217),
    .Q(\mem[0][12] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][13]$_DFFE_PP_  (.D(_0020_),
    .DE(net217),
    .Q(\mem[0][13] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][14]$_DFFE_PP_  (.D(_0021_),
    .DE(net217),
    .Q(\mem[0][14] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][15]$_DFFE_PP_  (.D(_0022_),
    .DE(net217),
    .Q(\mem[0][15] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][16]$_DFFE_PP_  (.D(_0023_),
    .DE(_0015_),
    .Q(\mem[0][16] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][17]$_DFFE_PP_  (.D(_0024_),
    .DE(net217),
    .Q(\mem[0][17] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][18]$_DFFE_PP_  (.D(_0025_),
    .DE(_0015_),
    .Q(\mem[0][18] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][19]$_DFFE_PP_  (.D(_0026_),
    .DE(_0015_),
    .Q(\mem[0][19] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][1]$_DFFE_PP_  (.D(_0027_),
    .DE(net217),
    .Q(\mem[0][1] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][20]$_DFFE_PP_  (.D(_0028_),
    .DE(_0015_),
    .Q(\mem[0][20] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][21]$_DFFE_PP_  (.D(_0029_),
    .DE(_0015_),
    .Q(\mem[0][21] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][22]$_DFFE_PP_  (.D(_0030_),
    .DE(_0015_),
    .Q(\mem[0][22] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][23]$_DFFE_PP_  (.D(_0031_),
    .DE(_0015_),
    .Q(\mem[0][23] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][24]$_DFFE_PP_  (.D(_0032_),
    .DE(net217),
    .Q(\mem[0][24] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][25]$_DFFE_PP_  (.D(_0033_),
    .DE(_0015_),
    .Q(\mem[0][25] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][26]$_DFFE_PP_  (.D(_0034_),
    .DE(_0015_),
    .Q(\mem[0][26] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][27]$_DFFE_PP_  (.D(_0035_),
    .DE(_0015_),
    .Q(\mem[0][27] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][28]$_DFFE_PP_  (.D(_0036_),
    .DE(_0015_),
    .Q(\mem[0][28] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][29]$_DFFE_PP_  (.D(_0037_),
    .DE(net217),
    .Q(\mem[0][29] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][2]$_DFFE_PP_  (.D(_0038_),
    .DE(net217),
    .Q(\mem[0][2] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][30]$_DFFE_PP_  (.D(_0039_),
    .DE(_0015_),
    .Q(\mem[0][30] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][31]$_DFFE_PP_  (.D(_0040_),
    .DE(_0015_),
    .Q(\mem[0][31] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][3]$_DFFE_PP_  (.D(_0041_),
    .DE(_0015_),
    .Q(\mem[0][3] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][4]$_DFFE_PP_  (.D(_0042_),
    .DE(net217),
    .Q(\mem[0][4] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][5]$_DFFE_PP_  (.D(_0043_),
    .DE(net217),
    .Q(\mem[0][5] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][6]$_DFFE_PP_  (.D(_0044_),
    .DE(net217),
    .Q(\mem[0][6] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][7]$_DFFE_PP_  (.D(_0045_),
    .DE(net217),
    .Q(\mem[0][7] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][8]$_DFFE_PP_  (.D(_0046_),
    .DE(net217),
    .Q(\mem[0][8] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][9]$_DFFE_PP_  (.D(_0047_),
    .DE(net217),
    .Q(\mem[0][9] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][0]$_DFFE_PP_  (.D(net179),
    .DE(net152),
    .Q(\mem[10][0] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][10]$_DFFE_PP_  (.D(net183),
    .DE(net152),
    .Q(\mem[10][10] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][11]$_DFFE_PP_  (.D(_0050_),
    .DE(net152),
    .Q(\mem[10][11] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][12]$_DFFE_PP_  (.D(_0051_),
    .DE(net152),
    .Q(\mem[10][12] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][13]$_DFFE_PP_  (.D(_0052_),
    .DE(net152),
    .Q(\mem[10][13] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][14]$_DFFE_PP_  (.D(_0053_),
    .DE(_0014_),
    .Q(\mem[10][14] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][15]$_DFFE_PP_  (.D(_0054_),
    .DE(net152),
    .Q(\mem[10][15] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][16]$_DFFE_PP_  (.D(_0055_),
    .DE(_0014_),
    .Q(\mem[10][16] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][17]$_DFFE_PP_  (.D(_0056_),
    .DE(_0014_),
    .Q(\mem[10][17] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][18]$_DFFE_PP_  (.D(_0057_),
    .DE(_0014_),
    .Q(\mem[10][18] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][19]$_DFFE_PP_  (.D(_0058_),
    .DE(_0014_),
    .Q(\mem[10][19] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][1]$_DFFE_PP_  (.D(_0059_),
    .DE(net152),
    .Q(\mem[10][1] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][20]$_DFFE_PP_  (.D(_0060_),
    .DE(_0014_),
    .Q(\mem[10][20] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][21]$_DFFE_PP_  (.D(_0061_),
    .DE(_0014_),
    .Q(\mem[10][21] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][22]$_DFFE_PP_  (.D(_0062_),
    .DE(_0014_),
    .Q(\mem[10][22] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][23]$_DFFE_PP_  (.D(_0063_),
    .DE(_0014_),
    .Q(\mem[10][23] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][24]$_DFFE_PP_  (.D(_0064_),
    .DE(net152),
    .Q(\mem[10][24] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][25]$_DFFE_PP_  (.D(_0065_),
    .DE(_0014_),
    .Q(\mem[10][25] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][26]$_DFFE_PP_  (.D(_0066_),
    .DE(_0014_),
    .Q(\mem[10][26] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][27]$_DFFE_PP_  (.D(_0067_),
    .DE(_0014_),
    .Q(\mem[10][27] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][28]$_DFFE_PP_  (.D(_0068_),
    .DE(_0014_),
    .Q(\mem[10][28] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][29]$_DFFE_PP_  (.D(_0069_),
    .DE(net152),
    .Q(\mem[10][29] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][2]$_DFFE_PP_  (.D(_0070_),
    .DE(_0014_),
    .Q(\mem[10][2] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][30]$_DFFE_PP_  (.D(_0071_),
    .DE(_0014_),
    .Q(\mem[10][30] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][31]$_DFFE_PP_  (.D(_0072_),
    .DE(_0014_),
    .Q(\mem[10][31] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][3]$_DFFE_PP_  (.D(net212),
    .DE(net152),
    .Q(\mem[10][3] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][4]$_DFFE_PP_  (.D(_0074_),
    .DE(net152),
    .Q(\mem[10][4] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][5]$_DFFE_PP_  (.D(_0075_),
    .DE(net152),
    .Q(\mem[10][5] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][6]$_DFFE_PP_  (.D(_0076_),
    .DE(net152),
    .Q(\mem[10][6] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][7]$_DFFE_PP_  (.D(_0077_),
    .DE(net152),
    .Q(\mem[10][7] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][8]$_DFFE_PP_  (.D(_0078_),
    .DE(net152),
    .Q(\mem[10][8] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][9]$_DFFE_PP_  (.D(_0079_),
    .DE(net152),
    .Q(\mem[10][9] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][0]$_DFFE_PP_  (.D(_0080_),
    .DE(net150),
    .Q(\mem[11][0] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][10]$_DFFE_PP_  (.D(_0081_),
    .DE(net150),
    .Q(\mem[11][10] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][11]$_DFFE_PP_  (.D(_0082_),
    .DE(net150),
    .Q(\mem[11][11] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][12]$_DFFE_PP_  (.D(_0083_),
    .DE(net150),
    .Q(\mem[11][12] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][13]$_DFFE_PP_  (.D(net186),
    .DE(net150),
    .Q(\mem[11][13] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][14]$_DFFE_PP_  (.D(_0085_),
    .DE(net149),
    .Q(\mem[11][14] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][15]$_DFFE_PP_  (.D(_0086_),
    .DE(net150),
    .Q(\mem[11][15] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][16]$_DFFE_PP_  (.D(_0087_),
    .DE(net149),
    .Q(\mem[11][16] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][17]$_DFFE_PP_  (.D(_0088_),
    .DE(net149),
    .Q(\mem[11][17] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][18]$_DFFE_PP_  (.D(_0089_),
    .DE(net149),
    .Q(\mem[11][18] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][19]$_DFFE_PP_  (.D(_0090_),
    .DE(net149),
    .Q(\mem[11][19] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][1]$_DFFE_PP_  (.D(_0091_),
    .DE(net150),
    .Q(\mem[11][1] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][20]$_DFFE_PP_  (.D(_0092_),
    .DE(net149),
    .Q(\mem[11][20] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][21]$_DFFE_PP_  (.D(net196),
    .DE(net149),
    .Q(\mem[11][21] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][22]$_DFFE_PP_  (.D(_0094_),
    .DE(net149),
    .Q(\mem[11][22] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][23]$_DFFE_PP_  (.D(_0095_),
    .DE(net149),
    .Q(\mem[11][23] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][24]$_DFFE_PP_  (.D(_0096_),
    .DE(_0013_),
    .Q(\mem[11][24] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][25]$_DFFE_PP_  (.D(_0097_),
    .DE(net149),
    .Q(\mem[11][25] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][26]$_DFFE_PP_  (.D(_0098_),
    .DE(net149),
    .Q(\mem[11][26] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][27]$_DFFE_PP_  (.D(_0099_),
    .DE(net149),
    .Q(\mem[11][27] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][28]$_DFFE_PP_  (.D(_0100_),
    .DE(net149),
    .Q(\mem[11][28] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][29]$_DFFE_PP_  (.D(_0101_),
    .DE(_0013_),
    .Q(\mem[11][29] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][2]$_DFFE_PP_  (.D(_0102_),
    .DE(net149),
    .Q(\mem[11][2] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][30]$_DFFE_PP_  (.D(_0103_),
    .DE(net149),
    .Q(\mem[11][30] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][31]$_DFFE_PP_  (.D(_0104_),
    .DE(net149),
    .Q(\mem[11][31] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][3]$_DFFE_PP_  (.D(_0105_),
    .DE(_0013_),
    .Q(\mem[11][3] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][4]$_DFFE_PP_  (.D(_0106_),
    .DE(net150),
    .Q(\mem[11][4] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][5]$_DFFE_PP_  (.D(_0107_),
    .DE(net150),
    .Q(\mem[11][5] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][6]$_DFFE_PP_  (.D(_0108_),
    .DE(net150),
    .Q(\mem[11][6] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][7]$_DFFE_PP_  (.D(_0109_),
    .DE(net150),
    .Q(\mem[11][7] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][8]$_DFFE_PP_  (.D(_0110_),
    .DE(net150),
    .Q(\mem[11][8] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][9]$_DFFE_PP_  (.D(_0111_),
    .DE(net150),
    .Q(\mem[11][9] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][0]$_DFFE_PP_  (.D(_0112_),
    .DE(net154),
    .Q(\mem[12][0] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][10]$_DFFE_PP_  (.D(_0113_),
    .DE(net154),
    .Q(\mem[12][10] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][11]$_DFFE_PP_  (.D(_0114_),
    .DE(net154),
    .Q(\mem[12][11] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][12]$_DFFE_PP_  (.D(_0115_),
    .DE(net154),
    .Q(\mem[12][12] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][13]$_DFFE_PP_  (.D(_0116_),
    .DE(net154),
    .Q(\mem[12][13] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][14]$_DFFE_PP_  (.D(_0117_),
    .DE(net153),
    .Q(\mem[12][14] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][15]$_DFFE_PP_  (.D(_0118_),
    .DE(net154),
    .Q(\mem[12][15] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][16]$_DFFE_PP_  (.D(_0119_),
    .DE(net153),
    .Q(\mem[12][16] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][17]$_DFFE_PP_  (.D(_0120_),
    .DE(net153),
    .Q(\mem[12][17] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][18]$_DFFE_PP_  (.D(_0121_),
    .DE(net153),
    .Q(\mem[12][18] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][19]$_DFFE_PP_  (.D(_0122_),
    .DE(net153),
    .Q(\mem[12][19] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][1]$_DFFE_PP_  (.D(_0123_),
    .DE(net154),
    .Q(\mem[12][1] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][20]$_DFFE_PP_  (.D(_0124_),
    .DE(net153),
    .Q(\mem[12][20] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][21]$_DFFE_PP_  (.D(_0125_),
    .DE(net153),
    .Q(\mem[12][21] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][22]$_DFFE_PP_  (.D(_0126_),
    .DE(net153),
    .Q(\mem[12][22] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][23]$_DFFE_PP_  (.D(_0127_),
    .DE(net153),
    .Q(\mem[12][23] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][24]$_DFFE_PP_  (.D(_0128_),
    .DE(_0012_),
    .Q(\mem[12][24] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][25]$_DFFE_PP_  (.D(_0129_),
    .DE(net153),
    .Q(\mem[12][25] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][26]$_DFFE_PP_  (.D(_0130_),
    .DE(net153),
    .Q(\mem[12][26] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][27]$_DFFE_PP_  (.D(_0131_),
    .DE(net153),
    .Q(\mem[12][27] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][28]$_DFFE_PP_  (.D(_0132_),
    .DE(net153),
    .Q(\mem[12][28] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][29]$_DFFE_PP_  (.D(_0133_),
    .DE(_0012_),
    .Q(\mem[12][29] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][2]$_DFFE_PP_  (.D(_0134_),
    .DE(net153),
    .Q(\mem[12][2] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][30]$_DFFE_PP_  (.D(net202),
    .DE(net153),
    .Q(\mem[12][30] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][31]$_DFFE_PP_  (.D(_0136_),
    .DE(net153),
    .Q(\mem[12][31] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][3]$_DFFE_PP_  (.D(_0137_),
    .DE(net153),
    .Q(\mem[12][3] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][4]$_DFFE_PP_  (.D(_0138_),
    .DE(net154),
    .Q(\mem[12][4] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][5]$_DFFE_PP_  (.D(_0139_),
    .DE(net154),
    .Q(\mem[12][5] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][6]$_DFFE_PP_  (.D(_0140_),
    .DE(net154),
    .Q(\mem[12][6] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][7]$_DFFE_PP_  (.D(_0141_),
    .DE(net154),
    .Q(\mem[12][7] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][8]$_DFFE_PP_  (.D(_0142_),
    .DE(net154),
    .Q(\mem[12][8] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][9]$_DFFE_PP_  (.D(_0143_),
    .DE(net154),
    .Q(\mem[12][9] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][0]$_DFFE_PP_  (.D(_0144_),
    .DE(net155),
    .Q(\mem[13][0] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][10]$_DFFE_PP_  (.D(_0145_),
    .DE(net155),
    .Q(\mem[13][10] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][11]$_DFFE_PP_  (.D(_0146_),
    .DE(net155),
    .Q(\mem[13][11] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][12]$_DFFE_PP_  (.D(_0147_),
    .DE(net155),
    .Q(\mem[13][12] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][13]$_DFFE_PP_  (.D(_0148_),
    .DE(net155),
    .Q(\mem[13][13] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][14]$_DFFE_PP_  (.D(_0149_),
    .DE(net155),
    .Q(\mem[13][14] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][15]$_DFFE_PP_  (.D(_0150_),
    .DE(net155),
    .Q(\mem[13][15] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][16]$_DFFE_PP_  (.D(_0151_),
    .DE(_0011_),
    .Q(\mem[13][16] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][17]$_DFFE_PP_  (.D(_0152_),
    .DE(_0011_),
    .Q(\mem[13][17] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][18]$_DFFE_PP_  (.D(_0153_),
    .DE(_0011_),
    .Q(\mem[13][18] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][19]$_DFFE_PP_  (.D(_0154_),
    .DE(_0011_),
    .Q(\mem[13][19] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][1]$_DFFE_PP_  (.D(_0155_),
    .DE(net155),
    .Q(\mem[13][1] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][20]$_DFFE_PP_  (.D(_0156_),
    .DE(_0011_),
    .Q(\mem[13][20] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][21]$_DFFE_PP_  (.D(_0157_),
    .DE(_0011_),
    .Q(\mem[13][21] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][22]$_DFFE_PP_  (.D(_0158_),
    .DE(_0011_),
    .Q(\mem[13][22] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][23]$_DFFE_PP_  (.D(_0159_),
    .DE(_0011_),
    .Q(\mem[13][23] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][24]$_DFFE_PP_  (.D(_0160_),
    .DE(net155),
    .Q(\mem[13][24] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][25]$_DFFE_PP_  (.D(net206),
    .DE(_0011_),
    .Q(\mem[13][25] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][26]$_DFFE_PP_  (.D(net175),
    .DE(_0011_),
    .Q(\mem[13][26] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][27]$_DFFE_PP_  (.D(_0163_),
    .DE(_0011_),
    .Q(\mem[13][27] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][28]$_DFFE_PP_  (.D(_0164_),
    .DE(_0011_),
    .Q(\mem[13][28] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][29]$_DFFE_PP_  (.D(_0165_),
    .DE(net155),
    .Q(\mem[13][29] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][2]$_DFFE_PP_  (.D(_0166_),
    .DE(_0011_),
    .Q(\mem[13][2] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][30]$_DFFE_PP_  (.D(_0167_),
    .DE(_0011_),
    .Q(\mem[13][30] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][31]$_DFFE_PP_  (.D(_0168_),
    .DE(_0011_),
    .Q(\mem[13][31] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][3]$_DFFE_PP_  (.D(_0169_),
    .DE(_0011_),
    .Q(\mem[13][3] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][4]$_DFFE_PP_  (.D(_0170_),
    .DE(net155),
    .Q(\mem[13][4] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][5]$_DFFE_PP_  (.D(_0171_),
    .DE(net155),
    .Q(\mem[13][5] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][6]$_DFFE_PP_  (.D(_0172_),
    .DE(net155),
    .Q(\mem[13][6] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][7]$_DFFE_PP_  (.D(_0173_),
    .DE(net155),
    .Q(\mem[13][7] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][8]$_DFFE_PP_  (.D(_0174_),
    .DE(net155),
    .Q(\mem[13][8] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][9]$_DFFE_PP_  (.D(_0175_),
    .DE(net155),
    .Q(\mem[13][9] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][0]$_DFFE_PP_  (.D(_0176_),
    .DE(net157),
    .Q(\mem[14][0] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][10]$_DFFE_PP_  (.D(_0177_),
    .DE(net157),
    .Q(\mem[14][10] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][11]$_DFFE_PP_  (.D(_0178_),
    .DE(net157),
    .Q(\mem[14][11] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][12]$_DFFE_PP_  (.D(_0179_),
    .DE(net157),
    .Q(\mem[14][12] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][13]$_DFFE_PP_  (.D(_0180_),
    .DE(net157),
    .Q(\mem[14][13] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][14]$_DFFE_PP_  (.D(_0181_),
    .DE(net156),
    .Q(\mem[14][14] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][15]$_DFFE_PP_  (.D(_0182_),
    .DE(net157),
    .Q(\mem[14][15] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][16]$_DFFE_PP_  (.D(_0183_),
    .DE(net156),
    .Q(\mem[14][16] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][17]$_DFFE_PP_  (.D(_0184_),
    .DE(net156),
    .Q(\mem[14][17] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][18]$_DFFE_PP_  (.D(_0185_),
    .DE(net156),
    .Q(\mem[14][18] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][19]$_DFFE_PP_  (.D(_0186_),
    .DE(net156),
    .Q(\mem[14][19] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][1]$_DFFE_PP_  (.D(_0187_),
    .DE(net157),
    .Q(\mem[14][1] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][20]$_DFFE_PP_  (.D(_0188_),
    .DE(net156),
    .Q(\mem[14][20] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][21]$_DFFE_PP_  (.D(_0189_),
    .DE(net156),
    .Q(\mem[14][21] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][22]$_DFFE_PP_  (.D(_0190_),
    .DE(net156),
    .Q(\mem[14][22] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][23]$_DFFE_PP_  (.D(_0191_),
    .DE(net156),
    .Q(\mem[14][23] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][24]$_DFFE_PP_  (.D(_0192_),
    .DE(_0010_),
    .Q(\mem[14][24] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][25]$_DFFE_PP_  (.D(_0193_),
    .DE(net156),
    .Q(\mem[14][25] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][26]$_DFFE_PP_  (.D(_0194_),
    .DE(net156),
    .Q(\mem[14][26] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][27]$_DFFE_PP_  (.D(_0195_),
    .DE(net156),
    .Q(\mem[14][27] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][28]$_DFFE_PP_  (.D(_0196_),
    .DE(net156),
    .Q(\mem[14][28] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][29]$_DFFE_PP_  (.D(_0197_),
    .DE(_0010_),
    .Q(\mem[14][29] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][2]$_DFFE_PP_  (.D(_0198_),
    .DE(net156),
    .Q(\mem[14][2] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][30]$_DFFE_PP_  (.D(_0199_),
    .DE(net156),
    .Q(\mem[14][30] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][31]$_DFFE_PP_  (.D(_0200_),
    .DE(net156),
    .Q(\mem[14][31] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][3]$_DFFE_PP_  (.D(_0201_),
    .DE(net156),
    .Q(\mem[14][3] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][4]$_DFFE_PP_  (.D(net190),
    .DE(net157),
    .Q(\mem[14][4] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][5]$_DFFE_PP_  (.D(_0203_),
    .DE(net157),
    .Q(\mem[14][5] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][6]$_DFFE_PP_  (.D(_0204_),
    .DE(net157),
    .Q(\mem[14][6] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][7]$_DFFE_PP_  (.D(_0205_),
    .DE(net157),
    .Q(\mem[14][7] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][8]$_DFFE_PP_  (.D(_0206_),
    .DE(net157),
    .Q(\mem[14][8] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][9]$_DFFE_PP_  (.D(_0207_),
    .DE(net157),
    .Q(\mem[14][9] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][0]$_DFFE_PP_  (.D(_0208_),
    .DE(_0009_),
    .Q(\mem[15][0] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][10]$_DFFE_PP_  (.D(_0209_),
    .DE(_0009_),
    .Q(\mem[15][10] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][11]$_DFFE_PP_  (.D(_0210_),
    .DE(_0009_),
    .Q(\mem[15][11] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][12]$_DFFE_PP_  (.D(_0211_),
    .DE(_0009_),
    .Q(\mem[15][12] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][13]$_DFFE_PP_  (.D(_0212_),
    .DE(_0009_),
    .Q(\mem[15][13] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][14]$_DFFE_PP_  (.D(_0213_),
    .DE(_0009_),
    .Q(\mem[15][14] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][15]$_DFFE_PP_  (.D(_0214_),
    .DE(_0009_),
    .Q(\mem[15][15] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][16]$_DFFE_PP_  (.D(_0215_),
    .DE(net158),
    .Q(\mem[15][16] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][17]$_DFFE_PP_  (.D(_0216_),
    .DE(net158),
    .Q(\mem[15][17] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][18]$_DFFE_PP_  (.D(_0217_),
    .DE(net158),
    .Q(\mem[15][18] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][19]$_DFFE_PP_  (.D(_0218_),
    .DE(net158),
    .Q(\mem[15][19] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][1]$_DFFE_PP_  (.D(_0219_),
    .DE(_0009_),
    .Q(\mem[15][1] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][20]$_DFFE_PP_  (.D(_0220_),
    .DE(net158),
    .Q(\mem[15][20] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][21]$_DFFE_PP_  (.D(_0221_),
    .DE(net158),
    .Q(\mem[15][21] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][22]$_DFFE_PP_  (.D(_0222_),
    .DE(net158),
    .Q(\mem[15][22] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][23]$_DFFE_PP_  (.D(_0223_),
    .DE(net158),
    .Q(\mem[15][23] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][24]$_DFFE_PP_  (.D(_0224_),
    .DE(net158),
    .Q(\mem[15][24] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][25]$_DFFE_PP_  (.D(_0225_),
    .DE(net158),
    .Q(\mem[15][25] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][26]$_DFFE_PP_  (.D(_0226_),
    .DE(net158),
    .Q(\mem[15][26] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][27]$_DFFE_PP_  (.D(_0227_),
    .DE(net158),
    .Q(\mem[15][27] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][28]$_DFFE_PP_  (.D(_0228_),
    .DE(net158),
    .Q(\mem[15][28] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][29]$_DFFE_PP_  (.D(_0229_),
    .DE(net158),
    .Q(\mem[15][29] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][2]$_DFFE_PP_  (.D(_0230_),
    .DE(net158),
    .Q(\mem[15][2] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][30]$_DFFE_PP_  (.D(_0231_),
    .DE(net158),
    .Q(\mem[15][30] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][31]$_DFFE_PP_  (.D(_0232_),
    .DE(net158),
    .Q(\mem[15][31] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][3]$_DFFE_PP_  (.D(_0233_),
    .DE(net158),
    .Q(\mem[15][3] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][4]$_DFFE_PP_  (.D(_0234_),
    .DE(_0009_),
    .Q(\mem[15][4] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][5]$_DFFE_PP_  (.D(_0235_),
    .DE(_0009_),
    .Q(\mem[15][5] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][6]$_DFFE_PP_  (.D(_0236_),
    .DE(_0009_),
    .Q(\mem[15][6] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][7]$_DFFE_PP_  (.D(_0237_),
    .DE(_0009_),
    .Q(\mem[15][7] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][8]$_DFFE_PP_  (.D(_0238_),
    .DE(_0009_),
    .Q(\mem[15][8] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][9]$_DFFE_PP_  (.D(_0239_),
    .DE(_0009_),
    .Q(\mem[15][9] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][0]$_DFFE_PP_  (.D(_0240_),
    .DE(_0008_),
    .Q(\mem[1][0] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][10]$_DFFE_PP_  (.D(_0241_),
    .DE(net162),
    .Q(\mem[1][10] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][11]$_DFFE_PP_  (.D(_0242_),
    .DE(net162),
    .Q(\mem[1][11] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][12]$_DFFE_PP_  (.D(_0243_),
    .DE(net162),
    .Q(\mem[1][12] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][13]$_DFFE_PP_  (.D(_0244_),
    .DE(net162),
    .Q(\mem[1][13] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][14]$_DFFE_PP_  (.D(_0245_),
    .DE(net162),
    .Q(\mem[1][14] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][15]$_DFFE_PP_  (.D(_0246_),
    .DE(net162),
    .Q(\mem[1][15] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][16]$_DFFE_PP_  (.D(_0247_),
    .DE(net162),
    .Q(\mem[1][16] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][17]$_DFFE_PP_  (.D(_0248_),
    .DE(net162),
    .Q(\mem[1][17] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][18]$_DFFE_PP_  (.D(_0249_),
    .DE(net162),
    .Q(\mem[1][18] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][19]$_DFFE_PP_  (.D(_0250_),
    .DE(net162),
    .Q(\mem[1][19] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][1]$_DFFE_PP_  (.D(_0251_),
    .DE(_0008_),
    .Q(\mem[1][1] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][20]$_DFFE_PP_  (.D(_0252_),
    .DE(net162),
    .Q(\mem[1][20] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][21]$_DFFE_PP_  (.D(_0253_),
    .DE(net162),
    .Q(\mem[1][21] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][22]$_DFFE_PP_  (.D(_0254_),
    .DE(net162),
    .Q(\mem[1][22] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][23]$_DFFE_PP_  (.D(_0255_),
    .DE(_0008_),
    .Q(\mem[1][23] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][24]$_DFFE_PP_  (.D(_0256_),
    .DE(net162),
    .Q(\mem[1][24] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][25]$_DFFE_PP_  (.D(_0257_),
    .DE(_0008_),
    .Q(\mem[1][25] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][26]$_DFFE_PP_  (.D(_0258_),
    .DE(_0008_),
    .Q(\mem[1][26] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][27]$_DFFE_PP_  (.D(_0259_),
    .DE(_0008_),
    .Q(\mem[1][27] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][28]$_DFFE_PP_  (.D(_0260_),
    .DE(_0008_),
    .Q(\mem[1][28] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][29]$_DFFE_PP_  (.D(_0261_),
    .DE(net162),
    .Q(\mem[1][29] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][2]$_DFFE_PP_  (.D(_0262_),
    .DE(net162),
    .Q(\mem[1][2] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][30]$_DFFE_PP_  (.D(_0263_),
    .DE(_0008_),
    .Q(\mem[1][30] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][31]$_DFFE_PP_  (.D(_0264_),
    .DE(_0008_),
    .Q(\mem[1][31] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][3]$_DFFE_PP_  (.D(_0265_),
    .DE(_0008_),
    .Q(\mem[1][3] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][4]$_DFFE_PP_  (.D(_0266_),
    .DE(_0008_),
    .Q(\mem[1][4] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][5]$_DFFE_PP_  (.D(_0267_),
    .DE(_0008_),
    .Q(\mem[1][5] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][6]$_DFFE_PP_  (.D(_0268_),
    .DE(_0008_),
    .Q(\mem[1][6] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][7]$_DFFE_PP_  (.D(_0269_),
    .DE(_0008_),
    .Q(\mem[1][7] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][8]$_DFFE_PP_  (.D(_0270_),
    .DE(_0008_),
    .Q(\mem[1][8] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][9]$_DFFE_PP_  (.D(_0271_),
    .DE(_0008_),
    .Q(\mem[1][9] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][0]$_DFFE_PP_  (.D(_0272_),
    .DE(net218),
    .Q(\mem[2][0] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][10]$_DFFE_PP_  (.D(_0273_),
    .DE(net218),
    .Q(\mem[2][10] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][11]$_DFFE_PP_  (.D(_0274_),
    .DE(net218),
    .Q(\mem[2][11] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][12]$_DFFE_PP_  (.D(_0275_),
    .DE(net218),
    .Q(\mem[2][12] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][13]$_DFFE_PP_  (.D(_0276_),
    .DE(net218),
    .Q(\mem[2][13] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][14]$_DFFE_PP_  (.D(_0277_),
    .DE(net218),
    .Q(\mem[2][14] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][15]$_DFFE_PP_  (.D(_0278_),
    .DE(net218),
    .Q(\mem[2][15] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][16]$_DFFE_PP_  (.D(_0279_),
    .DE(_0007_),
    .Q(\mem[2][16] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][17]$_DFFE_PP_  (.D(_0280_),
    .DE(net218),
    .Q(\mem[2][17] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][18]$_DFFE_PP_  (.D(_0281_),
    .DE(_0007_),
    .Q(\mem[2][18] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][19]$_DFFE_PP_  (.D(_0282_),
    .DE(_0007_),
    .Q(\mem[2][19] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][1]$_DFFE_PP_  (.D(_0283_),
    .DE(net218),
    .Q(\mem[2][1] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][20]$_DFFE_PP_  (.D(_0284_),
    .DE(_0007_),
    .Q(\mem[2][20] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][21]$_DFFE_PP_  (.D(_0285_),
    .DE(_0007_),
    .Q(\mem[2][21] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][22]$_DFFE_PP_  (.D(_0286_),
    .DE(_0007_),
    .Q(\mem[2][22] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][23]$_DFFE_PP_  (.D(_0287_),
    .DE(_0007_),
    .Q(\mem[2][23] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][24]$_DFFE_PP_  (.D(_0288_),
    .DE(net218),
    .Q(\mem[2][24] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][25]$_DFFE_PP_  (.D(_0289_),
    .DE(_0007_),
    .Q(\mem[2][25] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][26]$_DFFE_PP_  (.D(_0290_),
    .DE(_0007_),
    .Q(\mem[2][26] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][27]$_DFFE_PP_  (.D(_0291_),
    .DE(_0007_),
    .Q(\mem[2][27] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][28]$_DFFE_PP_  (.D(_0292_),
    .DE(_0007_),
    .Q(\mem[2][28] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][29]$_DFFE_PP_  (.D(_0293_),
    .DE(net218),
    .Q(\mem[2][29] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][2]$_DFFE_PP_  (.D(_0294_),
    .DE(net218),
    .Q(\mem[2][2] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][30]$_DFFE_PP_  (.D(_0295_),
    .DE(_0007_),
    .Q(\mem[2][30] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][31]$_DFFE_PP_  (.D(_0296_),
    .DE(_0007_),
    .Q(\mem[2][31] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][3]$_DFFE_PP_  (.D(_0297_),
    .DE(_0007_),
    .Q(\mem[2][3] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][4]$_DFFE_PP_  (.D(_0298_),
    .DE(net218),
    .Q(\mem[2][4] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][5]$_DFFE_PP_  (.D(_0299_),
    .DE(net218),
    .Q(\mem[2][5] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][6]$_DFFE_PP_  (.D(_0300_),
    .DE(_0007_),
    .Q(\mem[2][6] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][7]$_DFFE_PP_  (.D(_0301_),
    .DE(net218),
    .Q(\mem[2][7] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][8]$_DFFE_PP_  (.D(_0302_),
    .DE(net218),
    .Q(\mem[2][8] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][9]$_DFFE_PP_  (.D(_0303_),
    .DE(net218),
    .Q(\mem[2][9] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][0]$_DFFE_PP_  (.D(_0304_),
    .DE(net160),
    .Q(\mem[3][0] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][10]$_DFFE_PP_  (.D(_0305_),
    .DE(net160),
    .Q(\mem[3][10] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][11]$_DFFE_PP_  (.D(_0306_),
    .DE(net160),
    .Q(\mem[3][11] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][12]$_DFFE_PP_  (.D(_0307_),
    .DE(net160),
    .Q(\mem[3][12] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][13]$_DFFE_PP_  (.D(_0308_),
    .DE(net159),
    .Q(\mem[3][13] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][14]$_DFFE_PP_  (.D(_0309_),
    .DE(net159),
    .Q(\mem[3][14] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][15]$_DFFE_PP_  (.D(_0310_),
    .DE(net160),
    .Q(\mem[3][15] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][16]$_DFFE_PP_  (.D(_0311_),
    .DE(net159),
    .Q(\mem[3][16] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][17]$_DFFE_PP_  (.D(_0312_),
    .DE(net159),
    .Q(\mem[3][17] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][18]$_DFFE_PP_  (.D(_0313_),
    .DE(net159),
    .Q(\mem[3][18] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][19]$_DFFE_PP_  (.D(_0314_),
    .DE(net159),
    .Q(\mem[3][19] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][1]$_DFFE_PP_  (.D(_0315_),
    .DE(net160),
    .Q(\mem[3][1] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][20]$_DFFE_PP_  (.D(_0316_),
    .DE(net159),
    .Q(\mem[3][20] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][21]$_DFFE_PP_  (.D(_0317_),
    .DE(net159),
    .Q(\mem[3][21] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][22]$_DFFE_PP_  (.D(_0318_),
    .DE(net159),
    .Q(\mem[3][22] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][23]$_DFFE_PP_  (.D(_0319_),
    .DE(_0006_),
    .Q(\mem[3][23] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][24]$_DFFE_PP_  (.D(_0320_),
    .DE(net159),
    .Q(\mem[3][24] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][25]$_DFFE_PP_  (.D(_0321_),
    .DE(_0006_),
    .Q(\mem[3][25] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][26]$_DFFE_PP_  (.D(_0322_),
    .DE(_0006_),
    .Q(\mem[3][26] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][27]$_DFFE_PP_  (.D(_0323_),
    .DE(_0006_),
    .Q(\mem[3][27] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][28]$_DFFE_PP_  (.D(_0324_),
    .DE(_0006_),
    .Q(\mem[3][28] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][29]$_DFFE_PP_  (.D(_0325_),
    .DE(net159),
    .Q(\mem[3][29] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][2]$_DFFE_PP_  (.D(_0326_),
    .DE(net159),
    .Q(\mem[3][2] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][30]$_DFFE_PP_  (.D(_0327_),
    .DE(_0006_),
    .Q(\mem[3][30] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][31]$_DFFE_PP_  (.D(_0328_),
    .DE(_0006_),
    .Q(\mem[3][31] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][3]$_DFFE_PP_  (.D(_0329_),
    .DE(_0006_),
    .Q(\mem[3][3] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][4]$_DFFE_PP_  (.D(_0330_),
    .DE(net160),
    .Q(\mem[3][4] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][5]$_DFFE_PP_  (.D(_0331_),
    .DE(net159),
    .Q(\mem[3][5] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][6]$_DFFE_PP_  (.D(_0332_),
    .DE(net160),
    .Q(\mem[3][6] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][7]$_DFFE_PP_  (.D(_0333_),
    .DE(net160),
    .Q(\mem[3][7] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][8]$_DFFE_PP_  (.D(_0334_),
    .DE(net160),
    .Q(\mem[3][8] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][9]$_DFFE_PP_  (.D(_0335_),
    .DE(net160),
    .Q(\mem[3][9] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][0]$_DFFE_PP_  (.D(_0336_),
    .DE(_0005_),
    .Q(\mem[4][0] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][10]$_DFFE_PP_  (.D(_0337_),
    .DE(_0005_),
    .Q(\mem[4][10] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][11]$_DFFE_PP_  (.D(_0338_),
    .DE(_0005_),
    .Q(\mem[4][11] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][12]$_DFFE_PP_  (.D(_0339_),
    .DE(_0005_),
    .Q(\mem[4][12] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][13]$_DFFE_PP_  (.D(_0340_),
    .DE(net148),
    .Q(\mem[4][13] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][14]$_DFFE_PP_  (.D(_0341_),
    .DE(net148),
    .Q(\mem[4][14] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][15]$_DFFE_PP_  (.D(_0342_),
    .DE(_0005_),
    .Q(\mem[4][15] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][16]$_DFFE_PP_  (.D(_0343_),
    .DE(net148),
    .Q(\mem[4][16] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][17]$_DFFE_PP_  (.D(_0344_),
    .DE(net148),
    .Q(\mem[4][17] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][18]$_DFFE_PP_  (.D(_0345_),
    .DE(net148),
    .Q(\mem[4][18] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][19]$_DFFE_PP_  (.D(_0346_),
    .DE(net148),
    .Q(\mem[4][19] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][1]$_DFFE_PP_  (.D(_0347_),
    .DE(_0005_),
    .Q(\mem[4][1] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][20]$_DFFE_PP_  (.D(_0348_),
    .DE(net148),
    .Q(\mem[4][20] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][21]$_DFFE_PP_  (.D(_0349_),
    .DE(net148),
    .Q(\mem[4][21] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][22]$_DFFE_PP_  (.D(_0350_),
    .DE(net148),
    .Q(\mem[4][22] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][23]$_DFFE_PP_  (.D(_0351_),
    .DE(net148),
    .Q(\mem[4][23] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][24]$_DFFE_PP_  (.D(_0352_),
    .DE(net148),
    .Q(\mem[4][24] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][25]$_DFFE_PP_  (.D(_0353_),
    .DE(net148),
    .Q(\mem[4][25] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][26]$_DFFE_PP_  (.D(_0354_),
    .DE(net148),
    .Q(\mem[4][26] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][27]$_DFFE_PP_  (.D(_0355_),
    .DE(net148),
    .Q(\mem[4][27] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][28]$_DFFE_PP_  (.D(_0356_),
    .DE(net148),
    .Q(\mem[4][28] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][29]$_DFFE_PP_  (.D(_0357_),
    .DE(_0005_),
    .Q(\mem[4][29] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][2]$_DFFE_PP_  (.D(_0358_),
    .DE(_0005_),
    .Q(\mem[4][2] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][30]$_DFFE_PP_  (.D(_0359_),
    .DE(net148),
    .Q(\mem[4][30] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][31]$_DFFE_PP_  (.D(_0360_),
    .DE(net148),
    .Q(\mem[4][31] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][3]$_DFFE_PP_  (.D(_0361_),
    .DE(_0005_),
    .Q(\mem[4][3] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][4]$_DFFE_PP_  (.D(_0362_),
    .DE(_0005_),
    .Q(\mem[4][4] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][5]$_DFFE_PP_  (.D(_0363_),
    .DE(_0005_),
    .Q(\mem[4][5] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][6]$_DFFE_PP_  (.D(_0364_),
    .DE(_0005_),
    .Q(\mem[4][6] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][7]$_DFFE_PP_  (.D(_0365_),
    .DE(_0005_),
    .Q(\mem[4][7] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][8]$_DFFE_PP_  (.D(_0366_),
    .DE(_0005_),
    .Q(\mem[4][8] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][9]$_DFFE_PP_  (.D(_0367_),
    .DE(_0005_),
    .Q(\mem[4][9] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][0]$_DFFE_PP_  (.D(_0368_),
    .DE(_0004_),
    .Q(\mem[5][0] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][10]$_DFFE_PP_  (.D(_0369_),
    .DE(_0004_),
    .Q(\mem[5][10] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][11]$_DFFE_PP_  (.D(_0370_),
    .DE(_0004_),
    .Q(\mem[5][11] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][12]$_DFFE_PP_  (.D(_0371_),
    .DE(_0004_),
    .Q(\mem[5][12] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][13]$_DFFE_PP_  (.D(_0372_),
    .DE(_0004_),
    .Q(\mem[5][13] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][14]$_DFFE_PP_  (.D(_0373_),
    .DE(net161),
    .Q(\mem[5][14] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][15]$_DFFE_PP_  (.D(_0374_),
    .DE(_0004_),
    .Q(\mem[5][15] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][16]$_DFFE_PP_  (.D(_0375_),
    .DE(net161),
    .Q(\mem[5][16] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][17]$_DFFE_PP_  (.D(_0376_),
    .DE(net161),
    .Q(\mem[5][17] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][18]$_DFFE_PP_  (.D(_0377_),
    .DE(net161),
    .Q(\mem[5][18] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][19]$_DFFE_PP_  (.D(_0378_),
    .DE(net161),
    .Q(\mem[5][19] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][1]$_DFFE_PP_  (.D(_0379_),
    .DE(_0004_),
    .Q(\mem[5][1] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][20]$_DFFE_PP_  (.D(_0380_),
    .DE(net161),
    .Q(\mem[5][20] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][21]$_DFFE_PP_  (.D(_0381_),
    .DE(net161),
    .Q(\mem[5][21] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][22]$_DFFE_PP_  (.D(_0382_),
    .DE(net161),
    .Q(\mem[5][22] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][23]$_DFFE_PP_  (.D(_0383_),
    .DE(net161),
    .Q(\mem[5][23] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][24]$_DFFE_PP_  (.D(_0384_),
    .DE(net161),
    .Q(\mem[5][24] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][25]$_DFFE_PP_  (.D(_0385_),
    .DE(net161),
    .Q(\mem[5][25] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][26]$_DFFE_PP_  (.D(_0386_),
    .DE(net161),
    .Q(\mem[5][26] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][27]$_DFFE_PP_  (.D(_0387_),
    .DE(net161),
    .Q(\mem[5][27] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][28]$_DFFE_PP_  (.D(_0388_),
    .DE(net161),
    .Q(\mem[5][28] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][29]$_DFFE_PP_  (.D(_0389_),
    .DE(net161),
    .Q(\mem[5][29] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][2]$_DFFE_PP_  (.D(_0390_),
    .DE(net161),
    .Q(\mem[5][2] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][30]$_DFFE_PP_  (.D(_0391_),
    .DE(net161),
    .Q(\mem[5][30] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][31]$_DFFE_PP_  (.D(_0392_),
    .DE(net161),
    .Q(\mem[5][31] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][3]$_DFFE_PP_  (.D(_0393_),
    .DE(net161),
    .Q(\mem[5][3] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][4]$_DFFE_PP_  (.D(_0394_),
    .DE(_0004_),
    .Q(\mem[5][4] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][5]$_DFFE_PP_  (.D(_0395_),
    .DE(_0004_),
    .Q(\mem[5][5] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][6]$_DFFE_PP_  (.D(_0396_),
    .DE(_0004_),
    .Q(\mem[5][6] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][7]$_DFFE_PP_  (.D(_0397_),
    .DE(_0004_),
    .Q(\mem[5][7] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][8]$_DFFE_PP_  (.D(_0398_),
    .DE(_0004_),
    .Q(\mem[5][8] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][9]$_DFFE_PP_  (.D(_0399_),
    .DE(_0004_),
    .Q(\mem[5][9] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][0]$_DFFE_PP_  (.D(_0400_),
    .DE(_0003_),
    .Q(\mem[6][0] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][10]$_DFFE_PP_  (.D(_0401_),
    .DE(_0003_),
    .Q(\mem[6][10] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][11]$_DFFE_PP_  (.D(_0402_),
    .DE(_0003_),
    .Q(\mem[6][11] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][12]$_DFFE_PP_  (.D(_0403_),
    .DE(_0003_),
    .Q(\mem[6][12] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][13]$_DFFE_PP_  (.D(_0404_),
    .DE(_0003_),
    .Q(\mem[6][13] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][14]$_DFFE_PP_  (.D(_0405_),
    .DE(net216),
    .Q(\mem[6][14] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][15]$_DFFE_PP_  (.D(_0406_),
    .DE(_0003_),
    .Q(\mem[6][15] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][16]$_DFFE_PP_  (.D(_0407_),
    .DE(net216),
    .Q(\mem[6][16] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][17]$_DFFE_PP_  (.D(_0408_),
    .DE(net216),
    .Q(\mem[6][17] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][18]$_DFFE_PP_  (.D(_0409_),
    .DE(net216),
    .Q(\mem[6][18] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][19]$_DFFE_PP_  (.D(_0410_),
    .DE(net216),
    .Q(\mem[6][19] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][1]$_DFFE_PP_  (.D(_0411_),
    .DE(_0003_),
    .Q(\mem[6][1] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][20]$_DFFE_PP_  (.D(_0412_),
    .DE(net216),
    .Q(\mem[6][20] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][21]$_DFFE_PP_  (.D(_0413_),
    .DE(net216),
    .Q(\mem[6][21] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][22]$_DFFE_PP_  (.D(_0414_),
    .DE(net216),
    .Q(\mem[6][22] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][23]$_DFFE_PP_  (.D(_0415_),
    .DE(net216),
    .Q(\mem[6][23] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][24]$_DFFE_PP_  (.D(_0416_),
    .DE(net216),
    .Q(\mem[6][24] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][25]$_DFFE_PP_  (.D(_0417_),
    .DE(net216),
    .Q(\mem[6][25] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][26]$_DFFE_PP_  (.D(_0418_),
    .DE(net216),
    .Q(\mem[6][26] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][27]$_DFFE_PP_  (.D(_0419_),
    .DE(net216),
    .Q(\mem[6][27] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][28]$_DFFE_PP_  (.D(_0420_),
    .DE(net216),
    .Q(\mem[6][28] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][29]$_DFFE_PP_  (.D(_0421_),
    .DE(_0003_),
    .Q(\mem[6][29] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][2]$_DFFE_PP_  (.D(_0422_),
    .DE(net216),
    .Q(\mem[6][2] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][30]$_DFFE_PP_  (.D(_0423_),
    .DE(net216),
    .Q(\mem[6][30] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][31]$_DFFE_PP_  (.D(_0424_),
    .DE(net216),
    .Q(\mem[6][31] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][3]$_DFFE_PP_  (.D(_0425_),
    .DE(net216),
    .Q(\mem[6][3] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][4]$_DFFE_PP_  (.D(_0426_),
    .DE(_0003_),
    .Q(\mem[6][4] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][5]$_DFFE_PP_  (.D(_0427_),
    .DE(_0003_),
    .Q(\mem[6][5] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][6]$_DFFE_PP_  (.D(_0428_),
    .DE(_0003_),
    .Q(\mem[6][6] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][7]$_DFFE_PP_  (.D(_0429_),
    .DE(_0003_),
    .Q(\mem[6][7] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][8]$_DFFE_PP_  (.D(_0430_),
    .DE(_0003_),
    .Q(\mem[6][8] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][9]$_DFFE_PP_  (.D(_0431_),
    .DE(_0003_),
    .Q(\mem[6][9] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][0]$_DFFE_PP_  (.D(_0432_),
    .DE(_0002_),
    .Q(\mem[7][0] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][10]$_DFFE_PP_  (.D(_0433_),
    .DE(_0002_),
    .Q(\mem[7][10] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][11]$_DFFE_PP_  (.D(_0434_),
    .DE(_0002_),
    .Q(\mem[7][11] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][12]$_DFFE_PP_  (.D(_0435_),
    .DE(_0002_),
    .Q(\mem[7][12] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][13]$_DFFE_PP_  (.D(_0436_),
    .DE(_0002_),
    .Q(\mem[7][13] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][14]$_DFFE_PP_  (.D(_0437_),
    .DE(net151),
    .Q(\mem[7][14] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][15]$_DFFE_PP_  (.D(_0438_),
    .DE(_0002_),
    .Q(\mem[7][15] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][16]$_DFFE_PP_  (.D(_0439_),
    .DE(net151),
    .Q(\mem[7][16] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][17]$_DFFE_PP_  (.D(_0440_),
    .DE(net151),
    .Q(\mem[7][17] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][18]$_DFFE_PP_  (.D(_0441_),
    .DE(net151),
    .Q(\mem[7][18] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][19]$_DFFE_PP_  (.D(_0442_),
    .DE(net151),
    .Q(\mem[7][19] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][1]$_DFFE_PP_  (.D(_0443_),
    .DE(_0002_),
    .Q(\mem[7][1] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][20]$_DFFE_PP_  (.D(_0444_),
    .DE(net151),
    .Q(\mem[7][20] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][21]$_DFFE_PP_  (.D(_0445_),
    .DE(net151),
    .Q(\mem[7][21] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][22]$_DFFE_PP_  (.D(_0446_),
    .DE(net151),
    .Q(\mem[7][22] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][23]$_DFFE_PP_  (.D(_0447_),
    .DE(net151),
    .Q(\mem[7][23] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][24]$_DFFE_PP_  (.D(_0448_),
    .DE(net151),
    .Q(\mem[7][24] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][25]$_DFFE_PP_  (.D(_0449_),
    .DE(net151),
    .Q(\mem[7][25] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][26]$_DFFE_PP_  (.D(_0450_),
    .DE(net151),
    .Q(\mem[7][26] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][27]$_DFFE_PP_  (.D(_0451_),
    .DE(net151),
    .Q(\mem[7][27] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][28]$_DFFE_PP_  (.D(_0452_),
    .DE(net151),
    .Q(\mem[7][28] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][29]$_DFFE_PP_  (.D(_0453_),
    .DE(net151),
    .Q(\mem[7][29] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][2]$_DFFE_PP_  (.D(_0454_),
    .DE(net151),
    .Q(\mem[7][2] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][30]$_DFFE_PP_  (.D(_0455_),
    .DE(net151),
    .Q(\mem[7][30] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][31]$_DFFE_PP_  (.D(_0456_),
    .DE(net151),
    .Q(\mem[7][31] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][3]$_DFFE_PP_  (.D(_0457_),
    .DE(net151),
    .Q(\mem[7][3] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][4]$_DFFE_PP_  (.D(_0458_),
    .DE(_0002_),
    .Q(\mem[7][4] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][5]$_DFFE_PP_  (.D(_0459_),
    .DE(_0002_),
    .Q(\mem[7][5] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][6]$_DFFE_PP_  (.D(_0460_),
    .DE(_0002_),
    .Q(\mem[7][6] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][7]$_DFFE_PP_  (.D(_0461_),
    .DE(_0002_),
    .Q(\mem[7][7] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][8]$_DFFE_PP_  (.D(_0462_),
    .DE(_0002_),
    .Q(\mem[7][8] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][9]$_DFFE_PP_  (.D(_0463_),
    .DE(_0002_),
    .Q(\mem[7][9] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][0]$_DFFE_PP_  (.D(_0464_),
    .DE(net147),
    .Q(\mem[8][0] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][10]$_DFFE_PP_  (.D(_0465_),
    .DE(net147),
    .Q(\mem[8][10] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][11]$_DFFE_PP_  (.D(_0466_),
    .DE(net147),
    .Q(\mem[8][11] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][12]$_DFFE_PP_  (.D(_0467_),
    .DE(net147),
    .Q(\mem[8][12] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][13]$_DFFE_PP_  (.D(_0468_),
    .DE(net147),
    .Q(\mem[8][13] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][14]$_DFFE_PP_  (.D(_0469_),
    .DE(_0001_),
    .Q(\mem[8][14] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][15]$_DFFE_PP_  (.D(_0470_),
    .DE(net147),
    .Q(\mem[8][15] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][16]$_DFFE_PP_  (.D(_0471_),
    .DE(_0001_),
    .Q(\mem[8][16] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][17]$_DFFE_PP_  (.D(_0472_),
    .DE(_0001_),
    .Q(\mem[8][17] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][18]$_DFFE_PP_  (.D(_0473_),
    .DE(_0001_),
    .Q(\mem[8][18] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][19]$_DFFE_PP_  (.D(_0474_),
    .DE(_0001_),
    .Q(\mem[8][19] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][1]$_DFFE_PP_  (.D(_0475_),
    .DE(net147),
    .Q(\mem[8][1] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][20]$_DFFE_PP_  (.D(_0476_),
    .DE(_0001_),
    .Q(\mem[8][20] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][21]$_DFFE_PP_  (.D(_0477_),
    .DE(_0001_),
    .Q(\mem[8][21] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][22]$_DFFE_PP_  (.D(_0478_),
    .DE(_0001_),
    .Q(\mem[8][22] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][23]$_DFFE_PP_  (.D(_0479_),
    .DE(_0001_),
    .Q(\mem[8][23] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][24]$_DFFE_PP_  (.D(_0480_),
    .DE(net147),
    .Q(\mem[8][24] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][25]$_DFFE_PP_  (.D(_0481_),
    .DE(_0001_),
    .Q(\mem[8][25] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][26]$_DFFE_PP_  (.D(_0482_),
    .DE(_0001_),
    .Q(\mem[8][26] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][27]$_DFFE_PP_  (.D(_0483_),
    .DE(_0001_),
    .Q(\mem[8][27] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][28]$_DFFE_PP_  (.D(_0484_),
    .DE(_0001_),
    .Q(\mem[8][28] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][29]$_DFFE_PP_  (.D(_0485_),
    .DE(net147),
    .Q(\mem[8][29] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][2]$_DFFE_PP_  (.D(_0486_),
    .DE(_0001_),
    .Q(\mem[8][2] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][30]$_DFFE_PP_  (.D(_0487_),
    .DE(_0001_),
    .Q(\mem[8][30] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][31]$_DFFE_PP_  (.D(_0488_),
    .DE(_0001_),
    .Q(\mem[8][31] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][3]$_DFFE_PP_  (.D(_0489_),
    .DE(_0001_),
    .Q(\mem[8][3] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][4]$_DFFE_PP_  (.D(_0490_),
    .DE(net147),
    .Q(\mem[8][4] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][5]$_DFFE_PP_  (.D(_0491_),
    .DE(net147),
    .Q(\mem[8][5] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][6]$_DFFE_PP_  (.D(_0492_),
    .DE(net147),
    .Q(\mem[8][6] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][7]$_DFFE_PP_  (.D(_0493_),
    .DE(net147),
    .Q(\mem[8][7] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][8]$_DFFE_PP_  (.D(_0494_),
    .DE(net147),
    .Q(\mem[8][8] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][9]$_DFFE_PP_  (.D(_0495_),
    .DE(net147),
    .Q(\mem[8][9] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][0]$_DFFE_PP_  (.D(_0496_),
    .DE(_0000_),
    .Q(\mem[9][0] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][10]$_DFFE_PP_  (.D(_0497_),
    .DE(_0000_),
    .Q(\mem[9][10] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][11]$_DFFE_PP_  (.D(_0498_),
    .DE(_0000_),
    .Q(\mem[9][11] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][12]$_DFFE_PP_  (.D(_0499_),
    .DE(_0000_),
    .Q(\mem[9][12] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][13]$_DFFE_PP_  (.D(_0500_),
    .DE(_0000_),
    .Q(\mem[9][13] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][14]$_DFFE_PP_  (.D(_0501_),
    .DE(net146),
    .Q(\mem[9][14] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][15]$_DFFE_PP_  (.D(_0502_),
    .DE(_0000_),
    .Q(\mem[9][15] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][16]$_DFFE_PP_  (.D(_0503_),
    .DE(net146),
    .Q(\mem[9][16] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][17]$_DFFE_PP_  (.D(_0504_),
    .DE(net146),
    .Q(\mem[9][17] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][18]$_DFFE_PP_  (.D(_0505_),
    .DE(net146),
    .Q(\mem[9][18] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][19]$_DFFE_PP_  (.D(_0506_),
    .DE(net146),
    .Q(\mem[9][19] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][1]$_DFFE_PP_  (.D(_0507_),
    .DE(_0000_),
    .Q(\mem[9][1] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][20]$_DFFE_PP_  (.D(_0508_),
    .DE(net146),
    .Q(\mem[9][20] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][21]$_DFFE_PP_  (.D(_0509_),
    .DE(net146),
    .Q(\mem[9][21] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][22]$_DFFE_PP_  (.D(_0510_),
    .DE(net146),
    .Q(\mem[9][22] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][23]$_DFFE_PP_  (.D(_0511_),
    .DE(net146),
    .Q(\mem[9][23] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][24]$_DFFE_PP_  (.D(_0512_),
    .DE(net146),
    .Q(\mem[9][24] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][25]$_DFFE_PP_  (.D(_0513_),
    .DE(net146),
    .Q(\mem[9][25] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][26]$_DFFE_PP_  (.D(_0514_),
    .DE(net146),
    .Q(\mem[9][26] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][27]$_DFFE_PP_  (.D(_0515_),
    .DE(net146),
    .Q(\mem[9][27] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][28]$_DFFE_PP_  (.D(_0516_),
    .DE(net146),
    .Q(\mem[9][28] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][29]$_DFFE_PP_  (.D(_0517_),
    .DE(net146),
    .Q(\mem[9][29] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][2]$_DFFE_PP_  (.D(_0518_),
    .DE(net146),
    .Q(\mem[9][2] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][30]$_DFFE_PP_  (.D(_0519_),
    .DE(net146),
    .Q(\mem[9][30] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][31]$_DFFE_PP_  (.D(_0520_),
    .DE(net146),
    .Q(\mem[9][31] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][3]$_DFFE_PP_  (.D(_0521_),
    .DE(net146),
    .Q(\mem[9][3] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][4]$_DFFE_PP_  (.D(_0522_),
    .DE(_0000_),
    .Q(\mem[9][4] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][5]$_DFFE_PP_  (.D(_0523_),
    .DE(_0000_),
    .Q(\mem[9][5] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][6]$_DFFE_PP_  (.D(_0524_),
    .DE(_0000_),
    .Q(\mem[9][6] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][7]$_DFFE_PP_  (.D(_0525_),
    .DE(_0000_),
    .Q(\mem[9][7] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][8]$_DFFE_PP_  (.D(_0526_),
    .DE(_0000_),
    .Q(\mem[9][8] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][9]$_DFFE_PP_  (.D(_0527_),
    .DE(_0000_),
    .Q(\mem[9][9] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][0]$_DFFE_PN0P_  (.D(_0535_),
    .Q(net78),
    .RESET_B(net1),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][10]$_DFFE_PN0P_  (.D(_0536_),
    .Q(net79),
    .RESET_B(net1),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][11]$_DFFE_PN0P_  (.D(_0537_),
    .Q(net80),
    .RESET_B(net1),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][12]$_DFFE_PN0P_  (.D(_0538_),
    .Q(net81),
    .RESET_B(net1),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][13]$_DFFE_PN0P_  (.D(_0539_),
    .Q(net82),
    .RESET_B(net1),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][14]$_DFFE_PN0P_  (.D(_0540_),
    .Q(net83),
    .RESET_B(net1),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][15]$_DFFE_PN0P_  (.D(_0541_),
    .Q(net84),
    .RESET_B(net1),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][16]$_DFFE_PN0P_  (.D(_0542_),
    .Q(net85),
    .RESET_B(net1),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][17]$_DFFE_PN0P_  (.D(_0543_),
    .Q(net86),
    .RESET_B(net1),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][18]$_DFFE_PN0P_  (.D(_0544_),
    .Q(net87),
    .RESET_B(net1),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][19]$_DFFE_PN0P_  (.D(_0545_),
    .Q(net88),
    .RESET_B(net1),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][1]$_DFFE_PN0P_  (.D(_0546_),
    .Q(net89),
    .RESET_B(net1),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][20]$_DFFE_PN0P_  (.D(_0547_),
    .Q(net90),
    .RESET_B(net1),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][21]$_DFFE_PN0P_  (.D(_0548_),
    .Q(net91),
    .RESET_B(net1),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][22]$_DFFE_PN0P_  (.D(_0549_),
    .Q(net92),
    .RESET_B(net1),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][23]$_DFFE_PN0P_  (.D(_0550_),
    .Q(net93),
    .RESET_B(net1),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][24]$_DFFE_PN0P_  (.D(_0551_),
    .Q(net94),
    .RESET_B(net1),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][25]$_DFFE_PN0P_  (.D(_0552_),
    .Q(net95),
    .RESET_B(net1),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][26]$_DFFE_PN0P_  (.D(_0553_),
    .Q(net96),
    .RESET_B(net1),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][27]$_DFFE_PN0P_  (.D(_0554_),
    .Q(net97),
    .RESET_B(net1),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][28]$_DFFE_PN0P_  (.D(_0555_),
    .Q(net98),
    .RESET_B(net1),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][29]$_DFFE_PN0P_  (.D(_0556_),
    .Q(net99),
    .RESET_B(net1),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][2]$_DFFE_PN0P_  (.D(_0557_),
    .Q(net100),
    .RESET_B(net1),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][30]$_DFFE_PN0P_  (.D(_0558_),
    .Q(net101),
    .RESET_B(net1),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][31]$_DFFE_PN0P_  (.D(_0559_),
    .Q(net102),
    .RESET_B(net1),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][3]$_DFFE_PN0P_  (.D(_0560_),
    .Q(net111),
    .RESET_B(net1),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][4]$_DFFE_PN0P_  (.D(_0561_),
    .Q(net122),
    .RESET_B(net1),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][5]$_DFFE_PN0P_  (.D(_0562_),
    .Q(net133),
    .RESET_B(net1),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][6]$_DFFE_PN0P_  (.D(_0563_),
    .Q(net138),
    .RESET_B(net1),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][7]$_DFFE_PN0P_  (.D(_0564_),
    .Q(net139),
    .RESET_B(net1),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][8]$_DFFE_PN0P_  (.D(_0565_),
    .Q(net140),
    .RESET_B(net1),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[0][9]$_DFFE_PN0P_  (.D(_0566_),
    .Q(net141),
    .RESET_B(net1),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][0]$_DFFE_PN0P_  (.D(_0567_),
    .Q(net103),
    .RESET_B(net1),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][10]$_DFFE_PN0P_  (.D(_0568_),
    .Q(net114),
    .RESET_B(net1),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][11]$_DFFE_PN0P_  (.D(_0569_),
    .Q(net115),
    .RESET_B(net1),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][12]$_DFFE_PN0P_  (.D(_0570_),
    .Q(net116),
    .RESET_B(net1),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][13]$_DFFE_PN0P_  (.D(_0571_),
    .Q(net117),
    .RESET_B(net1),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][14]$_DFFE_PN0P_  (.D(_0572_),
    .Q(net118),
    .RESET_B(net1),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][15]$_DFFE_PN0P_  (.D(_0573_),
    .Q(net119),
    .RESET_B(net1),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][16]$_DFFE_PN0P_  (.D(_0574_),
    .Q(net120),
    .RESET_B(net1),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][17]$_DFFE_PN0P_  (.D(_0575_),
    .Q(net121),
    .RESET_B(net1),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][18]$_DFFE_PN0P_  (.D(_0576_),
    .Q(net123),
    .RESET_B(net1),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][19]$_DFFE_PN0P_  (.D(_0577_),
    .Q(net124),
    .RESET_B(net1),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][1]$_DFFE_PN0P_  (.D(_0578_),
    .Q(net104),
    .RESET_B(net1),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][20]$_DFFE_PN0P_  (.D(_0579_),
    .Q(net125),
    .RESET_B(net1),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][21]$_DFFE_PN0P_  (.D(_0580_),
    .Q(net126),
    .RESET_B(net1),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][22]$_DFFE_PN0P_  (.D(_0581_),
    .Q(net127),
    .RESET_B(net1),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][23]$_DFFE_PN0P_  (.D(_0582_),
    .Q(net128),
    .RESET_B(net1),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_2 \rd_data_regs[1][24]$_DFFE_PN0P_  (.D(_0583_),
    .Q(net129),
    .RESET_B(net1),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][25]$_DFFE_PN0P_  (.D(_0584_),
    .Q(net130),
    .RESET_B(net1),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][26]$_DFFE_PN0P_  (.D(_0585_),
    .Q(net131),
    .RESET_B(net1),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][27]$_DFFE_PN0P_  (.D(_0586_),
    .Q(net132),
    .RESET_B(net1),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][28]$_DFFE_PN0P_  (.D(_0587_),
    .Q(net134),
    .RESET_B(net1),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_2 \rd_data_regs[1][29]$_DFFE_PN0P_  (.D(_0588_),
    .Q(net135),
    .RESET_B(net1),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][2]$_DFFE_PN0P_  (.D(_0589_),
    .Q(net105),
    .RESET_B(net1),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][30]$_DFFE_PN0P_  (.D(_0590_),
    .Q(net136),
    .RESET_B(net1),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][31]$_DFFE_PN0P_  (.D(_0591_),
    .Q(net137),
    .RESET_B(net1),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][3]$_DFFE_PN0P_  (.D(_0592_),
    .Q(net106),
    .RESET_B(net1),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][4]$_DFFE_PN0P_  (.D(_0593_),
    .Q(net107),
    .RESET_B(net1),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][5]$_DFFE_PN0P_  (.D(_0594_),
    .Q(net108),
    .RESET_B(net1),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][6]$_DFFE_PN0P_  (.D(_0595_),
    .Q(net109),
    .RESET_B(net1),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][7]$_DFFE_PN0P_  (.D(_0596_),
    .Q(net110),
    .RESET_B(net1),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][8]$_DFFE_PN0P_  (.D(_0597_),
    .Q(net112),
    .RESET_B(net1),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_regs[1][9]$_DFFE_PN0P_  (.D(_0598_),
    .Q(net113),
    .RESET_B(net1),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[0]$_DFFE_PN0N_  (.D(_0599_),
    .Q(\rd_ptr[0] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[1]$_DFFE_PN0N_  (.D(_0600_),
    .Q(\rd_ptr[1] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[2]$_DFFE_PN0N_  (.D(_0601_),
    .Q(\rd_ptr[2] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[3]$_DFFE_PN0N_  (.D(_0602_),
    .Q(\rd_ptr[3] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_valid_regs[0]$_DFF_PN0_  (.D(_0529_),
    .Q(net142),
    .RESET_B(net1),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_valid_regs[1]$_DFF_PN0_  (.D(_2537_),
    .Q(net143),
    .RESET_B(net1),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_4 \wr_ptr[0]$_DFFE_PN0N_  (.D(_0603_),
    .Q(\wr_ptr[0] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[1]$_DFFE_PN0N_  (.D(_0604_),
    .Q(\wr_ptr[1] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[2]$_DFFE_PN0N_  (.D(_0605_),
    .Q(\wr_ptr[2] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[3]$_DFFE_PN0N_  (.D(_0606_),
    .Q(\wr_ptr[3] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__buf_16 hold1 (.A(net171),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_872 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(rd_en[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(net178),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(net182),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(wr_data[11]),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(wr_data[12]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(net185),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(net184),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(wr_data[15]),
    .X(net9));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(wr_data[16]),
    .X(net10));
 sky130_fd_sc_hd__dlymetal6s2s_1 input10 (.A(wr_data[17]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(net172),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(wr_data[19]),
    .X(net13));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(wr_data[1]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input14 (.A(wr_data[20]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(net195),
    .X(net16));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(wr_data[22]),
    .X(net17));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(wr_data[23]),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input18 (.A(net210),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(net205),
    .X(net20));
 sky130_fd_sc_hd__dlymetal6s2s_1 input20 (.A(net176),
    .X(net21));
 sky130_fd_sc_hd__dlymetal6s2s_1 input21 (.A(wr_data[27]),
    .X(net22));
 sky130_fd_sc_hd__dlymetal6s2s_1 input22 (.A(wr_data[28]),
    .X(net23));
 sky130_fd_sc_hd__buf_2 input23 (.A(net215),
    .X(net24));
 sky130_fd_sc_hd__dlymetal6s2s_1 input24 (.A(wr_data[2]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(net208),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 input26 (.A(wr_data[31]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(net181),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(net204),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(net209),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(net211),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(net192),
    .X(net32));
 sky130_fd_sc_hd__dlymetal6s2s_1 input32 (.A(wr_data[37]),
    .X(net33));
 sky130_fd_sc_hd__dlymetal6s2s_1 input33 (.A(wr_data[38]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(net177),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(net214),
    .X(net36));
 sky130_fd_sc_hd__dlymetal6s2s_1 input36 (.A(wr_data[40]),
    .X(net37));
 sky130_fd_sc_hd__dlymetal6s2s_1 input37 (.A(wr_data[41]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(net187),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(net203),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(net193),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(net191),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(net188),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(net199),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(net180),
    .X(net45));
 sky130_fd_sc_hd__dlymetal6s2s_1 input45 (.A(wr_data[49]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(net189),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(net173),
    .X(net48));
 sky130_fd_sc_hd__dlymetal6s2s_1 input48 (.A(wr_data[51]),
    .X(net49));
 sky130_fd_sc_hd__dlymetal6s2s_1 input49 (.A(wr_data[52]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(net197),
    .X(net51));
 sky130_fd_sc_hd__dlymetal6s2s_1 input51 (.A(wr_data[54]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(net200),
    .X(net53));
 sky130_fd_sc_hd__buf_2 input53 (.A(net213),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(net207),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(net174),
    .X(net56));
 sky130_fd_sc_hd__dlymetal6s2s_1 input56 (.A(wr_data[59]),
    .X(net57));
 sky130_fd_sc_hd__dlymetal6s2s_1 input57 (.A(wr_data[5]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(net198),
    .X(net59));
 sky130_fd_sc_hd__buf_2 input59 (.A(wr_data[61]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(net201),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(net194),
    .X(net62));
 sky130_fd_sc_hd__dlymetal6s2s_1 input62 (.A(wr_data[6]),
    .X(net63));
 sky130_fd_sc_hd__dlymetal6s2s_1 input63 (.A(wr_data[7]),
    .X(net64));
 sky130_fd_sc_hd__dlymetal6s2s_1 input64 (.A(wr_data[8]),
    .X(net65));
 sky130_fd_sc_hd__dlymetal6s2s_1 input65 (.A(wr_data[9]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(wr_en[0]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(wr_en[1]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net69),
    .X(almost_empty));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(net70),
    .X(almost_full));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net71),
    .X(data_count[0]));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(net72),
    .X(data_count[1]));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(net73),
    .X(data_count[2]));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(net74),
    .X(data_count[3]));
 sky130_fd_sc_hd__clkbuf_1 output74 (.A(net223),
    .X(data_count[4]));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(net76),
    .X(empty));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(net77),
    .X(full));
 sky130_fd_sc_hd__clkbuf_1 output77 (.A(net78),
    .X(rd_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(net79),
    .X(rd_data[10]));
 sky130_fd_sc_hd__clkbuf_1 output79 (.A(net80),
    .X(rd_data[11]));
 sky130_fd_sc_hd__clkbuf_1 output80 (.A(net81),
    .X(rd_data[12]));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(net82),
    .X(rd_data[13]));
 sky130_fd_sc_hd__clkbuf_1 output82 (.A(net83),
    .X(rd_data[14]));
 sky130_fd_sc_hd__clkbuf_1 output83 (.A(net84),
    .X(rd_data[15]));
 sky130_fd_sc_hd__clkbuf_1 output84 (.A(net85),
    .X(rd_data[16]));
 sky130_fd_sc_hd__clkbuf_1 output85 (.A(net86),
    .X(rd_data[17]));
 sky130_fd_sc_hd__clkbuf_1 output86 (.A(net87),
    .X(rd_data[18]));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(net88),
    .X(rd_data[19]));
 sky130_fd_sc_hd__clkbuf_1 output88 (.A(net89),
    .X(rd_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(net90),
    .X(rd_data[20]));
 sky130_fd_sc_hd__clkbuf_1 output90 (.A(net91),
    .X(rd_data[21]));
 sky130_fd_sc_hd__clkbuf_1 output91 (.A(net92),
    .X(rd_data[22]));
 sky130_fd_sc_hd__clkbuf_1 output92 (.A(net93),
    .X(rd_data[23]));
 sky130_fd_sc_hd__clkbuf_1 output93 (.A(net94),
    .X(rd_data[24]));
 sky130_fd_sc_hd__clkbuf_1 output94 (.A(net95),
    .X(rd_data[25]));
 sky130_fd_sc_hd__clkbuf_1 output95 (.A(net96),
    .X(rd_data[26]));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(net97),
    .X(rd_data[27]));
 sky130_fd_sc_hd__clkbuf_1 output97 (.A(net98),
    .X(rd_data[28]));
 sky130_fd_sc_hd__clkbuf_1 output98 (.A(net99),
    .X(rd_data[29]));
 sky130_fd_sc_hd__clkbuf_1 output99 (.A(net100),
    .X(rd_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output100 (.A(net101),
    .X(rd_data[30]));
 sky130_fd_sc_hd__clkbuf_1 output101 (.A(net102),
    .X(rd_data[31]));
 sky130_fd_sc_hd__clkbuf_1 output102 (.A(net103),
    .X(rd_data[32]));
 sky130_fd_sc_hd__clkbuf_1 output103 (.A(net104),
    .X(rd_data[33]));
 sky130_fd_sc_hd__clkbuf_1 output104 (.A(net105),
    .X(rd_data[34]));
 sky130_fd_sc_hd__clkbuf_1 output105 (.A(net106),
    .X(rd_data[35]));
 sky130_fd_sc_hd__clkbuf_1 output106 (.A(net107),
    .X(rd_data[36]));
 sky130_fd_sc_hd__clkbuf_1 output107 (.A(net108),
    .X(rd_data[37]));
 sky130_fd_sc_hd__clkbuf_1 output108 (.A(net109),
    .X(rd_data[38]));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(net110),
    .X(rd_data[39]));
 sky130_fd_sc_hd__clkbuf_1 output110 (.A(net111),
    .X(rd_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output111 (.A(net112),
    .X(rd_data[40]));
 sky130_fd_sc_hd__clkbuf_1 output112 (.A(net113),
    .X(rd_data[41]));
 sky130_fd_sc_hd__clkbuf_1 output113 (.A(net114),
    .X(rd_data[42]));
 sky130_fd_sc_hd__clkbuf_1 output114 (.A(net115),
    .X(rd_data[43]));
 sky130_fd_sc_hd__clkbuf_1 output115 (.A(net116),
    .X(rd_data[44]));
 sky130_fd_sc_hd__clkbuf_1 output116 (.A(net117),
    .X(rd_data[45]));
 sky130_fd_sc_hd__clkbuf_1 output117 (.A(net118),
    .X(rd_data[46]));
 sky130_fd_sc_hd__clkbuf_1 output118 (.A(net119),
    .X(rd_data[47]));
 sky130_fd_sc_hd__clkbuf_1 output119 (.A(net120),
    .X(rd_data[48]));
 sky130_fd_sc_hd__clkbuf_1 output120 (.A(net121),
    .X(rd_data[49]));
 sky130_fd_sc_hd__clkbuf_1 output121 (.A(net122),
    .X(rd_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output122 (.A(net123),
    .X(rd_data[50]));
 sky130_fd_sc_hd__clkbuf_1 output123 (.A(net124),
    .X(rd_data[51]));
 sky130_fd_sc_hd__clkbuf_1 output124 (.A(net125),
    .X(rd_data[52]));
 sky130_fd_sc_hd__clkbuf_1 output125 (.A(net126),
    .X(rd_data[53]));
 sky130_fd_sc_hd__clkbuf_1 output126 (.A(net127),
    .X(rd_data[54]));
 sky130_fd_sc_hd__clkbuf_1 output127 (.A(net128),
    .X(rd_data[55]));
 sky130_fd_sc_hd__clkbuf_1 output128 (.A(net129),
    .X(rd_data[56]));
 sky130_fd_sc_hd__clkbuf_1 output129 (.A(net130),
    .X(rd_data[57]));
 sky130_fd_sc_hd__clkbuf_1 output130 (.A(net131),
    .X(rd_data[58]));
 sky130_fd_sc_hd__clkbuf_1 output131 (.A(net132),
    .X(rd_data[59]));
 sky130_fd_sc_hd__clkbuf_1 output132 (.A(net133),
    .X(rd_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output133 (.A(net134),
    .X(rd_data[60]));
 sky130_fd_sc_hd__clkbuf_1 output134 (.A(net135),
    .X(rd_data[61]));
 sky130_fd_sc_hd__clkbuf_1 output135 (.A(net136),
    .X(rd_data[62]));
 sky130_fd_sc_hd__clkbuf_1 output136 (.A(net137),
    .X(rd_data[63]));
 sky130_fd_sc_hd__clkbuf_1 output137 (.A(net138),
    .X(rd_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output138 (.A(net139),
    .X(rd_data[7]));
 sky130_fd_sc_hd__clkbuf_1 output139 (.A(net140),
    .X(rd_data[8]));
 sky130_fd_sc_hd__clkbuf_1 output140 (.A(net141),
    .X(rd_data[9]));
 sky130_fd_sc_hd__clkbuf_1 output141 (.A(net142),
    .X(rd_valid[0]));
 sky130_fd_sc_hd__clkbuf_1 output142 (.A(net143),
    .X(rd_valid[1]));
 sky130_fd_sc_hd__clkbuf_1 output143 (.A(net144),
    .X(wr_ready[0]));
 sky130_fd_sc_hd__clkbuf_1 output144 (.A(net145),
    .X(wr_ready[1]));
 sky130_fd_sc_hd__buf_12 max_cap145 (.A(_0000_),
    .X(net146));
 sky130_fd_sc_hd__buf_16 max_cap146 (.A(_0001_),
    .X(net147));
 sky130_fd_sc_hd__buf_16 load_slew147 (.A(_0005_),
    .X(net148));
 sky130_fd_sc_hd__buf_16 load_slew148 (.A(_0013_),
    .X(net149));
 sky130_fd_sc_hd__buf_16 load_slew149 (.A(_0013_),
    .X(net150));
 sky130_fd_sc_hd__buf_12 max_cap150 (.A(_0002_),
    .X(net151));
 sky130_fd_sc_hd__buf_12 max_cap151 (.A(_0014_),
    .X(net152));
 sky130_fd_sc_hd__buf_16 load_slew152 (.A(_0012_),
    .X(net153));
 sky130_fd_sc_hd__buf_16 load_slew153 (.A(_0012_),
    .X(net154));
 sky130_fd_sc_hd__buf_12 wire154 (.A(_0011_),
    .X(net155));
 sky130_fd_sc_hd__buf_16 load_slew155 (.A(_0010_),
    .X(net156));
 sky130_fd_sc_hd__buf_16 load_slew156 (.A(_0010_),
    .X(net157));
 sky130_fd_sc_hd__buf_12 wire157 (.A(_0009_),
    .X(net158));
 sky130_fd_sc_hd__buf_16 load_slew158 (.A(net160),
    .X(net159));
 sky130_fd_sc_hd__buf_16 load_slew159 (.A(_0006_),
    .X(net160));
 sky130_fd_sc_hd__buf_16 max_cap160 (.A(_0004_),
    .X(net161));
 sky130_fd_sc_hd__buf_16 load_slew161 (.A(_0008_),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload0 (.A(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload1 (.A(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkinv_8 clkload2 (.A(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload3 (.A(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload4 (.A(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload5 (.A(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload6 (.A(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload7 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload8 (.A(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload9 (.A(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload10 (.A(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkinv_1 clkload11 (.A(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkinv_2 clkload12 (.A(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload13 (.A(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkinv_2 clkload14 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload15 (.A(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload16 (.A(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkinv_2 clkload17 (.A(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload18 (.A(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload19 (.A(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkinv_2 clkload20 (.A(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkinv_2 clkload21 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload22 (.A(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkinv_2 clkload23 (.A(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkinv_1 clkload24 (.A(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkinv_2 clkload25 (.A(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload26 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload27 (.A(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload28 (.A(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload29 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload30 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload31 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkinv_2 clkload32 (.A(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload33 (.A(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload34 (.A(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload35 (.A(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload36 (.A(clknet_leaf_48_clk));
 sky130_fd_sc_hd__bufinv_16 clkload37 (.A(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload38 (.A(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkinv_2 clkload39 (.A(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload40 (.A(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkinv_1 clkload41 (.A(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkinv_2 clkload42 (.A(clknet_leaf_41_clk));
 sky130_fd_sc_hd__bufinv_16 clkload43 (.A(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload44 (.A(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload45 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload46 (.A(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload47 (.A(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload48 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload49 (.A(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload50 (.A(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload51 (.A(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload52 (.A(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload53 (.A(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload54 (.A(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkinv_2 clkload55 (.A(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkinv_2 clkload56 (.A(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload57 (.A(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clone1 (.A(net165),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(_0720_),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net164),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(_2547_),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net223),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net74),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net169),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(rst_n),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(wr_data[18]),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(wr_data[50]),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(wr_data[58]),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_0162_),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(wr_data[26]),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(wr_data[39]),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(wr_data[0]),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(_0048_),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(wr_data[48]),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(wr_data[32]),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(wr_data[10]),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_0049_),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(wr_data[14]),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(wr_data[13]),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_0084_),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(wr_data[42]),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(wr_data[46]),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(wr_data[4]),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_0202_),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(wr_data[45]),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(wr_data[36]),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(wr_data[44]),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(wr_data[63]),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(wr_data[21]),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0093_),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(wr_data[53]),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(wr_data[60]),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(wr_data[47]),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(wr_data[55]),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(wr_data[62]),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_0135_),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(wr_data[43]),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(wr_data[33]),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(wr_data[25]),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_0161_),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(wr_data[57]),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(wr_data[30]),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(wr_data[34]),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(wr_data[24]),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(wr_data[35]),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_0073_),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(wr_data[56]),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(wr_data[3]),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(wr_data[29]),
    .X(net215));
 sky130_fd_sc_hd__buf_16 load_slew1 (.A(_0003_),
    .X(net216));
 sky130_fd_sc_hd__buf_16 load_slew2 (.A(_0015_),
    .X(net217));
 sky130_fd_sc_hd__buf_16 load_slew3 (.A(_0007_),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(_0712_),
    .X(net219));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer10 (.A(net219),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(_0714_),
    .X(net221));
 sky130_fd_sc_hd__buf_6 rebuffer12 (.A(_0529_),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net75),
    .X(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_1279_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_1365_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_2494_));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_432 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_552 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_42 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_216 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_87 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_420 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_332 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_72 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_300 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_410 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_563 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_488 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_282 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_438 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_504 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_383 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_534 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_542 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_550 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_102 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_440 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_501 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_486 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_44 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_532 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_396 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_550 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_70 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_240 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_194 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_364 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_500 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_532 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_564 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_524 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_260 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_348 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_36 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_380 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_500 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_514 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_290 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_510 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_294 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_353 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_70 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_350 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_460 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_173 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_460 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_194 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_354 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_563 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_468 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_320 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_390 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_468 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_72 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_503 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_397 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_540 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_44 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_498 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_552 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_380 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_484 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_21 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_34 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_314 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_83 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_526 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_92 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_396 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_19 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_564 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_44 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_214 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_469 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_554 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_280 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_413 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_294 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_320 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_430 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_468 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_477 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_87 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_210 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_563 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_283 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_354 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_64 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_514 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_555 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_74 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_468 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_476 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_542 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_550 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_170 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_194 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_390 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_147 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_260 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_66 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_72 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_464 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_552 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_396 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_260 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_438 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_480 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_380 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_557 ();
endmodule
