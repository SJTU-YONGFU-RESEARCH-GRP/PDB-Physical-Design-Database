module axi_lite_master (arready,
    arvalid,
    awready,
    awvalid,
    bready,
    bvalid,
    clk,
    read_done,
    read_req,
    rready,
    rst_n,
    rvalid,
    wready,
    write_done,
    write_req,
    wvalid,
    araddr,
    awaddr,
    bresp,
    rdata,
    read_addr,
    read_data,
    rresp,
    wdata,
    write_addr,
    write_data,
    write_strb,
    wstrb);
 input arready;
 output arvalid;
 input awready;
 output awvalid;
 output bready;
 input bvalid;
 input clk;
 output read_done;
 input read_req;
 output rready;
 input rst_n;
 input rvalid;
 input wready;
 output write_done;
 input write_req;
 output wvalid;
 output [31:0] araddr;
 output [31:0] awaddr;
 input [1:0] bresp;
 input [31:0] rdata;
 input [31:0] read_addr;
 output [31:0] read_data;
 input [1:0] rresp;
 output [31:0] wdata;
 input [31:0] write_addr;
 input [31:0] write_data;
 input [3:0] write_strb;
 output [3:0] wstrb;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire net15;
 wire net14;
 wire net13;
 wire _149_;
 wire net12;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire net11;
 wire net10;
 wire net9;
 wire net8;
 wire net7;
 wire net6;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire net5;
 wire net4;
 wire net3;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire net2;
 wire net1;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire \state_r[0] ;
 wire \state_r[1] ;
 wire \state_r[2] ;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net283;
 wire net285;
 wire clknet_0_clk;
 wire net284;
 wire net286;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net287;

 gf180mcu_fd_sc_mcu9t5v0__inv_4 _203_ (.I(\state_r[1] ),
    .ZN(_142_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _204_ (.I(\state_r[0] ),
    .ZN(_143_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _205_ (.A1(_142_),
    .A2(_143_),
    .A3(net68),
    .ZN(_144_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _206_ (.A1(\state_r[2] ),
    .A2(_144_),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input15 (.I(rdata[1]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _208_ (.I0(net141),
    .I1(net36),
    .S(net283),
    .Z(_000_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _209_ (.I0(net142),
    .I1(net37),
    .S(net283),
    .Z(_001_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _210_ (.I0(net143),
    .I1(net38),
    .S(net283),
    .Z(_002_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _211_ (.I0(net144),
    .I1(net39),
    .S(net283),
    .Z(_003_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _212_ (.I0(net145),
    .I1(net40),
    .S(net283),
    .Z(_004_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _213_ (.I0(net146),
    .I1(net41),
    .S(net283),
    .Z(_005_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _214_ (.I0(net147),
    .I1(net42),
    .S(net283),
    .Z(_006_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _215_ (.I0(net148),
    .I1(net43),
    .S(net283),
    .Z(_007_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _216_ (.I0(net149),
    .I1(net44),
    .S(net283),
    .Z(_008_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _217_ (.I0(net150),
    .I1(net45),
    .S(net283),
    .Z(_009_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input14 (.I(rdata[19]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _219_ (.I0(net151),
    .I1(net46),
    .S(net283),
    .Z(_010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _220_ (.I0(net152),
    .I1(net47),
    .S(net283),
    .Z(_011_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _221_ (.I0(net153),
    .I1(net48),
    .S(_145_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _222_ (.I0(net154),
    .I1(net49),
    .S(net283),
    .Z(_013_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _223_ (.I0(net155),
    .I1(net50),
    .S(net283),
    .Z(_014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _224_ (.I0(net156),
    .I1(net51),
    .S(_145_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _225_ (.I0(net157),
    .I1(net52),
    .S(net283),
    .Z(_016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _226_ (.I0(net158),
    .I1(net53),
    .S(net283),
    .Z(_017_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _227_ (.I0(net159),
    .I1(net54),
    .S(net283),
    .Z(_018_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _228_ (.I0(net160),
    .I1(net55),
    .S(_145_),
    .Z(_019_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input13 (.I(rdata[18]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _230_ (.I0(net161),
    .I1(net56),
    .S(_145_),
    .Z(_020_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _231_ (.I0(net162),
    .I1(net57),
    .S(_145_),
    .Z(_021_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _232_ (.I0(net163),
    .I1(net58),
    .S(_145_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _233_ (.I0(net164),
    .I1(net59),
    .S(_145_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _234_ (.I0(net165),
    .I1(net60),
    .S(_145_),
    .Z(_024_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _235_ (.I0(net166),
    .I1(net61),
    .S(_145_),
    .Z(_025_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _236_ (.I0(net167),
    .I1(net62),
    .S(_145_),
    .Z(_026_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _237_ (.I0(net168),
    .I1(net63),
    .S(_145_),
    .Z(_027_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _238_ (.I0(net169),
    .I1(net64),
    .S(_145_),
    .Z(_028_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _239_ (.I0(net170),
    .I1(net65),
    .S(_145_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _240_ (.I0(net171),
    .I1(net66),
    .S(net283),
    .Z(_030_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _241_ (.I0(net172),
    .I1(net67),
    .S(net283),
    .Z(_031_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _242_ (.I(net173),
    .ZN(_149_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input12 (.I(rdata[17]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _244_ (.A1(_149_),
    .A2(_144_),
    .B(\state_r[2] ),
    .ZN(_151_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _245_ (.A1(_143_),
    .A2(net1),
    .B(_149_),
    .C(\state_r[1] ),
    .ZN(_152_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _246_ (.A1(_151_),
    .A2(_152_),
    .Z(_032_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _247_ (.A1(\state_r[2] ),
    .A2(\state_r[0] ),
    .ZN(_153_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _248_ (.A1(_142_),
    .A2(net136),
    .A3(_153_),
    .Z(_154_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input11 (.I(rdata[16]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(rdata[15]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(rdata[14]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _252_ (.I0(net174),
    .I1(net72),
    .S(net284),
    .Z(_033_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _253_ (.I0(net175),
    .I1(net73),
    .S(net284),
    .Z(_034_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _254_ (.I0(net176),
    .I1(net74),
    .S(net284),
    .Z(_035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _255_ (.I0(net177),
    .I1(net75),
    .S(net284),
    .Z(_036_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _256_ (.I0(net178),
    .I1(net76),
    .S(net284),
    .Z(_037_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _257_ (.I0(net179),
    .I1(net77),
    .S(net284),
    .Z(_038_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _258_ (.I0(net180),
    .I1(net78),
    .S(net284),
    .Z(_039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _259_ (.I0(net181),
    .I1(net79),
    .S(net284),
    .Z(_040_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _260_ (.I0(net182),
    .I1(net80),
    .S(net284),
    .Z(_041_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(rdata[13]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _262_ (.I0(net183),
    .I1(net81),
    .S(net284),
    .Z(_042_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _263_ (.I0(net184),
    .I1(net82),
    .S(net284),
    .Z(_043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _264_ (.I0(net185),
    .I1(net83),
    .S(net284),
    .Z(_044_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _265_ (.I0(net186),
    .I1(net84),
    .S(net284),
    .Z(_045_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _266_ (.I0(net187),
    .I1(net85),
    .S(net284),
    .Z(_046_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _267_ (.I0(net188),
    .I1(net86),
    .S(net284),
    .Z(_047_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _268_ (.I0(net189),
    .I1(net87),
    .S(net284),
    .Z(_048_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _269_ (.I0(net190),
    .I1(net88),
    .S(net284),
    .Z(_049_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _270_ (.I0(net191),
    .I1(net89),
    .S(net284),
    .Z(_050_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _271_ (.I0(net192),
    .I1(net90),
    .S(net284),
    .Z(_051_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(rdata[12]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _273_ (.I0(net193),
    .I1(net91),
    .S(_154_),
    .Z(_052_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _274_ (.I0(net194),
    .I1(net92),
    .S(_154_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _275_ (.I0(net195),
    .I1(net93),
    .S(_154_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _276_ (.I0(net196),
    .I1(net94),
    .S(_154_),
    .Z(_055_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _277_ (.I0(net197),
    .I1(net95),
    .S(_154_),
    .Z(_056_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _278_ (.I0(net198),
    .I1(net96),
    .S(_154_),
    .Z(_057_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _279_ (.I0(net199),
    .I1(net97),
    .S(_154_),
    .Z(_058_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _280_ (.I0(net200),
    .I1(net98),
    .S(_154_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _281_ (.I0(net201),
    .I1(net99),
    .S(_154_),
    .Z(_060_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _282_ (.I0(net202),
    .I1(net100),
    .S(_154_),
    .Z(_061_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(rdata[11]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _284_ (.I0(net203),
    .I1(net101),
    .S(net284),
    .Z(_062_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _285_ (.I0(net204),
    .I1(net102),
    .S(net284),
    .Z(_063_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _286_ (.I0(net205),
    .I1(net103),
    .S(net284),
    .Z(_064_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _287_ (.I(\state_r[2] ),
    .ZN(_161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _288_ (.A1(_161_),
    .A2(net206),
    .ZN(_162_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _289_ (.A1(_142_),
    .A2(\state_r[0] ),
    .Z(_163_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _290_ (.A1(net2),
    .A2(_163_),
    .Z(_164_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _291_ (.A1(\state_r[2] ),
    .A2(net206),
    .B1(net136),
    .B2(_153_),
    .ZN(_165_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _292_ (.A1(_162_),
    .A2(_164_),
    .B1(_165_),
    .B2(\state_r[1] ),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _293_ (.I(net207),
    .ZN(_166_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _294_ (.A1(_166_),
    .A2(net3),
    .B(\state_r[0] ),
    .ZN(_167_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _295_ (.A1(_161_),
    .A2(_167_),
    .ZN(_168_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _296_ (.A1(net279),
    .A2(net71),
    .Z(_169_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _297_ (.A1(\state_r[1] ),
    .A2(_169_),
    .B(net207),
    .ZN(_170_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _298_ (.A1(\state_r[1] ),
    .A2(_168_),
    .B(_170_),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _299_ (.A1(net241),
    .A2(net70),
    .Z(_171_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _300_ (.A1(\state_r[2] ),
    .A2(_163_),
    .A3(_171_),
    .Z(_172_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(rdata[10]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _302_ (.I0(net208),
    .I1(net4),
    .S(_172_),
    .Z(_067_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _303_ (.I0(net209),
    .I1(net5),
    .S(_172_),
    .Z(_068_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _304_ (.I0(net210),
    .I1(net6),
    .S(_172_),
    .Z(_069_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _305_ (.I0(net211),
    .I1(net7),
    .S(_172_),
    .Z(_070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _306_ (.I0(net212),
    .I1(net8),
    .S(_172_),
    .Z(_071_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _307_ (.I0(net213),
    .I1(net9),
    .S(_172_),
    .Z(_072_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _308_ (.I0(net214),
    .I1(net10),
    .S(_172_),
    .Z(_073_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _309_ (.I0(net215),
    .I1(net11),
    .S(_172_),
    .Z(_074_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _310_ (.I0(net216),
    .I1(net12),
    .S(_172_),
    .Z(_075_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _311_ (.I0(net217),
    .I1(net13),
    .S(_172_),
    .Z(_076_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(rdata[0]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _313_ (.I0(net218),
    .I1(net14),
    .S(_172_),
    .Z(_077_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _314_ (.I0(net219),
    .I1(net15),
    .S(_172_),
    .Z(_078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _315_ (.I0(net220),
    .I1(net16),
    .S(_172_),
    .Z(_079_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _316_ (.I0(net221),
    .I1(net17),
    .S(_172_),
    .Z(_080_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _317_ (.I0(net222),
    .I1(net18),
    .S(_172_),
    .Z(_081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _318_ (.I0(net223),
    .I1(net19),
    .S(_172_),
    .Z(_082_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _319_ (.I0(net224),
    .I1(net20),
    .S(_172_),
    .Z(_083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _320_ (.I0(net225),
    .I1(net21),
    .S(_172_),
    .Z(_084_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _321_ (.I0(net226),
    .I1(net22),
    .S(_172_),
    .Z(_085_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _322_ (.I0(net227),
    .I1(net23),
    .S(_172_),
    .Z(_086_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(bvalid),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _324_ (.I0(net228),
    .I1(net24),
    .S(_172_),
    .Z(_087_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _325_ (.I0(net229),
    .I1(net25),
    .S(_172_),
    .Z(_088_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _326_ (.I0(net230),
    .I1(net26),
    .S(_172_),
    .Z(_089_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _327_ (.I0(net231),
    .I1(net27),
    .S(_172_),
    .Z(_090_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _328_ (.I0(net232),
    .I1(net28),
    .S(_172_),
    .Z(_091_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _329_ (.I0(net233),
    .I1(net29),
    .S(_172_),
    .Z(_092_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _330_ (.I0(net234),
    .I1(net30),
    .S(_172_),
    .Z(_093_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _331_ (.I0(net235),
    .I1(net31),
    .S(_172_),
    .Z(_094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _332_ (.I0(net236),
    .I1(net32),
    .S(_172_),
    .Z(_095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _333_ (.I0(net237),
    .I1(net33),
    .S(_172_),
    .Z(_096_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _334_ (.I0(net238),
    .I1(net34),
    .S(_172_),
    .Z(_097_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _335_ (.I0(net239),
    .I1(net35),
    .S(_172_),
    .Z(_098_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _336_ (.A1(_163_),
    .A2(_171_),
    .B(net240),
    .ZN(_176_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _337_ (.A1(\state_r[1] ),
    .A2(\state_r[0] ),
    .B(net240),
    .ZN(_177_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _338_ (.A1(_161_),
    .A2(_176_),
    .B(_177_),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _339_ (.I(net241),
    .ZN(_178_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _340_ (.A1(\state_r[2] ),
    .A2(_143_),
    .A3(net173),
    .A4(net1),
    .Z(_179_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _341_ (.A1(\state_r[0] ),
    .A2(net70),
    .B(_178_),
    .ZN(_180_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _342_ (.A1(_179_),
    .A2(_180_),
    .B(_142_),
    .ZN(_181_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _343_ (.A1(\state_r[2] ),
    .A2(_178_),
    .B(_181_),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _344_ (.I(net284),
    .ZN(_182_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _345_ (.A1(net206),
    .A2(net2),
    .Z(_183_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _346_ (.A1(\state_r[2] ),
    .A2(_143_),
    .A3(_183_),
    .ZN(_184_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _347_ (.A1(_161_),
    .A2(_143_),
    .A3(_171_),
    .ZN(_185_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _348_ (.A1(_179_),
    .A2(_184_),
    .A3(_185_),
    .B(_142_),
    .ZN(_186_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _349_ (.A1(\state_r[0] ),
    .A2(net207),
    .A3(net3),
    .ZN(_187_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _350_ (.A1(\state_r[0] ),
    .A2(_169_),
    .B(_187_),
    .ZN(_188_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _351_ (.A1(\state_r[2] ),
    .A2(_142_),
    .A3(_188_),
    .Z(_189_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _352_ (.A1(_182_),
    .A2(_186_),
    .A3(_189_),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _353_ (.A1(_163_),
    .A2(_183_),
    .B1(_187_),
    .B2(\state_r[1] ),
    .ZN(_190_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _354_ (.A1(\state_r[2] ),
    .A2(_190_),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _355_ (.A1(_143_),
    .A2(net68),
    .ZN(_191_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _356_ (.A1(\state_r[0] ),
    .A2(_171_),
    .Z(_192_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _357_ (.A1(net136),
    .A2(_191_),
    .B1(_192_),
    .B2(_161_),
    .ZN(_193_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _358_ (.A1(_142_),
    .A2(_193_),
    .Z(_103_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _359_ (.I0(net242),
    .I1(net104),
    .S(net284),
    .Z(_104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _360_ (.I0(net243),
    .I1(net105),
    .S(net284),
    .Z(_105_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _361_ (.I0(net244),
    .I1(net106),
    .S(net284),
    .Z(_106_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _362_ (.I0(net245),
    .I1(net107),
    .S(net284),
    .Z(_107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _363_ (.I0(net246),
    .I1(net108),
    .S(net284),
    .Z(_108_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _364_ (.I0(net247),
    .I1(net109),
    .S(net284),
    .Z(_109_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _365_ (.I0(net248),
    .I1(net110),
    .S(net284),
    .Z(_110_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(awready),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _367_ (.I0(net249),
    .I1(net111),
    .S(net284),
    .Z(_111_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _368_ (.I0(net250),
    .I1(net112),
    .S(net284),
    .Z(_112_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _369_ (.I0(net251),
    .I1(net113),
    .S(net284),
    .Z(_113_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _370_ (.I0(net252),
    .I1(net114),
    .S(net284),
    .Z(_114_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _371_ (.I0(net253),
    .I1(net115),
    .S(net284),
    .Z(_115_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _372_ (.I0(net254),
    .I1(net116),
    .S(net284),
    .Z(_116_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _373_ (.I0(net255),
    .I1(net117),
    .S(net284),
    .Z(_117_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _374_ (.I0(net256),
    .I1(net118),
    .S(net284),
    .Z(_118_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _375_ (.I0(net257),
    .I1(net119),
    .S(net284),
    .Z(_119_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _376_ (.I0(net258),
    .I1(net120),
    .S(net284),
    .Z(_120_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input1 (.I(arready),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _378_ (.I0(net259),
    .I1(net121),
    .S(_154_),
    .Z(_121_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _379_ (.I0(net260),
    .I1(net122),
    .S(_154_),
    .Z(_122_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _380_ (.I0(net261),
    .I1(net123),
    .S(_154_),
    .Z(_123_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _381_ (.I0(net262),
    .I1(net124),
    .S(_154_),
    .Z(_124_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _382_ (.I0(net263),
    .I1(net125),
    .S(_154_),
    .Z(_125_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _383_ (.I0(net264),
    .I1(net126),
    .S(_154_),
    .Z(_126_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _384_ (.I0(net265),
    .I1(net127),
    .S(_154_),
    .Z(_127_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _385_ (.I0(net266),
    .I1(net128),
    .S(_154_),
    .Z(_128_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _386_ (.I0(net267),
    .I1(net129),
    .S(_154_),
    .Z(_129_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _387_ (.I0(net268),
    .I1(net130),
    .S(_154_),
    .Z(_130_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _388_ (.I0(net269),
    .I1(net131),
    .S(net284),
    .Z(_131_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _389_ (.I0(net270),
    .I1(net132),
    .S(net284),
    .Z(_132_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _390_ (.I0(net271),
    .I1(net133),
    .S(net284),
    .Z(_133_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _391_ (.I0(net272),
    .I1(net134),
    .S(net284),
    .Z(_134_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _392_ (.I0(net273),
    .I1(net135),
    .S(net284),
    .Z(_135_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _393_ (.I(net274),
    .ZN(_196_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _394_ (.A1(\state_r[2] ),
    .A2(_187_),
    .B(_196_),
    .ZN(_197_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _395_ (.A1(\state_r[1] ),
    .A2(_197_),
    .ZN(_198_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _396_ (.A1(_196_),
    .A2(_153_),
    .B(_198_),
    .ZN(_136_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _397_ (.I0(net275),
    .I1(net137),
    .S(net284),
    .Z(_137_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _398_ (.I0(net276),
    .I1(net138),
    .S(net284),
    .Z(_138_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _399_ (.I0(net277),
    .I1(net139),
    .S(net284),
    .Z(_139_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _400_ (.I0(net278),
    .I1(net140),
    .S(net284),
    .Z(_140_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _401_ (.A1(_143_),
    .A2(net71),
    .ZN(_199_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _402_ (.A1(_161_),
    .A2(net279),
    .A3(_199_),
    .ZN(_200_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _403_ (.A1(_161_),
    .A2(\state_r[0] ),
    .A3(_183_),
    .Z(_201_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _404_ (.A1(net279),
    .A2(_201_),
    .B(_142_),
    .ZN(_202_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _405_ (.A1(_200_),
    .A2(_202_),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[0]$_DFFE_PN0P_  (.D(_000_),
    .RN(net285),
    .CLK(clknet_4_2_0_clk),
    .Q(net141));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[10]$_DFFE_PN0P_  (.D(_001_),
    .RN(net285),
    .CLK(clknet_4_8_0_clk),
    .Q(net142));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[11]$_DFFE_PN0P_  (.D(_002_),
    .RN(net285),
    .CLK(clknet_4_8_0_clk),
    .Q(net143));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[12]$_DFFE_PN0P_  (.D(_003_),
    .RN(net285),
    .CLK(clknet_4_8_0_clk),
    .Q(net144));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[13]$_DFFE_PN0P_  (.D(_004_),
    .RN(net285),
    .CLK(clknet_4_2_0_clk),
    .Q(net145));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[14]$_DFFE_PN0P_  (.D(_005_),
    .RN(net285),
    .CLK(clknet_4_8_0_clk),
    .Q(net146));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[15]$_DFFE_PN0P_  (.D(_006_),
    .RN(net285),
    .CLK(clknet_4_2_0_clk),
    .Q(net147));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[16]$_DFFE_PN0P_  (.D(_007_),
    .RN(net285),
    .CLK(clknet_4_8_0_clk),
    .Q(net148));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[17]$_DFFE_PN0P_  (.D(_008_),
    .RN(net285),
    .CLK(clknet_4_8_0_clk),
    .Q(net149));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[18]$_DFFE_PN0P_  (.D(_009_),
    .RN(net285),
    .CLK(clknet_4_8_0_clk),
    .Q(net150));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[19]$_DFFE_PN0P_  (.D(_010_),
    .RN(net286),
    .CLK(clknet_4_10_0_clk),
    .Q(net151));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[1]$_DFFE_PN0P_  (.D(_011_),
    .RN(net286),
    .CLK(clknet_4_10_0_clk),
    .Q(net152));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[20]$_DFFE_PN0P_  (.D(_012_),
    .RN(net286),
    .CLK(clknet_4_10_0_clk),
    .Q(net153));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[21]$_DFFE_PN0P_  (.D(_013_),
    .RN(net286),
    .CLK(clknet_4_10_0_clk),
    .Q(net154));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[22]$_DFFE_PN0P_  (.D(_014_),
    .RN(net286),
    .CLK(clknet_4_8_0_clk),
    .Q(net155));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[23]$_DFFE_PN0P_  (.D(_015_),
    .RN(net286),
    .CLK(clknet_4_10_0_clk),
    .Q(net156));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[24]$_DFFE_PN0P_  (.D(_016_),
    .RN(net286),
    .CLK(clknet_4_10_0_clk),
    .Q(net157));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[25]$_DFFE_PN0P_  (.D(_017_),
    .RN(net286),
    .CLK(clknet_4_10_0_clk),
    .Q(net158));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[26]$_DFFE_PN0P_  (.D(_018_),
    .RN(net286),
    .CLK(clknet_4_10_0_clk),
    .Q(net159));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[27]$_DFFE_PN0P_  (.D(_019_),
    .RN(net286),
    .CLK(clknet_4_10_0_clk),
    .Q(net160));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[28]$_DFFE_PN0P_  (.D(_020_),
    .RN(net286),
    .CLK(clknet_4_11_0_clk),
    .Q(net161));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[29]$_DFFE_PN0P_  (.D(_021_),
    .RN(net286),
    .CLK(clknet_4_9_0_clk),
    .Q(net162));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[2]$_DFFE_PN0P_  (.D(_022_),
    .RN(net286),
    .CLK(clknet_4_11_0_clk),
    .Q(net163));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[30]$_DFFE_PN0P_  (.D(_023_),
    .RN(net286),
    .CLK(clknet_4_11_0_clk),
    .Q(net164));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[31]$_DFFE_PN0P_  (.D(_024_),
    .RN(net286),
    .CLK(clknet_4_11_0_clk),
    .Q(net165));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[3]$_DFFE_PN0P_  (.D(_025_),
    .RN(net286),
    .CLK(clknet_4_11_0_clk),
    .Q(net166));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[4]$_DFFE_PN0P_  (.D(_026_),
    .RN(net286),
    .CLK(clknet_4_9_0_clk),
    .Q(net167));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[5]$_DFFE_PN0P_  (.D(_027_),
    .RN(net286),
    .CLK(clknet_4_11_0_clk),
    .Q(net168));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[6]$_DFFE_PN0P_  (.D(_028_),
    .RN(net286),
    .CLK(clknet_4_10_0_clk),
    .Q(net169));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[7]$_DFFE_PN0P_  (.D(_029_),
    .RN(net286),
    .CLK(clknet_4_11_0_clk),
    .Q(net170));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[8]$_DFFE_PN0P_  (.D(_030_),
    .RN(net285),
    .CLK(clknet_4_8_0_clk),
    .Q(net171));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \araddr[9]$_DFFE_PN0P_  (.D(_031_),
    .RN(net285),
    .CLK(clknet_4_8_0_clk),
    .Q(net172));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \arvalid$_DFFE_PN0P_  (.D(_032_),
    .RN(net286),
    .CLK(clknet_4_9_0_clk),
    .Q(net173));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[0]$_DFFE_PN0P_  (.D(_033_),
    .RN(net285),
    .CLK(clknet_4_2_0_clk),
    .Q(net174));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[10]$_DFFE_PN0P_  (.D(_034_),
    .RN(net285),
    .CLK(clknet_4_2_0_clk),
    .Q(net175));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[11]$_DFFE_PN0P_  (.D(_035_),
    .RN(net285),
    .CLK(clknet_4_2_0_clk),
    .Q(net176));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[12]$_DFFE_PN0P_  (.D(_036_),
    .RN(net285),
    .CLK(clknet_4_0_0_clk),
    .Q(net177));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[13]$_DFFE_PN0P_  (.D(_037_),
    .RN(net285),
    .CLK(clknet_4_2_0_clk),
    .Q(net178));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[14]$_DFFE_PN0P_  (.D(_038_),
    .RN(net285),
    .CLK(clknet_4_0_0_clk),
    .Q(net179));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[15]$_DFFE_PN0P_  (.D(_039_),
    .RN(net285),
    .CLK(clknet_4_2_0_clk),
    .Q(net180));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[16]$_DFFE_PN0P_  (.D(_040_),
    .RN(net285),
    .CLK(clknet_4_0_0_clk),
    .Q(net181));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[17]$_DFFE_PN0P_  (.D(_041_),
    .RN(net285),
    .CLK(clknet_4_2_0_clk),
    .Q(net182));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[18]$_DFFE_PN0P_  (.D(_042_),
    .RN(net285),
    .CLK(clknet_4_5_0_clk),
    .Q(net183));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[19]$_DFFE_PN0P_  (.D(_043_),
    .RN(net285),
    .CLK(clknet_4_5_0_clk),
    .Q(net184));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[1]$_DFFE_PN0P_  (.D(_044_),
    .RN(net285),
    .CLK(clknet_4_5_0_clk),
    .Q(net185));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[20]$_DFFE_PN0P_  (.D(_045_),
    .RN(net285),
    .CLK(clknet_4_5_0_clk),
    .Q(net186));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[21]$_DFFE_PN0P_  (.D(_046_),
    .RN(net69),
    .CLK(clknet_4_5_0_clk),
    .Q(net187));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[22]$_DFFE_PN0P_  (.D(_047_),
    .RN(net69),
    .CLK(clknet_4_5_0_clk),
    .Q(net188));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[23]$_DFFE_PN0P_  (.D(_048_),
    .RN(net285),
    .CLK(clknet_4_5_0_clk),
    .Q(net189));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[24]$_DFFE_PN0P_  (.D(_049_),
    .RN(net285),
    .CLK(clknet_4_5_0_clk),
    .Q(net190));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[25]$_DFFE_PN0P_  (.D(_050_),
    .RN(net285),
    .CLK(clknet_4_5_0_clk),
    .Q(net191));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[26]$_DFFE_PN0P_  (.D(_051_),
    .RN(net69),
    .CLK(clknet_4_5_0_clk),
    .Q(net192));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[27]$_DFFE_PN0P_  (.D(_052_),
    .RN(net286),
    .CLK(clknet_4_12_0_clk),
    .Q(net193));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[28]$_DFFE_PN0P_  (.D(_053_),
    .RN(net286),
    .CLK(clknet_4_14_0_clk),
    .Q(net194));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[29]$_DFFE_PN0P_  (.D(_054_),
    .RN(net286),
    .CLK(clknet_4_9_0_clk),
    .Q(net195));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[2]$_DFFE_PN0P_  (.D(_055_),
    .RN(net286),
    .CLK(clknet_4_9_0_clk),
    .Q(net196));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[30]$_DFFE_PN0P_  (.D(_056_),
    .RN(net286),
    .CLK(clknet_4_14_0_clk),
    .Q(net197));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[31]$_DFFE_PN0P_  (.D(_057_),
    .RN(net286),
    .CLK(clknet_4_14_0_clk),
    .Q(net198));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[3]$_DFFE_PN0P_  (.D(_058_),
    .RN(net286),
    .CLK(clknet_4_14_0_clk),
    .Q(net199));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[4]$_DFFE_PN0P_  (.D(_059_),
    .RN(net286),
    .CLK(clknet_4_11_0_clk),
    .Q(net200));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[5]$_DFFE_PN0P_  (.D(_060_),
    .RN(net286),
    .CLK(clknet_4_11_0_clk),
    .Q(net201));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[6]$_DFFE_PN0P_  (.D(_061_),
    .RN(net286),
    .CLK(clknet_4_14_0_clk),
    .Q(net202));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[7]$_DFFE_PN0P_  (.D(_062_),
    .RN(net286),
    .CLK(clknet_4_6_0_clk),
    .Q(net203));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[8]$_DFFE_PN0P_  (.D(_063_),
    .RN(net285),
    .CLK(clknet_4_4_0_clk),
    .Q(net204));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awaddr[9]$_DFFE_PN0P_  (.D(_064_),
    .RN(net285),
    .CLK(clknet_4_4_0_clk),
    .Q(net205));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \awvalid$_DFFE_PN0P_  (.D(_065_),
    .RN(net286),
    .CLK(clknet_4_12_0_clk),
    .Q(net206));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bready$_DFFE_PN0P_  (.D(_066_),
    .RN(net285),
    .CLK(clknet_4_3_0_clk),
    .Q(net207));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[0]$_DFFE_PN0P_  (.D(_067_),
    .RN(net69),
    .CLK(clknet_4_15_0_clk),
    .Q(net208));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[10]$_DFFE_PN0P_  (.D(_068_),
    .RN(net286),
    .CLK(clknet_4_12_0_clk),
    .Q(net209));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[11]$_DFFE_PN0P_  (.D(_069_),
    .RN(net69),
    .CLK(clknet_4_12_0_clk),
    .Q(net210));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[12]$_DFFE_PN0P_  (.D(_070_),
    .RN(net286),
    .CLK(clknet_4_14_0_clk),
    .Q(net211));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[13]$_DFFE_PN0P_  (.D(_071_),
    .RN(net69),
    .CLK(clknet_4_15_0_clk),
    .Q(net212));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[14]$_DFFE_PN0P_  (.D(_072_),
    .RN(net69),
    .CLK(clknet_4_14_0_clk),
    .Q(net213));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[15]$_DFFE_PN0P_  (.D(_073_),
    .RN(net286),
    .CLK(clknet_4_12_0_clk),
    .Q(net214));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[16]$_DFFE_PN0P_  (.D(_074_),
    .RN(net69),
    .CLK(clknet_4_15_0_clk),
    .Q(net215));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[17]$_DFFE_PN0P_  (.D(_075_),
    .RN(net286),
    .CLK(clknet_4_14_0_clk),
    .Q(net216));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[18]$_DFFE_PN0P_  (.D(_076_),
    .RN(net286),
    .CLK(clknet_4_12_0_clk),
    .Q(net217));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[19]$_DFFE_PN0P_  (.D(_077_),
    .RN(net69),
    .CLK(clknet_4_7_0_clk),
    .Q(net218));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[1]$_DFFE_PN0P_  (.D(_078_),
    .RN(net69),
    .CLK(clknet_4_7_0_clk),
    .Q(net219));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[20]$_DFFE_PN0P_  (.D(_079_),
    .RN(net69),
    .CLK(clknet_4_7_0_clk),
    .Q(net220));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[21]$_DFFE_PN0P_  (.D(_080_),
    .RN(net69),
    .CLK(clknet_4_7_0_clk),
    .Q(net221));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[22]$_DFFE_PN0P_  (.D(_081_),
    .RN(net286),
    .CLK(clknet_4_6_0_clk),
    .Q(net222));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[23]$_DFFE_PN0P_  (.D(_082_),
    .RN(net69),
    .CLK(clknet_4_7_0_clk),
    .Q(net223));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[24]$_DFFE_PN0P_  (.D(_083_),
    .RN(net69),
    .CLK(clknet_4_6_0_clk),
    .Q(net224));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[25]$_DFFE_PN0P_  (.D(_084_),
    .RN(net69),
    .CLK(clknet_4_7_0_clk),
    .Q(net225));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[26]$_DFFE_PN0P_  (.D(_085_),
    .RN(net69),
    .CLK(clknet_4_7_0_clk),
    .Q(net226));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[27]$_DFFE_PN0P_  (.D(_086_),
    .RN(net69),
    .CLK(clknet_4_7_0_clk),
    .Q(net227));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[28]$_DFFE_PN0P_  (.D(_087_),
    .RN(net286),
    .CLK(clknet_4_13_0_clk),
    .Q(net228));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[29]$_DFFE_PN0P_  (.D(_088_),
    .RN(net69),
    .CLK(clknet_4_13_0_clk),
    .Q(net229));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[2]$_DFFE_PN0P_  (.D(_089_),
    .RN(net69),
    .CLK(clknet_4_13_0_clk),
    .Q(net230));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[30]$_DFFE_PN0P_  (.D(_090_),
    .RN(net286),
    .CLK(clknet_4_12_0_clk),
    .Q(net231));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[31]$_DFFE_PN0P_  (.D(_091_),
    .RN(net69),
    .CLK(clknet_4_12_0_clk),
    .Q(net232));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[3]$_DFFE_PN0P_  (.D(_092_),
    .RN(net69),
    .CLK(clknet_4_13_0_clk),
    .Q(net233));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[4]$_DFFE_PN0P_  (.D(_093_),
    .RN(net69),
    .CLK(clknet_4_13_0_clk),
    .Q(net234));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[5]$_DFFE_PN0P_  (.D(_094_),
    .RN(net69),
    .CLK(clknet_4_13_0_clk),
    .Q(net235));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[6]$_DFFE_PN0P_  (.D(_095_),
    .RN(net69),
    .CLK(clknet_4_13_0_clk),
    .Q(net236));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[7]$_DFFE_PN0P_  (.D(_096_),
    .RN(net69),
    .CLK(clknet_4_13_0_clk),
    .Q(net237));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[8]$_DFFE_PN0P_  (.D(_097_),
    .RN(net286),
    .CLK(clknet_4_7_0_clk),
    .Q(net238));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[9]$_DFFE_PN0P_  (.D(_098_),
    .RN(net286),
    .CLK(clknet_4_13_0_clk),
    .Q(net239));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_done_r$_DFFE_PN0P_  (.D(_099_),
    .RN(net286),
    .CLK(clknet_4_6_0_clk),
    .Q(net240));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rready$_DFFE_PN0P_  (.D(_100_),
    .RN(net286),
    .CLK(clknet_4_9_0_clk),
    .Q(net241));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \state_r[0]$_DFFE_PN0P_  (.D(_101_),
    .RN(net285),
    .CLK(clknet_4_3_0_clk),
    .Q(\state_r[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \state_r[1]$_DFFE_PN0P_  (.D(_102_),
    .RN(net285),
    .CLK(clknet_4_3_0_clk),
    .Q(\state_r[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \state_r[2]$_DFFE_PN0P_  (.D(_103_),
    .RN(net286),
    .CLK(clknet_4_9_0_clk),
    .Q(\state_r[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[0]$_DFFE_PN0P_  (.D(_104_),
    .RN(net285),
    .CLK(clknet_4_4_0_clk),
    .Q(net242));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[10]$_DFFE_PN0P_  (.D(_105_),
    .RN(net286),
    .CLK(clknet_4_6_0_clk),
    .Q(net243));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[11]$_DFFE_PN0P_  (.D(_106_),
    .RN(net285),
    .CLK(clknet_4_4_0_clk),
    .Q(net244));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[12]$_DFFE_PN0P_  (.D(_107_),
    .RN(net285),
    .CLK(clknet_4_4_0_clk),
    .Q(net245));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[13]$_DFFE_PN0P_  (.D(_108_),
    .RN(net285),
    .CLK(clknet_4_6_0_clk),
    .Q(net246));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[14]$_DFFE_PN0P_  (.D(_109_),
    .RN(net285),
    .CLK(clknet_4_1_0_clk),
    .Q(net247));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[15]$_DFFE_PN0P_  (.D(_110_),
    .RN(net286),
    .CLK(clknet_4_7_0_clk),
    .Q(net248));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[16]$_DFFE_PN0P_  (.D(_111_),
    .RN(net285),
    .CLK(clknet_4_1_0_clk),
    .Q(net249));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[17]$_DFFE_PN0P_  (.D(_112_),
    .RN(net285),
    .CLK(clknet_4_1_0_clk),
    .Q(net250));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[18]$_DFFE_PN0P_  (.D(_113_),
    .RN(net285),
    .CLK(clknet_4_6_0_clk),
    .Q(net251));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[19]$_DFFE_PN0P_  (.D(_114_),
    .RN(net285),
    .CLK(clknet_4_1_0_clk),
    .Q(net252));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[1]$_DFFE_PN0P_  (.D(_115_),
    .RN(net285),
    .CLK(clknet_4_6_0_clk),
    .Q(net253));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[20]$_DFFE_PN0P_  (.D(_116_),
    .RN(net285),
    .CLK(clknet_4_1_0_clk),
    .Q(net254));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[21]$_DFFE_PN0P_  (.D(_117_),
    .RN(net285),
    .CLK(clknet_4_1_0_clk),
    .Q(net255));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[22]$_DFFE_PN0P_  (.D(_118_),
    .RN(net285),
    .CLK(clknet_4_4_0_clk),
    .Q(net256));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[23]$_DFFE_PN0P_  (.D(_119_),
    .RN(net285),
    .CLK(clknet_4_4_0_clk),
    .Q(net257));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[24]$_DFFE_PN0P_  (.D(_120_),
    .RN(net285),
    .CLK(clknet_4_1_0_clk),
    .Q(net258));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[25]$_DFFE_PN0P_  (.D(_121_),
    .RN(net69),
    .CLK(clknet_4_15_0_clk),
    .Q(net259));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[26]$_DFFE_PN0P_  (.D(_122_),
    .RN(net69),
    .CLK(clknet_4_15_0_clk),
    .Q(net260));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[27]$_DFFE_PN0P_  (.D(_123_),
    .RN(net286),
    .CLK(clknet_4_15_0_clk),
    .Q(net261));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[28]$_DFFE_PN0P_  (.D(_124_),
    .RN(net69),
    .CLK(clknet_4_13_0_clk),
    .Q(net262));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[29]$_DFFE_PN0P_  (.D(_125_),
    .RN(net69),
    .CLK(clknet_4_15_0_clk),
    .Q(net263));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[2]$_DFFE_PN0P_  (.D(_126_),
    .RN(net69),
    .CLK(clknet_4_15_0_clk),
    .Q(net264));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[30]$_DFFE_PN0P_  (.D(_127_),
    .RN(net69),
    .CLK(clknet_4_15_0_clk),
    .Q(net265));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[31]$_DFFE_PN0P_  (.D(_128_),
    .RN(net69),
    .CLK(clknet_4_15_0_clk),
    .Q(net266));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[3]$_DFFE_PN0P_  (.D(_129_),
    .RN(net69),
    .CLK(clknet_4_15_0_clk),
    .Q(net267));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[4]$_DFFE_PN0P_  (.D(_130_),
    .RN(net286),
    .CLK(clknet_4_15_0_clk),
    .Q(net268));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[5]$_DFFE_PN0P_  (.D(_131_),
    .RN(net285),
    .CLK(clknet_4_1_0_clk),
    .Q(net269));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[6]$_DFFE_PN0P_  (.D(_132_),
    .RN(net285),
    .CLK(clknet_4_2_0_clk),
    .Q(net270));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[7]$_DFFE_PN0P_  (.D(_133_),
    .RN(net285),
    .CLK(clknet_4_0_0_clk),
    .Q(net271));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[8]$_DFFE_PN0P_  (.D(_134_),
    .RN(net285),
    .CLK(clknet_4_0_0_clk),
    .Q(net272));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wdata[9]$_DFFE_PN0P_  (.D(_135_),
    .RN(net285),
    .CLK(clknet_4_0_0_clk),
    .Q(net273));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \write_done_r$_DFFE_PN0P_  (.D(_136_),
    .RN(net285),
    .CLK(clknet_4_3_0_clk),
    .Q(net274));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wstrb[0]$_DFFE_PN0P_  (.D(_137_),
    .RN(net285),
    .CLK(clknet_4_0_0_clk),
    .Q(net275));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wstrb[1]$_DFFE_PN0P_  (.D(_138_),
    .RN(net285),
    .CLK(clknet_4_0_0_clk),
    .Q(net276));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wstrb[2]$_DFFE_PN0P_  (.D(_139_),
    .RN(net285),
    .CLK(clknet_4_0_0_clk),
    .Q(net277));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wstrb[3]$_DFFE_PN0P_  (.D(_140_),
    .RN(net285),
    .CLK(clknet_4_0_0_clk),
    .Q(net278));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wvalid$_DFFE_PN0P_  (.D(_141_),
    .RN(net285),
    .CLK(clknet_4_3_0_clk),
    .Q(net279));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input16 (.I(rdata[20]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input17 (.I(rdata[21]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input18 (.I(rdata[22]),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input19 (.I(rdata[23]),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input20 (.I(rdata[24]),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input21 (.I(rdata[25]),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input22 (.I(rdata[26]),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input23 (.I(rdata[27]),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input24 (.I(rdata[28]),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input25 (.I(rdata[29]),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input26 (.I(rdata[2]),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input27 (.I(rdata[30]),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input28 (.I(rdata[31]),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input29 (.I(rdata[3]),
    .Z(net29));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input30 (.I(rdata[4]),
    .Z(net30));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input31 (.I(rdata[5]),
    .Z(net31));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input32 (.I(rdata[6]),
    .Z(net32));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input33 (.I(rdata[7]),
    .Z(net33));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input34 (.I(rdata[8]),
    .Z(net34));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input35 (.I(rdata[9]),
    .Z(net35));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input36 (.I(read_addr[0]),
    .Z(net36));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input37 (.I(read_addr[10]),
    .Z(net37));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input38 (.I(read_addr[11]),
    .Z(net38));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input39 (.I(read_addr[12]),
    .Z(net39));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input40 (.I(read_addr[13]),
    .Z(net40));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input41 (.I(read_addr[14]),
    .Z(net41));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input42 (.I(read_addr[15]),
    .Z(net42));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input43 (.I(read_addr[16]),
    .Z(net43));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input44 (.I(read_addr[17]),
    .Z(net44));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input45 (.I(read_addr[18]),
    .Z(net45));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input46 (.I(read_addr[19]),
    .Z(net46));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input47 (.I(read_addr[1]),
    .Z(net47));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input48 (.I(read_addr[20]),
    .Z(net48));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input49 (.I(read_addr[21]),
    .Z(net49));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input50 (.I(read_addr[22]),
    .Z(net50));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input51 (.I(read_addr[23]),
    .Z(net51));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input52 (.I(read_addr[24]),
    .Z(net52));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input53 (.I(read_addr[25]),
    .Z(net53));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input54 (.I(read_addr[26]),
    .Z(net54));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input55 (.I(read_addr[27]),
    .Z(net55));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input56 (.I(read_addr[28]),
    .Z(net56));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input57 (.I(read_addr[29]),
    .Z(net57));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input58 (.I(read_addr[2]),
    .Z(net58));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input59 (.I(read_addr[30]),
    .Z(net59));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input60 (.I(read_addr[31]),
    .Z(net60));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input61 (.I(read_addr[3]),
    .Z(net61));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input62 (.I(read_addr[4]),
    .Z(net62));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input63 (.I(read_addr[5]),
    .Z(net63));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input64 (.I(read_addr[6]),
    .Z(net64));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input65 (.I(read_addr[7]),
    .Z(net65));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input66 (.I(read_addr[8]),
    .Z(net66));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input67 (.I(read_addr[9]),
    .Z(net67));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input68 (.I(read_req),
    .Z(net68));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input69 (.I(net287),
    .Z(net69));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input70 (.I(rvalid),
    .Z(net70));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input71 (.I(wready),
    .Z(net71));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input72 (.I(write_addr[0]),
    .Z(net72));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input73 (.I(write_addr[10]),
    .Z(net73));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input74 (.I(write_addr[11]),
    .Z(net74));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input75 (.I(write_addr[12]),
    .Z(net75));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input76 (.I(write_addr[13]),
    .Z(net76));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input77 (.I(write_addr[14]),
    .Z(net77));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input78 (.I(write_addr[15]),
    .Z(net78));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input79 (.I(write_addr[16]),
    .Z(net79));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input80 (.I(write_addr[17]),
    .Z(net80));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input81 (.I(write_addr[18]),
    .Z(net81));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input82 (.I(write_addr[19]),
    .Z(net82));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input83 (.I(write_addr[1]),
    .Z(net83));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input84 (.I(write_addr[20]),
    .Z(net84));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input85 (.I(write_addr[21]),
    .Z(net85));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input86 (.I(write_addr[22]),
    .Z(net86));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input87 (.I(write_addr[23]),
    .Z(net87));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input88 (.I(write_addr[24]),
    .Z(net88));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input89 (.I(write_addr[25]),
    .Z(net89));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input90 (.I(write_addr[26]),
    .Z(net90));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input91 (.I(write_addr[27]),
    .Z(net91));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input92 (.I(write_addr[28]),
    .Z(net92));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input93 (.I(write_addr[29]),
    .Z(net93));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input94 (.I(write_addr[2]),
    .Z(net94));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input95 (.I(write_addr[30]),
    .Z(net95));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input96 (.I(write_addr[31]),
    .Z(net96));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input97 (.I(write_addr[3]),
    .Z(net97));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input98 (.I(write_addr[4]),
    .Z(net98));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input99 (.I(write_addr[5]),
    .Z(net99));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input100 (.I(write_addr[6]),
    .Z(net100));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input101 (.I(write_addr[7]),
    .Z(net101));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input102 (.I(write_addr[8]),
    .Z(net102));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input103 (.I(write_addr[9]),
    .Z(net103));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input104 (.I(write_data[0]),
    .Z(net104));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input105 (.I(write_data[10]),
    .Z(net105));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input106 (.I(write_data[11]),
    .Z(net106));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input107 (.I(write_data[12]),
    .Z(net107));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input108 (.I(write_data[13]),
    .Z(net108));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input109 (.I(write_data[14]),
    .Z(net109));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input110 (.I(write_data[15]),
    .Z(net110));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input111 (.I(write_data[16]),
    .Z(net111));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input112 (.I(write_data[17]),
    .Z(net112));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input113 (.I(write_data[18]),
    .Z(net113));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input114 (.I(write_data[19]),
    .Z(net114));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input115 (.I(write_data[1]),
    .Z(net115));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input116 (.I(write_data[20]),
    .Z(net116));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input117 (.I(write_data[21]),
    .Z(net117));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input118 (.I(write_data[22]),
    .Z(net118));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input119 (.I(write_data[23]),
    .Z(net119));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input120 (.I(write_data[24]),
    .Z(net120));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input121 (.I(write_data[25]),
    .Z(net121));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input122 (.I(write_data[26]),
    .Z(net122));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input123 (.I(write_data[27]),
    .Z(net123));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input124 (.I(write_data[28]),
    .Z(net124));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input125 (.I(write_data[29]),
    .Z(net125));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input126 (.I(write_data[2]),
    .Z(net126));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input127 (.I(write_data[30]),
    .Z(net127));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input128 (.I(write_data[31]),
    .Z(net128));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input129 (.I(write_data[3]),
    .Z(net129));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input130 (.I(write_data[4]),
    .Z(net130));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input131 (.I(write_data[5]),
    .Z(net131));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input132 (.I(write_data[6]),
    .Z(net132));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input133 (.I(write_data[7]),
    .Z(net133));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input134 (.I(write_data[8]),
    .Z(net134));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input135 (.I(write_data[9]),
    .Z(net135));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input136 (.I(write_req),
    .Z(net136));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input137 (.I(write_strb[0]),
    .Z(net137));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input138 (.I(write_strb[1]),
    .Z(net138));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input139 (.I(write_strb[2]),
    .Z(net139));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input140 (.I(write_strb[3]),
    .Z(net140));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output141 (.I(net141),
    .Z(araddr[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output142 (.I(net142),
    .Z(araddr[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output143 (.I(net143),
    .Z(araddr[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output144 (.I(net144),
    .Z(araddr[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output145 (.I(net145),
    .Z(araddr[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output146 (.I(net146),
    .Z(araddr[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output147 (.I(net147),
    .Z(araddr[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output148 (.I(net148),
    .Z(araddr[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output149 (.I(net149),
    .Z(araddr[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output150 (.I(net150),
    .Z(araddr[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output151 (.I(net151),
    .Z(araddr[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output152 (.I(net152),
    .Z(araddr[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output153 (.I(net153),
    .Z(araddr[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output154 (.I(net154),
    .Z(araddr[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output155 (.I(net155),
    .Z(araddr[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output156 (.I(net156),
    .Z(araddr[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output157 (.I(net157),
    .Z(araddr[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output158 (.I(net158),
    .Z(araddr[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output159 (.I(net159),
    .Z(araddr[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output160 (.I(net160),
    .Z(araddr[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output161 (.I(net161),
    .Z(araddr[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output162 (.I(net162),
    .Z(araddr[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output163 (.I(net163),
    .Z(araddr[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output164 (.I(net164),
    .Z(araddr[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output165 (.I(net165),
    .Z(araddr[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output166 (.I(net166),
    .Z(araddr[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output167 (.I(net167),
    .Z(araddr[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output168 (.I(net168),
    .Z(araddr[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output169 (.I(net169),
    .Z(araddr[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output170 (.I(net170),
    .Z(araddr[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output171 (.I(net171),
    .Z(araddr[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output172 (.I(net172),
    .Z(araddr[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output173 (.I(net173),
    .Z(arvalid));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output174 (.I(net174),
    .Z(awaddr[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output175 (.I(net175),
    .Z(awaddr[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output176 (.I(net176),
    .Z(awaddr[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output177 (.I(net177),
    .Z(awaddr[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output178 (.I(net178),
    .Z(awaddr[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output179 (.I(net179),
    .Z(awaddr[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output180 (.I(net180),
    .Z(awaddr[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output181 (.I(net181),
    .Z(awaddr[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output182 (.I(net182),
    .Z(awaddr[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output183 (.I(net183),
    .Z(awaddr[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output184 (.I(net184),
    .Z(awaddr[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output185 (.I(net185),
    .Z(awaddr[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output186 (.I(net186),
    .Z(awaddr[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output187 (.I(net187),
    .Z(awaddr[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output188 (.I(net188),
    .Z(awaddr[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output189 (.I(net189),
    .Z(awaddr[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output190 (.I(net190),
    .Z(awaddr[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output191 (.I(net191),
    .Z(awaddr[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output192 (.I(net192),
    .Z(awaddr[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output193 (.I(net193),
    .Z(awaddr[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output194 (.I(net194),
    .Z(awaddr[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output195 (.I(net195),
    .Z(awaddr[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output196 (.I(net196),
    .Z(awaddr[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output197 (.I(net197),
    .Z(awaddr[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output198 (.I(net198),
    .Z(awaddr[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output199 (.I(net199),
    .Z(awaddr[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output200 (.I(net200),
    .Z(awaddr[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output201 (.I(net201),
    .Z(awaddr[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output202 (.I(net202),
    .Z(awaddr[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output203 (.I(net203),
    .Z(awaddr[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output204 (.I(net204),
    .Z(awaddr[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output205 (.I(net205),
    .Z(awaddr[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output206 (.I(net206),
    .Z(awvalid));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output207 (.I(net207),
    .Z(bready));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output208 (.I(net208),
    .Z(read_data[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output209 (.I(net209),
    .Z(read_data[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output210 (.I(net210),
    .Z(read_data[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output211 (.I(net211),
    .Z(read_data[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output212 (.I(net212),
    .Z(read_data[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output213 (.I(net213),
    .Z(read_data[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output214 (.I(net214),
    .Z(read_data[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output215 (.I(net215),
    .Z(read_data[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output216 (.I(net216),
    .Z(read_data[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output217 (.I(net217),
    .Z(read_data[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output218 (.I(net218),
    .Z(read_data[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output219 (.I(net219),
    .Z(read_data[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output220 (.I(net220),
    .Z(read_data[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output221 (.I(net221),
    .Z(read_data[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output222 (.I(net222),
    .Z(read_data[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output223 (.I(net223),
    .Z(read_data[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output224 (.I(net224),
    .Z(read_data[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output225 (.I(net225),
    .Z(read_data[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output226 (.I(net226),
    .Z(read_data[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output227 (.I(net227),
    .Z(read_data[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output228 (.I(net228),
    .Z(read_data[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output229 (.I(net229),
    .Z(read_data[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output230 (.I(net230),
    .Z(read_data[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output231 (.I(net231),
    .Z(read_data[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output232 (.I(net232),
    .Z(read_data[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output233 (.I(net233),
    .Z(read_data[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output234 (.I(net234),
    .Z(read_data[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output235 (.I(net235),
    .Z(read_data[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output236 (.I(net236),
    .Z(read_data[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output237 (.I(net237),
    .Z(read_data[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output238 (.I(net238),
    .Z(read_data[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output239 (.I(net239),
    .Z(read_data[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output240 (.I(net240),
    .Z(read_done));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output241 (.I(net241),
    .Z(rready));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output242 (.I(net242),
    .Z(wdata[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output243 (.I(net243),
    .Z(wdata[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output244 (.I(net244),
    .Z(wdata[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output245 (.I(net245),
    .Z(wdata[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output246 (.I(net246),
    .Z(wdata[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output247 (.I(net247),
    .Z(wdata[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output248 (.I(net248),
    .Z(wdata[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output249 (.I(net249),
    .Z(wdata[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output250 (.I(net250),
    .Z(wdata[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output251 (.I(net251),
    .Z(wdata[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output252 (.I(net252),
    .Z(wdata[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output253 (.I(net253),
    .Z(wdata[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output254 (.I(net254),
    .Z(wdata[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output255 (.I(net255),
    .Z(wdata[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output256 (.I(net256),
    .Z(wdata[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output257 (.I(net257),
    .Z(wdata[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output258 (.I(net258),
    .Z(wdata[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output259 (.I(net259),
    .Z(wdata[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output260 (.I(net260),
    .Z(wdata[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output261 (.I(net261),
    .Z(wdata[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output262 (.I(net262),
    .Z(wdata[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output263 (.I(net263),
    .Z(wdata[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output264 (.I(net264),
    .Z(wdata[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output265 (.I(net265),
    .Z(wdata[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output266 (.I(net266),
    .Z(wdata[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output267 (.I(net267),
    .Z(wdata[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output268 (.I(net268),
    .Z(wdata[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output269 (.I(net269),
    .Z(wdata[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output270 (.I(net270),
    .Z(wdata[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output271 (.I(net271),
    .Z(wdata[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output272 (.I(net272),
    .Z(wdata[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output273 (.I(net273),
    .Z(wdata[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output274 (.I(net274),
    .Z(write_done));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output275 (.I(net275),
    .Z(wstrb[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output276 (.I(net276),
    .Z(wstrb[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output277 (.I(net277),
    .Z(wstrb[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output278 (.I(net278),
    .Z(wstrb[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output279 (.I(net279),
    .Z(wvalid));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place283 (.I(_145_),
    .Z(net283));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place285 (.I(net69),
    .Z(net285));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place284 (.I(_154_),
    .Z(net284));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place286 (.I(net285),
    .Z(net286));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_0_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_1_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_2_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_3_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_4_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_5_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_6_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_7_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_8_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_9_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_10_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_11_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_12_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_13_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_14_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_15_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload0 (.I(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload1 (.I(clknet_4_1_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload2 (.I(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload3 (.I(clknet_4_3_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload4 (.I(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload5 (.I(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload6 (.I(clknet_4_6_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload7 (.I(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload8 (.I(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload9 (.I(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload10 (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload11 (.I(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload12 (.I(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload13 (.I(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload14 (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold287 (.I(rst_n),
    .Z(net287));
endmodule
