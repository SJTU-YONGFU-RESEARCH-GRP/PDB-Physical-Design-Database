module multi_phase_pwm_controller (clk,
    enable,
    rst_n,
    deadtime,
    duty,
    pwm_n_out,
    pwm_p_out);
 input clk;
 input enable;
 input rst_n;
 input [5:0] deadtime;
 input [7:0] duty;
 output [2:0] pwm_n_out;
 output [2:0] pwm_p_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 INV_X1 _0563_ (.A(_0361_),
    .ZN(_0321_));
 CLKBUF_X3 _0564_ (.A(_0330_),
    .Z(_0014_));
 XNOR2_X2 _0565_ (.A(_0014_),
    .B(_0326_),
    .ZN(_0388_));
 BUF_X1 _0566_ (.A(\counter[7] ),
    .Z(_0015_));
 INV_X1 _0567_ (.A(_0337_),
    .ZN(_0016_));
 INV_X1 _0568_ (.A(_0345_),
    .ZN(_0017_));
 BUF_X2 _0569_ (.A(\counter[6] ),
    .Z(_0018_));
 INV_X2 _0570_ (.A(\counter[5] ),
    .ZN(_0019_));
 NOR2_X1 _0571_ (.A1(_0018_),
    .A2(_0019_),
    .ZN(_0020_));
 NAND2_X1 _0572_ (.A1(\counter[0] ),
    .A2(_0485_),
    .ZN(_0021_));
 NAND2_X2 _0573_ (.A1(_0353_),
    .A2(_0021_),
    .ZN(_0022_));
 BUF_X2 _0574_ (.A(\counter[4] ),
    .Z(_0023_));
 BUF_X4 _0575_ (.A(\counter[3] ),
    .Z(_0024_));
 INV_X4 _0576_ (.A(_0024_),
    .ZN(_0025_));
 NOR4_X2 _0577_ (.A1(_0018_),
    .A2(_0019_),
    .A3(_0023_),
    .A4(_0025_),
    .ZN(_0026_));
 AOI221_X2 _0578_ (.A(_0016_),
    .B1(_0017_),
    .B2(_0020_),
    .C1(_0022_),
    .C2(_0026_),
    .ZN(_0027_));
 XNOR2_X1 _0579_ (.A(_0015_),
    .B(_0027_),
    .ZN(_0028_));
 INV_X1 _0580_ (.A(_0028_),
    .ZN(_0415_));
 INV_X2 _0581_ (.A(_0023_),
    .ZN(_0029_));
 CLKBUF_X2 _0582_ (.A(\counter[2] ),
    .Z(_0030_));
 OAI21_X2 _0583_ (.A(_0024_),
    .B1(_0030_),
    .B2(_0433_),
    .ZN(_0031_));
 AOI21_X2 _0584_ (.A(_0019_),
    .B1(_0029_),
    .B2(_0031_),
    .ZN(_0032_));
 XNOR2_X2 _0585_ (.A(_0016_),
    .B(_0032_),
    .ZN(_0033_));
 INV_X2 _0586_ (.A(_0033_),
    .ZN(_0418_));
 NAND2_X1 _0587_ (.A1(_0029_),
    .A2(_0024_),
    .ZN(_0034_));
 AOI21_X1 _0588_ (.A(_0030_),
    .B1(_0485_),
    .B2(\counter[0] ),
    .ZN(_0035_));
 OAI21_X1 _0589_ (.A(_0345_),
    .B1(_0034_),
    .B2(_0035_),
    .ZN(_0036_));
 XNOR2_X2 _0590_ (.A(_0019_),
    .B(_0036_),
    .ZN(_0450_));
 INV_X2 _0591_ (.A(_0450_),
    .ZN(_0421_));
 XNOR2_X2 _0592_ (.A(_0345_),
    .B(_0031_),
    .ZN(_0453_));
 INV_X2 _0593_ (.A(_0453_),
    .ZN(_0424_));
 XNOR2_X2 _0594_ (.A(_0025_),
    .B(_0022_),
    .ZN(_0444_));
 INV_X2 _0595_ (.A(_0444_),
    .ZN(_0427_));
 XOR2_X2 _0596_ (.A(_0353_),
    .B(_0433_),
    .Z(_0447_));
 INV_X2 _0597_ (.A(_0447_),
    .ZN(_0430_));
 INV_X1 _0598_ (.A(_0018_),
    .ZN(_0037_));
 OAI21_X2 _0599_ (.A(_0023_),
    .B1(_0024_),
    .B2(_0487_),
    .ZN(_0038_));
 AOI21_X2 _0600_ (.A(_0037_),
    .B1(_0019_),
    .B2(_0038_),
    .ZN(_0039_));
 XNOR2_X2 _0601_ (.A(_0333_),
    .B(_0039_),
    .ZN(_0470_));
 NAND2_X1 _0602_ (.A1(_0019_),
    .A2(_0023_),
    .ZN(_0040_));
 AOI21_X1 _0603_ (.A(_0024_),
    .B1(_0030_),
    .B2(\counter[1] ),
    .ZN(_0041_));
 OAI21_X1 _0604_ (.A(_0341_),
    .B1(_0040_),
    .B2(_0041_),
    .ZN(_0042_));
 XNOR2_X2 _0605_ (.A(_0018_),
    .B(_0042_),
    .ZN(_0473_));
 XNOR2_X2 _0606_ (.A(_0341_),
    .B(_0038_),
    .ZN(_0499_));
 INV_X2 _0607_ (.A(_0499_),
    .ZN(_0476_));
 NAND2_X1 _0608_ (.A1(_0030_),
    .A2(\counter[1] ),
    .ZN(_0043_));
 OAI21_X1 _0609_ (.A(_0349_),
    .B1(_0043_),
    .B2(_0024_),
    .ZN(_0044_));
 XNOR2_X2 _0610_ (.A(_0029_),
    .B(_0044_),
    .ZN(_0502_));
 INV_X2 _0611_ (.A(_0502_),
    .ZN(_0479_));
 XOR2_X2 _0612_ (.A(_0349_),
    .B(_0487_),
    .Z(_0493_));
 INV_X2 _0613_ (.A(_0493_),
    .ZN(_0482_));
 INV_X1 _0614_ (.A(net8),
    .ZN(_0324_));
 INV_X1 _0615_ (.A(_0363_),
    .ZN(_0325_));
 INV_X1 _0616_ (.A(_0327_),
    .ZN(_0375_));
 INV_X1 _0617_ (.A(_0486_),
    .ZN(_0496_));
 INV_X2 _0618_ (.A(net6),
    .ZN(_0391_));
 INV_X2 _0619_ (.A(net5),
    .ZN(_0396_));
 INV_X2 _0620_ (.A(net4),
    .ZN(_0380_));
 INV_X2 _0621_ (.A(net3),
    .ZN(_0328_));
 INV_X1 _0622_ (.A(_0362_),
    .ZN(_0366_));
 BUF_X2 _0623_ (.A(net13),
    .Z(_0045_));
 NOR2_X1 _0624_ (.A1(_0045_),
    .A2(_0392_),
    .ZN(_0046_));
 INV_X1 _0625_ (.A(_0381_),
    .ZN(_0047_));
 INV_X1 _0626_ (.A(_0371_),
    .ZN(_0048_));
 INV_X1 _0627_ (.A(_0357_),
    .ZN(_0049_));
 OAI21_X1 _0628_ (.A(_0048_),
    .B1(_0361_),
    .B2(_0049_),
    .ZN(_0050_));
 AOI21_X2 _0629_ (.A(_0329_),
    .B1(_0050_),
    .B2(_0014_),
    .ZN(_0051_));
 BUF_X2 _0630_ (.A(_0382_),
    .Z(_0052_));
 INV_X2 _0631_ (.A(_0052_),
    .ZN(_0053_));
 OAI21_X1 _0632_ (.A(_0047_),
    .B1(_0051_),
    .B2(_0053_),
    .ZN(_0054_));
 BUF_X2 _0633_ (.A(_0398_),
    .Z(_0055_));
 AOI21_X2 _0634_ (.A(_0397_),
    .B1(_0054_),
    .B2(_0055_),
    .ZN(_0056_));
 BUF_X2 _0635_ (.A(_0393_),
    .Z(_0057_));
 INV_X1 _0636_ (.A(_0057_),
    .ZN(_0058_));
 OAI21_X1 _0637_ (.A(_0046_),
    .B1(_0056_),
    .B2(_0058_),
    .ZN(_0059_));
 XNOR2_X2 _0638_ (.A(net14),
    .B(_0059_),
    .ZN(_0334_));
 INV_X1 _0639_ (.A(_0392_),
    .ZN(_0060_));
 AOI21_X1 _0640_ (.A(_0329_),
    .B1(_0322_),
    .B2(_0014_),
    .ZN(_0061_));
 OAI21_X2 _0641_ (.A(_0047_),
    .B1(_0061_),
    .B2(_0053_),
    .ZN(_0062_));
 AOI21_X1 _0642_ (.A(_0397_),
    .B1(_0062_),
    .B2(_0055_),
    .ZN(_0063_));
 OAI21_X1 _0643_ (.A(_0060_),
    .B1(_0063_),
    .B2(_0058_),
    .ZN(_0064_));
 XNOR2_X2 _0644_ (.A(_0045_),
    .B(_0064_),
    .ZN(_0338_));
 XNOR2_X2 _0645_ (.A(_0057_),
    .B(_0056_),
    .ZN(_0342_));
 INV_X2 _0646_ (.A(_0055_),
    .ZN(_0065_));
 XNOR2_X2 _0647_ (.A(_0065_),
    .B(_0062_),
    .ZN(_0346_));
 XNOR2_X2 _0648_ (.A(_0052_),
    .B(_0051_),
    .ZN(_0350_));
 XOR2_X2 _0649_ (.A(_0014_),
    .B(_0322_),
    .Z(_0354_));
 INV_X1 _0650_ (.A(_0331_),
    .ZN(_0066_));
 AOI21_X2 _0651_ (.A(_0372_),
    .B1(_0049_),
    .B2(_0363_),
    .ZN(_0067_));
 OAI21_X1 _0652_ (.A(_0066_),
    .B1(_0067_),
    .B2(_0014_),
    .ZN(_0068_));
 XNOR2_X2 _0653_ (.A(_0053_),
    .B(_0068_),
    .ZN(_0385_));
 INV_X1 _0654_ (.A(_0399_),
    .ZN(_0069_));
 INV_X1 _0655_ (.A(_0383_),
    .ZN(_0070_));
 OAI21_X2 _0656_ (.A(_0070_),
    .B1(_0052_),
    .B2(_0066_),
    .ZN(_0071_));
 NOR3_X2 _0657_ (.A1(_0014_),
    .A2(_0052_),
    .A3(_0055_),
    .ZN(_0072_));
 INV_X1 _0658_ (.A(_0372_),
    .ZN(_0073_));
 OAI21_X2 _0659_ (.A(_0073_),
    .B1(_0357_),
    .B2(_0325_),
    .ZN(_0074_));
 AOI22_X4 _0660_ (.A1(_0065_),
    .A2(_0071_),
    .B1(_0072_),
    .B2(_0074_),
    .ZN(_0075_));
 NAND2_X1 _0661_ (.A1(_0069_),
    .A2(_0075_),
    .ZN(_0076_));
 XNOR2_X2 _0662_ (.A(_0058_),
    .B(_0076_),
    .ZN(_0401_));
 NOR2_X1 _0663_ (.A1(_0014_),
    .A2(_0326_),
    .ZN(_0077_));
 OAI21_X1 _0664_ (.A(_0053_),
    .B1(_0077_),
    .B2(_0331_),
    .ZN(_0078_));
 NAND2_X1 _0665_ (.A1(_0070_),
    .A2(_0078_),
    .ZN(_0079_));
 XNOR2_X2 _0666_ (.A(_0065_),
    .B(_0079_),
    .ZN(_0404_));
 INV_X2 _0667_ (.A(net2),
    .ZN(_0320_));
 INV_X1 _0668_ (.A(net7),
    .ZN(_0360_));
 INV_X2 _0669_ (.A(_0434_),
    .ZN(_0435_));
 INV_X2 _0670_ (.A(net15),
    .ZN(_0080_));
 BUF_X4 _0671_ (.A(enable),
    .Z(_0081_));
 INV_X4 _0672_ (.A(_0081_),
    .ZN(_0082_));
 NAND2_X1 _0673_ (.A1(_0082_),
    .A2(\counter[0] ),
    .ZN(_0083_));
 AND3_X1 _0674_ (.A1(_0024_),
    .A2(_0030_),
    .A3(_0433_),
    .ZN(_0084_));
 AND3_X1 _0675_ (.A1(\counter[5] ),
    .A2(_0023_),
    .A3(_0084_),
    .ZN(_0085_));
 NAND2_X1 _0676_ (.A1(_0015_),
    .A2(_0018_),
    .ZN(_0086_));
 INV_X1 _0677_ (.A(_0086_),
    .ZN(_0087_));
 NAND2_X2 _0678_ (.A1(_0085_),
    .A2(_0087_),
    .ZN(_0088_));
 NAND3_X1 _0679_ (.A1(_0081_),
    .A2(_0365_),
    .A3(_0088_),
    .ZN(_0089_));
 AOI21_X1 _0680_ (.A(_0080_),
    .B1(_0083_),
    .B2(_0089_),
    .ZN(_0000_));
 NAND2_X1 _0681_ (.A1(_0082_),
    .A2(\counter[1] ),
    .ZN(_0090_));
 NAND3_X1 _0682_ (.A1(_0081_),
    .A2(_0434_),
    .A3(_0088_),
    .ZN(_0091_));
 AOI21_X1 _0683_ (.A(_0080_),
    .B1(_0090_),
    .B2(_0091_),
    .ZN(_0001_));
 NAND2_X1 _0684_ (.A1(_0082_),
    .A2(_0030_),
    .ZN(_0092_));
 NAND3_X1 _0685_ (.A1(_0081_),
    .A2(_0430_),
    .A3(_0088_),
    .ZN(_0093_));
 AOI21_X1 _0686_ (.A(_0080_),
    .B1(_0092_),
    .B2(_0093_),
    .ZN(_0002_));
 AND2_X1 _0687_ (.A1(\counter[0] ),
    .A2(_0487_),
    .ZN(_0094_));
 NAND3_X1 _0688_ (.A1(_0081_),
    .A2(_0025_),
    .A3(_0094_),
    .ZN(_0095_));
 OAI21_X1 _0689_ (.A(_0095_),
    .B1(_0094_),
    .B2(_0025_),
    .ZN(_0096_));
 AOI22_X1 _0690_ (.A1(_0082_),
    .A2(_0024_),
    .B1(_0088_),
    .B2(_0096_),
    .ZN(_0097_));
 NOR2_X1 _0691_ (.A1(_0080_),
    .A2(_0097_),
    .ZN(_0003_));
 NAND2_X1 _0692_ (.A1(_0081_),
    .A2(_0084_),
    .ZN(_0098_));
 XNOR2_X1 _0693_ (.A(_0029_),
    .B(_0098_),
    .ZN(_0099_));
 NOR2_X1 _0694_ (.A1(_0080_),
    .A2(_0099_),
    .ZN(_0004_));
 NAND2_X1 _0695_ (.A1(_0082_),
    .A2(\counter[5] ),
    .ZN(_0100_));
 NAND3_X1 _0696_ (.A1(_0023_),
    .A2(_0024_),
    .A3(_0094_),
    .ZN(_0101_));
 XOR2_X1 _0697_ (.A(_0341_),
    .B(_0101_),
    .Z(_0102_));
 NAND3_X1 _0698_ (.A1(_0081_),
    .A2(_0088_),
    .A3(_0102_),
    .ZN(_0103_));
 AOI21_X1 _0699_ (.A(_0080_),
    .B1(_0100_),
    .B2(_0103_),
    .ZN(_0005_));
 NAND2_X1 _0700_ (.A1(_0082_),
    .A2(_0018_),
    .ZN(_0104_));
 NAND3_X1 _0701_ (.A1(_0337_),
    .A2(_0085_),
    .A3(_0086_),
    .ZN(_0105_));
 OAI21_X1 _0702_ (.A(_0105_),
    .B1(_0085_),
    .B2(_0337_),
    .ZN(_0106_));
 NAND2_X1 _0703_ (.A1(_0081_),
    .A2(_0106_),
    .ZN(_0107_));
 AOI21_X1 _0704_ (.A(_0080_),
    .B1(_0104_),
    .B2(_0107_),
    .ZN(_0006_));
 NAND2_X1 _0705_ (.A1(_0082_),
    .A2(_0015_),
    .ZN(_0108_));
 NOR3_X1 _0706_ (.A1(_0037_),
    .A2(_0019_),
    .A3(_0101_),
    .ZN(_0109_));
 XNOR2_X1 _0707_ (.A(_0333_),
    .B(_0109_),
    .ZN(_0110_));
 NAND3_X1 _0708_ (.A1(_0081_),
    .A2(_0088_),
    .A3(_0110_),
    .ZN(_0111_));
 AOI21_X1 _0709_ (.A(_0080_),
    .B1(_0108_),
    .B2(_0111_),
    .ZN(_0007_));
 NAND2_X4 _0710_ (.A1(net15),
    .A2(_0081_),
    .ZN(_0112_));
 INV_X1 _0711_ (.A(_0015_),
    .ZN(_0113_));
 NAND3_X1 _0712_ (.A1(_0412_),
    .A2(_0408_),
    .A3(_0410_),
    .ZN(_0114_));
 NAND2_X1 _0713_ (.A1(_0514_),
    .A2(_0414_),
    .ZN(_0115_));
 INV_X1 _0714_ (.A(_0468_),
    .ZN(_0116_));
 NAND3_X1 _0715_ (.A1(_0116_),
    .A2(_0514_),
    .A3(_0414_),
    .ZN(_0117_));
 AOI21_X1 _0716_ (.A(_0413_),
    .B1(_0513_),
    .B2(_0414_),
    .ZN(_0118_));
 AOI21_X1 _0717_ (.A(_0114_),
    .B1(_0117_),
    .B2(_0118_),
    .ZN(_0119_));
 INV_X1 _0718_ (.A(_0408_),
    .ZN(_0120_));
 AOI21_X1 _0719_ (.A(_0409_),
    .B1(_0410_),
    .B2(_0411_),
    .ZN(_0121_));
 NOR2_X1 _0720_ (.A1(_0120_),
    .A2(_0121_),
    .ZN(_0122_));
 OAI33_X1 _0721_ (.A1(_0467_),
    .A2(_0114_),
    .A3(_0115_),
    .B1(_0119_),
    .B2(_0122_),
    .B3(_0407_),
    .ZN(_0123_));
 AOI21_X1 _0722_ (.A(_0113_),
    .B1(_0018_),
    .B2(_0123_),
    .ZN(_0124_));
 INV_X1 _0723_ (.A(_0394_),
    .ZN(_0125_));
 AND3_X1 _0724_ (.A1(net14),
    .A2(_0069_),
    .A3(_0125_),
    .ZN(_0126_));
 OR3_X1 _0725_ (.A1(_0014_),
    .A2(_0052_),
    .A3(_0055_),
    .ZN(_0127_));
 AOI21_X1 _0726_ (.A(_0383_),
    .B1(_0053_),
    .B2(_0331_),
    .ZN(_0128_));
 OAI221_X2 _0727_ (.A(_0126_),
    .B1(_0127_),
    .B2(_0067_),
    .C1(_0055_),
    .C2(_0128_),
    .ZN(_0129_));
 INV_X1 _0728_ (.A(_0045_),
    .ZN(_0130_));
 NOR2_X1 _0729_ (.A1(net14),
    .A2(_0130_),
    .ZN(_0131_));
 NAND2_X1 _0730_ (.A1(_0058_),
    .A2(_0131_),
    .ZN(_0132_));
 OR2_X1 _0731_ (.A1(_0075_),
    .A2(_0132_),
    .ZN(_0133_));
 OAI21_X1 _0732_ (.A(_0125_),
    .B1(_0069_),
    .B2(_0057_),
    .ZN(_0134_));
 OAI21_X1 _0733_ (.A(_0045_),
    .B1(_0058_),
    .B2(_0394_),
    .ZN(_0135_));
 AOI22_X2 _0734_ (.A1(_0131_),
    .A2(_0134_),
    .B1(_0135_),
    .B2(net14),
    .ZN(_0136_));
 AND3_X1 _0735_ (.A1(_0129_),
    .A2(_0133_),
    .A3(_0136_),
    .ZN(_0137_));
 OR2_X1 _0736_ (.A1(_0045_),
    .A2(_0057_),
    .ZN(_0138_));
 NAND3_X1 _0737_ (.A1(_0045_),
    .A2(_0069_),
    .A3(_0125_),
    .ZN(_0139_));
 OR2_X1 _0738_ (.A1(_0331_),
    .A2(_0383_),
    .ZN(_0140_));
 OAI221_X2 _0739_ (.A(_0065_),
    .B1(_0077_),
    .B2(_0140_),
    .C1(_0383_),
    .C2(_0053_),
    .ZN(_0141_));
 MUX2_X2 _0740_ (.A(_0138_),
    .B(_0139_),
    .S(_0141_),
    .Z(_0142_));
 NAND2_X1 _0741_ (.A1(_0045_),
    .A2(_0057_),
    .ZN(_0143_));
 OAI22_X2 _0742_ (.A1(_0069_),
    .A2(_0138_),
    .B1(_0143_),
    .B2(_0394_),
    .ZN(_0144_));
 AOI21_X4 _0743_ (.A(_0144_),
    .B1(_0394_),
    .B2(_0130_),
    .ZN(_0145_));
 NAND3_X1 _0744_ (.A1(_0387_),
    .A2(_0406_),
    .A3(_0403_),
    .ZN(_0146_));
 AOI21_X1 _0745_ (.A(_0389_),
    .B1(_0378_),
    .B2(_0390_),
    .ZN(_0147_));
 INV_X1 _0746_ (.A(_0377_),
    .ZN(_0148_));
 INV_X1 _0747_ (.A(_0367_),
    .ZN(_0149_));
 OAI211_X2 _0748_ (.A(_0148_),
    .B(_0390_),
    .C1(_0368_),
    .C2(_0149_),
    .ZN(_0150_));
 AOI21_X2 _0749_ (.A(_0146_),
    .B1(_0147_),
    .B2(_0150_),
    .ZN(_0151_));
 AOI21_X1 _0750_ (.A(_0402_),
    .B1(_0405_),
    .B2(_0403_),
    .ZN(_0152_));
 NAND3_X1 _0751_ (.A1(_0406_),
    .A2(_0403_),
    .A3(_0386_),
    .ZN(_0153_));
 NAND2_X1 _0752_ (.A1(_0152_),
    .A2(_0153_),
    .ZN(_0154_));
 OAI211_X2 _0753_ (.A(_0142_),
    .B(_0145_),
    .C1(_0151_),
    .C2(_0154_),
    .ZN(_0155_));
 AOI211_X2 _0754_ (.A(_0151_),
    .B(_0154_),
    .C1(_0142_),
    .C2(_0145_),
    .ZN(_0156_));
 OAI21_X1 _0755_ (.A(_0155_),
    .B1(_0156_),
    .B2(_0337_),
    .ZN(_0157_));
 OAI21_X1 _0756_ (.A(_0124_),
    .B1(_0137_),
    .B2(_0157_),
    .ZN(_0158_));
 NAND3_X1 _0757_ (.A1(_0336_),
    .A2(_0340_),
    .A3(_0344_),
    .ZN(_0159_));
 NOR2_X1 _0758_ (.A1(_0359_),
    .A2(_0439_),
    .ZN(_0160_));
 NAND4_X1 _0759_ (.A1(_0352_),
    .A2(_0348_),
    .A3(_0356_),
    .A4(_0160_),
    .ZN(_0161_));
 OR2_X1 _0760_ (.A1(_0159_),
    .A2(_0161_),
    .ZN(_0162_));
 AOI21_X1 _0761_ (.A(_0339_),
    .B1(_0343_),
    .B2(_0340_),
    .ZN(_0163_));
 INV_X1 _0762_ (.A(_0163_),
    .ZN(_0164_));
 AOI21_X1 _0763_ (.A(_0335_),
    .B1(_0164_),
    .B2(_0336_),
    .ZN(_0165_));
 OAI21_X1 _0764_ (.A(_0348_),
    .B1(_0351_),
    .B2(_0352_),
    .ZN(_0166_));
 NOR2_X1 _0765_ (.A1(_0351_),
    .A2(_0355_),
    .ZN(_0167_));
 NOR2_X1 _0766_ (.A1(_0440_),
    .A2(_0359_),
    .ZN(_0168_));
 OAI21_X1 _0767_ (.A(_0356_),
    .B1(_0491_),
    .B2(_0168_),
    .ZN(_0169_));
 AOI21_X1 _0768_ (.A(_0166_),
    .B1(_0167_),
    .B2(_0169_),
    .ZN(_0170_));
 NOR2_X1 _0769_ (.A1(_0347_),
    .A2(_0170_),
    .ZN(_0171_));
 OAI21_X1 _0770_ (.A(_0165_),
    .B1(_0171_),
    .B2(_0159_),
    .ZN(_0172_));
 OAI211_X2 _0771_ (.A(_0129_),
    .B(_0136_),
    .C1(_0132_),
    .C2(_0075_),
    .ZN(_0173_));
 AOI21_X1 _0772_ (.A(_0173_),
    .B1(_0123_),
    .B2(_0087_),
    .ZN(_0174_));
 AOI22_X1 _0773_ (.A1(_0162_),
    .A2(_0172_),
    .B1(_0157_),
    .B2(_0174_),
    .ZN(_0175_));
 AOI21_X1 _0774_ (.A(_0112_),
    .B1(_0158_),
    .B2(_0175_),
    .ZN(_0008_));
 NAND3_X1 _0775_ (.A1(_0461_),
    .A2(_0459_),
    .A3(_0463_),
    .ZN(_0176_));
 NAND3_X1 _0776_ (.A1(_0467_),
    .A2(_0457_),
    .A3(_0465_),
    .ZN(_0177_));
 INV_X1 _0777_ (.A(_0458_),
    .ZN(_0178_));
 INV_X1 _0778_ (.A(_0466_),
    .ZN(_0179_));
 AOI21_X1 _0779_ (.A(_0464_),
    .B1(_0465_),
    .B2(_0179_),
    .ZN(_0180_));
 OAI21_X1 _0780_ (.A(_0178_),
    .B1(_0176_),
    .B2(_0180_),
    .ZN(_0181_));
 INV_X1 _0781_ (.A(_0456_),
    .ZN(_0182_));
 AOI21_X1 _0782_ (.A(_0460_),
    .B1(_0462_),
    .B2(_0461_),
    .ZN(_0183_));
 INV_X1 _0783_ (.A(_0459_),
    .ZN(_0184_));
 OAI21_X1 _0784_ (.A(_0182_),
    .B1(_0183_),
    .B2(_0184_),
    .ZN(_0185_));
 OAI222_X2 _0785_ (.A1(_0457_),
    .A2(_0456_),
    .B1(_0176_),
    .B2(_0177_),
    .C1(_0181_),
    .C2(_0185_),
    .ZN(_0186_));
 INV_X1 _0786_ (.A(_0445_),
    .ZN(_0187_));
 OAI21_X1 _0787_ (.A(_0446_),
    .B1(_0449_),
    .B2(_0448_),
    .ZN(_0188_));
 OR2_X1 _0788_ (.A1(_0442_),
    .A2(_0448_),
    .ZN(_0189_));
 NAND2_X1 _0789_ (.A1(_0368_),
    .A2(_0369_),
    .ZN(_0190_));
 AOI21_X1 _0790_ (.A(_0189_),
    .B1(_0190_),
    .B2(_0443_),
    .ZN(_0191_));
 OAI21_X1 _0791_ (.A(_0187_),
    .B1(_0188_),
    .B2(_0191_),
    .ZN(_0192_));
 NAND2_X1 _0792_ (.A1(_0455_),
    .A2(_0452_),
    .ZN(_0193_));
 INV_X1 _0793_ (.A(_0193_),
    .ZN(_0194_));
 AOI221_X2 _0794_ (.A(_0451_),
    .B1(_0192_),
    .B2(_0194_),
    .C1(_0454_),
    .C2(_0452_),
    .ZN(_0195_));
 NAND2_X2 _0795_ (.A1(_0142_),
    .A2(_0145_),
    .ZN(_0196_));
 AOI21_X1 _0796_ (.A(_0186_),
    .B1(_0195_),
    .B2(_0196_),
    .ZN(_0197_));
 NOR2_X2 _0797_ (.A1(_0080_),
    .A2(_0082_),
    .ZN(_0198_));
 NAND2_X1 _0798_ (.A1(_0113_),
    .A2(_0198_),
    .ZN(_0199_));
 NAND2_X1 _0799_ (.A1(_0015_),
    .A2(_0198_),
    .ZN(_0200_));
 MUX2_X1 _0800_ (.A(_0199_),
    .B(_0200_),
    .S(_0027_),
    .Z(_0201_));
 NOR2_X1 _0801_ (.A1(_0418_),
    .A2(_0201_),
    .ZN(_0202_));
 NOR2_X1 _0802_ (.A1(_0033_),
    .A2(_0196_),
    .ZN(_0203_));
 NOR2_X1 _0803_ (.A1(_0201_),
    .A2(_0195_),
    .ZN(_0204_));
 AOI221_X2 _0804_ (.A(_0137_),
    .B1(_0197_),
    .B2(_0202_),
    .C1(_0203_),
    .C2(_0204_),
    .ZN(_0205_));
 AOI21_X1 _0805_ (.A(_0033_),
    .B1(_0142_),
    .B2(_0145_),
    .ZN(_0206_));
 AOI221_X1 _0806_ (.A(_0201_),
    .B1(_0186_),
    .B2(_0033_),
    .C1(_0206_),
    .C2(_0173_),
    .ZN(_0207_));
 NOR3_X1 _0807_ (.A1(_0028_),
    .A2(_0112_),
    .A3(_0206_),
    .ZN(_0208_));
 OAI21_X1 _0808_ (.A(_0195_),
    .B1(_0196_),
    .B2(_0418_),
    .ZN(_0209_));
 AOI21_X1 _0809_ (.A(_0207_),
    .B1(_0208_),
    .B2(_0209_),
    .ZN(_0210_));
 AND3_X1 _0810_ (.A1(_0417_),
    .A2(_0420_),
    .A3(_0423_),
    .ZN(_0211_));
 INV_X1 _0811_ (.A(_0425_),
    .ZN(_0212_));
 INV_X1 _0812_ (.A(_0426_),
    .ZN(_0213_));
 INV_X1 _0813_ (.A(_0431_),
    .ZN(_0214_));
 INV_X1 _0814_ (.A(_0438_),
    .ZN(_0215_));
 AOI21_X1 _0815_ (.A(_0436_),
    .B1(_0215_),
    .B2(_0437_),
    .ZN(_0216_));
 INV_X1 _0816_ (.A(_0432_),
    .ZN(_0217_));
 OAI21_X1 _0817_ (.A(_0214_),
    .B1(_0216_),
    .B2(_0217_),
    .ZN(_0218_));
 AOI21_X1 _0818_ (.A(_0428_),
    .B1(_0218_),
    .B2(_0429_),
    .ZN(_0219_));
 OAI21_X1 _0819_ (.A(_0212_),
    .B1(_0213_),
    .B2(_0219_),
    .ZN(_0220_));
 AOI21_X1 _0820_ (.A(_0419_),
    .B1(_0422_),
    .B2(_0420_),
    .ZN(_0221_));
 INV_X1 _0821_ (.A(_0221_),
    .ZN(_0222_));
 AOI221_X2 _0822_ (.A(_0416_),
    .B1(_0211_),
    .B2(_0220_),
    .C1(_0222_),
    .C2(_0417_),
    .ZN(_0223_));
 NAND2_X1 _0823_ (.A1(_0439_),
    .A2(_0437_),
    .ZN(_0224_));
 NAND4_X1 _0824_ (.A1(_0429_),
    .A2(_0426_),
    .A3(_0432_),
    .A4(_0211_),
    .ZN(_0225_));
 OAI21_X1 _0825_ (.A(_0198_),
    .B1(_0224_),
    .B2(_0225_),
    .ZN(_0226_));
 OAI22_X1 _0826_ (.A1(_0205_),
    .A2(_0210_),
    .B1(_0223_),
    .B2(_0226_),
    .ZN(_0009_));
 INV_X1 _0827_ (.A(_0495_),
    .ZN(_0227_));
 OAI21_X1 _0828_ (.A(_0501_),
    .B1(_0503_),
    .B2(_0504_),
    .ZN(_0228_));
 OR2_X1 _0829_ (.A1(_0227_),
    .A2(_0228_),
    .ZN(_0229_));
 AOI21_X1 _0830_ (.A(_0497_),
    .B1(_0376_),
    .B2(_0498_),
    .ZN(_0230_));
 AND2_X1 _0831_ (.A1(_0377_),
    .A2(_0498_),
    .ZN(_0231_));
 OAI21_X1 _0832_ (.A(_0231_),
    .B1(_0149_),
    .B2(_0368_),
    .ZN(_0232_));
 AOI21_X1 _0833_ (.A(_0229_),
    .B1(_0230_),
    .B2(_0232_),
    .ZN(_0233_));
 NOR2_X1 _0834_ (.A1(_0494_),
    .A2(_0503_),
    .ZN(_0234_));
 NOR2_X1 _0835_ (.A1(_0228_),
    .A2(_0234_),
    .ZN(_0235_));
 NOR3_X1 _0836_ (.A1(_0500_),
    .A2(_0233_),
    .A3(_0235_),
    .ZN(_0236_));
 NAND2_X1 _0837_ (.A1(_0196_),
    .A2(_0236_),
    .ZN(_0237_));
 OAI21_X1 _0838_ (.A(_0473_),
    .B1(_0196_),
    .B2(_0236_),
    .ZN(_0238_));
 AND2_X1 _0839_ (.A1(_0470_),
    .A2(_0198_),
    .ZN(_0239_));
 NAND4_X1 _0840_ (.A1(_0137_),
    .A2(_0237_),
    .A3(_0238_),
    .A4(_0239_),
    .ZN(_0240_));
 AOI21_X1 _0841_ (.A(_0137_),
    .B1(_0237_),
    .B2(_0238_),
    .ZN(_0241_));
 NOR2_X1 _0842_ (.A1(_0470_),
    .A2(_0112_),
    .ZN(_0242_));
 INV_X1 _0843_ (.A(_0505_),
    .ZN(_0243_));
 AND3_X1 _0844_ (.A1(_0510_),
    .A2(_0508_),
    .A3(_0512_),
    .ZN(_0244_));
 NOR2_X1 _0845_ (.A1(_0468_),
    .A2(_0514_),
    .ZN(_0245_));
 OAI21_X1 _0846_ (.A(_0244_),
    .B1(_0245_),
    .B2(_0515_),
    .ZN(_0246_));
 AOI21_X1 _0847_ (.A(_0509_),
    .B1(_0511_),
    .B2(_0510_),
    .ZN(_0247_));
 INV_X1 _0848_ (.A(_0508_),
    .ZN(_0248_));
 OAI21_X1 _0849_ (.A(_0246_),
    .B1(_0247_),
    .B2(_0248_),
    .ZN(_0249_));
 OAI21_X1 _0850_ (.A(_0506_),
    .B1(_0249_),
    .B2(_0507_),
    .ZN(_0250_));
 INV_X1 _0851_ (.A(_0506_),
    .ZN(_0251_));
 NOR3_X1 _0852_ (.A1(_0467_),
    .A2(_0514_),
    .A3(_0251_),
    .ZN(_0252_));
 AOI22_X1 _0853_ (.A1(_0243_),
    .A2(_0250_),
    .B1(_0252_),
    .B2(_0244_),
    .ZN(_0253_));
 OAI21_X1 _0854_ (.A(_0242_),
    .B1(_0253_),
    .B2(_0473_),
    .ZN(_0254_));
 INV_X1 _0855_ (.A(_0439_),
    .ZN(_0255_));
 NAND2_X1 _0856_ (.A1(_0255_),
    .A2(_0490_),
    .ZN(_0256_));
 INV_X1 _0857_ (.A(_0492_),
    .ZN(_0257_));
 AND3_X1 _0858_ (.A1(_0472_),
    .A2(_0475_),
    .A3(_0478_),
    .ZN(_0258_));
 NAND4_X1 _0859_ (.A1(_0484_),
    .A2(_0257_),
    .A3(_0481_),
    .A4(_0258_),
    .ZN(_0259_));
 OAI21_X1 _0860_ (.A(_0198_),
    .B1(_0256_),
    .B2(_0259_),
    .ZN(_0260_));
 INV_X1 _0861_ (.A(_0480_),
    .ZN(_0261_));
 INV_X1 _0862_ (.A(_0484_),
    .ZN(_0262_));
 INV_X1 _0863_ (.A(_0489_),
    .ZN(_0263_));
 NOR2_X1 _0864_ (.A1(_0440_),
    .A2(_0492_),
    .ZN(_0264_));
 OAI21_X1 _0865_ (.A(_0490_),
    .B1(_0358_),
    .B2(_0264_),
    .ZN(_0265_));
 AOI21_X1 _0866_ (.A(_0262_),
    .B1(_0263_),
    .B2(_0265_),
    .ZN(_0266_));
 OAI21_X1 _0867_ (.A(_0481_),
    .B1(_0483_),
    .B2(_0266_),
    .ZN(_0267_));
 NAND2_X1 _0868_ (.A1(_0261_),
    .A2(_0267_),
    .ZN(_0268_));
 AOI21_X1 _0869_ (.A(_0474_),
    .B1(_0477_),
    .B2(_0475_),
    .ZN(_0269_));
 INV_X1 _0870_ (.A(_0269_),
    .ZN(_0270_));
 AOI221_X2 _0871_ (.A(_0471_),
    .B1(_0268_),
    .B2(_0258_),
    .C1(_0270_),
    .C2(_0472_),
    .ZN(_0271_));
 OAI221_X1 _0872_ (.A(_0240_),
    .B1(_0241_),
    .B2(_0254_),
    .C1(_0260_),
    .C2(_0271_),
    .ZN(_0010_));
 AND4_X1 _0873_ (.A1(_0548_),
    .A2(_0550_),
    .A3(_0552_),
    .A4(_0554_),
    .ZN(_0272_));
 INV_X1 _0874_ (.A(_0544_),
    .ZN(_0273_));
 AND4_X1 _0875_ (.A1(_0560_),
    .A2(_0273_),
    .A3(_0556_),
    .A4(_0558_),
    .ZN(_0274_));
 INV_X1 _0876_ (.A(_0556_),
    .ZN(_0275_));
 INV_X1 _0877_ (.A(_0559_),
    .ZN(_0276_));
 INV_X1 _0878_ (.A(_0560_),
    .ZN(_0277_));
 OAI21_X1 _0879_ (.A(_0276_),
    .B1(_0277_),
    .B2(_0545_),
    .ZN(_0278_));
 AOI21_X1 _0880_ (.A(_0557_),
    .B1(_0278_),
    .B2(_0558_),
    .ZN(_0279_));
 NOR2_X1 _0881_ (.A1(_0275_),
    .A2(_0279_),
    .ZN(_0280_));
 OAI21_X1 _0882_ (.A(_0272_),
    .B1(_0280_),
    .B2(_0555_),
    .ZN(_0281_));
 INV_X1 _0883_ (.A(_0549_),
    .ZN(_0282_));
 AOI21_X1 _0884_ (.A(_0551_),
    .B1(_0552_),
    .B2(_0553_),
    .ZN(_0283_));
 INV_X1 _0885_ (.A(_0550_),
    .ZN(_0284_));
 OAI21_X1 _0886_ (.A(_0282_),
    .B1(_0283_),
    .B2(_0284_),
    .ZN(_0285_));
 AOI21_X1 _0887_ (.A(_0547_),
    .B1(_0285_),
    .B2(_0548_),
    .ZN(_0286_));
 AOI221_X1 _0888_ (.A(_0112_),
    .B1(_0272_),
    .B2(_0274_),
    .C1(_0281_),
    .C2(_0286_),
    .ZN(_0011_));
 AND4_X1 _0889_ (.A1(_0530_),
    .A2(_0534_),
    .A3(_0536_),
    .A4(_0532_),
    .ZN(_0287_));
 AND4_X1 _0890_ (.A1(_0544_),
    .A2(_0538_),
    .A3(_0540_),
    .A4(_0542_),
    .ZN(_0288_));
 INV_X1 _0891_ (.A(_0538_),
    .ZN(_0289_));
 INV_X1 _0892_ (.A(_0541_),
    .ZN(_0290_));
 INV_X1 _0893_ (.A(_0542_),
    .ZN(_0291_));
 OAI21_X1 _0894_ (.A(_0290_),
    .B1(_0543_),
    .B2(_0291_),
    .ZN(_0292_));
 AOI21_X1 _0895_ (.A(_0539_),
    .B1(_0292_),
    .B2(_0540_),
    .ZN(_0293_));
 NOR2_X1 _0896_ (.A1(_0289_),
    .A2(_0293_),
    .ZN(_0294_));
 OAI21_X1 _0897_ (.A(_0287_),
    .B1(_0294_),
    .B2(_0537_),
    .ZN(_0295_));
 INV_X1 _0898_ (.A(_0531_),
    .ZN(_0296_));
 AOI21_X1 _0899_ (.A(_0533_),
    .B1(_0535_),
    .B2(_0534_),
    .ZN(_0297_));
 INV_X1 _0900_ (.A(_0532_),
    .ZN(_0298_));
 OAI21_X1 _0901_ (.A(_0296_),
    .B1(_0297_),
    .B2(_0298_),
    .ZN(_0299_));
 AOI21_X1 _0902_ (.A(_0529_),
    .B1(_0299_),
    .B2(_0530_),
    .ZN(_0300_));
 AOI221_X2 _0903_ (.A(_0112_),
    .B1(_0287_),
    .B2(_0288_),
    .C1(_0295_),
    .C2(_0300_),
    .ZN(_0012_));
 AND4_X1 _0904_ (.A1(_0518_),
    .A2(_0520_),
    .A3(_0522_),
    .A4(_0524_),
    .ZN(_0301_));
 AND4_X1 _0905_ (.A1(_0526_),
    .A2(_0277_),
    .A3(_0273_),
    .A4(_0528_),
    .ZN(_0302_));
 INV_X1 _0906_ (.A(_0526_),
    .ZN(_0303_));
 INV_X1 _0907_ (.A(_0527_),
    .ZN(_0304_));
 NOR2_X1 _0908_ (.A1(_0545_),
    .A2(_0560_),
    .ZN(_0305_));
 OAI21_X1 _0909_ (.A(_0528_),
    .B1(_0561_),
    .B2(_0305_),
    .ZN(_0306_));
 AOI21_X1 _0910_ (.A(_0303_),
    .B1(_0304_),
    .B2(_0306_),
    .ZN(_0307_));
 OAI21_X1 _0911_ (.A(_0301_),
    .B1(_0307_),
    .B2(_0525_),
    .ZN(_0308_));
 INV_X1 _0912_ (.A(_0519_),
    .ZN(_0309_));
 AOI21_X1 _0913_ (.A(_0521_),
    .B1(_0522_),
    .B2(_0523_),
    .ZN(_0310_));
 INV_X1 _0914_ (.A(_0520_),
    .ZN(_0311_));
 OAI21_X1 _0915_ (.A(_0309_),
    .B1(_0310_),
    .B2(_0311_),
    .ZN(_0312_));
 AOI21_X1 _0916_ (.A(_0517_),
    .B1(_0312_),
    .B2(_0518_),
    .ZN(_0313_));
 AOI221_X1 _0917_ (.A(_0112_),
    .B1(_0301_),
    .B2(_0302_),
    .C1(_0308_),
    .C2(_0313_),
    .ZN(_0013_));
 FA_X1 _0918_ (.A(_0320_),
    .B(net8),
    .CI(_0321_),
    .CO(_0322_),
    .S(_0323_));
 FA_X1 _0919_ (.A(_0320_),
    .B(_0324_),
    .CI(_0325_),
    .CO(_0326_),
    .S(_0327_));
 HA_X1 _0920_ (.A(_0328_),
    .B(net9),
    .CO(_0329_),
    .S(_0330_));
 HA_X1 _0921_ (.A(net3),
    .B(net9),
    .CO(_0331_),
    .S(_0332_));
 HA_X1 _0922_ (.A(_0333_),
    .B(_0334_),
    .CO(_0335_),
    .S(_0336_));
 HA_X1 _0923_ (.A(_0337_),
    .B(_0338_),
    .CO(_0339_),
    .S(_0340_));
 HA_X1 _0924_ (.A(_0341_),
    .B(_0342_),
    .CO(_0343_),
    .S(_0344_));
 HA_X1 _0925_ (.A(_0345_),
    .B(_0346_),
    .CO(_0347_),
    .S(_0348_));
 HA_X1 _0926_ (.A(_0349_),
    .B(_0350_),
    .CO(_0351_),
    .S(_0352_));
 HA_X1 _0927_ (.A(_0353_),
    .B(_0354_),
    .CO(_0355_),
    .S(_0356_));
 HA_X1 _0928_ (.A(_0323_),
    .B(\counter[1] ),
    .CO(_0358_),
    .S(_0359_));
 HA_X1 _0929_ (.A(net1),
    .B(_0360_),
    .CO(_0361_),
    .S(_0362_));
 HA_X1 _0930_ (.A(net1),
    .B(net7),
    .CO(_0363_),
    .S(_0364_));
 HA_X1 _0931_ (.A(_0365_),
    .B(_0366_),
    .CO(_0367_),
    .S(_0368_));
 HA_X1 _0932_ (.A(\counter[0] ),
    .B(_0366_),
    .CO(_0369_),
    .S(_0370_));
 HA_X1 _0933_ (.A(_0320_),
    .B(net8),
    .CO(_0371_),
    .S(_0357_));
 HA_X1 _0934_ (.A(net2),
    .B(net8),
    .CO(_0372_),
    .S(_0373_));
 HA_X1 _0935_ (.A(_0374_),
    .B(_0375_),
    .CO(_0376_),
    .S(_0377_));
 HA_X1 _0936_ (.A(\counter[1] ),
    .B(_0375_),
    .CO(_0378_),
    .S(_0379_));
 HA_X1 _0937_ (.A(_0380_),
    .B(net10),
    .CO(_0381_),
    .S(_0382_));
 HA_X1 _0938_ (.A(net4),
    .B(net10),
    .CO(_0383_),
    .S(_0384_));
 HA_X1 _0939_ (.A(\counter[3] ),
    .B(_0385_),
    .CO(_0386_),
    .S(_0387_));
 HA_X1 _0940_ (.A(\counter[2] ),
    .B(_0388_),
    .CO(_0389_),
    .S(_0390_));
 HA_X1 _0941_ (.A(_0391_),
    .B(net12),
    .CO(_0392_),
    .S(_0393_));
 HA_X1 _0942_ (.A(net6),
    .B(net12),
    .CO(_0394_),
    .S(_0395_));
 HA_X1 _0943_ (.A(_0396_),
    .B(net11),
    .CO(_0397_),
    .S(_0398_));
 HA_X1 _0944_ (.A(net5),
    .B(net11),
    .CO(_0399_),
    .S(_0400_));
 HA_X1 _0945_ (.A(\counter[5] ),
    .B(_0401_),
    .CO(_0402_),
    .S(_0403_));
 HA_X1 _0946_ (.A(\counter[4] ),
    .B(_0404_),
    .CO(_0405_),
    .S(_0406_));
 HA_X1 _0947_ (.A(_0341_),
    .B(_0391_),
    .CO(_0407_),
    .S(_0408_));
 HA_X1 _0948_ (.A(_0345_),
    .B(_0396_),
    .CO(_0409_),
    .S(_0410_));
 HA_X1 _0949_ (.A(_0349_),
    .B(_0380_),
    .CO(_0411_),
    .S(_0412_));
 HA_X1 _0950_ (.A(_0353_),
    .B(_0328_),
    .CO(_0413_),
    .S(_0414_));
 HA_X1 _0951_ (.A(_0334_),
    .B(_0415_),
    .CO(_0416_),
    .S(_0417_));
 HA_X1 _0952_ (.A(_0338_),
    .B(_0418_),
    .CO(_0419_),
    .S(_0420_));
 HA_X1 _0953_ (.A(_0342_),
    .B(_0421_),
    .CO(_0422_),
    .S(_0423_));
 HA_X1 _0954_ (.A(_0346_),
    .B(_0424_),
    .CO(_0425_),
    .S(_0426_));
 HA_X1 _0955_ (.A(_0350_),
    .B(_0427_),
    .CO(_0428_),
    .S(_0429_));
 HA_X1 _0956_ (.A(_0354_),
    .B(_0430_),
    .CO(_0431_),
    .S(_0432_));
 HA_X1 _0957_ (.A(\counter[0] ),
    .B(\counter[1] ),
    .CO(_0433_),
    .S(_0434_));
 HA_X1 _0958_ (.A(_0323_),
    .B(_0435_),
    .CO(_0436_),
    .S(_0437_));
 HA_X1 _0959_ (.A(_0365_),
    .B(_0362_),
    .CO(_0438_),
    .S(_0439_));
 HA_X1 _0960_ (.A(\counter[0] ),
    .B(_0362_),
    .CO(_0440_),
    .S(_0441_));
 HA_X1 _0961_ (.A(_0375_),
    .B(_0434_),
    .CO(_0442_),
    .S(_0443_));
 HA_X1 _0962_ (.A(_0385_),
    .B(_0444_),
    .CO(_0445_),
    .S(_0446_));
 HA_X1 _0963_ (.A(_0388_),
    .B(_0447_),
    .CO(_0448_),
    .S(_0449_));
 HA_X1 _0964_ (.A(_0401_),
    .B(_0450_),
    .CO(_0451_),
    .S(_0452_));
 HA_X1 _0965_ (.A(_0404_),
    .B(_0453_),
    .CO(_0454_),
    .S(_0455_));
 HA_X1 _0966_ (.A(_0391_),
    .B(_0421_),
    .CO(_0456_),
    .S(_0457_));
 HA_X1 _0967_ (.A(_0396_),
    .B(_0424_),
    .CO(_0458_),
    .S(_0459_));
 HA_X1 _0968_ (.A(_0380_),
    .B(_0427_),
    .CO(_0460_),
    .S(_0461_));
 HA_X1 _0969_ (.A(_0328_),
    .B(_0430_),
    .CO(_0462_),
    .S(_0463_));
 HA_X1 _0970_ (.A(_0320_),
    .B(_0435_),
    .CO(_0464_),
    .S(_0465_));
 HA_X1 _0971_ (.A(_0365_),
    .B(net1),
    .CO(_0466_),
    .S(_0467_));
 HA_X1 _0972_ (.A(\counter[0] ),
    .B(net1),
    .CO(_0468_),
    .S(_0469_));
 HA_X1 _0973_ (.A(_0470_),
    .B(_0334_),
    .CO(_0471_),
    .S(_0472_));
 HA_X1 _0974_ (.A(_0473_),
    .B(_0338_),
    .CO(_0474_),
    .S(_0475_));
 HA_X1 _0975_ (.A(_0476_),
    .B(_0342_),
    .CO(_0477_),
    .S(_0478_));
 HA_X1 _0976_ (.A(_0479_),
    .B(_0346_),
    .CO(_0480_),
    .S(_0481_));
 HA_X1 _0977_ (.A(_0482_),
    .B(_0350_),
    .CO(_0483_),
    .S(_0484_));
 HA_X1 _0978_ (.A(\counter[1] ),
    .B(_0353_),
    .CO(_0485_),
    .S(_0486_));
 HA_X1 _0979_ (.A(\counter[1] ),
    .B(\counter[2] ),
    .CO(_0487_),
    .S(_0488_));
 HA_X1 _0980_ (.A(_0486_),
    .B(_0354_),
    .CO(_0489_),
    .S(_0490_));
 HA_X1 _0981_ (.A(_0374_),
    .B(_0323_),
    .CO(_0491_),
    .S(_0492_));
 HA_X1 _0982_ (.A(_0493_),
    .B(_0385_),
    .CO(_0494_),
    .S(_0495_));
 HA_X1 _0983_ (.A(_0496_),
    .B(_0388_),
    .CO(_0497_),
    .S(_0498_));
 HA_X1 _0984_ (.A(_0499_),
    .B(_0401_),
    .CO(_0500_),
    .S(_0501_));
 HA_X1 _0985_ (.A(_0502_),
    .B(_0404_),
    .CO(_0503_),
    .S(_0504_));
 HA_X1 _0986_ (.A(_0391_),
    .B(_0476_),
    .CO(_0505_),
    .S(_0506_));
 HA_X1 _0987_ (.A(_0396_),
    .B(_0479_),
    .CO(_0507_),
    .S(_0508_));
 HA_X1 _0988_ (.A(_0380_),
    .B(_0482_),
    .CO(_0509_),
    .S(_0510_));
 HA_X1 _0989_ (.A(_0328_),
    .B(_0486_),
    .CO(_0511_),
    .S(_0512_));
 HA_X1 _0990_ (.A(_0374_),
    .B(_0320_),
    .CO(_0513_),
    .S(_0514_));
 HA_X1 _0991_ (.A(\counter[1] ),
    .B(_0320_),
    .CO(_0515_),
    .S(_0516_));
 HA_X1 _0992_ (.A(net14),
    .B(_0470_),
    .CO(_0517_),
    .S(_0518_));
 HA_X1 _0993_ (.A(net13),
    .B(_0473_),
    .CO(_0519_),
    .S(_0520_));
 HA_X1 _0994_ (.A(net12),
    .B(_0476_),
    .CO(_0521_),
    .S(_0522_));
 HA_X1 _0995_ (.A(net11),
    .B(_0479_),
    .CO(_0523_),
    .S(_0524_));
 HA_X1 _0996_ (.A(net10),
    .B(_0482_),
    .CO(_0525_),
    .S(_0526_));
 HA_X1 _0997_ (.A(net9),
    .B(_0486_),
    .CO(_0527_),
    .S(_0528_));
 HA_X1 _0998_ (.A(net14),
    .B(_0415_),
    .CO(_0529_),
    .S(_0530_));
 HA_X1 _0999_ (.A(net13),
    .B(_0418_),
    .CO(_0531_),
    .S(_0532_));
 HA_X1 _1000_ (.A(net12),
    .B(_0421_),
    .CO(_0533_),
    .S(_0534_));
 HA_X1 _1001_ (.A(net11),
    .B(_0424_),
    .CO(_0535_),
    .S(_0536_));
 HA_X1 _1002_ (.A(net10),
    .B(_0427_),
    .CO(_0537_),
    .S(_0538_));
 HA_X1 _1003_ (.A(net9),
    .B(_0430_),
    .CO(_0539_),
    .S(_0540_));
 HA_X1 _1004_ (.A(net8),
    .B(_0435_),
    .CO(_0541_),
    .S(_0542_));
 HA_X1 _1005_ (.A(_0365_),
    .B(_0360_),
    .CO(_0543_),
    .S(_0544_));
 HA_X1 _1006_ (.A(\counter[0] ),
    .B(_0360_),
    .CO(_0545_),
    .S(_0546_));
 HA_X1 _1007_ (.A(_0333_),
    .B(net14),
    .CO(_0547_),
    .S(_0548_));
 HA_X1 _1008_ (.A(_0337_),
    .B(net13),
    .CO(_0549_),
    .S(_0550_));
 HA_X1 _1009_ (.A(_0341_),
    .B(net12),
    .CO(_0551_),
    .S(_0552_));
 HA_X1 _1010_ (.A(_0345_),
    .B(net11),
    .CO(_0553_),
    .S(_0554_));
 HA_X1 _1011_ (.A(_0349_),
    .B(net10),
    .CO(_0555_),
    .S(_0556_));
 HA_X1 _1012_ (.A(_0353_),
    .B(net9),
    .CO(_0557_),
    .S(_0558_));
 HA_X1 _1013_ (.A(_0374_),
    .B(net8),
    .CO(_0559_),
    .S(_0560_));
 HA_X1 _1014_ (.A(\counter[1] ),
    .B(net8),
    .CO(_0561_),
    .S(_0562_));
 DFF_X2 \counter[0]$_SDFFE_PN0P_  (.D(_0000_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[0] ),
    .QN(_0365_));
 DFF_X2 \counter[1]$_SDFFE_PN0P_  (.D(_0001_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[1] ),
    .QN(_0374_));
 DFF_X2 \counter[2]$_SDFFE_PN0P_  (.D(_0002_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[2] ),
    .QN(_0353_));
 DFF_X2 \counter[3]$_SDFFE_PN0P_  (.D(_0003_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[3] ),
    .QN(_0349_));
 DFF_X2 \counter[4]$_SDFFE_PN0P_  (.D(_0004_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[4] ),
    .QN(_0345_));
 DFF_X2 \counter[5]$_SDFFE_PN0P_  (.D(_0005_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[5] ),
    .QN(_0341_));
 DFF_X2 \counter[6]$_SDFFE_PN0P_  (.D(_0006_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[6] ),
    .QN(_0337_));
 DFF_X2 \counter[7]$_SDFFE_PN0P_  (.D(_0007_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\counter[7] ),
    .QN(_0333_));
 DFF_X1 \pwm_n_reg[0]$_SDFF_PN0_  (.D(_0008_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net16),
    .QN(_0319_));
 DFF_X1 \pwm_n_reg[1]$_SDFF_PN0_  (.D(_0009_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net17),
    .QN(_0318_));
 DFF_X1 \pwm_n_reg[2]$_SDFF_PN0_  (.D(_0010_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net18),
    .QN(_0317_));
 DFF_X1 \pwm_p_reg[0]$_SDFF_PN0_  (.D(_0011_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net19),
    .QN(_0316_));
 DFF_X1 \pwm_p_reg[1]$_SDFF_PN0_  (.D(_0012_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net20),
    .QN(_0315_));
 DFF_X1 \pwm_p_reg[2]$_SDFF_PN0_  (.D(_0013_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net21),
    .QN(_0314_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_95 ();
 BUF_X2 input1 (.A(deadtime[0]),
    .Z(net1));
 BUF_X1 input2 (.A(deadtime[1]),
    .Z(net2));
 BUF_X1 input3 (.A(deadtime[2]),
    .Z(net3));
 BUF_X1 input4 (.A(deadtime[3]),
    .Z(net4));
 BUF_X1 input5 (.A(deadtime[4]),
    .Z(net5));
 BUF_X1 input6 (.A(deadtime[5]),
    .Z(net6));
 BUF_X1 input7 (.A(duty[0]),
    .Z(net7));
 BUF_X4 input8 (.A(duty[1]),
    .Z(net8));
 CLKBUF_X3 input9 (.A(duty[2]),
    .Z(net9));
 CLKBUF_X3 input10 (.A(duty[3]),
    .Z(net10));
 CLKBUF_X3 input11 (.A(duty[4]),
    .Z(net11));
 CLKBUF_X3 input12 (.A(duty[5]),
    .Z(net12));
 BUF_X2 input13 (.A(duty[6]),
    .Z(net13));
 CLKBUF_X3 input14 (.A(duty[7]),
    .Z(net14));
 CLKBUF_X2 input15 (.A(rst_n),
    .Z(net15));
 BUF_X1 output16 (.A(net16),
    .Z(pwm_n_out[0]));
 BUF_X1 output17 (.A(net17),
    .Z(pwm_n_out[1]));
 BUF_X1 output18 (.A(net18),
    .Z(pwm_n_out[2]));
 BUF_X1 output19 (.A(net19),
    .Z(pwm_p_out[0]));
 BUF_X1 output20 (.A(net20),
    .Z(pwm_p_out[1]));
 BUF_X1 output21 (.A(net21),
    .Z(pwm_p_out[2]));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 INV_X1 clkload0 (.A(clknet_1_0__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X16 FILLER_0_97 ();
 FILLCELL_X4 FILLER_0_113 ();
 FILLCELL_X1 FILLER_0_117 ();
 FILLCELL_X16 FILLER_0_123 ();
 FILLCELL_X8 FILLER_0_139 ();
 FILLCELL_X2 FILLER_0_147 ();
 FILLCELL_X1 FILLER_0_149 ();
 FILLCELL_X16 FILLER_0_155 ();
 FILLCELL_X8 FILLER_0_171 ();
 FILLCELL_X4 FILLER_0_179 ();
 FILLCELL_X4 FILLER_0_186 ();
 FILLCELL_X2 FILLER_0_190 ();
 FILLCELL_X8 FILLER_0_195 ();
 FILLCELL_X4 FILLER_0_203 ();
 FILLCELL_X8 FILLER_0_210 ();
 FILLCELL_X4 FILLER_0_218 ();
 FILLCELL_X2 FILLER_0_222 ();
 FILLCELL_X32 FILLER_0_236 ();
 FILLCELL_X32 FILLER_0_268 ();
 FILLCELL_X32 FILLER_0_300 ();
 FILLCELL_X16 FILLER_0_332 ();
 FILLCELL_X8 FILLER_0_348 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X16 FILLER_1_129 ();
 FILLCELL_X4 FILLER_1_145 ();
 FILLCELL_X1 FILLER_1_149 ();
 FILLCELL_X32 FILLER_1_153 ();
 FILLCELL_X4 FILLER_1_185 ();
 FILLCELL_X2 FILLER_1_189 ();
 FILLCELL_X8 FILLER_1_208 ();
 FILLCELL_X2 FILLER_1_216 ();
 FILLCELL_X32 FILLER_1_223 ();
 FILLCELL_X32 FILLER_1_255 ();
 FILLCELL_X32 FILLER_1_287 ();
 FILLCELL_X32 FILLER_1_319 ();
 FILLCELL_X4 FILLER_1_351 ();
 FILLCELL_X1 FILLER_1_355 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X16 FILLER_2_129 ();
 FILLCELL_X2 FILLER_2_145 ();
 FILLCELL_X1 FILLER_2_147 ();
 FILLCELL_X4 FILLER_2_161 ();
 FILLCELL_X2 FILLER_2_165 ();
 FILLCELL_X32 FILLER_2_184 ();
 FILLCELL_X32 FILLER_2_216 ();
 FILLCELL_X32 FILLER_2_248 ();
 FILLCELL_X32 FILLER_2_280 ();
 FILLCELL_X32 FILLER_2_312 ();
 FILLCELL_X8 FILLER_2_344 ();
 FILLCELL_X4 FILLER_2_352 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X16 FILLER_3_97 ();
 FILLCELL_X8 FILLER_3_113 ();
 FILLCELL_X1 FILLER_3_121 ();
 FILLCELL_X1 FILLER_3_136 ();
 FILLCELL_X2 FILLER_3_142 ();
 FILLCELL_X16 FILLER_3_154 ();
 FILLCELL_X4 FILLER_3_170 ();
 FILLCELL_X16 FILLER_3_191 ();
 FILLCELL_X4 FILLER_3_207 ();
 FILLCELL_X2 FILLER_3_211 ();
 FILLCELL_X32 FILLER_3_226 ();
 FILLCELL_X32 FILLER_3_258 ();
 FILLCELL_X32 FILLER_3_290 ();
 FILLCELL_X32 FILLER_3_322 ();
 FILLCELL_X2 FILLER_3_354 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X4 FILLER_4_97 ();
 FILLCELL_X2 FILLER_4_101 ();
 FILLCELL_X1 FILLER_4_103 ();
 FILLCELL_X2 FILLER_4_108 ();
 FILLCELL_X2 FILLER_4_112 ();
 FILLCELL_X1 FILLER_4_120 ();
 FILLCELL_X4 FILLER_4_123 ();
 FILLCELL_X8 FILLER_4_133 ();
 FILLCELL_X4 FILLER_4_151 ();
 FILLCELL_X4 FILLER_4_159 ();
 FILLCELL_X32 FILLER_4_179 ();
 FILLCELL_X8 FILLER_4_211 ();
 FILLCELL_X4 FILLER_4_219 ();
 FILLCELL_X32 FILLER_4_249 ();
 FILLCELL_X32 FILLER_4_281 ();
 FILLCELL_X32 FILLER_4_313 ();
 FILLCELL_X8 FILLER_4_345 ();
 FILLCELL_X2 FILLER_4_353 ();
 FILLCELL_X1 FILLER_4_355 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X2 FILLER_5_97 ();
 FILLCELL_X1 FILLER_5_99 ();
 FILLCELL_X1 FILLER_5_107 ();
 FILLCELL_X16 FILLER_5_124 ();
 FILLCELL_X8 FILLER_5_140 ();
 FILLCELL_X4 FILLER_5_148 ();
 FILLCELL_X1 FILLER_5_152 ();
 FILLCELL_X4 FILLER_5_163 ();
 FILLCELL_X16 FILLER_5_177 ();
 FILLCELL_X8 FILLER_5_193 ();
 FILLCELL_X2 FILLER_5_201 ();
 FILLCELL_X4 FILLER_5_209 ();
 FILLCELL_X8 FILLER_5_217 ();
 FILLCELL_X1 FILLER_5_225 ();
 FILLCELL_X1 FILLER_5_236 ();
 FILLCELL_X1 FILLER_5_247 ();
 FILLCELL_X32 FILLER_5_250 ();
 FILLCELL_X32 FILLER_5_282 ();
 FILLCELL_X32 FILLER_5_314 ();
 FILLCELL_X8 FILLER_5_346 ();
 FILLCELL_X2 FILLER_5_354 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X16 FILLER_6_65 ();
 FILLCELL_X8 FILLER_6_81 ();
 FILLCELL_X4 FILLER_6_89 ();
 FILLCELL_X2 FILLER_6_93 ();
 FILLCELL_X1 FILLER_6_95 ();
 FILLCELL_X4 FILLER_6_108 ();
 FILLCELL_X2 FILLER_6_112 ();
 FILLCELL_X1 FILLER_6_114 ();
 FILLCELL_X32 FILLER_6_117 ();
 FILLCELL_X8 FILLER_6_149 ();
 FILLCELL_X2 FILLER_6_157 ();
 FILLCELL_X1 FILLER_6_159 ();
 FILLCELL_X32 FILLER_6_168 ();
 FILLCELL_X32 FILLER_6_236 ();
 FILLCELL_X32 FILLER_6_268 ();
 FILLCELL_X32 FILLER_6_300 ();
 FILLCELL_X16 FILLER_6_332 ();
 FILLCELL_X8 FILLER_6_348 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X16 FILLER_7_65 ();
 FILLCELL_X8 FILLER_7_81 ();
 FILLCELL_X4 FILLER_7_89 ();
 FILLCELL_X2 FILLER_7_93 ();
 FILLCELL_X32 FILLER_7_105 ();
 FILLCELL_X16 FILLER_7_137 ();
 FILLCELL_X4 FILLER_7_153 ();
 FILLCELL_X2 FILLER_7_157 ();
 FILLCELL_X1 FILLER_7_159 ();
 FILLCELL_X32 FILLER_7_165 ();
 FILLCELL_X8 FILLER_7_197 ();
 FILLCELL_X4 FILLER_7_205 ();
 FILLCELL_X2 FILLER_7_209 ();
 FILLCELL_X4 FILLER_7_221 ();
 FILLCELL_X2 FILLER_7_225 ();
 FILLCELL_X1 FILLER_7_227 ();
 FILLCELL_X32 FILLER_7_238 ();
 FILLCELL_X32 FILLER_7_270 ();
 FILLCELL_X32 FILLER_7_302 ();
 FILLCELL_X16 FILLER_7_334 ();
 FILLCELL_X4 FILLER_7_350 ();
 FILLCELL_X2 FILLER_7_354 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X16 FILLER_8_97 ();
 FILLCELL_X8 FILLER_8_113 ();
 FILLCELL_X4 FILLER_8_121 ();
 FILLCELL_X8 FILLER_8_154 ();
 FILLCELL_X4 FILLER_8_162 ();
 FILLCELL_X1 FILLER_8_166 ();
 FILLCELL_X16 FILLER_8_187 ();
 FILLCELL_X2 FILLER_8_203 ();
 FILLCELL_X1 FILLER_8_205 ();
 FILLCELL_X32 FILLER_8_216 ();
 FILLCELL_X32 FILLER_8_248 ();
 FILLCELL_X32 FILLER_8_280 ();
 FILLCELL_X4 FILLER_8_312 ();
 FILLCELL_X2 FILLER_8_316 ();
 FILLCELL_X32 FILLER_8_323 ();
 FILLCELL_X1 FILLER_8_355 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X16 FILLER_9_97 ();
 FILLCELL_X8 FILLER_9_113 ();
 FILLCELL_X1 FILLER_9_121 ();
 FILLCELL_X2 FILLER_9_132 ();
 FILLCELL_X2 FILLER_9_138 ();
 FILLCELL_X1 FILLER_9_157 ();
 FILLCELL_X4 FILLER_9_165 ();
 FILLCELL_X1 FILLER_9_169 ();
 FILLCELL_X4 FILLER_9_180 ();
 FILLCELL_X1 FILLER_9_184 ();
 FILLCELL_X1 FILLER_9_187 ();
 FILLCELL_X32 FILLER_9_198 ();
 FILLCELL_X32 FILLER_9_230 ();
 FILLCELL_X32 FILLER_9_262 ();
 FILLCELL_X32 FILLER_9_294 ();
 FILLCELL_X16 FILLER_9_326 ();
 FILLCELL_X8 FILLER_9_342 ();
 FILLCELL_X4 FILLER_9_350 ();
 FILLCELL_X2 FILLER_9_354 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X8 FILLER_10_65 ();
 FILLCELL_X4 FILLER_10_73 ();
 FILLCELL_X2 FILLER_10_77 ();
 FILLCELL_X4 FILLER_10_113 ();
 FILLCELL_X2 FILLER_10_117 ();
 FILLCELL_X1 FILLER_10_119 ();
 FILLCELL_X16 FILLER_10_127 ();
 FILLCELL_X4 FILLER_10_143 ();
 FILLCELL_X16 FILLER_10_149 ();
 FILLCELL_X4 FILLER_10_165 ();
 FILLCELL_X2 FILLER_10_169 ();
 FILLCELL_X16 FILLER_10_176 ();
 FILLCELL_X8 FILLER_10_192 ();
 FILLCELL_X4 FILLER_10_200 ();
 FILLCELL_X2 FILLER_10_204 ();
 FILLCELL_X8 FILLER_10_209 ();
 FILLCELL_X4 FILLER_10_217 ();
 FILLCELL_X4 FILLER_10_241 ();
 FILLCELL_X2 FILLER_10_245 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X32 FILLER_10_289 ();
 FILLCELL_X32 FILLER_10_321 ();
 FILLCELL_X2 FILLER_10_353 ();
 FILLCELL_X1 FILLER_10_355 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X8 FILLER_11_65 ();
 FILLCELL_X4 FILLER_11_83 ();
 FILLCELL_X2 FILLER_11_87 ();
 FILLCELL_X1 FILLER_11_89 ();
 FILLCELL_X8 FILLER_11_94 ();
 FILLCELL_X1 FILLER_11_102 ();
 FILLCELL_X2 FILLER_11_107 ();
 FILLCELL_X1 FILLER_11_109 ();
 FILLCELL_X16 FILLER_11_121 ();
 FILLCELL_X4 FILLER_11_137 ();
 FILLCELL_X2 FILLER_11_141 ();
 FILLCELL_X2 FILLER_11_153 ();
 FILLCELL_X1 FILLER_11_155 ();
 FILLCELL_X32 FILLER_11_160 ();
 FILLCELL_X1 FILLER_11_203 ();
 FILLCELL_X8 FILLER_11_208 ();
 FILLCELL_X4 FILLER_11_216 ();
 FILLCELL_X32 FILLER_11_252 ();
 FILLCELL_X32 FILLER_11_284 ();
 FILLCELL_X32 FILLER_11_316 ();
 FILLCELL_X8 FILLER_11_348 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X8 FILLER_12_65 ();
 FILLCELL_X4 FILLER_12_73 ();
 FILLCELL_X8 FILLER_12_87 ();
 FILLCELL_X4 FILLER_12_95 ();
 FILLCELL_X1 FILLER_12_99 ();
 FILLCELL_X16 FILLER_12_120 ();
 FILLCELL_X4 FILLER_12_136 ();
 FILLCELL_X2 FILLER_12_140 ();
 FILLCELL_X8 FILLER_12_152 ();
 FILLCELL_X4 FILLER_12_160 ();
 FILLCELL_X1 FILLER_12_164 ();
 FILLCELL_X32 FILLER_12_175 ();
 FILLCELL_X16 FILLER_12_207 ();
 FILLCELL_X2 FILLER_12_223 ();
 FILLCELL_X1 FILLER_12_227 ();
 FILLCELL_X32 FILLER_12_232 ();
 FILLCELL_X32 FILLER_12_264 ();
 FILLCELL_X32 FILLER_12_296 ();
 FILLCELL_X16 FILLER_12_328 ();
 FILLCELL_X8 FILLER_12_344 ();
 FILLCELL_X4 FILLER_12_352 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X8 FILLER_13_65 ();
 FILLCELL_X4 FILLER_13_73 ();
 FILLCELL_X1 FILLER_13_77 ();
 FILLCELL_X2 FILLER_13_88 ();
 FILLCELL_X1 FILLER_13_90 ();
 FILLCELL_X1 FILLER_13_93 ();
 FILLCELL_X16 FILLER_13_108 ();
 FILLCELL_X4 FILLER_13_124 ();
 FILLCELL_X2 FILLER_13_128 ();
 FILLCELL_X4 FILLER_13_154 ();
 FILLCELL_X2 FILLER_13_158 ();
 FILLCELL_X1 FILLER_13_174 ();
 FILLCELL_X4 FILLER_13_179 ();
 FILLCELL_X2 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_205 ();
 FILLCELL_X32 FILLER_13_237 ();
 FILLCELL_X32 FILLER_13_269 ();
 FILLCELL_X32 FILLER_13_301 ();
 FILLCELL_X16 FILLER_13_333 ();
 FILLCELL_X4 FILLER_13_349 ();
 FILLCELL_X2 FILLER_13_353 ();
 FILLCELL_X1 FILLER_13_355 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X16 FILLER_14_129 ();
 FILLCELL_X1 FILLER_14_145 ();
 FILLCELL_X16 FILLER_14_148 ();
 FILLCELL_X4 FILLER_14_164 ();
 FILLCELL_X2 FILLER_14_168 ();
 FILLCELL_X16 FILLER_14_188 ();
 FILLCELL_X8 FILLER_14_204 ();
 FILLCELL_X4 FILLER_14_212 ();
 FILLCELL_X4 FILLER_14_226 ();
 FILLCELL_X1 FILLER_14_230 ();
 FILLCELL_X2 FILLER_14_234 ();
 FILLCELL_X32 FILLER_14_246 ();
 FILLCELL_X32 FILLER_14_278 ();
 FILLCELL_X4 FILLER_14_310 ();
 FILLCELL_X2 FILLER_14_314 ();
 FILLCELL_X1 FILLER_14_316 ();
 FILLCELL_X32 FILLER_14_320 ();
 FILLCELL_X4 FILLER_14_352 ();
 FILLCELL_X16 FILLER_15_1 ();
 FILLCELL_X8 FILLER_15_17 ();
 FILLCELL_X4 FILLER_15_25 ();
 FILLCELL_X1 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_37 ();
 FILLCELL_X32 FILLER_15_69 ();
 FILLCELL_X32 FILLER_15_101 ();
 FILLCELL_X8 FILLER_15_133 ();
 FILLCELL_X32 FILLER_15_145 ();
 FILLCELL_X16 FILLER_15_177 ();
 FILLCELL_X2 FILLER_15_193 ();
 FILLCELL_X16 FILLER_15_199 ();
 FILLCELL_X2 FILLER_15_215 ();
 FILLCELL_X2 FILLER_15_221 ();
 FILLCELL_X2 FILLER_15_228 ();
 FILLCELL_X1 FILLER_15_230 ();
 FILLCELL_X32 FILLER_15_236 ();
 FILLCELL_X32 FILLER_15_268 ();
 FILLCELL_X32 FILLER_15_300 ();
 FILLCELL_X16 FILLER_15_332 ();
 FILLCELL_X8 FILLER_15_348 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X16 FILLER_16_33 ();
 FILLCELL_X8 FILLER_16_61 ();
 FILLCELL_X4 FILLER_16_69 ();
 FILLCELL_X16 FILLER_16_83 ();
 FILLCELL_X8 FILLER_16_99 ();
 FILLCELL_X8 FILLER_16_130 ();
 FILLCELL_X4 FILLER_16_138 ();
 FILLCELL_X1 FILLER_16_142 ();
 FILLCELL_X4 FILLER_16_154 ();
 FILLCELL_X1 FILLER_16_158 ();
 FILLCELL_X32 FILLER_16_164 ();
 FILLCELL_X16 FILLER_16_196 ();
 FILLCELL_X4 FILLER_16_212 ();
 FILLCELL_X1 FILLER_16_218 ();
 FILLCELL_X32 FILLER_16_243 ();
 FILLCELL_X32 FILLER_16_275 ();
 FILLCELL_X32 FILLER_16_307 ();
 FILLCELL_X16 FILLER_16_339 ();
 FILLCELL_X1 FILLER_16_355 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X16 FILLER_17_33 ();
 FILLCELL_X4 FILLER_17_49 ();
 FILLCELL_X2 FILLER_17_53 ();
 FILLCELL_X1 FILLER_17_55 ();
 FILLCELL_X2 FILLER_17_79 ();
 FILLCELL_X16 FILLER_17_85 ();
 FILLCELL_X8 FILLER_17_101 ();
 FILLCELL_X4 FILLER_17_109 ();
 FILLCELL_X2 FILLER_17_113 ();
 FILLCELL_X1 FILLER_17_115 ();
 FILLCELL_X16 FILLER_17_123 ();
 FILLCELL_X2 FILLER_17_139 ();
 FILLCELL_X2 FILLER_17_152 ();
 FILLCELL_X1 FILLER_17_161 ();
 FILLCELL_X16 FILLER_17_176 ();
 FILLCELL_X4 FILLER_17_192 ();
 FILLCELL_X2 FILLER_17_196 ();
 FILLCELL_X1 FILLER_17_209 ();
 FILLCELL_X32 FILLER_17_252 ();
 FILLCELL_X32 FILLER_17_284 ();
 FILLCELL_X32 FILLER_17_316 ();
 FILLCELL_X8 FILLER_17_348 ();
 FILLCELL_X8 FILLER_18_1 ();
 FILLCELL_X2 FILLER_18_9 ();
 FILLCELL_X32 FILLER_18_14 ();
 FILLCELL_X8 FILLER_18_46 ();
 FILLCELL_X2 FILLER_18_54 ();
 FILLCELL_X2 FILLER_18_58 ();
 FILLCELL_X16 FILLER_18_85 ();
 FILLCELL_X8 FILLER_18_101 ();
 FILLCELL_X8 FILLER_18_121 ();
 FILLCELL_X4 FILLER_18_129 ();
 FILLCELL_X1 FILLER_18_133 ();
 FILLCELL_X16 FILLER_18_172 ();
 FILLCELL_X2 FILLER_18_188 ();
 FILLCELL_X4 FILLER_18_214 ();
 FILLCELL_X2 FILLER_18_218 ();
 FILLCELL_X1 FILLER_18_220 ();
 FILLCELL_X32 FILLER_18_246 ();
 FILLCELL_X32 FILLER_18_278 ();
 FILLCELL_X32 FILLER_18_310 ();
 FILLCELL_X8 FILLER_18_342 ();
 FILLCELL_X4 FILLER_18_350 ();
 FILLCELL_X2 FILLER_18_354 ();
 FILLCELL_X2 FILLER_19_1 ();
 FILLCELL_X1 FILLER_19_3 ();
 FILLCELL_X32 FILLER_19_7 ();
 FILLCELL_X8 FILLER_19_39 ();
 FILLCELL_X2 FILLER_19_47 ();
 FILLCELL_X2 FILLER_19_59 ();
 FILLCELL_X1 FILLER_19_61 ();
 FILLCELL_X8 FILLER_19_65 ();
 FILLCELL_X2 FILLER_19_73 ();
 FILLCELL_X2 FILLER_19_77 ();
 FILLCELL_X1 FILLER_19_79 ();
 FILLCELL_X4 FILLER_19_96 ();
 FILLCELL_X2 FILLER_19_110 ();
 FILLCELL_X1 FILLER_19_112 ();
 FILLCELL_X4 FILLER_19_122 ();
 FILLCELL_X2 FILLER_19_126 ();
 FILLCELL_X1 FILLER_19_151 ();
 FILLCELL_X4 FILLER_19_161 ();
 FILLCELL_X2 FILLER_19_165 ();
 FILLCELL_X1 FILLER_19_167 ();
 FILLCELL_X8 FILLER_19_178 ();
 FILLCELL_X8 FILLER_19_196 ();
 FILLCELL_X4 FILLER_19_204 ();
 FILLCELL_X1 FILLER_19_208 ();
 FILLCELL_X8 FILLER_19_229 ();
 FILLCELL_X2 FILLER_19_237 ();
 FILLCELL_X32 FILLER_19_253 ();
 FILLCELL_X32 FILLER_19_285 ();
 FILLCELL_X32 FILLER_19_317 ();
 FILLCELL_X4 FILLER_19_349 ();
 FILLCELL_X2 FILLER_19_353 ();
 FILLCELL_X1 FILLER_19_355 ();
 FILLCELL_X16 FILLER_20_1 ();
 FILLCELL_X4 FILLER_20_17 ();
 FILLCELL_X1 FILLER_20_21 ();
 FILLCELL_X32 FILLER_20_29 ();
 FILLCELL_X32 FILLER_20_61 ();
 FILLCELL_X32 FILLER_20_93 ();
 FILLCELL_X16 FILLER_20_125 ();
 FILLCELL_X4 FILLER_20_141 ();
 FILLCELL_X2 FILLER_20_145 ();
 FILLCELL_X1 FILLER_20_147 ();
 FILLCELL_X32 FILLER_20_158 ();
 FILLCELL_X32 FILLER_20_190 ();
 FILLCELL_X16 FILLER_20_222 ();
 FILLCELL_X2 FILLER_20_238 ();
 FILLCELL_X1 FILLER_20_240 ();
 FILLCELL_X32 FILLER_20_253 ();
 FILLCELL_X32 FILLER_20_285 ();
 FILLCELL_X32 FILLER_20_317 ();
 FILLCELL_X4 FILLER_20_349 ();
 FILLCELL_X2 FILLER_20_353 ();
 FILLCELL_X1 FILLER_20_355 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X32 FILLER_21_193 ();
 FILLCELL_X16 FILLER_21_225 ();
 FILLCELL_X1 FILLER_21_241 ();
 FILLCELL_X32 FILLER_21_256 ();
 FILLCELL_X32 FILLER_21_288 ();
 FILLCELL_X32 FILLER_21_320 ();
 FILLCELL_X4 FILLER_21_352 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X1 FILLER_22_97 ();
 FILLCELL_X8 FILLER_22_108 ();
 FILLCELL_X4 FILLER_22_116 ();
 FILLCELL_X32 FILLER_22_130 ();
 FILLCELL_X2 FILLER_22_162 ();
 FILLCELL_X1 FILLER_22_174 ();
 FILLCELL_X8 FILLER_22_177 ();
 FILLCELL_X4 FILLER_22_185 ();
 FILLCELL_X1 FILLER_22_189 ();
 FILLCELL_X16 FILLER_22_195 ();
 FILLCELL_X1 FILLER_22_221 ();
 FILLCELL_X4 FILLER_22_232 ();
 FILLCELL_X2 FILLER_22_236 ();
 FILLCELL_X32 FILLER_22_262 ();
 FILLCELL_X32 FILLER_22_294 ();
 FILLCELL_X16 FILLER_22_326 ();
 FILLCELL_X8 FILLER_22_342 ();
 FILLCELL_X4 FILLER_22_350 ();
 FILLCELL_X2 FILLER_22_354 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X8 FILLER_23_65 ();
 FILLCELL_X2 FILLER_23_73 ();
 FILLCELL_X4 FILLER_23_85 ();
 FILLCELL_X1 FILLER_23_89 ();
 FILLCELL_X1 FILLER_23_107 ();
 FILLCELL_X2 FILLER_23_118 ();
 FILLCELL_X1 FILLER_23_120 ();
 FILLCELL_X8 FILLER_23_123 ();
 FILLCELL_X1 FILLER_23_131 ();
 FILLCELL_X4 FILLER_23_170 ();
 FILLCELL_X2 FILLER_23_174 ();
 FILLCELL_X1 FILLER_23_176 ();
 FILLCELL_X16 FILLER_23_190 ();
 FILLCELL_X1 FILLER_23_225 ();
 FILLCELL_X8 FILLER_23_228 ();
 FILLCELL_X4 FILLER_23_241 ();
 FILLCELL_X32 FILLER_23_259 ();
 FILLCELL_X32 FILLER_23_291 ();
 FILLCELL_X32 FILLER_23_323 ();
 FILLCELL_X1 FILLER_23_355 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X16 FILLER_24_65 ();
 FILLCELL_X4 FILLER_24_91 ();
 FILLCELL_X1 FILLER_24_110 ();
 FILLCELL_X4 FILLER_24_113 ();
 FILLCELL_X1 FILLER_24_117 ();
 FILLCELL_X1 FILLER_24_128 ();
 FILLCELL_X2 FILLER_24_135 ();
 FILLCELL_X1 FILLER_24_137 ();
 FILLCELL_X4 FILLER_24_155 ();
 FILLCELL_X8 FILLER_24_164 ();
 FILLCELL_X1 FILLER_24_172 ();
 FILLCELL_X16 FILLER_24_186 ();
 FILLCELL_X4 FILLER_24_202 ();
 FILLCELL_X1 FILLER_24_206 ();
 FILLCELL_X16 FILLER_24_218 ();
 FILLCELL_X8 FILLER_24_234 ();
 FILLCELL_X1 FILLER_24_242 ();
 FILLCELL_X32 FILLER_24_260 ();
 FILLCELL_X16 FILLER_24_292 ();
 FILLCELL_X8 FILLER_24_308 ();
 FILLCELL_X2 FILLER_24_316 ();
 FILLCELL_X32 FILLER_24_321 ();
 FILLCELL_X2 FILLER_24_353 ();
 FILLCELL_X1 FILLER_24_355 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X8 FILLER_25_65 ();
 FILLCELL_X4 FILLER_25_73 ();
 FILLCELL_X4 FILLER_25_93 ();
 FILLCELL_X2 FILLER_25_97 ();
 FILLCELL_X16 FILLER_25_102 ();
 FILLCELL_X8 FILLER_25_118 ();
 FILLCELL_X1 FILLER_25_126 ();
 FILLCELL_X8 FILLER_25_133 ();
 FILLCELL_X4 FILLER_25_141 ();
 FILLCELL_X2 FILLER_25_145 ();
 FILLCELL_X1 FILLER_25_147 ();
 FILLCELL_X2 FILLER_25_162 ();
 FILLCELL_X1 FILLER_25_164 ();
 FILLCELL_X2 FILLER_25_168 ();
 FILLCELL_X4 FILLER_25_174 ();
 FILLCELL_X2 FILLER_25_178 ();
 FILLCELL_X16 FILLER_25_184 ();
 FILLCELL_X8 FILLER_25_200 ();
 FILLCELL_X2 FILLER_25_208 ();
 FILLCELL_X16 FILLER_25_216 ();
 FILLCELL_X8 FILLER_25_232 ();
 FILLCELL_X1 FILLER_25_240 ();
 FILLCELL_X16 FILLER_25_245 ();
 FILLCELL_X8 FILLER_25_261 ();
 FILLCELL_X2 FILLER_25_269 ();
 FILLCELL_X32 FILLER_25_288 ();
 FILLCELL_X32 FILLER_25_320 ();
 FILLCELL_X4 FILLER_25_352 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X8 FILLER_26_65 ();
 FILLCELL_X4 FILLER_26_73 ();
 FILLCELL_X1 FILLER_26_77 ();
 FILLCELL_X8 FILLER_26_80 ();
 FILLCELL_X32 FILLER_26_91 ();
 FILLCELL_X32 FILLER_26_123 ();
 FILLCELL_X32 FILLER_26_155 ();
 FILLCELL_X1 FILLER_26_187 ();
 FILLCELL_X8 FILLER_26_191 ();
 FILLCELL_X4 FILLER_26_199 ();
 FILLCELL_X2 FILLER_26_203 ();
 FILLCELL_X1 FILLER_26_205 ();
 FILLCELL_X16 FILLER_26_219 ();
 FILLCELL_X8 FILLER_26_235 ();
 FILLCELL_X2 FILLER_26_243 ();
 FILLCELL_X1 FILLER_26_245 ();
 FILLCELL_X32 FILLER_26_248 ();
 FILLCELL_X32 FILLER_26_280 ();
 FILLCELL_X32 FILLER_26_312 ();
 FILLCELL_X8 FILLER_26_344 ();
 FILLCELL_X4 FILLER_26_352 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X16 FILLER_27_65 ();
 FILLCELL_X2 FILLER_27_81 ();
 FILLCELL_X32 FILLER_27_85 ();
 FILLCELL_X16 FILLER_27_117 ();
 FILLCELL_X8 FILLER_27_133 ();
 FILLCELL_X4 FILLER_27_141 ();
 FILLCELL_X32 FILLER_27_148 ();
 FILLCELL_X16 FILLER_27_180 ();
 FILLCELL_X8 FILLER_27_196 ();
 FILLCELL_X4 FILLER_27_204 ();
 FILLCELL_X2 FILLER_27_208 ();
 FILLCELL_X32 FILLER_27_217 ();
 FILLCELL_X2 FILLER_27_249 ();
 FILLCELL_X1 FILLER_27_251 ();
 FILLCELL_X8 FILLER_27_257 ();
 FILLCELL_X4 FILLER_27_265 ();
 FILLCELL_X2 FILLER_27_269 ();
 FILLCELL_X32 FILLER_27_288 ();
 FILLCELL_X32 FILLER_27_320 ();
 FILLCELL_X4 FILLER_27_352 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X4 FILLER_28_97 ();
 FILLCELL_X2 FILLER_28_101 ();
 FILLCELL_X1 FILLER_28_103 ();
 FILLCELL_X32 FILLER_28_116 ();
 FILLCELL_X8 FILLER_28_148 ();
 FILLCELL_X4 FILLER_28_156 ();
 FILLCELL_X1 FILLER_28_160 ();
 FILLCELL_X8 FILLER_28_171 ();
 FILLCELL_X2 FILLER_28_179 ();
 FILLCELL_X1 FILLER_28_181 ();
 FILLCELL_X8 FILLER_28_185 ();
 FILLCELL_X1 FILLER_28_193 ();
 FILLCELL_X32 FILLER_28_197 ();
 FILLCELL_X4 FILLER_28_229 ();
 FILLCELL_X8 FILLER_28_238 ();
 FILLCELL_X1 FILLER_28_246 ();
 FILLCELL_X32 FILLER_28_255 ();
 FILLCELL_X16 FILLER_28_287 ();
 FILLCELL_X8 FILLER_28_303 ();
 FILLCELL_X4 FILLER_28_311 ();
 FILLCELL_X2 FILLER_28_315 ();
 FILLCELL_X32 FILLER_28_320 ();
 FILLCELL_X4 FILLER_28_352 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X4 FILLER_29_65 ();
 FILLCELL_X1 FILLER_29_69 ();
 FILLCELL_X1 FILLER_29_96 ();
 FILLCELL_X16 FILLER_29_111 ();
 FILLCELL_X8 FILLER_29_131 ();
 FILLCELL_X4 FILLER_29_139 ();
 FILLCELL_X1 FILLER_29_155 ();
 FILLCELL_X1 FILLER_29_166 ();
 FILLCELL_X4 FILLER_29_171 ();
 FILLCELL_X2 FILLER_29_175 ();
 FILLCELL_X1 FILLER_29_177 ();
 FILLCELL_X32 FILLER_29_202 ();
 FILLCELL_X2 FILLER_29_234 ();
 FILLCELL_X1 FILLER_29_236 ();
 FILLCELL_X32 FILLER_29_261 ();
 FILLCELL_X32 FILLER_29_293 ();
 FILLCELL_X16 FILLER_29_325 ();
 FILLCELL_X8 FILLER_29_341 ();
 FILLCELL_X4 FILLER_29_349 ();
 FILLCELL_X2 FILLER_29_353 ();
 FILLCELL_X1 FILLER_29_355 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X8 FILLER_30_65 ();
 FILLCELL_X2 FILLER_30_73 ();
 FILLCELL_X1 FILLER_30_75 ();
 FILLCELL_X2 FILLER_30_79 ();
 FILLCELL_X4 FILLER_30_107 ();
 FILLCELL_X1 FILLER_30_111 ();
 FILLCELL_X1 FILLER_30_122 ();
 FILLCELL_X2 FILLER_30_143 ();
 FILLCELL_X16 FILLER_30_148 ();
 FILLCELL_X8 FILLER_30_164 ();
 FILLCELL_X4 FILLER_30_172 ();
 FILLCELL_X1 FILLER_30_176 ();
 FILLCELL_X1 FILLER_30_192 ();
 FILLCELL_X32 FILLER_30_204 ();
 FILLCELL_X4 FILLER_30_236 ();
 FILLCELL_X2 FILLER_30_240 ();
 FILLCELL_X1 FILLER_30_242 ();
 FILLCELL_X32 FILLER_30_260 ();
 FILLCELL_X32 FILLER_30_292 ();
 FILLCELL_X32 FILLER_30_324 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X8 FILLER_31_65 ();
 FILLCELL_X4 FILLER_31_73 ();
 FILLCELL_X2 FILLER_31_77 ();
 FILLCELL_X1 FILLER_31_79 ();
 FILLCELL_X2 FILLER_31_84 ();
 FILLCELL_X2 FILLER_31_90 ();
 FILLCELL_X16 FILLER_31_122 ();
 FILLCELL_X4 FILLER_31_138 ();
 FILLCELL_X2 FILLER_31_142 ();
 FILLCELL_X1 FILLER_31_144 ();
 FILLCELL_X2 FILLER_31_159 ();
 FILLCELL_X2 FILLER_31_165 ();
 FILLCELL_X16 FILLER_31_199 ();
 FILLCELL_X8 FILLER_31_215 ();
 FILLCELL_X4 FILLER_31_223 ();
 FILLCELL_X1 FILLER_31_227 ();
 FILLCELL_X32 FILLER_31_250 ();
 FILLCELL_X32 FILLER_31_282 ();
 FILLCELL_X32 FILLER_31_314 ();
 FILLCELL_X8 FILLER_31_346 ();
 FILLCELL_X2 FILLER_31_354 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X8 FILLER_32_225 ();
 FILLCELL_X4 FILLER_32_233 ();
 FILLCELL_X32 FILLER_32_254 ();
 FILLCELL_X8 FILLER_32_303 ();
 FILLCELL_X4 FILLER_32_311 ();
 FILLCELL_X2 FILLER_32_315 ();
 FILLCELL_X32 FILLER_32_320 ();
 FILLCELL_X4 FILLER_32_352 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X16 FILLER_33_97 ();
 FILLCELL_X4 FILLER_33_113 ();
 FILLCELL_X32 FILLER_33_120 ();
 FILLCELL_X32 FILLER_33_152 ();
 FILLCELL_X32 FILLER_33_184 ();
 FILLCELL_X16 FILLER_33_216 ();
 FILLCELL_X2 FILLER_33_232 ();
 FILLCELL_X1 FILLER_33_234 ();
 FILLCELL_X32 FILLER_33_239 ();
 FILLCELL_X32 FILLER_33_271 ();
 FILLCELL_X32 FILLER_33_303 ();
 FILLCELL_X16 FILLER_33_335 ();
 FILLCELL_X4 FILLER_33_351 ();
 FILLCELL_X1 FILLER_33_355 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X16 FILLER_34_65 ();
 FILLCELL_X4 FILLER_34_81 ();
 FILLCELL_X1 FILLER_34_85 ();
 FILLCELL_X8 FILLER_34_105 ();
 FILLCELL_X2 FILLER_34_113 ();
 FILLCELL_X1 FILLER_34_115 ();
 FILLCELL_X2 FILLER_34_125 ();
 FILLCELL_X2 FILLER_34_137 ();
 FILLCELL_X1 FILLER_34_139 ();
 FILLCELL_X32 FILLER_34_149 ();
 FILLCELL_X2 FILLER_34_181 ();
 FILLCELL_X4 FILLER_34_193 ();
 FILLCELL_X2 FILLER_34_197 ();
 FILLCELL_X16 FILLER_34_209 ();
 FILLCELL_X8 FILLER_34_225 ();
 FILLCELL_X1 FILLER_34_238 ();
 FILLCELL_X1 FILLER_34_242 ();
 FILLCELL_X32 FILLER_34_249 ();
 FILLCELL_X32 FILLER_34_281 ();
 FILLCELL_X32 FILLER_34_313 ();
 FILLCELL_X8 FILLER_34_345 ();
 FILLCELL_X2 FILLER_34_353 ();
 FILLCELL_X1 FILLER_34_355 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X16 FILLER_35_107 ();
 FILLCELL_X4 FILLER_35_123 ();
 FILLCELL_X4 FILLER_35_131 ();
 FILLCELL_X1 FILLER_35_135 ();
 FILLCELL_X2 FILLER_35_139 ();
 FILLCELL_X1 FILLER_35_141 ();
 FILLCELL_X2 FILLER_35_146 ();
 FILLCELL_X8 FILLER_35_159 ();
 FILLCELL_X8 FILLER_35_195 ();
 FILLCELL_X4 FILLER_35_215 ();
 FILLCELL_X2 FILLER_35_219 ();
 FILLCELL_X1 FILLER_35_221 ();
 FILLCELL_X1 FILLER_35_232 ();
 FILLCELL_X1 FILLER_35_235 ();
 FILLCELL_X32 FILLER_35_243 ();
 FILLCELL_X32 FILLER_35_275 ();
 FILLCELL_X32 FILLER_35_307 ();
 FILLCELL_X16 FILLER_35_339 ();
 FILLCELL_X1 FILLER_35_355 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X16 FILLER_36_65 ();
 FILLCELL_X8 FILLER_36_81 ();
 FILLCELL_X1 FILLER_36_89 ();
 FILLCELL_X2 FILLER_36_98 ();
 FILLCELL_X1 FILLER_36_135 ();
 FILLCELL_X2 FILLER_36_169 ();
 FILLCELL_X1 FILLER_36_171 ();
 FILLCELL_X2 FILLER_36_189 ();
 FILLCELL_X1 FILLER_36_194 ();
 FILLCELL_X2 FILLER_36_205 ();
 FILLCELL_X8 FILLER_36_221 ();
 FILLCELL_X1 FILLER_36_229 ();
 FILLCELL_X1 FILLER_36_235 ();
 FILLCELL_X4 FILLER_36_241 ();
 FILLCELL_X2 FILLER_36_245 ();
 FILLCELL_X1 FILLER_36_247 ();
 FILLCELL_X32 FILLER_36_252 ();
 FILLCELL_X32 FILLER_36_284 ();
 FILLCELL_X32 FILLER_36_316 ();
 FILLCELL_X8 FILLER_36_348 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X8 FILLER_37_65 ();
 FILLCELL_X1 FILLER_37_73 ();
 FILLCELL_X1 FILLER_37_101 ();
 FILLCELL_X8 FILLER_37_105 ();
 FILLCELL_X4 FILLER_37_113 ();
 FILLCELL_X16 FILLER_37_125 ();
 FILLCELL_X1 FILLER_37_141 ();
 FILLCELL_X4 FILLER_37_146 ();
 FILLCELL_X1 FILLER_37_150 ();
 FILLCELL_X16 FILLER_37_155 ();
 FILLCELL_X8 FILLER_37_171 ();
 FILLCELL_X4 FILLER_37_179 ();
 FILLCELL_X2 FILLER_37_183 ();
 FILLCELL_X16 FILLER_37_201 ();
 FILLCELL_X4 FILLER_37_217 ();
 FILLCELL_X2 FILLER_37_221 ();
 FILLCELL_X1 FILLER_37_223 ();
 FILLCELL_X2 FILLER_37_229 ();
 FILLCELL_X32 FILLER_37_261 ();
 FILLCELL_X32 FILLER_37_293 ();
 FILLCELL_X16 FILLER_37_325 ();
 FILLCELL_X8 FILLER_37_341 ();
 FILLCELL_X4 FILLER_37_349 ();
 FILLCELL_X2 FILLER_37_353 ();
 FILLCELL_X1 FILLER_37_355 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X2 FILLER_38_161 ();
 FILLCELL_X1 FILLER_38_163 ();
 FILLCELL_X8 FILLER_38_167 ();
 FILLCELL_X2 FILLER_38_175 ();
 FILLCELL_X32 FILLER_38_180 ();
 FILLCELL_X16 FILLER_38_212 ();
 FILLCELL_X4 FILLER_38_228 ();
 FILLCELL_X2 FILLER_38_232 ();
 FILLCELL_X1 FILLER_38_234 ();
 FILLCELL_X32 FILLER_38_242 ();
 FILLCELL_X32 FILLER_38_274 ();
 FILLCELL_X32 FILLER_38_306 ();
 FILLCELL_X16 FILLER_38_338 ();
 FILLCELL_X2 FILLER_38_354 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X8 FILLER_39_129 ();
 FILLCELL_X4 FILLER_39_137 ();
 FILLCELL_X2 FILLER_39_141 ();
 FILLCELL_X4 FILLER_39_151 ();
 FILLCELL_X2 FILLER_39_155 ();
 FILLCELL_X1 FILLER_39_157 ();
 FILLCELL_X4 FILLER_39_169 ();
 FILLCELL_X2 FILLER_39_177 ();
 FILLCELL_X1 FILLER_39_179 ();
 FILLCELL_X8 FILLER_39_184 ();
 FILLCELL_X4 FILLER_39_192 ();
 FILLCELL_X1 FILLER_39_196 ();
 FILLCELL_X4 FILLER_39_201 ();
 FILLCELL_X2 FILLER_39_205 ();
 FILLCELL_X1 FILLER_39_207 ();
 FILLCELL_X8 FILLER_39_214 ();
 FILLCELL_X4 FILLER_39_222 ();
 FILLCELL_X1 FILLER_39_226 ();
 FILLCELL_X2 FILLER_39_246 ();
 FILLCELL_X32 FILLER_39_251 ();
 FILLCELL_X32 FILLER_39_283 ();
 FILLCELL_X32 FILLER_39_315 ();
 FILLCELL_X8 FILLER_39_347 ();
 FILLCELL_X1 FILLER_39_355 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X2 FILLER_40_129 ();
 FILLCELL_X2 FILLER_40_136 ();
 FILLCELL_X1 FILLER_40_138 ();
 FILLCELL_X4 FILLER_40_147 ();
 FILLCELL_X8 FILLER_40_158 ();
 FILLCELL_X2 FILLER_40_166 ();
 FILLCELL_X1 FILLER_40_168 ();
 FILLCELL_X8 FILLER_40_172 ();
 FILLCELL_X2 FILLER_40_180 ();
 FILLCELL_X2 FILLER_40_188 ();
 FILLCELL_X1 FILLER_40_190 ();
 FILLCELL_X8 FILLER_40_210 ();
 FILLCELL_X4 FILLER_40_218 ();
 FILLCELL_X2 FILLER_40_226 ();
 FILLCELL_X32 FILLER_40_235 ();
 FILLCELL_X32 FILLER_40_267 ();
 FILLCELL_X32 FILLER_40_299 ();
 FILLCELL_X16 FILLER_40_331 ();
 FILLCELL_X8 FILLER_40_347 ();
 FILLCELL_X1 FILLER_40_355 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X16 FILLER_41_148 ();
 FILLCELL_X2 FILLER_41_164 ();
 FILLCELL_X1 FILLER_41_166 ();
 FILLCELL_X1 FILLER_41_190 ();
 FILLCELL_X32 FILLER_41_198 ();
 FILLCELL_X2 FILLER_41_230 ();
 FILLCELL_X32 FILLER_41_244 ();
 FILLCELL_X32 FILLER_41_276 ();
 FILLCELL_X32 FILLER_41_308 ();
 FILLCELL_X16 FILLER_41_340 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X32 FILLER_42_129 ();
 FILLCELL_X32 FILLER_42_161 ();
 FILLCELL_X32 FILLER_42_193 ();
 FILLCELL_X32 FILLER_42_225 ();
 FILLCELL_X32 FILLER_42_257 ();
 FILLCELL_X32 FILLER_42_289 ();
 FILLCELL_X32 FILLER_42_321 ();
 FILLCELL_X2 FILLER_42_353 ();
 FILLCELL_X1 FILLER_42_355 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X4 FILLER_43_97 ();
 FILLCELL_X2 FILLER_43_101 ();
 FILLCELL_X32 FILLER_43_110 ();
 FILLCELL_X32 FILLER_43_142 ();
 FILLCELL_X32 FILLER_43_174 ();
 FILLCELL_X32 FILLER_43_206 ();
 FILLCELL_X32 FILLER_43_238 ();
 FILLCELL_X32 FILLER_43_270 ();
 FILLCELL_X32 FILLER_43_302 ();
 FILLCELL_X16 FILLER_43_334 ();
 FILLCELL_X4 FILLER_43_350 ();
 FILLCELL_X2 FILLER_43_354 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X32 FILLER_44_65 ();
 FILLCELL_X32 FILLER_44_97 ();
 FILLCELL_X32 FILLER_44_129 ();
 FILLCELL_X32 FILLER_44_161 ();
 FILLCELL_X32 FILLER_44_193 ();
 FILLCELL_X32 FILLER_44_225 ();
 FILLCELL_X32 FILLER_44_257 ();
 FILLCELL_X32 FILLER_44_289 ();
 FILLCELL_X32 FILLER_44_321 ();
 FILLCELL_X2 FILLER_44_353 ();
 FILLCELL_X1 FILLER_44_355 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X32 FILLER_45_65 ();
 FILLCELL_X32 FILLER_45_97 ();
 FILLCELL_X32 FILLER_45_129 ();
 FILLCELL_X32 FILLER_45_161 ();
 FILLCELL_X32 FILLER_45_193 ();
 FILLCELL_X32 FILLER_45_225 ();
 FILLCELL_X32 FILLER_45_257 ();
 FILLCELL_X32 FILLER_45_289 ();
 FILLCELL_X32 FILLER_45_321 ();
 FILLCELL_X2 FILLER_45_353 ();
 FILLCELL_X1 FILLER_45_355 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X32 FILLER_46_33 ();
 FILLCELL_X32 FILLER_46_65 ();
 FILLCELL_X32 FILLER_46_97 ();
 FILLCELL_X32 FILLER_46_129 ();
 FILLCELL_X32 FILLER_46_161 ();
 FILLCELL_X32 FILLER_46_193 ();
 FILLCELL_X32 FILLER_46_225 ();
 FILLCELL_X32 FILLER_46_257 ();
 FILLCELL_X32 FILLER_46_289 ();
 FILLCELL_X32 FILLER_46_321 ();
 FILLCELL_X2 FILLER_46_353 ();
 FILLCELL_X1 FILLER_46_355 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X32 FILLER_47_33 ();
 FILLCELL_X32 FILLER_47_65 ();
 FILLCELL_X32 FILLER_47_97 ();
 FILLCELL_X32 FILLER_47_129 ();
 FILLCELL_X32 FILLER_47_161 ();
 FILLCELL_X32 FILLER_47_193 ();
 FILLCELL_X8 FILLER_47_225 ();
 FILLCELL_X2 FILLER_47_233 ();
 FILLCELL_X1 FILLER_47_235 ();
 FILLCELL_X32 FILLER_47_240 ();
 FILLCELL_X32 FILLER_47_272 ();
 FILLCELL_X32 FILLER_47_304 ();
 FILLCELL_X16 FILLER_47_336 ();
 FILLCELL_X4 FILLER_47_352 ();
endmodule
