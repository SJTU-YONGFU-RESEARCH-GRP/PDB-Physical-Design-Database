module dma_controller (clk,
    debug_has_active_channels,
    rst_n,
    channel_busy,
    channel_done,
    channel_dst_addr,
    channel_enable,
    channel_error,
    channel_length,
    channel_mode,
    channel_src_addr,
    channel_start,
    debug_active_channels,
    debug_channel_state,
    debug_transfer_count,
    dst_addr,
    dst_wdata,
    dst_wready,
    dst_write,
    dst_wstrb,
    src_addr,
    src_rdata,
    src_read,
    src_rready,
    src_rvalid);
 input clk;
 output debug_has_active_channels;
 input rst_n;
 output [3:0] channel_busy;
 output [3:0] channel_done;
 input [127:0] channel_dst_addr;
 input [3:0] channel_enable;
 output [3:0] channel_error;
 input [127:0] channel_length;
 input [7:0] channel_mode;
 input [127:0] channel_src_addr;
 input [3:0] channel_start;
 output [3:0] debug_active_channels;
 output [11:0] debug_channel_state;
 output [127:0] debug_transfer_count;
 output [127:0] dst_addr;
 output [127:0] dst_wdata;
 input [3:0] dst_wready;
 output [3:0] dst_write;
 output [15:0] dst_wstrb;
 output [127:0] src_addr;
 input [127:0] src_rdata;
 output [3:0] src_read;
 output [3:0] src_rready;
 input [3:0] src_rvalid;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire clknet_0_clk;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire \active_channel_count[0] ;
 wire \active_channel_count[1] ;
 wire \active_channel_count[2] ;
 wire \active_channel_count[3] ;
 wire \channel_state[0][0] ;
 wire \channel_state[0][1] ;
 wire \channel_state[0][2] ;
 wire \channel_state[1][0] ;
 wire \channel_state[1][1] ;
 wire \channel_state[1][2] ;
 wire \channel_state[2][0] ;
 wire \channel_state[2][1] ;
 wire \channel_state[2][2] ;
 wire \channel_state[3][0] ;
 wire \channel_state[3][1] ;
 wire \channel_state[3][2] ;
 wire \transfer_count[0][0] ;
 wire \transfer_count[0][10] ;
 wire \transfer_count[0][11] ;
 wire \transfer_count[0][12] ;
 wire \transfer_count[0][13] ;
 wire \transfer_count[0][14] ;
 wire \transfer_count[0][15] ;
 wire \transfer_count[0][16] ;
 wire \transfer_count[0][17] ;
 wire \transfer_count[0][18] ;
 wire \transfer_count[0][19] ;
 wire \transfer_count[0][1] ;
 wire \transfer_count[0][20] ;
 wire \transfer_count[0][21] ;
 wire \transfer_count[0][22] ;
 wire \transfer_count[0][23] ;
 wire \transfer_count[0][24] ;
 wire \transfer_count[0][25] ;
 wire \transfer_count[0][26] ;
 wire \transfer_count[0][27] ;
 wire \transfer_count[0][28] ;
 wire \transfer_count[0][29] ;
 wire \transfer_count[0][2] ;
 wire \transfer_count[0][30] ;
 wire \transfer_count[0][31] ;
 wire \transfer_count[0][3] ;
 wire \transfer_count[0][4] ;
 wire \transfer_count[0][5] ;
 wire \transfer_count[0][6] ;
 wire \transfer_count[0][7] ;
 wire \transfer_count[0][8] ;
 wire \transfer_count[0][9] ;
 wire \transfer_count[1][0] ;
 wire \transfer_count[1][10] ;
 wire \transfer_count[1][11] ;
 wire \transfer_count[1][12] ;
 wire \transfer_count[1][13] ;
 wire \transfer_count[1][14] ;
 wire \transfer_count[1][15] ;
 wire \transfer_count[1][16] ;
 wire \transfer_count[1][17] ;
 wire \transfer_count[1][18] ;
 wire \transfer_count[1][19] ;
 wire \transfer_count[1][1] ;
 wire \transfer_count[1][20] ;
 wire \transfer_count[1][21] ;
 wire \transfer_count[1][22] ;
 wire \transfer_count[1][23] ;
 wire \transfer_count[1][24] ;
 wire \transfer_count[1][25] ;
 wire \transfer_count[1][26] ;
 wire \transfer_count[1][27] ;
 wire \transfer_count[1][28] ;
 wire \transfer_count[1][29] ;
 wire \transfer_count[1][2] ;
 wire \transfer_count[1][30] ;
 wire \transfer_count[1][31] ;
 wire \transfer_count[1][3] ;
 wire \transfer_count[1][4] ;
 wire \transfer_count[1][5] ;
 wire \transfer_count[1][6] ;
 wire \transfer_count[1][7] ;
 wire \transfer_count[1][8] ;
 wire \transfer_count[1][9] ;
 wire \transfer_count[2][0] ;
 wire \transfer_count[2][10] ;
 wire \transfer_count[2][11] ;
 wire \transfer_count[2][12] ;
 wire \transfer_count[2][13] ;
 wire \transfer_count[2][14] ;
 wire \transfer_count[2][15] ;
 wire \transfer_count[2][16] ;
 wire \transfer_count[2][17] ;
 wire \transfer_count[2][18] ;
 wire \transfer_count[2][19] ;
 wire \transfer_count[2][1] ;
 wire \transfer_count[2][20] ;
 wire \transfer_count[2][21] ;
 wire \transfer_count[2][22] ;
 wire \transfer_count[2][23] ;
 wire \transfer_count[2][24] ;
 wire \transfer_count[2][25] ;
 wire \transfer_count[2][26] ;
 wire \transfer_count[2][27] ;
 wire \transfer_count[2][28] ;
 wire \transfer_count[2][29] ;
 wire \transfer_count[2][2] ;
 wire \transfer_count[2][30] ;
 wire \transfer_count[2][31] ;
 wire \transfer_count[2][3] ;
 wire \transfer_count[2][4] ;
 wire \transfer_count[2][5] ;
 wire \transfer_count[2][6] ;
 wire \transfer_count[2][7] ;
 wire \transfer_count[2][8] ;
 wire \transfer_count[2][9] ;
 wire \transfer_count[3][0] ;
 wire \transfer_count[3][10] ;
 wire \transfer_count[3][11] ;
 wire \transfer_count[3][12] ;
 wire \transfer_count[3][13] ;
 wire \transfer_count[3][14] ;
 wire \transfer_count[3][15] ;
 wire \transfer_count[3][16] ;
 wire \transfer_count[3][17] ;
 wire \transfer_count[3][18] ;
 wire \transfer_count[3][19] ;
 wire \transfer_count[3][1] ;
 wire \transfer_count[3][20] ;
 wire \transfer_count[3][21] ;
 wire \transfer_count[3][22] ;
 wire \transfer_count[3][23] ;
 wire \transfer_count[3][24] ;
 wire \transfer_count[3][25] ;
 wire \transfer_count[3][26] ;
 wire \transfer_count[3][27] ;
 wire \transfer_count[3][28] ;
 wire \transfer_count[3][29] ;
 wire \transfer_count[3][2] ;
 wire \transfer_count[3][30] ;
 wire \transfer_count[3][31] ;
 wire \transfer_count[3][3] ;
 wire \transfer_count[3][4] ;
 wire \transfer_count[3][5] ;
 wire \transfer_count[3][6] ;
 wire \transfer_count[3][7] ;
 wire \transfer_count[3][8] ;
 wire \transfer_count[3][9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net715;
 wire net716;
 wire net717;

 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1392_ (.A1(\transfer_count[1][0] ),
    .A2(\transfer_count[1][1] ),
    .A3(\transfer_count[1][4] ),
    .A4(\transfer_count[1][5] ),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1393_ (.A1(\transfer_count[1][2] ),
    .A2(\transfer_count[1][3] ),
    .A3(_0747_),
    .Z(_0748_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _1394_ (.A1(\transfer_count[1][7] ),
    .A2(\transfer_count[1][6] ),
    .A3(_0748_),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1395_ (.A1(\transfer_count[1][10] ),
    .A2(\transfer_count[1][9] ),
    .A3(\transfer_count[1][8] ),
    .Z(_0750_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _1396_ (.A1(\transfer_count[1][12] ),
    .A2(\transfer_count[1][11] ),
    .A3(_0749_),
    .A4(_0750_),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1397_ (.A1(\transfer_count[1][13] ),
    .A2(_0751_),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1398_ (.A1(\transfer_count[1][8] ),
    .A2(_0749_),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1399_ (.A1(\transfer_count[1][9] ),
    .A2(_0752_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1400_ (.A1(\transfer_count[1][28] ),
    .A2(\transfer_count[1][27] ),
    .A3(\transfer_count[1][26] ),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1401_ (.A1(\transfer_count[1][13] ),
    .A2(\transfer_count[1][12] ),
    .A3(\transfer_count[1][11] ),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1402_ (.A1(\transfer_count[1][14] ),
    .A2(\transfer_count[1][15] ),
    .Z(_0755_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1403_ (.A1(\transfer_count[1][16] ),
    .A2(_0750_),
    .A3(_0754_),
    .A4(_0755_),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1404_ (.A1(\transfer_count[1][19] ),
    .A2(\transfer_count[1][18] ),
    .A3(\transfer_count[1][17] ),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1405_ (.A1(\transfer_count[1][20] ),
    .A2(_0757_),
    .Z(_0758_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1406_ (.A1(\transfer_count[1][22] ),
    .A2(\transfer_count[1][21] ),
    .A3(_0756_),
    .A4(_0758_),
    .Z(_0759_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1407_ (.A1(\transfer_count[1][25] ),
    .A2(\transfer_count[1][24] ),
    .A3(\transfer_count[1][23] ),
    .Z(_0760_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1408_ (.A1(_0749_),
    .A2(_0753_),
    .A3(_0759_),
    .A4(_0760_),
    .Z(_0761_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1409_ (.A1(\transfer_count[1][29] ),
    .A2(_0761_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1410_ (.A1(_0749_),
    .A2(_0759_),
    .Z(_0762_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1411_ (.A1(\transfer_count[1][24] ),
    .A2(\transfer_count[1][23] ),
    .A3(_0762_),
    .Z(_0763_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1412_ (.A1(\transfer_count[1][25] ),
    .A2(_0763_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1413_ (.A1(_0749_),
    .A2(_0756_),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1414_ (.A1(_0758_),
    .A2(_0764_),
    .Z(_0765_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1415_ (.A1(\transfer_count[1][21] ),
    .A2(_0765_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1416_ (.A1(\transfer_count[1][17] ),
    .A2(_0764_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _1417_ (.A1(\channel_state[1][0] ),
    .A2(\channel_state[1][1] ),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1418_ (.A1(net139),
    .A2(\channel_state[1][2] ),
    .Z(_0767_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1419_ (.A1(_0766_),
    .A2(_0767_),
    .Z(_0768_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1420_ (.I(_0768_),
    .Z(_0769_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1421_ (.A1(_1002_),
    .A2(_0993_),
    .A3(_0999_),
    .A4(_1005_),
    .Z(_0770_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1422_ (.A1(_0984_),
    .A2(_0990_),
    .A3(_0987_),
    .Z(_0771_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1423_ (.A1(_0996_),
    .A2(_0770_),
    .A3(_0771_),
    .Z(_0772_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1424_ (.A1(_1374_),
    .A2(_1380_),
    .A3(_1377_),
    .A4(_1383_),
    .Z(_0773_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1425_ (.A1(_0772_),
    .A2(_0773_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1426_ (.I(_1365_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1427_ (.I(_1364_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1428_ (.A1(_0775_),
    .A2(_1359_),
    .B(_0776_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1429_ (.A1(_1368_),
    .A2(_1371_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1430_ (.A1(_1368_),
    .A2(_1370_),
    .B1(_0777_),
    .B2(_0778_),
    .C(_1367_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1431_ (.A1(_1374_),
    .A2(_1377_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1432_ (.A1(_1380_),
    .A2(_1382_),
    .B(_1379_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1433_ (.A1(_1374_),
    .A2(_1376_),
    .B(_1373_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1434_ (.A1(_0780_),
    .A2(_0781_),
    .B(_0782_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1435_ (.A1(_0772_),
    .A2(_0783_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1436_ (.A1(_0774_),
    .A2(_0779_),
    .B(_0784_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _1437_ (.A1(_1002_),
    .A2(_1004_),
    .B(_1001_),
    .C(_0998_),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1438_ (.A1(_0999_),
    .A2(_0998_),
    .B(_0996_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1439_ (.A1(_0992_),
    .A2(_0995_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1440_ (.A1(_0786_),
    .A2(_0787_),
    .B(_0788_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _1441_ (.A1(_0993_),
    .A2(_0992_),
    .B(_0771_),
    .C(_0789_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1442_ (.A1(_0987_),
    .A2(_0989_),
    .Z(_0791_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1443_ (.A1(_0986_),
    .A2(_0791_),
    .Z(_0792_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1444_ (.A1(_0984_),
    .A2(_0792_),
    .B(_0983_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1445_ (.A1(_0790_),
    .A2(_0793_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1446_ (.A1(_1035_),
    .A2(_1037_),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1447_ (.A1(_1034_),
    .A2(_0795_),
    .Z(_0796_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _1448_ (.A1(_1050_),
    .A2(_1052_),
    .B(_1049_),
    .C(_1046_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1449_ (.A1(_1047_),
    .A2(_1046_),
    .B(_1044_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1450_ (.A1(_1040_),
    .A2(_1043_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1451_ (.A1(_0797_),
    .A2(_0798_),
    .B(_0799_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1452_ (.A1(_1041_),
    .A2(_1040_),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1453_ (.A1(_1032_),
    .A2(_1038_),
    .A3(_1035_),
    .A4(_0801_),
    .Z(_0802_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1454_ (.A1(_1032_),
    .A2(_0796_),
    .B1(_0800_),
    .B2(_0802_),
    .C(_1031_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1455_ (.A1(_1008_),
    .A2(_1014_),
    .A3(_1011_),
    .A4(_1017_),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1456_ (.A1(_1026_),
    .A2(_1028_),
    .B(_1025_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1457_ (.A1(_1020_),
    .A2(_1023_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1458_ (.A1(_1020_),
    .A2(_1022_),
    .B(_1019_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1459_ (.A1(_0805_),
    .A2(_0806_),
    .B(_0807_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1460_ (.A1(_1008_),
    .A2(_1011_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1461_ (.A1(_1014_),
    .A2(_1016_),
    .B(_1013_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1462_ (.A1(_1008_),
    .A2(_1010_),
    .B(_1007_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1463_ (.A1(_0809_),
    .A2(_0810_),
    .B(_0811_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1464_ (.A1(_0804_),
    .A2(_0808_),
    .B(_0812_),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1465_ (.A1(_0803_),
    .A2(_0813_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _1466_ (.A1(_1032_),
    .A2(_1038_),
    .A3(_1050_),
    .A4(_1035_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _1467_ (.A1(_1044_),
    .A2(_1041_),
    .A3(_1047_),
    .A4(_1053_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _1468_ (.A1(_0809_),
    .A2(_0810_),
    .B1(_0815_),
    .B2(_0816_),
    .C(_0811_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1469_ (.A1(_0804_),
    .A2(_0808_),
    .B(_0817_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1470_ (.A1(_1020_),
    .A2(_1026_),
    .A3(_1023_),
    .A4(_1029_),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1471_ (.A1(_0804_),
    .A2(_0819_),
    .Z(_0820_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _1472_ (.A1(_0804_),
    .A2(_0808_),
    .B(_0812_),
    .C(_0820_),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _1473_ (.A1(_1368_),
    .A2(_1365_),
    .A3(_1360_),
    .A4(_1371_),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _1474_ (.A1(_0815_),
    .A2(_0816_),
    .A3(_0822_),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1475_ (.A1(_0820_),
    .A2(_0772_),
    .A3(_0773_),
    .A4(_0823_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _1476_ (.A1(_0803_),
    .A2(_0818_),
    .B(_0821_),
    .C(_0824_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _1477_ (.A1(_0785_),
    .A2(_0794_),
    .A3(_0814_),
    .B(_0825_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _1478_ (.I(\channel_state[1][2] ),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1479_ (.A1(net3),
    .A2(_0827_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1480_ (.A1(net135),
    .A2(_0828_),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1481_ (.A1(_0766_),
    .A2(_0829_),
    .B(net147),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1482_ (.A1(_0769_),
    .A2(_0826_),
    .B(_0830_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1483_ (.A1(\transfer_count[3][27] ),
    .A2(\transfer_count[3][26] ),
    .A3(\transfer_count[3][25] ),
    .A4(\transfer_count[3][24] ),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1484_ (.A1(\transfer_count[3][28] ),
    .A2(_0831_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1485_ (.A1(\transfer_count[3][19] ),
    .A2(\transfer_count[3][18] ),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1486_ (.A1(\transfer_count[3][22] ),
    .A2(\transfer_count[3][21] ),
    .A3(\transfer_count[3][20] ),
    .A4(_0833_),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1487_ (.A1(\transfer_count[3][17] ),
    .A2(\transfer_count[3][16] ),
    .A3(\transfer_count[3][15] ),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1488_ (.A1(\transfer_count[3][14] ),
    .A2(\transfer_count[3][13] ),
    .A3(\transfer_count[3][12] ),
    .A4(\transfer_count[3][11] ),
    .Z(_0836_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1489_ (.A1(_0835_),
    .A2(_0836_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1490_ (.A1(\transfer_count[3][10] ),
    .A2(\transfer_count[3][9] ),
    .A3(\transfer_count[3][8] ),
    .A4(\transfer_count[3][7] ),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1491_ (.A1(\transfer_count[3][5] ),
    .A2(\transfer_count[3][4] ),
    .A3(\transfer_count[3][3] ),
    .A4(\transfer_count[3][2] ),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1492_ (.A1(\transfer_count[3][1] ),
    .A2(\transfer_count[3][0] ),
    .Z(_0840_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1493_ (.A1(\transfer_count[3][6] ),
    .A2(_0838_),
    .A3(_0839_),
    .A4(_0840_),
    .Z(_0841_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1494_ (.A1(\transfer_count[3][23] ),
    .A2(_0834_),
    .A3(_0837_),
    .A4(_0841_),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1495_ (.A1(_0832_),
    .A2(_0842_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1496_ (.A1(\transfer_count[3][29] ),
    .A2(_0843_),
    .Z(_1060_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _1497_ (.A1(\transfer_count[3][26] ),
    .A2(\transfer_count[3][25] ),
    .A3(\transfer_count[3][24] ),
    .A4(_0842_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1498_ (.A1(\transfer_count[3][27] ),
    .A2(_0844_),
    .Z(_1066_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1499_ (.A1(\transfer_count[3][24] ),
    .A2(_0842_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1500_ (.A1(\transfer_count[3][25] ),
    .A2(_0845_),
    .Z(_1072_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1501_ (.A1(_0837_),
    .A2(_0841_),
    .Z(_0846_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1502_ (.A1(_0834_),
    .A2(_0846_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1503_ (.A1(\transfer_count[3][23] ),
    .A2(_0847_),
    .Z(_1078_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1504_ (.A1(_0836_),
    .A2(_0841_),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _1505_ (.A1(\transfer_count[3][20] ),
    .A2(_0833_),
    .A3(_0835_),
    .A4(_0848_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1506_ (.A1(\transfer_count[3][21] ),
    .A2(_0849_),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1507_ (.A1(\transfer_count[3][18] ),
    .A2(_0846_),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1508_ (.A1(\transfer_count[3][19] ),
    .A2(_0850_),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1509_ (.A1(\transfer_count[3][15] ),
    .A2(_0848_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1510_ (.A1(\transfer_count[3][12] ),
    .A2(\transfer_count[3][11] ),
    .A3(_0841_),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1511_ (.A1(\transfer_count[3][13] ),
    .A2(_0851_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1512_ (.A1(\transfer_count[3][11] ),
    .A2(_0841_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1513_ (.A1(\transfer_count[3][6] ),
    .A2(_0839_),
    .A3(_0840_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1514_ (.A1(\transfer_count[3][8] ),
    .A2(\transfer_count[3][7] ),
    .A3(_0852_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1515_ (.A1(\transfer_count[3][9] ),
    .A2(_0853_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1516_ (.A1(\transfer_count[3][7] ),
    .A2(_0852_),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1517_ (.A1(\transfer_count[3][4] ),
    .A2(\transfer_count[3][3] ),
    .A3(\transfer_count[3][2] ),
    .A4(_0840_),
    .Z(_0854_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1518_ (.A1(\transfer_count[3][5] ),
    .A2(_0854_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1519_ (.A1(\transfer_count[3][2] ),
    .A2(_0840_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1520_ (.A1(\transfer_count[3][3] ),
    .A2(_0855_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1521_ (.A1(_1116_),
    .A2(_1113_),
    .Z(_0856_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1522_ (.A1(_1107_),
    .A2(_1119_),
    .A3(_1125_),
    .A4(_1110_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1523_ (.A1(_1104_),
    .A2(_1122_),
    .A3(_0856_),
    .A4(_0857_),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _1524_ (.A1(_1128_),
    .A2(_1131_),
    .A3(_1137_),
    .A4(_1134_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1525_ (.I(_1148_),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1526_ (.I(_1147_),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1527_ (.A1(_0860_),
    .A2(_1151_),
    .B(_0861_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1528_ (.A1(_1140_),
    .A2(_1143_),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _1529_ (.A1(_1140_),
    .A2(_1142_),
    .B1(_0862_),
    .B2(_0863_),
    .C(_1139_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1530_ (.A1(_1136_),
    .A2(_1131_),
    .A3(_1134_),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1531_ (.A1(_1131_),
    .A2(_1133_),
    .Z(_0866_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _1532_ (.A1(_1130_),
    .A2(_0865_),
    .A3(_0866_),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1533_ (.A1(_1128_),
    .A2(_0867_),
    .B(_1127_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1534_ (.A1(_0859_),
    .A2(_0864_),
    .B(_0868_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1535_ (.A1(_1124_),
    .A2(_1119_),
    .A3(_1122_),
    .Z(_0870_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1536_ (.A1(_1119_),
    .A2(_1121_),
    .Z(_0871_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _1537_ (.A1(_1118_),
    .A2(_0870_),
    .A3(_0871_),
    .B(_0856_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1538_ (.A1(_1112_),
    .A2(_1109_),
    .Z(_0873_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1539_ (.A1(_1104_),
    .A2(_1106_),
    .B1(_1115_),
    .B2(_1113_),
    .C(_0873_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1540_ (.I(_1104_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1541_ (.A1(_1110_),
    .A2(_1109_),
    .Z(_0876_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1542_ (.A1(_1107_),
    .A2(_0876_),
    .B(_1106_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _1543_ (.A1(_0872_),
    .A2(_0874_),
    .B(_0875_),
    .C(_0877_),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _1544_ (.A1(_0858_),
    .A2(_0869_),
    .B(_0878_),
    .C(_1103_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _1545_ (.A1(_1140_),
    .A2(_1148_),
    .A3(_1152_),
    .A4(_1143_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1546_ (.A1(_0859_),
    .A2(_0880_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1547_ (.A1(_0858_),
    .A2(_0881_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1548_ (.A1(_1056_),
    .A2(_1059_),
    .A3(_1065_),
    .A4(_1062_),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1549_ (.A1(_1068_),
    .A2(_1071_),
    .A3(_1077_),
    .A4(_1074_),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1550_ (.A1(_1080_),
    .A2(_1083_),
    .A3(_0883_),
    .A4(_0884_),
    .Z(_0885_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1551_ (.A1(_1095_),
    .A2(_1098_),
    .A3(_1101_),
    .A4(_1086_),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _1552_ (.A1(_1092_),
    .A2(_1089_),
    .A3(_0885_),
    .A4(_0886_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1553_ (.A1(_0882_),
    .A2(_0887_),
    .Z(_0888_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1554_ (.I(_0882_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1555_ (.I(_0883_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1556_ (.A1(_1080_),
    .A2(_1082_),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1557_ (.A1(_1079_),
    .A2(_0891_),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1558_ (.A1(_1076_),
    .A2(_1071_),
    .A3(_1074_),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1559_ (.A1(_1071_),
    .A2(_1073_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _1560_ (.A1(_1070_),
    .A2(_0893_),
    .A3(_0894_),
    .Z(_0895_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1561_ (.A1(_0884_),
    .A2(_0892_),
    .B1(_0895_),
    .B2(_1068_),
    .C(_1067_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1562_ (.A1(_1100_),
    .A2(_1098_),
    .B(_1097_),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1563_ (.A1(_1092_),
    .A2(_1095_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1564_ (.A1(_0897_),
    .A2(_0898_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1565_ (.A1(_1092_),
    .A2(_1094_),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _1566_ (.A1(_1088_),
    .A2(_1085_),
    .A3(_1091_),
    .A4(_0900_),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1567_ (.A1(_1080_),
    .A2(_1083_),
    .A3(_0883_),
    .A4(_0884_),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1568_ (.I(_1085_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1569_ (.A1(_1088_),
    .A2(_1089_),
    .B(_1086_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1570_ (.A1(_0903_),
    .A2(_0904_),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _1571_ (.A1(_0899_),
    .A2(_0901_),
    .B(_0902_),
    .C(_0905_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1572_ (.A1(_1064_),
    .A2(_1062_),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _1573_ (.A1(_1061_),
    .A2(_0907_),
    .B(_1056_),
    .C(_1059_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1574_ (.A1(_1056_),
    .A2(_1058_),
    .B(_1055_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1575_ (.A1(_0908_),
    .A2(_0909_),
    .Z(_0910_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _1576_ (.A1(_0890_),
    .A2(_0896_),
    .B(_0906_),
    .C(_0910_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1577_ (.A1(_0889_),
    .A2(_0887_),
    .B(_0911_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1578_ (.A1(\channel_state[3][0] ),
    .A2(\channel_state[3][1] ),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1579_ (.A1(\channel_state[3][2] ),
    .A2(_0913_),
    .Z(_0914_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _1580_ (.A1(net141),
    .A2(_0914_),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1581_ (.I(_0915_),
    .Z(_0916_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _1582_ (.A1(_0879_),
    .A2(_0888_),
    .B(_0912_),
    .C(_0916_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _1583_ (.I(\channel_state[3][2] ),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1584_ (.A1(net5),
    .A2(_0918_),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1585_ (.A1(net137),
    .A2(_0913_),
    .A3(_0919_),
    .Z(_0920_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1586_ (.A1(net149),
    .A2(_0920_),
    .Z(_0921_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1587_ (.A1(_0917_),
    .A2(_0921_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1588_ (.I(\channel_state[0][2] ),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1589_ (.A1(net134),
    .A2(_0922_),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _1590_ (.A1(net134),
    .A2(net2),
    .A3(_0922_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1591_ (.I(\channel_state[0][1] ),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1592_ (.I0(_0923_),
    .I1(_0924_),
    .S(_0925_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1593_ (.A1(\channel_state[0][0] ),
    .A2(_0926_),
    .Z(_0927_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1594_ (.A1(net154),
    .A2(_0927_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1595_ (.A1(\transfer_count[0][2] ),
    .A2(\transfer_count[0][1] ),
    .A3(\transfer_count[0][0] ),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1596_ (.A1(\transfer_count[0][3] ),
    .A2(\transfer_count[0][4] ),
    .A3(_0928_),
    .Z(_0929_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1597_ (.A1(\transfer_count[0][5] ),
    .A2(_0929_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1598_ (.A1(\transfer_count[0][12] ),
    .A2(\transfer_count[0][11] ),
    .Z(_0930_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1599_ (.A1(\transfer_count[0][10] ),
    .A2(\transfer_count[0][9] ),
    .A3(\transfer_count[0][8] ),
    .Z(_0931_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1600_ (.A1(\transfer_count[0][3] ),
    .A2(\transfer_count[0][5] ),
    .A3(\transfer_count[0][4] ),
    .Z(_0932_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1601_ (.A1(\transfer_count[0][6] ),
    .A2(\transfer_count[0][7] ),
    .A3(_0928_),
    .A4(_0932_),
    .Z(_0933_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _1602_ (.A1(_0930_),
    .A2(_0931_),
    .A3(_0933_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1603_ (.A1(\transfer_count[0][13] ),
    .A2(_0934_),
    .Z(_1186_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1604_ (.A1(\transfer_count[0][6] ),
    .A2(_0928_),
    .A3(_0932_),
    .Z(_0935_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1605_ (.A1(\transfer_count[0][7] ),
    .A2(_0935_),
    .Z(_0936_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1606_ (.A1(\transfer_count[0][8] ),
    .A2(_0936_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1607_ (.A1(\transfer_count[0][9] ),
    .A2(_0937_),
    .Z(_1198_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1608_ (.A1(\transfer_count[0][25] ),
    .A2(\transfer_count[0][24] ),
    .A3(\transfer_count[0][23] ),
    .A4(\transfer_count[0][22] ),
    .Z(_0938_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1609_ (.A1(\transfer_count[0][28] ),
    .A2(\transfer_count[0][27] ),
    .A3(\transfer_count[0][26] ),
    .A4(_0938_),
    .Z(_0939_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1610_ (.A1(\transfer_count[0][19] ),
    .A2(\transfer_count[0][18] ),
    .A3(\transfer_count[0][17] ),
    .A4(\transfer_count[0][16] ),
    .Z(_0940_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1611_ (.A1(\transfer_count[0][21] ),
    .A2(\transfer_count[0][20] ),
    .A3(_0940_),
    .Z(_0941_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1612_ (.A1(\transfer_count[0][14] ),
    .A2(\transfer_count[0][13] ),
    .A3(_0930_),
    .A4(_0931_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1613_ (.A1(\transfer_count[0][15] ),
    .A2(_0933_),
    .A3(_0942_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1614_ (.A1(_0939_),
    .A2(_0941_),
    .A3(_0943_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1615_ (.A1(\transfer_count[0][29] ),
    .A2(_0944_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1616_ (.A1(\transfer_count[0][15] ),
    .A2(_0933_),
    .A3(_0941_),
    .A4(_0942_),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1617_ (.A1(\transfer_count[0][24] ),
    .A2(\transfer_count[0][23] ),
    .A3(\transfer_count[0][22] ),
    .A4(_0945_),
    .Z(_0946_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1618_ (.A1(\transfer_count[0][25] ),
    .A2(_0946_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1619_ (.A1(\transfer_count[0][20] ),
    .A2(_0940_),
    .A3(_0943_),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1620_ (.A1(\transfer_count[0][21] ),
    .A2(_0947_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1621_ (.A1(\transfer_count[0][16] ),
    .A2(_0943_),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1622_ (.A1(\transfer_count[0][17] ),
    .A2(_0948_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1623_ (.I(\channel_state[0][0] ),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1624_ (.A1(_0949_),
    .A2(_0925_),
    .Z(_0950_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _1625_ (.A1(net138),
    .A2(\channel_state[0][2] ),
    .A3(_0950_),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1626_ (.I(_0951_),
    .Z(_0952_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1627_ (.A1(_1164_),
    .A2(_1167_),
    .A3(_1179_),
    .Z(_0953_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1628_ (.I(_1161_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1629_ (.I(_1160_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1630_ (.A1(_0954_),
    .A2(_1155_),
    .B(_0955_),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1631_ (.I(_1179_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1632_ (.A1(_1164_),
    .A2(_1166_),
    .B(_1163_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1633_ (.A1(_0957_),
    .A2(_0958_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1634_ (.I(_1170_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1635_ (.A1(_1173_),
    .A2(_1175_),
    .B(_1172_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1636_ (.A1(_1169_),
    .A2(_1178_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1637_ (.A1(_0960_),
    .A2(_0961_),
    .B(_0962_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _1638_ (.A1(_0953_),
    .A2(_0956_),
    .B(_0959_),
    .C(_0963_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1639_ (.I(_1172_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1640_ (.A1(_1176_),
    .A2(_1175_),
    .B(_1173_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1641_ (.A1(_0965_),
    .A2(_0146_),
    .B(_0960_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1642_ (.A1(_1182_),
    .A2(_1188_),
    .A3(_1185_),
    .Z(_0148_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1643_ (.A1(_1194_),
    .A2(_1200_),
    .A3(_1191_),
    .A4(_1197_),
    .Z(_0149_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1644_ (.A1(_1203_),
    .A2(_0148_),
    .A3(_0149_),
    .Z(_0150_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1645_ (.A1(_1169_),
    .A2(_0147_),
    .B(_0150_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1646_ (.A1(_1185_),
    .A2(_1187_),
    .Z(_0152_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1647_ (.A1(_1184_),
    .A2(_0152_),
    .Z(_0153_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1648_ (.A1(_1182_),
    .A2(_0153_),
    .B(_1181_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _1649_ (.A1(_0964_),
    .A2(_0151_),
    .B(_0154_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _1650_ (.A1(_1230_),
    .A2(_1233_),
    .A3(_1235_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1651_ (.A1(_1230_),
    .A2(_1232_),
    .B(_1229_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _1652_ (.A1(_1206_),
    .A2(_1212_),
    .A3(_1209_),
    .A4(_1215_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _1653_ (.A1(_1218_),
    .A2(_1224_),
    .A3(_1221_),
    .A4(_1227_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _1654_ (.A1(_0156_),
    .A2(_0157_),
    .B(_0158_),
    .C(_0159_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _1655_ (.A1(_1212_),
    .A2(_1214_),
    .B(_1211_),
    .C(_1208_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1656_ (.A1(_1209_),
    .A2(_1208_),
    .B(_1206_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1657_ (.I(_1205_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1658_ (.A1(_0161_),
    .A2(_0162_),
    .B(_0163_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1659_ (.A1(_0160_),
    .A2(_0164_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _1660_ (.A1(_1200_),
    .A2(_1202_),
    .B(_1199_),
    .C(_1196_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1661_ (.A1(_1197_),
    .A2(_1196_),
    .B(_1194_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1662_ (.A1(_1190_),
    .A2(_1193_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1663_ (.A1(_0166_),
    .A2(_0167_),
    .B(_0168_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _1664_ (.A1(_1191_),
    .A2(_1190_),
    .B(_0148_),
    .C(_0169_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _1665_ (.A1(_1230_),
    .A2(_1236_),
    .A3(_1233_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _1666_ (.A1(_0158_),
    .A2(_0159_),
    .A3(_0171_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _1667_ (.A1(_1242_),
    .A2(_1239_),
    .A3(_1245_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1668_ (.A1(_1248_),
    .A2(_1250_),
    .B(_1247_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1669_ (.A1(_1239_),
    .A2(_1241_),
    .B(_1238_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _1670_ (.A1(_1242_),
    .A2(_1239_),
    .A3(_1244_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _1671_ (.A1(_0173_),
    .A2(_0174_),
    .B(_0175_),
    .C(_0176_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1672_ (.A1(_1224_),
    .A2(_1226_),
    .B(_1223_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1673_ (.A1(_1218_),
    .A2(_1221_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1674_ (.A1(_1218_),
    .A2(_1220_),
    .B(_1217_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1675_ (.A1(_0178_),
    .A2(_0179_),
    .B(_0180_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1676_ (.A1(_1206_),
    .A2(_1212_),
    .A3(_1209_),
    .A4(_1215_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _1677_ (.A1(_0172_),
    .A2(_0177_),
    .B1(_0181_),
    .B2(_0182_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _1678_ (.A1(_0165_),
    .A2(_0170_),
    .A3(_0183_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1679_ (.A1(_1248_),
    .A2(_1251_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1680_ (.A1(_0173_),
    .A2(_0185_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _1681_ (.A1(_0172_),
    .A2(_0186_),
    .B(_0160_),
    .C(_0164_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1682_ (.A1(_1156_),
    .A2(_1170_),
    .A3(_1176_),
    .A4(_1173_),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1683_ (.A1(_1161_),
    .A2(_0953_),
    .A3(_0188_),
    .Z(_0189_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1684_ (.A1(_0172_),
    .A2(_0186_),
    .A3(_0189_),
    .A4(_0150_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1685_ (.A1(_0183_),
    .A2(_0187_),
    .B(_0190_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1686_ (.A1(_0155_),
    .A2(_0184_),
    .B(_0191_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _1687_ (.A1(\channel_state[0][0] ),
    .A2(\channel_state[0][1] ),
    .A3(_0924_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1688_ (.I(net146),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _1689_ (.A1(_0952_),
    .A2(_0192_),
    .B1(_0193_),
    .B2(_0194_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1690_ (.I(\transfer_count[3][0] ),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _1691_ (.A1(_0915_),
    .A2(_0920_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1692_ (.I0(_0916_),
    .I1(_0195_),
    .S(\transfer_count[3][0] ),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1693_ (.I(_0195_),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _1694_ (.A1(_1145_),
    .A2(_0916_),
    .B1(_0196_),
    .B2(\transfer_count[3][1] ),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1695_ (.I(_0197_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1696_ (.A1(_1144_),
    .A2(_0916_),
    .Z(_0198_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _1697_ (.A1(net141),
    .A2(_0914_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1698_ (.I(_0199_),
    .Z(_0200_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1699_ (.A1(_0915_),
    .A2(_0920_),
    .Z(_0201_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1700_ (.I(_0201_),
    .Z(_0202_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1701_ (.A1(_1144_),
    .A2(_0200_),
    .B(_0202_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1702_ (.I0(_0198_),
    .I1(_0203_),
    .S(\transfer_count[3][2] ),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1703_ (.I(_0199_),
    .Z(_0204_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1704_ (.I(_0204_),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1705_ (.A1(\transfer_count[3][3] ),
    .A2(_0196_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1706_ (.A1(_1138_),
    .A2(_0205_),
    .B(_0206_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1707_ (.A1(\transfer_count[3][3] ),
    .A2(\transfer_count[3][2] ),
    .A3(_1144_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1708_ (.A1(\transfer_count[3][4] ),
    .A2(_0207_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1709_ (.A1(\transfer_count[3][4] ),
    .A2(_0196_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1710_ (.A1(_0205_),
    .A2(_1135_),
    .B(_0208_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1711_ (.A1(\transfer_count[3][5] ),
    .A2(_0196_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1712_ (.A1(_1132_),
    .A2(_0205_),
    .B(_0209_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1713_ (.A1(_1144_),
    .A2(_0839_),
    .Z(_0210_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1714_ (.A1(_0916_),
    .A2(_0210_),
    .Z(_0211_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1715_ (.A1(_0204_),
    .A2(_0210_),
    .B(_0202_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1716_ (.I0(_0211_),
    .I1(_0212_),
    .S(\transfer_count[3][6] ),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1717_ (.I(_0915_),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1718_ (.A1(_0852_),
    .A2(_0213_),
    .Z(_0214_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1719_ (.A1(_0852_),
    .A2(_0200_),
    .B(_0202_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1720_ (.I0(_0214_),
    .I1(_0215_),
    .S(\transfer_count[3][7] ),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1721_ (.A1(\transfer_count[3][6] ),
    .A2(_1144_),
    .Z(_0216_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1722_ (.A1(_0839_),
    .A2(_0216_),
    .Z(_0217_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1723_ (.A1(\transfer_count[3][7] ),
    .A2(_0217_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1724_ (.A1(\transfer_count[3][8] ),
    .A2(_0218_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1725_ (.A1(\transfer_count[3][8] ),
    .A2(_0196_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1726_ (.A1(_0205_),
    .A2(_1123_),
    .B(_0219_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1727_ (.A1(\transfer_count[3][9] ),
    .A2(_0196_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1728_ (.A1(_1120_),
    .A2(_0205_),
    .B(_0220_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1729_ (.A1(\transfer_count[3][9] ),
    .A2(\transfer_count[3][8] ),
    .A3(\transfer_count[3][7] ),
    .A4(_0217_),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1730_ (.A1(\transfer_count[3][10] ),
    .A2(_0221_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1731_ (.A1(\transfer_count[3][10] ),
    .A2(_0196_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1732_ (.A1(_0205_),
    .A2(_1117_),
    .B(_0222_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1733_ (.A1(_0841_),
    .A2(_0213_),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1734_ (.A1(_0841_),
    .A2(_0200_),
    .B(_0202_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1735_ (.I0(_0223_),
    .I1(_0224_),
    .S(\transfer_count[3][11] ),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1736_ (.A1(_0838_),
    .A2(_0839_),
    .A3(_0216_),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1737_ (.A1(\transfer_count[3][11] ),
    .A2(_0225_),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1738_ (.A1(\transfer_count[3][12] ),
    .A2(_0226_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1739_ (.A1(\transfer_count[3][12] ),
    .A2(_0196_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1740_ (.A1(_0205_),
    .A2(_1111_),
    .B(_0227_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1741_ (.A1(_0851_),
    .A2(_0213_),
    .Z(_0228_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1742_ (.A1(_0851_),
    .A2(_0200_),
    .B(_0202_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1743_ (.I0(_0228_),
    .I1(_0229_),
    .S(\transfer_count[3][13] ),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1744_ (.A1(\transfer_count[3][13] ),
    .A2(\transfer_count[3][12] ),
    .A3(\transfer_count[3][11] ),
    .A4(_0225_),
    .Z(_0230_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1745_ (.A1(_0916_),
    .A2(_0230_),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1746_ (.A1(_0204_),
    .A2(_0230_),
    .B(_0201_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1747_ (.I0(_0231_),
    .I1(_0232_),
    .S(\transfer_count[3][14] ),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1748_ (.A1(_0836_),
    .A2(_0838_),
    .A3(_0852_),
    .A4(_0915_),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1749_ (.A1(_0848_),
    .A2(_0200_),
    .B(_0201_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1750_ (.I0(_0233_),
    .I1(_0234_),
    .S(\transfer_count[3][15] ),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _1751_ (.A1(\transfer_count[3][15] ),
    .A2(\transfer_count[3][14] ),
    .A3(_0230_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1752_ (.A1(_0213_),
    .A2(_0235_),
    .Z(_0236_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1753_ (.A1(_0195_),
    .A2(_0236_),
    .B(\transfer_count[3][16] ),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _1754_ (.A1(\transfer_count[3][16] ),
    .A2(_0205_),
    .A3(_0235_),
    .B(_0237_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _1755_ (.A1(\transfer_count[3][16] ),
    .A2(\transfer_count[3][15] ),
    .A3(_0848_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1756_ (.A1(_0213_),
    .A2(_0238_),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1757_ (.A1(_0195_),
    .A2(_0239_),
    .B(\transfer_count[3][17] ),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _1758_ (.A1(\transfer_count[3][17] ),
    .A2(_0205_),
    .A3(_0238_),
    .B(_0240_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1759_ (.A1(_0837_),
    .A2(_0915_),
    .A3(_0225_),
    .Z(_0241_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1760_ (.A1(_0835_),
    .A2(_0836_),
    .A3(_0838_),
    .Z(_0242_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1761_ (.A1(_0242_),
    .A2(_0217_),
    .Z(_0243_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1762_ (.A1(_0200_),
    .A2(_0243_),
    .B(_0201_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1763_ (.I0(_0241_),
    .I1(_0244_),
    .S(\transfer_count[3][18] ),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1764_ (.A1(\transfer_count[3][19] ),
    .A2(_0196_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1765_ (.A1(_1090_),
    .A2(_0205_),
    .B(_0245_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1766_ (.A1(_0833_),
    .A2(_0837_),
    .A3(_0915_),
    .A4(_0225_),
    .Z(_0246_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1767_ (.A1(_0833_),
    .A2(_0243_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1768_ (.A1(_0200_),
    .A2(_0247_),
    .B(_0201_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1769_ (.I0(_0246_),
    .I1(_0248_),
    .S(\transfer_count[3][20] ),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1770_ (.A1(_0849_),
    .A2(_0213_),
    .Z(_0249_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1771_ (.A1(_0195_),
    .A2(_0249_),
    .B(\transfer_count[3][21] ),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _1772_ (.A1(\transfer_count[3][21] ),
    .A2(_0849_),
    .A3(_0204_),
    .B(_0250_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1773_ (.A1(\transfer_count[3][21] ),
    .A2(\transfer_count[3][20] ),
    .A3(_0833_),
    .A4(_0243_),
    .Z(_0251_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1774_ (.A1(_0916_),
    .A2(_0251_),
    .B(\transfer_count[3][22] ),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1775_ (.A1(_0200_),
    .A2(_0251_),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1776_ (.A1(\transfer_count[3][22] ),
    .A2(_0202_),
    .A3(_0253_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1777_ (.A1(_0252_),
    .A2(_0254_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1778_ (.A1(_0847_),
    .A2(_0213_),
    .Z(_0255_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1779_ (.A1(_0195_),
    .A2(_0255_),
    .B(\transfer_count[3][23] ),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _1780_ (.A1(\transfer_count[3][23] ),
    .A2(_0847_),
    .A3(_0204_),
    .B(_0256_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1781_ (.A1(\transfer_count[3][23] ),
    .A2(_0834_),
    .A3(_0242_),
    .A4(_0217_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1782_ (.I(_0257_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1783_ (.A1(_0200_),
    .A2(_0257_),
    .B(_0202_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1784_ (.A1(\transfer_count[3][24] ),
    .A2(_0259_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _1785_ (.A1(\transfer_count[3][24] ),
    .A2(_0204_),
    .A3(_0258_),
    .B(_0260_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1786_ (.A1(_0845_),
    .A2(_0213_),
    .Z(_0261_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1787_ (.A1(_0195_),
    .A2(_0261_),
    .B(\transfer_count[3][25] ),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _1788_ (.A1(\transfer_count[3][25] ),
    .A2(_0845_),
    .A3(_0204_),
    .B(_0262_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1789_ (.A1(\transfer_count[3][25] ),
    .A2(\transfer_count[3][24] ),
    .A3(_0257_),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1790_ (.A1(_0916_),
    .A2(_0263_),
    .B(\transfer_count[3][26] ),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1791_ (.A1(_0200_),
    .A2(_0263_),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1792_ (.A1(\transfer_count[3][26] ),
    .A2(_0202_),
    .A3(_0265_),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1793_ (.A1(_0264_),
    .A2(_0266_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1794_ (.A1(_0844_),
    .A2(_0213_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1795_ (.A1(_0195_),
    .A2(_0267_),
    .B(\transfer_count[3][27] ),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _1796_ (.A1(\transfer_count[3][27] ),
    .A2(_0844_),
    .A3(_0204_),
    .B(_0268_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1797_ (.A1(_0831_),
    .A2(_0257_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1798_ (.A1(_0916_),
    .A2(_0269_),
    .B(\transfer_count[3][28] ),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1799_ (.A1(_0199_),
    .A2(_0269_),
    .Z(_0271_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1800_ (.A1(\transfer_count[3][28] ),
    .A2(_0202_),
    .A3(_0271_),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1801_ (.A1(_0270_),
    .A2(_0272_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1802_ (.A1(_0843_),
    .A2(_0915_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1803_ (.A1(_0195_),
    .A2(_0273_),
    .B(\transfer_count[3][29] ),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _1804_ (.A1(\transfer_count[3][29] ),
    .A2(_0843_),
    .A3(_0204_),
    .B(_0274_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1805_ (.A1(\transfer_count[3][29] ),
    .A2(_0832_),
    .Z(_0275_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1806_ (.A1(_0257_),
    .A2(_0275_),
    .Z(_0276_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1807_ (.A1(_0916_),
    .A2(_0276_),
    .B(\transfer_count[3][30] ),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1808_ (.A1(_0199_),
    .A2(_0276_),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1809_ (.A1(\transfer_count[3][30] ),
    .A2(_0202_),
    .A3(_0278_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1810_ (.A1(_0277_),
    .A2(_0279_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _1811_ (.A1(\transfer_count[3][30] ),
    .A2(_0842_),
    .A3(_0275_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1812_ (.A1(_0213_),
    .A2(_0280_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1813_ (.A1(_0195_),
    .A2(_0281_),
    .B(\transfer_count[3][31] ),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _1814_ (.A1(\transfer_count[3][31] ),
    .A2(_0204_),
    .A3(_0280_),
    .B(_0282_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1815_ (.I(\transfer_count[2][0] ),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1816_ (.I(\channel_state[2][0] ),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1817_ (.A1(\channel_state[2][2] ),
    .A2(_0283_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1818_ (.A1(\channel_state[2][1] ),
    .A2(_0284_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1819_ (.A1(net140),
    .A2(_0285_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1820_ (.I(_0286_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _1821_ (.A1(net140),
    .A2(_0285_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1822_ (.I(net4),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1823_ (.I(net136),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _1824_ (.A1(_0289_),
    .A2(\channel_state[2][2] ),
    .A3(\channel_state[2][0] ),
    .A4(_0290_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1825_ (.A1(\channel_state[2][1] ),
    .A2(_0291_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1826_ (.A1(_0288_),
    .A2(_0292_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1827_ (.I0(_0287_),
    .I1(_0293_),
    .S(\transfer_count[2][0] ),
    .Z(_0077_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _1828_ (.A1(_1349_),
    .A2(_0287_),
    .B1(_0293_),
    .B2(\transfer_count[2][1] ),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1829_ (.I(_0294_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1830_ (.I(_0286_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1831_ (.A1(_1348_),
    .A2(_0295_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1832_ (.I(_0288_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _1833_ (.A1(_0288_),
    .A2(_0292_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1834_ (.I(_0298_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1835_ (.A1(_1348_),
    .A2(_0297_),
    .B(_0299_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1836_ (.I0(_0296_),
    .I1(_0300_),
    .S(\transfer_count[2][2] ),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1837_ (.A1(\transfer_count[2][0] ),
    .A2(\transfer_count[2][1] ),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1838_ (.A1(\transfer_count[2][2] ),
    .A2(_0301_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1839_ (.A1(\transfer_count[2][3] ),
    .A2(_0302_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1840_ (.I(_0288_),
    .Z(_0303_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1841_ (.A1(\transfer_count[2][3] ),
    .A2(_0293_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1842_ (.A1(_0303_),
    .A2(_1342_),
    .B(_0304_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1843_ (.A1(\transfer_count[2][2] ),
    .A2(\transfer_count[2][3] ),
    .A3(_1348_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1844_ (.A1(\transfer_count[2][4] ),
    .A2(_0305_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1845_ (.A1(\transfer_count[2][4] ),
    .A2(_0293_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1846_ (.A1(_0303_),
    .A2(_1339_),
    .B(_0306_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1847_ (.A1(\transfer_count[2][2] ),
    .A2(\transfer_count[2][3] ),
    .Z(_0307_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1848_ (.A1(\transfer_count[2][4] ),
    .A2(_0301_),
    .A3(_0307_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1849_ (.A1(\transfer_count[2][5] ),
    .A2(_0308_),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1850_ (.A1(_0287_),
    .A2(_0308_),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1851_ (.A1(_0303_),
    .A2(_0308_),
    .B(_0299_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1852_ (.I0(_0309_),
    .I1(_0310_),
    .S(\transfer_count[2][5] ),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1853_ (.A1(\transfer_count[2][4] ),
    .A2(\transfer_count[2][5] ),
    .A3(_0305_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1854_ (.A1(_0287_),
    .A2(_0311_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1855_ (.A1(_0303_),
    .A2(_0311_),
    .B(_0299_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1856_ (.I0(_0312_),
    .I1(_0313_),
    .S(\transfer_count[2][6] ),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1857_ (.A1(\transfer_count[2][5] ),
    .A2(\transfer_count[2][6] ),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1858_ (.A1(\transfer_count[2][4] ),
    .A2(_0301_),
    .A3(_0307_),
    .A4(_0314_),
    .Z(_0315_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1859_ (.A1(\transfer_count[2][7] ),
    .A2(_0315_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1860_ (.A1(_0287_),
    .A2(_0315_),
    .Z(_0316_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1861_ (.A1(_0303_),
    .A2(_0315_),
    .B(_0299_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1862_ (.I0(_0316_),
    .I1(_0317_),
    .S(\transfer_count[2][7] ),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1863_ (.A1(\transfer_count[2][6] ),
    .A2(\transfer_count[2][7] ),
    .A3(_0311_),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1864_ (.A1(_0287_),
    .A2(_0318_),
    .Z(_0319_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1865_ (.A1(_0303_),
    .A2(_0318_),
    .B(_0299_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1866_ (.I0(_0319_),
    .I1(_0320_),
    .S(\transfer_count[2][8] ),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1867_ (.A1(\transfer_count[2][7] ),
    .A2(\transfer_count[2][8] ),
    .A3(_0315_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1868_ (.A1(\transfer_count[2][9] ),
    .A2(_0321_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1869_ (.A1(_0287_),
    .A2(_0321_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1870_ (.I(_0288_),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1871_ (.A1(_0323_),
    .A2(_0321_),
    .B(_0299_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1872_ (.I0(_0322_),
    .I1(_0324_),
    .S(\transfer_count[2][9] ),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1873_ (.A1(\transfer_count[2][7] ),
    .A2(\transfer_count[2][8] ),
    .A3(\transfer_count[2][9] ),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1874_ (.A1(\transfer_count[2][4] ),
    .A2(_0305_),
    .A3(_0314_),
    .A4(_0325_),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1875_ (.A1(_0287_),
    .A2(_0326_),
    .Z(_0327_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1876_ (.A1(_0323_),
    .A2(_0326_),
    .B(_0299_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1877_ (.I0(_0327_),
    .I1(_0328_),
    .S(\transfer_count[2][10] ),
    .Z(_0078_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1878_ (.A1(\transfer_count[2][10] ),
    .A2(_0315_),
    .A3(_0325_),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1879_ (.A1(\transfer_count[2][11] ),
    .A2(_0329_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1880_ (.A1(_0287_),
    .A2(_0329_),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1881_ (.A1(_0323_),
    .A2(_0329_),
    .B(_0299_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1882_ (.I0(_0330_),
    .I1(_0331_),
    .S(\transfer_count[2][11] ),
    .Z(_0079_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _1883_ (.I(_0286_),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1884_ (.A1(\transfer_count[2][10] ),
    .A2(\transfer_count[2][11] ),
    .A3(_0326_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1885_ (.A1(_0332_),
    .A2(_0333_),
    .Z(_0334_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1886_ (.A1(_0323_),
    .A2(_0333_),
    .B(_0299_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1887_ (.I0(_0334_),
    .I1(_0335_),
    .S(\transfer_count[2][12] ),
    .Z(_0080_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _1888_ (.A1(\transfer_count[2][11] ),
    .A2(\transfer_count[2][12] ),
    .A3(_0329_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1889_ (.A1(\transfer_count[2][13] ),
    .A2(_0336_),
    .Z(_1312_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1890_ (.A1(_0303_),
    .A2(_0336_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1891_ (.I0(_0292_),
    .I1(_0336_),
    .S(_0295_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1892_ (.I0(_0337_),
    .I1(_0338_),
    .S(\transfer_count[2][13] ),
    .Z(_0081_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _1893_ (.A1(\transfer_count[2][12] ),
    .A2(\transfer_count[2][13] ),
    .A3(_0333_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1894_ (.A1(_0295_),
    .A2(_0339_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1895_ (.A1(_0293_),
    .A2(_0340_),
    .B(\transfer_count[2][14] ),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _1896_ (.A1(\transfer_count[2][14] ),
    .A2(_0303_),
    .A3(_0339_),
    .B(_0341_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1897_ (.A1(\transfer_count[2][10] ),
    .A2(\transfer_count[2][11] ),
    .A3(\transfer_count[2][12] ),
    .A4(\transfer_count[2][13] ),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1898_ (.A1(\transfer_count[2][14] ),
    .A2(_0342_),
    .Z(_0343_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1899_ (.A1(_0315_),
    .A2(_0325_),
    .A3(_0343_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1900_ (.A1(\transfer_count[2][15] ),
    .A2(_0344_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1901_ (.A1(_0332_),
    .A2(_0344_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1902_ (.I(_0298_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1903_ (.A1(_0323_),
    .A2(_0344_),
    .B(_0346_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1904_ (.I0(_0345_),
    .I1(_0347_),
    .S(\transfer_count[2][15] ),
    .Z(_0083_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1905_ (.A1(_0326_),
    .A2(_0343_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1906_ (.A1(\transfer_count[2][15] ),
    .A2(_0348_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1907_ (.A1(_0332_),
    .A2(_0349_),
    .Z(_0350_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1908_ (.A1(_0323_),
    .A2(_0349_),
    .B(_0346_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1909_ (.I0(_0350_),
    .I1(_0351_),
    .S(\transfer_count[2][16] ),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1910_ (.A1(\transfer_count[2][15] ),
    .A2(\transfer_count[2][16] ),
    .A3(_0344_),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1911_ (.A1(_0332_),
    .A2(_0352_),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1912_ (.A1(_0323_),
    .A2(_0352_),
    .B(_0346_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1913_ (.I0(_0353_),
    .I1(_0354_),
    .S(\transfer_count[2][17] ),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1914_ (.A1(\transfer_count[2][15] ),
    .A2(\transfer_count[2][16] ),
    .A3(\transfer_count[2][17] ),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1915_ (.A1(_0348_),
    .A2(_0355_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1916_ (.A1(_0332_),
    .A2(_0356_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1917_ (.A1(_0323_),
    .A2(_0356_),
    .B(_0346_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1918_ (.I0(_0357_),
    .I1(_0358_),
    .S(\transfer_count[2][18] ),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1919_ (.A1(\transfer_count[2][18] ),
    .A2(_0344_),
    .A3(_0355_),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1920_ (.A1(\transfer_count[2][19] ),
    .A2(_0359_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1921_ (.A1(_0332_),
    .A2(_0359_),
    .Z(_0360_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1922_ (.A1(_0323_),
    .A2(_0359_),
    .B(_0346_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1923_ (.I0(_0360_),
    .I1(_0361_),
    .S(\transfer_count[2][19] ),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1924_ (.A1(\transfer_count[2][18] ),
    .A2(\transfer_count[2][19] ),
    .A3(_0356_),
    .Z(_0362_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1925_ (.A1(_0332_),
    .A2(_0362_),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1926_ (.A1(_0323_),
    .A2(_0362_),
    .B(_0346_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1927_ (.I0(_0363_),
    .I1(_0364_),
    .S(\transfer_count[2][20] ),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1928_ (.A1(\transfer_count[2][18] ),
    .A2(\transfer_count[2][19] ),
    .A3(\transfer_count[2][20] ),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1929_ (.A1(_0355_),
    .A2(_0365_),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1930_ (.A1(_0344_),
    .A2(_0366_),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1931_ (.A1(\transfer_count[2][21] ),
    .A2(_0367_),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1932_ (.A1(_0332_),
    .A2(_0367_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1933_ (.A1(_0297_),
    .A2(_0367_),
    .B(_0346_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1934_ (.I0(_0368_),
    .I1(_0369_),
    .S(\transfer_count[2][21] ),
    .Z(_0090_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1935_ (.A1(\transfer_count[2][21] ),
    .A2(_0348_),
    .A3(_0366_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1936_ (.A1(_0332_),
    .A2(_0370_),
    .Z(_0371_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1937_ (.A1(_0297_),
    .A2(_0370_),
    .B(_0346_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1938_ (.I0(_0371_),
    .I1(_0372_),
    .S(\transfer_count[2][22] ),
    .Z(_0091_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1939_ (.A1(\transfer_count[2][21] ),
    .A2(\transfer_count[2][22] ),
    .A3(_0355_),
    .A4(_0365_),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1940_ (.A1(_0344_),
    .A2(_0373_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1941_ (.A1(\transfer_count[2][23] ),
    .A2(_0374_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1942_ (.A1(_0332_),
    .A2(_0374_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1943_ (.A1(_0297_),
    .A2(_0374_),
    .B(_0346_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1944_ (.I0(_0375_),
    .I1(_0376_),
    .S(\transfer_count[2][23] ),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1945_ (.A1(_0326_),
    .A2(_0343_),
    .A3(_0373_),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1946_ (.A1(\transfer_count[2][23] ),
    .A2(_0377_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1947_ (.A1(_0295_),
    .A2(_0378_),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1948_ (.A1(_0297_),
    .A2(_0378_),
    .B(_0346_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1949_ (.I0(_0379_),
    .I1(_0380_),
    .S(\transfer_count[2][24] ),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1950_ (.A1(\transfer_count[2][23] ),
    .A2(\transfer_count[2][24] ),
    .A3(_0374_),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1951_ (.A1(\transfer_count[2][25] ),
    .A2(_0381_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1952_ (.A1(_0295_),
    .A2(_0381_),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1953_ (.A1(_0297_),
    .A2(_0381_),
    .B(_0298_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1954_ (.I0(_0382_),
    .I1(_0383_),
    .S(\transfer_count[2][25] ),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1955_ (.A1(\transfer_count[2][23] ),
    .A2(\transfer_count[2][24] ),
    .A3(\transfer_count[2][25] ),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1956_ (.A1(_0377_),
    .A2(_0384_),
    .Z(_0385_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1957_ (.A1(_0295_),
    .A2(_0385_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1958_ (.A1(_0297_),
    .A2(_0385_),
    .B(_0298_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1959_ (.I0(_0386_),
    .I1(_0387_),
    .S(\transfer_count[2][26] ),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1960_ (.A1(\transfer_count[2][26] ),
    .A2(_0374_),
    .A3(_0384_),
    .Z(_0388_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1961_ (.A1(\transfer_count[2][27] ),
    .A2(_0388_),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1962_ (.A1(_0295_),
    .A2(_0388_),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1963_ (.A1(_0297_),
    .A2(_0388_),
    .B(_0298_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1964_ (.I0(_0389_),
    .I1(_0390_),
    .S(\transfer_count[2][27] ),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1965_ (.A1(\transfer_count[2][26] ),
    .A2(\transfer_count[2][27] ),
    .A3(_0384_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1966_ (.A1(_0377_),
    .A2(_0391_),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1967_ (.A1(_0295_),
    .A2(_0392_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1968_ (.A1(_0297_),
    .A2(_0392_),
    .B(_0298_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1969_ (.I0(_0393_),
    .I1(_0394_),
    .S(\transfer_count[2][28] ),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1970_ (.A1(\transfer_count[2][28] ),
    .A2(_0374_),
    .A3(_0391_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1971_ (.A1(\transfer_count[2][29] ),
    .A2(_0395_),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1972_ (.A1(_0295_),
    .A2(_0395_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1973_ (.A1(_0297_),
    .A2(_0395_),
    .B(_0298_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1974_ (.I0(_0396_),
    .I1(_0397_),
    .S(\transfer_count[2][29] ),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1975_ (.A1(\transfer_count[2][28] ),
    .A2(\transfer_count[2][29] ),
    .A3(_0391_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1976_ (.A1(_0377_),
    .A2(_0398_),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1977_ (.A1(_0287_),
    .A2(_0399_),
    .B(\transfer_count[2][30] ),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1978_ (.A1(_0288_),
    .A2(_0399_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1979_ (.A1(\transfer_count[2][30] ),
    .A2(_0299_),
    .A3(_0401_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1980_ (.A1(_0400_),
    .A2(_0402_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _1981_ (.A1(\transfer_count[2][30] ),
    .A2(_0374_),
    .A3(_0398_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1982_ (.A1(_0303_),
    .A2(_0403_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1983_ (.I0(_0292_),
    .I1(_0403_),
    .S(_0295_),
    .Z(_0405_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1984_ (.I0(_0404_),
    .I1(_0405_),
    .S(\transfer_count[2][31] ),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1985_ (.I(\transfer_count[1][0] ),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _1986_ (.A1(_0767_),
    .A2(_0829_),
    .B(_0766_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1987_ (.I0(_0769_),
    .I1(_0406_),
    .S(\transfer_count[1][0] ),
    .Z(_0045_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1988_ (.I(_0406_),
    .Z(_0407_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _1989_ (.A1(_1362_),
    .A2(_0769_),
    .B1(_0407_),
    .B2(\transfer_count[1][1] ),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1990_ (.I(_0408_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _1991_ (.I(_0768_),
    .Z(_0409_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1992_ (.A1(_1361_),
    .A2(_0409_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _1993_ (.A1(_0766_),
    .A2(_0767_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1994_ (.I(_0411_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1995_ (.A1(net139),
    .A2(\channel_state[1][2] ),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1996_ (.A1(net135),
    .A2(_0828_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _1997_ (.A1(_0413_),
    .A2(_0414_),
    .B(\channel_state[1][0] ),
    .C(\channel_state[1][1] ),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1998_ (.I(_0415_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1999_ (.A1(_1361_),
    .A2(_0412_),
    .B(_0416_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2000_ (.I0(_0410_),
    .I1(_0417_),
    .S(\transfer_count[1][2] ),
    .Z(_0067_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2001_ (.A1(\transfer_count[1][0] ),
    .A2(\transfer_count[1][1] ),
    .A3(\transfer_count[1][2] ),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2002_ (.A1(_0769_),
    .A2(_0418_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2003_ (.I(_0411_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2004_ (.A1(_0420_),
    .A2(_0418_),
    .B(_0416_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2005_ (.I0(_0419_),
    .I1(_0421_),
    .S(\transfer_count[1][3] ),
    .Z(_0070_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2006_ (.I(_0420_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2007_ (.A1(_1361_),
    .A2(\transfer_count[1][2] ),
    .A3(\transfer_count[1][3] ),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2008_ (.A1(\transfer_count[1][4] ),
    .A2(_0423_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2009_ (.A1(\transfer_count[1][4] ),
    .A2(_0407_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2010_ (.A1(_0422_),
    .A2(_1381_),
    .B(_0424_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2011_ (.A1(\transfer_count[1][3] ),
    .A2(\transfer_count[1][4] ),
    .A3(_0418_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2012_ (.A1(\transfer_count[1][5] ),
    .A2(_0425_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2013_ (.A1(\transfer_count[1][5] ),
    .A2(_0407_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2014_ (.A1(_0422_),
    .A2(_1378_),
    .B(_0426_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2015_ (.A1(\transfer_count[1][4] ),
    .A2(\transfer_count[1][5] ),
    .A3(_0423_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2016_ (.A1(_0769_),
    .A2(_0427_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2017_ (.A1(_0420_),
    .A2(_0427_),
    .B(_0416_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2018_ (.I0(_0428_),
    .I1(_0429_),
    .S(\transfer_count[1][6] ),
    .Z(_0073_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2019_ (.A1(\transfer_count[1][6] ),
    .A2(_0748_),
    .Z(_0430_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2020_ (.A1(_0769_),
    .A2(_0430_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2021_ (.A1(_0420_),
    .A2(_0430_),
    .B(_0416_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2022_ (.I0(_0431_),
    .I1(_0432_),
    .S(\transfer_count[1][7] ),
    .Z(_0074_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2023_ (.A1(\transfer_count[1][7] ),
    .A2(\transfer_count[1][6] ),
    .A3(_0427_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _2024_ (.I(_0433_),
    .Z(_0434_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2025_ (.A1(_0769_),
    .A2(_0434_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2026_ (.A1(_0420_),
    .A2(_0434_),
    .B(_0416_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2027_ (.I0(_0435_),
    .I1(_0436_),
    .S(\transfer_count[1][8] ),
    .Z(_0075_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2028_ (.A1(\transfer_count[1][9] ),
    .A2(_0407_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2029_ (.A1(_1000_),
    .A2(_0422_),
    .B(_0437_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2030_ (.A1(\transfer_count[1][9] ),
    .A2(\transfer_count[1][8] ),
    .A3(_0434_),
    .Z(_0438_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2031_ (.A1(\transfer_count[1][10] ),
    .A2(_0438_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2032_ (.A1(\transfer_count[1][10] ),
    .A2(_0407_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2033_ (.A1(_0422_),
    .A2(_0997_),
    .B(_0439_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2034_ (.A1(_0749_),
    .A2(_0750_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2035_ (.A1(\transfer_count[1][11] ),
    .A2(_0440_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2036_ (.A1(\transfer_count[1][11] ),
    .A2(_0407_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2037_ (.A1(_0422_),
    .A2(_0994_),
    .B(_0441_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2038_ (.A1(\transfer_count[1][11] ),
    .A2(_0750_),
    .A3(_0433_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2039_ (.A1(\transfer_count[1][12] ),
    .A2(_0442_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2040_ (.A1(\transfer_count[1][12] ),
    .A2(_0407_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2041_ (.A1(_0422_),
    .A2(_0991_),
    .B(_0443_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2042_ (.A1(_0751_),
    .A2(_0768_),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2043_ (.A1(_0406_),
    .A2(_0444_),
    .B(\transfer_count[1][13] ),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2044_ (.A1(\transfer_count[1][13] ),
    .A2(_0751_),
    .A3(_0420_),
    .B(_0445_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2045_ (.A1(_0750_),
    .A2(_0754_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2046_ (.A1(_0446_),
    .A2(_0434_),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2047_ (.A1(\transfer_count[1][14] ),
    .A2(_0447_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2048_ (.A1(\transfer_count[1][14] ),
    .A2(_0407_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2049_ (.A1(_0422_),
    .A2(_0985_),
    .B(_0448_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2050_ (.A1(\transfer_count[1][14] ),
    .A2(_0749_),
    .A3(_0446_),
    .Z(_0449_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2051_ (.A1(\transfer_count[1][15] ),
    .A2(_0449_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2052_ (.A1(\transfer_count[1][15] ),
    .A2(_0407_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2053_ (.A1(_0422_),
    .A2(_0982_),
    .B(_0450_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2054_ (.A1(_0446_),
    .A2(_0755_),
    .A3(_0434_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2055_ (.A1(_0768_),
    .A2(_0451_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2056_ (.A1(_0406_),
    .A2(_0452_),
    .B(\transfer_count[1][16] ),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2057_ (.A1(\transfer_count[1][16] ),
    .A2(_0422_),
    .A3(_0451_),
    .B(_0453_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2058_ (.A1(_0764_),
    .A2(_0409_),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2059_ (.A1(_0764_),
    .A2(_0412_),
    .B(_0416_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2060_ (.I0(_0454_),
    .I1(_0455_),
    .S(\transfer_count[1][17] ),
    .Z(_0053_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2061_ (.A1(_0756_),
    .A2(_0433_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2062_ (.A1(\transfer_count[1][17] ),
    .A2(_0456_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2063_ (.A1(_0769_),
    .A2(_0457_),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2064_ (.A1(_0420_),
    .A2(_0457_),
    .B(_0416_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2065_ (.I0(_0458_),
    .I1(_0459_),
    .S(\transfer_count[1][18] ),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2066_ (.A1(\transfer_count[1][18] ),
    .A2(\transfer_count[1][17] ),
    .A3(_0764_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2067_ (.A1(_0460_),
    .A2(_0409_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2068_ (.A1(_0460_),
    .A2(_0412_),
    .B(_0416_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2069_ (.I0(_0461_),
    .I1(_0462_),
    .S(\transfer_count[1][19] ),
    .Z(_0055_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2070_ (.A1(_0757_),
    .A2(_0456_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2071_ (.A1(_0769_),
    .A2(_0463_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2072_ (.A1(_0420_),
    .A2(_0463_),
    .B(_0416_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2073_ (.I0(_0464_),
    .I1(_0465_),
    .S(\transfer_count[1][20] ),
    .Z(_0057_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2074_ (.A1(\transfer_count[1][20] ),
    .A2(\transfer_count[1][19] ),
    .A3(_0460_),
    .A4(_0768_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2075_ (.A1(_0765_),
    .A2(_0412_),
    .B(_0416_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2076_ (.I0(_0466_),
    .I1(_0467_),
    .S(\transfer_count[1][21] ),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2077_ (.A1(\transfer_count[1][21] ),
    .A2(\transfer_count[1][20] ),
    .A3(_0757_),
    .A4(_0456_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2078_ (.A1(_0409_),
    .A2(_0468_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2079_ (.A1(_0420_),
    .A2(_0468_),
    .B(_0415_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2080_ (.I0(_0469_),
    .I1(_0470_),
    .S(\transfer_count[1][22] ),
    .Z(_0059_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2081_ (.A1(_0762_),
    .A2(_0409_),
    .Z(_0471_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2082_ (.A1(_0762_),
    .A2(_0412_),
    .B(_0415_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2083_ (.I0(_0471_),
    .I1(_0472_),
    .S(\transfer_count[1][23] ),
    .Z(_0060_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2084_ (.A1(\transfer_count[1][23] ),
    .A2(_0759_),
    .A3(_0434_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2085_ (.A1(_0409_),
    .A2(_0473_),
    .Z(_0474_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2086_ (.A1(_0420_),
    .A2(_0473_),
    .B(_0415_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2087_ (.I0(_0474_),
    .I1(_0475_),
    .S(\transfer_count[1][24] ),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2088_ (.A1(_0763_),
    .A2(_0768_),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2089_ (.A1(_0763_),
    .A2(_0412_),
    .B(_0415_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2090_ (.I0(_0476_),
    .I1(_0477_),
    .S(\transfer_count[1][25] ),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2091_ (.A1(_0759_),
    .A2(_0760_),
    .A3(_0434_),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2092_ (.A1(_0409_),
    .A2(_0478_),
    .Z(_0479_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2093_ (.A1(_0412_),
    .A2(_0478_),
    .B(_0415_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2094_ (.I0(_0479_),
    .I1(_0480_),
    .S(\transfer_count[1][26] ),
    .Z(_0063_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _2095_ (.A1(\transfer_count[1][26] ),
    .A2(_0749_),
    .A3(_0759_),
    .A4(_0760_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2096_ (.A1(_0768_),
    .A2(_0481_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2097_ (.A1(_0406_),
    .A2(_0482_),
    .B(\transfer_count[1][27] ),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2098_ (.A1(\transfer_count[1][27] ),
    .A2(_0422_),
    .A3(_0481_),
    .B(_0483_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2099_ (.A1(\transfer_count[1][27] ),
    .A2(\transfer_count[1][26] ),
    .A3(\transfer_count[1][24] ),
    .A4(\transfer_count[1][23] ),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2100_ (.A1(\transfer_count[1][25] ),
    .A2(_0759_),
    .A3(_0434_),
    .A4(_0484_),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2101_ (.A1(_0409_),
    .A2(_0485_),
    .Z(_0486_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2102_ (.A1(_0412_),
    .A2(_0485_),
    .B(_0415_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2103_ (.I0(_0486_),
    .I1(_0487_),
    .S(\transfer_count[1][28] ),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2104_ (.A1(_0761_),
    .A2(_0768_),
    .Z(_0488_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2105_ (.A1(_0761_),
    .A2(_0411_),
    .B(_0415_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2106_ (.I0(_0488_),
    .I1(_0489_),
    .S(\transfer_count[1][29] ),
    .Z(_0066_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2107_ (.A1(\transfer_count[1][29] ),
    .A2(_0753_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2108_ (.A1(_0759_),
    .A2(_0760_),
    .A3(_0434_),
    .A4(_0490_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2109_ (.A1(_0409_),
    .A2(_0491_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2110_ (.A1(_0412_),
    .A2(_0491_),
    .B(_0415_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2111_ (.I0(_0492_),
    .I1(_0493_),
    .S(\transfer_count[1][30] ),
    .Z(_0068_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2112_ (.A1(\transfer_count[1][30] ),
    .A2(\transfer_count[1][29] ),
    .A3(_0761_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2113_ (.A1(_0409_),
    .A2(_0494_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2114_ (.A1(_0412_),
    .A2(_0494_),
    .B(_0415_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2115_ (.I0(_0495_),
    .I1(_0496_),
    .S(\transfer_count[1][31] ),
    .Z(_0069_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2116_ (.I(\transfer_count[0][0] ),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2117_ (.A1(net138),
    .A2(\channel_state[0][2] ),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2118_ (.A1(\channel_state[0][0] ),
    .A2(\channel_state[0][1] ),
    .A3(_0497_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2119_ (.I(_0498_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _2120_ (.A1(_0499_),
    .A2(_0193_),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2121_ (.I0(_0952_),
    .I1(_0500_),
    .S(\transfer_count[0][0] ),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2122_ (.A1(\transfer_count[0][1] ),
    .A2(_0193_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2123_ (.I(_0499_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2124_ (.I0(_1158_),
    .I1(_0501_),
    .S(_0502_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _2125_ (.I(_0951_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2126_ (.A1(_1157_),
    .A2(_0503_),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2127_ (.I(_0499_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2128_ (.A1(_0499_),
    .A2(_0193_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2129_ (.I(_0506_),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2130_ (.A1(_1157_),
    .A2(_0505_),
    .B(_0507_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2131_ (.I0(_0504_),
    .I1(_0508_),
    .S(\transfer_count[0][2] ),
    .Z(_0035_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2132_ (.A1(_0928_),
    .A2(_0503_),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2133_ (.A1(_0928_),
    .A2(_0505_),
    .B(_0507_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2134_ (.I0(_0509_),
    .I1(_0510_),
    .S(\transfer_count[0][3] ),
    .Z(_0038_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2135_ (.A1(\transfer_count[0][2] ),
    .A2(\transfer_count[0][3] ),
    .A3(_1157_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2136_ (.A1(\transfer_count[0][4] ),
    .A2(_0511_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2137_ (.A1(\transfer_count[0][4] ),
    .A2(_0502_),
    .A3(_0193_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2138_ (.A1(_0502_),
    .A2(_1177_),
    .B(_0512_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2139_ (.A1(\transfer_count[0][5] ),
    .A2(_0500_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2140_ (.A1(_1174_),
    .A2(_0502_),
    .B(_0513_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2141_ (.A1(\transfer_count[0][2] ),
    .A2(_1157_),
    .A3(_0932_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2142_ (.A1(_0952_),
    .A2(_0514_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2143_ (.I(_0499_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2144_ (.A1(_0516_),
    .A2(_0514_),
    .B(_0507_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2145_ (.I0(_0515_),
    .I1(_0517_),
    .S(\transfer_count[0][6] ),
    .Z(_0041_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2146_ (.A1(_0935_),
    .A2(_0503_),
    .Z(_0518_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2147_ (.A1(_0935_),
    .A2(_0505_),
    .B(_0507_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2148_ (.I0(_0518_),
    .I1(_0519_),
    .S(\transfer_count[0][7] ),
    .Z(_0042_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2149_ (.A1(\transfer_count[0][6] ),
    .A2(\transfer_count[0][7] ),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2150_ (.A1(\transfer_count[0][2] ),
    .A2(_1157_),
    .A3(_0932_),
    .A4(_0520_),
    .Z(_0521_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2151_ (.A1(_0952_),
    .A2(_0521_),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2152_ (.A1(_0516_),
    .A2(_0521_),
    .B(_0507_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2153_ (.I0(_0522_),
    .I1(_0523_),
    .S(\transfer_count[0][8] ),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2154_ (.A1(_0937_),
    .A2(_0516_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2155_ (.I0(_0937_),
    .I1(_0193_),
    .S(_0499_),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2156_ (.I0(_0524_),
    .I1(_0525_),
    .S(\transfer_count[0][9] ),
    .Z(_0044_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2157_ (.A1(\transfer_count[0][9] ),
    .A2(\transfer_count[0][8] ),
    .A3(_0521_),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2158_ (.A1(\transfer_count[0][10] ),
    .A2(_0526_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2159_ (.A1(\transfer_count[0][10] ),
    .A2(_0500_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2160_ (.A1(_0502_),
    .A2(_1195_),
    .B(_0527_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2161_ (.A1(_0931_),
    .A2(_0936_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2162_ (.A1(_0528_),
    .A2(_0516_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2163_ (.I0(_0528_),
    .I1(_0193_),
    .S(_0499_),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2164_ (.I0(_0529_),
    .I1(_0530_),
    .S(\transfer_count[0][11] ),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2165_ (.A1(\transfer_count[0][11] ),
    .A2(_0931_),
    .A3(_0521_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2166_ (.A1(\transfer_count[0][12] ),
    .A2(_0531_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2167_ (.A1(\transfer_count[0][12] ),
    .A2(_0500_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2168_ (.A1(_0502_),
    .A2(_1189_),
    .B(_0532_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2169_ (.A1(_0934_),
    .A2(_0951_),
    .Z(_0533_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2170_ (.A1(_0500_),
    .A2(_0533_),
    .B(\transfer_count[0][13] ),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2171_ (.A1(\transfer_count[0][13] ),
    .A2(_0934_),
    .A3(_0502_),
    .B(_0534_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2172_ (.A1(\transfer_count[0][13] ),
    .A2(_0930_),
    .A3(_0931_),
    .A4(_0521_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2173_ (.A1(\transfer_count[0][14] ),
    .A2(_0535_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2174_ (.A1(\transfer_count[0][14] ),
    .A2(_0500_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2175_ (.A1(_0502_),
    .A2(_1183_),
    .B(_0536_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2176_ (.A1(_0933_),
    .A2(_0942_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2177_ (.A1(_0537_),
    .A2(_0951_),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2178_ (.A1(_0500_),
    .A2(_0538_),
    .B(\transfer_count[0][15] ),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2179_ (.A1(\transfer_count[0][15] ),
    .A2(_0537_),
    .A3(_0502_),
    .B(_0539_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2180_ (.A1(\transfer_count[0][15] ),
    .A2(_0942_),
    .A3(_0521_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2181_ (.A1(_0952_),
    .A2(_0540_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2182_ (.A1(_0516_),
    .A2(_0540_),
    .B(_0507_),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2183_ (.I0(_0541_),
    .I1(_0542_),
    .S(\transfer_count[0][16] ),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2184_ (.A1(_0948_),
    .A2(_0503_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2185_ (.A1(_0948_),
    .A2(_0505_),
    .B(_0507_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2186_ (.I0(_0543_),
    .I1(_0544_),
    .S(\transfer_count[0][17] ),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2187_ (.A1(\transfer_count[0][17] ),
    .A2(\transfer_count[0][16] ),
    .A3(_0540_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2188_ (.A1(_0952_),
    .A2(_0545_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2189_ (.A1(_0516_),
    .A2(_0545_),
    .B(_0507_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2190_ (.I0(_0546_),
    .I1(_0547_),
    .S(\transfer_count[0][18] ),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2191_ (.A1(\transfer_count[0][18] ),
    .A2(\transfer_count[0][17] ),
    .A3(\transfer_count[0][16] ),
    .A4(_0943_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2192_ (.A1(_0952_),
    .A2(_0548_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2193_ (.A1(_0516_),
    .A2(_0548_),
    .B(_0507_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2194_ (.I0(_0549_),
    .I1(_0550_),
    .S(\transfer_count[0][19] ),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2195_ (.A1(_0940_),
    .A2(_0540_),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2196_ (.A1(_0952_),
    .A2(_0551_),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2197_ (.I(_0506_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2198_ (.A1(_0516_),
    .A2(_0551_),
    .B(_0553_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2199_ (.I0(_0552_),
    .I1(_0554_),
    .S(\transfer_count[0][20] ),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2200_ (.A1(_0947_),
    .A2(_0951_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2201_ (.A1(_0947_),
    .A2(_0505_),
    .B(_0553_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2202_ (.I0(_0555_),
    .I1(_0556_),
    .S(\transfer_count[0][21] ),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2203_ (.A1(_0941_),
    .A2(_0540_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2204_ (.A1(_0952_),
    .A2(_0557_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2205_ (.A1(_0516_),
    .A2(_0557_),
    .B(_0553_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2206_ (.I0(_0558_),
    .I1(_0559_),
    .S(\transfer_count[0][22] ),
    .Z(_0027_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2207_ (.A1(\transfer_count[0][22] ),
    .A2(_0945_),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2208_ (.A1(_0503_),
    .A2(_0560_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2209_ (.A1(_0516_),
    .A2(_0560_),
    .B(_0553_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2210_ (.I0(_0561_),
    .I1(_0562_),
    .S(\transfer_count[0][23] ),
    .Z(_0028_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2211_ (.A1(\transfer_count[0][23] ),
    .A2(\transfer_count[0][22] ),
    .A3(_0557_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2212_ (.A1(_0503_),
    .A2(_0563_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2213_ (.A1(_0505_),
    .A2(_0563_),
    .B(_0553_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2214_ (.I0(_0564_),
    .I1(_0565_),
    .S(\transfer_count[0][24] ),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2215_ (.A1(_0946_),
    .A2(_0951_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2216_ (.A1(_0946_),
    .A2(_0499_),
    .B(_0553_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2217_ (.I0(_0566_),
    .I1(_0567_),
    .S(\transfer_count[0][25] ),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2218_ (.A1(_0938_),
    .A2(_0557_),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2219_ (.A1(_0503_),
    .A2(_0568_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2220_ (.A1(_0505_),
    .A2(_0568_),
    .B(_0553_),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2221_ (.I0(_0569_),
    .I1(_0570_),
    .S(\transfer_count[0][26] ),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2222_ (.A1(\transfer_count[0][26] ),
    .A2(_0938_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2223_ (.A1(_0571_),
    .A2(_0941_),
    .A3(_0943_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2224_ (.A1(_0503_),
    .A2(_0572_),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2225_ (.A1(_0505_),
    .A2(_0572_),
    .B(_0553_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2226_ (.I0(_0573_),
    .I1(_0574_),
    .S(\transfer_count[0][27] ),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2227_ (.A1(\transfer_count[0][27] ),
    .A2(_0571_),
    .A3(_0557_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2228_ (.A1(_0503_),
    .A2(_0575_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2229_ (.A1(_0505_),
    .A2(_0575_),
    .B(_0553_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2230_ (.I0(_0576_),
    .I1(_0577_),
    .S(\transfer_count[0][28] ),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2231_ (.A1(_0944_),
    .A2(_0951_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2232_ (.A1(_0944_),
    .A2(_0499_),
    .B(_0553_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2233_ (.I0(_0578_),
    .I1(_0579_),
    .S(\transfer_count[0][29] ),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2234_ (.A1(\transfer_count[0][29] ),
    .A2(_0939_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2235_ (.A1(_0557_),
    .A2(_0580_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2236_ (.A1(_0503_),
    .A2(_0581_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2237_ (.A1(_0505_),
    .A2(_0581_),
    .B(_0506_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2238_ (.I0(_0582_),
    .I1(_0583_),
    .S(\transfer_count[0][30] ),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2239_ (.A1(\transfer_count[0][30] ),
    .A2(_0945_),
    .A3(_0580_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2240_ (.A1(_0951_),
    .A2(_0584_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2241_ (.A1(_0500_),
    .A2(_0585_),
    .B(\transfer_count[0][31] ),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2242_ (.A1(\transfer_count[0][31] ),
    .A2(_0502_),
    .A3(_0584_),
    .B(_0586_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2243_ (.I(\active_channel_count[0] ),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2244_ (.A1(_0949_),
    .A2(\channel_state[0][1] ),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2245_ (.A1(\channel_state[0][0] ),
    .A2(_0925_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2246_ (.A1(_0587_),
    .A2(_0588_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2247_ (.A1(\channel_state[0][2] ),
    .A2(_0589_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2248_ (.A1(net2),
    .A2(net146),
    .A3(_0590_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2249_ (.I(\channel_state[1][1] ),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2250_ (.A1(\channel_state[1][0] ),
    .A2(_0592_),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2251_ (.A1(\channel_state[1][0] ),
    .A2(_0592_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2252_ (.A1(_0593_),
    .A2(_0594_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2253_ (.A1(\channel_state[1][2] ),
    .A2(_0595_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2254_ (.A1(net147),
    .A2(net3),
    .A3(_0596_),
    .Z(_0597_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2255_ (.I(\channel_state[3][0] ),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2256_ (.A1(_0598_),
    .A2(\channel_state[3][1] ),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _2257_ (.I(\channel_state[3][1] ),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2258_ (.A1(\channel_state[3][0] ),
    .A2(_0600_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2259_ (.A1(_0599_),
    .A2(_0601_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2260_ (.A1(\channel_state[3][2] ),
    .A2(_0602_),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2261_ (.A1(net149),
    .A2(net5),
    .A3(_0603_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2262_ (.A1(_0283_),
    .A2(\channel_state[2][1] ),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _2263_ (.I(\channel_state[2][1] ),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2264_ (.A1(\channel_state[2][0] ),
    .A2(_0606_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2265_ (.A1(_0605_),
    .A2(_0607_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2266_ (.I(net148),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _2267_ (.A1(\channel_state[2][2] ),
    .A2(_0608_),
    .B(_0609_),
    .C(_0289_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2268_ (.A1(_0591_),
    .A2(_0597_),
    .A3(_0604_),
    .A4(_0610_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2269_ (.A1(_1252_),
    .A2(_0611_),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2270_ (.A1(_1255_),
    .A2(_0611_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2271_ (.A1(_1256_),
    .A2(\active_channel_count[2] ),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2272_ (.A1(_0611_),
    .A2(_0612_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2273_ (.A1(\active_channel_count[0] ),
    .A2(\active_channel_count[2] ),
    .A3(\active_channel_count[1] ),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2274_ (.A1(\active_channel_count[3] ),
    .A2(_0613_),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2275_ (.A1(_0611_),
    .A2(_0614_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2276_ (.A1(net134),
    .A2(\channel_state[0][0] ),
    .A3(_0925_),
    .A4(\channel_state[0][2] ),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2277_ (.A1(_0949_),
    .A2(\channel_state[0][1] ),
    .A3(_0922_),
    .A4(net142),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2278_ (.A1(_0507_),
    .A2(_0615_),
    .A3(_0616_),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2279_ (.A1(\channel_state[0][2] ),
    .A2(_0588_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2280_ (.A1(_0949_),
    .A2(\channel_state[0][1] ),
    .A3(_0923_),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2281_ (.A1(_0968_),
    .A2(_0617_),
    .Z(_0980_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2282_ (.A1(\channel_state[0][0] ),
    .A2(\channel_state[0][1] ),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2283_ (.A1(net134),
    .A2(_0950_),
    .B(_0618_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2284_ (.I0(_0618_),
    .I1(_0619_),
    .S(\channel_state[0][2] ),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2285_ (.A1(net134),
    .A2(_0589_),
    .B(_0192_),
    .C(_0497_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2286_ (.A1(_0620_),
    .A2(_0621_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2287_ (.A1(_0827_),
    .A2(net143),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2288_ (.I(net135),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2289_ (.A1(\channel_state[1][2] ),
    .A2(\channel_state[1][0] ),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2290_ (.A1(_0623_),
    .A2(\channel_state[1][1] ),
    .A3(_0624_),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2291_ (.A1(_0593_),
    .A2(_0622_),
    .B(_0625_),
    .C(_0407_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2292_ (.A1(\channel_state[1][2] ),
    .A2(_0594_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2293_ (.A1(_0827_),
    .A2(_0595_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2294_ (.A1(_0623_),
    .A2(_0593_),
    .B(_0626_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2295_ (.I(net139),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2296_ (.A1(_0623_),
    .A2(_0624_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2297_ (.A1(_0627_),
    .A2(\channel_state[1][1] ),
    .A3(_0826_),
    .A4(_0628_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2298_ (.A1(\channel_state[1][0] ),
    .A2(\channel_state[1][1] ),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2299_ (.A1(net135),
    .A2(_0592_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2300_ (.A1(_0623_),
    .A2(\channel_state[1][1] ),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2301_ (.A1(\channel_state[1][0] ),
    .A2(_0632_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2302_ (.A1(_0631_),
    .A2(_0633_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2303_ (.I0(_0630_),
    .I1(_0634_),
    .S(\channel_state[1][2] ),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2304_ (.A1(_0629_),
    .A2(_0635_),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2305_ (.A1(net136),
    .A2(_0606_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2306_ (.A1(\channel_state[2][2] ),
    .A2(\channel_state[2][0] ),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2307_ (.I(\channel_state[2][2] ),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2308_ (.A1(_0638_),
    .A2(net144),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _2309_ (.A1(_0636_),
    .A2(_0637_),
    .B1(_0639_),
    .B2(_0605_),
    .C(_0293_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _2310_ (.A1(\channel_state[2][2] ),
    .A2(_0607_),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2311_ (.A1(_0638_),
    .A2(_0608_),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2312_ (.A1(_0290_),
    .A2(_0605_),
    .B(_0640_),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2313_ (.A1(net136),
    .A2(_0606_),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2314_ (.I0(\channel_state[2][1] ),
    .I1(_0641_),
    .S(\channel_state[2][2] ),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2315_ (.A1(_0290_),
    .A2(\channel_state[2][1] ),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2316_ (.A1(net140),
    .A2(_0606_),
    .B(_0284_),
    .C(_0643_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2317_ (.A1(\channel_state[2][0] ),
    .A2(_0642_),
    .B(_0644_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2318_ (.A1(\channel_state[2][0] ),
    .A2(_0643_),
    .B(_0636_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2319_ (.A1(_0638_),
    .A2(\channel_state[2][0] ),
    .A3(\channel_state[2][1] ),
    .Z(_0647_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2320_ (.A1(\channel_state[2][2] ),
    .A2(_0646_),
    .B(_0647_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2321_ (.I(_1299_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2322_ (.A1(_1304_),
    .A2(_1302_),
    .B(_1301_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2323_ (.A1(_0649_),
    .A2(_0650_),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2324_ (.A1(_1298_),
    .A2(_0651_),
    .B(_1296_),
    .C(_1293_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2325_ (.A1(_1293_),
    .A2(_1295_),
    .B(_1289_),
    .C(_1292_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2326_ (.A1(_0652_),
    .A2(_0653_),
    .Z(_0654_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2327_ (.A1(_1269_),
    .A2(_1275_),
    .A3(_1281_),
    .A4(_1278_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2328_ (.A1(_1260_),
    .A2(_1272_),
    .A3(_1263_),
    .A4(_1266_),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2329_ (.A1(_1284_),
    .A2(_1287_),
    .A3(_0655_),
    .A4(_0656_),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2330_ (.A1(_1290_),
    .A2(_1289_),
    .B(_0657_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2331_ (.A1(_1260_),
    .A2(_1263_),
    .A3(_1266_),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2332_ (.A1(_1280_),
    .A2(_1278_),
    .B(_1274_),
    .C(_1277_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2333_ (.A1(_1275_),
    .A2(_1274_),
    .B(_1272_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2334_ (.A1(_0660_),
    .A2(_0661_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2335_ (.A1(_1268_),
    .A2(_1271_),
    .A3(_0662_),
    .Z(_0663_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _2336_ (.A1(_1268_),
    .A2(_1269_),
    .B(_0659_),
    .C(_0663_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2337_ (.I(_1259_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2338_ (.A1(_1263_),
    .A2(_1265_),
    .Z(_0666_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2339_ (.A1(_1262_),
    .A2(_0666_),
    .B(_1260_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2340_ (.A1(_1284_),
    .A2(_1286_),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2341_ (.A1(_1283_),
    .A2(_0668_),
    .B(_0655_),
    .C(_0656_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2342_ (.A1(_0665_),
    .A2(_0667_),
    .A3(_0669_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _2343_ (.A1(_0654_),
    .A2(_0658_),
    .B(_0664_),
    .C(_0670_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2344_ (.I(_1323_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2345_ (.A1(_1328_),
    .A2(_1326_),
    .B(_1325_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2346_ (.A1(_0672_),
    .A2(_0673_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2347_ (.A1(_1322_),
    .A2(_0674_),
    .B(_1320_),
    .C(_1317_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2348_ (.A1(_1317_),
    .A2(_1319_),
    .B(_1313_),
    .C(_1316_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2349_ (.A1(_0675_),
    .A2(_0676_),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2350_ (.A1(_1314_),
    .A2(_1313_),
    .B(_1308_),
    .C(_1311_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2351_ (.A1(_1296_),
    .A2(_1293_),
    .A3(_1305_),
    .A4(_1290_),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2352_ (.A1(_1299_),
    .A2(_1302_),
    .A3(_0679_),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2353_ (.A1(_0657_),
    .A2(_0680_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2354_ (.A1(_1308_),
    .A2(_1310_),
    .B(_1307_),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2355_ (.A1(_1317_),
    .A2(_1323_),
    .A3(_1329_),
    .A4(_1314_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2356_ (.A1(_1308_),
    .A2(_1320_),
    .A3(_1311_),
    .A4(_1326_),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2357_ (.A1(_0683_),
    .A2(_0684_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2358_ (.A1(_0682_),
    .A2(_0685_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2359_ (.A1(_0657_),
    .A2(_0686_),
    .A3(_0680_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2360_ (.A1(_1332_),
    .A2(_1335_),
    .A3(_1341_),
    .A4(_1338_),
    .Z(_0688_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2361_ (.I(_1355_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2362_ (.A1(_1352_),
    .A2(_0689_),
    .B(_1351_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2363_ (.A1(_1344_),
    .A2(_1347_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2364_ (.A1(_1344_),
    .A2(_1346_),
    .B(_1343_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2365_ (.A1(_0690_),
    .A2(_0691_),
    .B(_0692_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2366_ (.A1(_1332_),
    .A2(_1335_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2367_ (.A1(_1340_),
    .A2(_1338_),
    .B(_1337_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2368_ (.A1(_1332_),
    .A2(_1334_),
    .B(_1331_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2369_ (.A1(_0694_),
    .A2(_0695_),
    .B(_0682_),
    .C(_0696_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2370_ (.A1(_0688_),
    .A2(_0693_),
    .B(_0697_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _2371_ (.A1(_0677_),
    .A2(_0678_),
    .A3(_0681_),
    .B1(_0687_),
    .B2(_0698_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2372_ (.A1(_0648_),
    .A2(_0671_),
    .A3(_0699_),
    .Z(_0700_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2373_ (.A1(_1344_),
    .A2(_1352_),
    .A3(_1356_),
    .A4(_1347_),
    .Z(_0701_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2374_ (.A1(_0688_),
    .A2(_0701_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2375_ (.A1(_0648_),
    .A2(_0685_),
    .A3(_0681_),
    .A4(_0702_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2376_ (.A1(_0645_),
    .A2(_0700_),
    .A3(_0703_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2377_ (.A1(\channel_state[3][2] ),
    .A2(_0601_),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2378_ (.A1(net137),
    .A2(_0600_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2379_ (.A1(\channel_state[3][2] ),
    .A2(\channel_state[3][0] ),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2380_ (.A1(_0918_),
    .A2(net145),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _2381_ (.A1(_0704_),
    .A2(_0705_),
    .B1(_0706_),
    .B2(_0599_),
    .C(_0196_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2382_ (.I(net137),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2383_ (.A1(_0918_),
    .A2(_0602_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2384_ (.A1(_0707_),
    .A2(_0599_),
    .B(_0708_),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2385_ (.A1(_0879_),
    .A2(_0888_),
    .B(_0912_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2386_ (.A1(_0707_),
    .A2(\channel_state[3][1] ),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2387_ (.A1(\channel_state[3][0] ),
    .A2(_0710_),
    .B(_0704_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2388_ (.A1(_0918_),
    .A2(\channel_state[3][0] ),
    .A3(\channel_state[3][1] ),
    .Z(_0712_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2389_ (.A1(\channel_state[3][2] ),
    .A2(_0711_),
    .B(_0712_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2390_ (.I0(_0600_),
    .I1(_0704_),
    .S(\channel_state[3][2] ),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2391_ (.A1(net141),
    .A2(_0600_),
    .Z(_0715_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2392_ (.A1(_0918_),
    .A2(\channel_state[3][0] ),
    .A3(_0710_),
    .A4(_0715_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _2393_ (.A1(_0709_),
    .A2(_0713_),
    .B1(_0714_),
    .B2(_0598_),
    .C(_0716_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2394_ (.A1(net142),
    .A2(_0587_),
    .B(_0588_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2395_ (.A1(_0922_),
    .A2(_0717_),
    .Z(_1391_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2396_ (.A1(_0952_),
    .A2(_0192_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2397_ (.I0(_0923_),
    .I1(_0924_),
    .S(_0949_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2398_ (.A1(\channel_state[0][1] ),
    .A2(_0719_),
    .B(net150),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2399_ (.A1(_0718_),
    .A2(_0720_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2400_ (.A1(net143),
    .A2(_0593_),
    .B(_0594_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2401_ (.A1(_0827_),
    .A2(_0721_),
    .Z(_1389_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2402_ (.A1(_0769_),
    .A2(_0826_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2403_ (.A1(\channel_state[1][0] ),
    .A2(_0414_),
    .B1(_0624_),
    .B2(net135),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2404_ (.A1(_0592_),
    .A2(_0723_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2405_ (.A1(net151),
    .A2(_0724_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2406_ (.A1(_0722_),
    .A2(_0725_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2407_ (.A1(_0598_),
    .A2(net137),
    .A3(_0919_),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2408_ (.A1(net137),
    .A2(_0705_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2409_ (.A1(_0726_),
    .A2(_0727_),
    .B(_0600_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2410_ (.A1(net153),
    .A2(_0728_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2411_ (.A1(_0917_),
    .A2(_0729_),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2412_ (.A1(net144),
    .A2(_0605_),
    .B(_0607_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2413_ (.A1(_0638_),
    .A2(_0730_),
    .Z(_1386_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2414_ (.A1(_0288_),
    .A2(_0685_),
    .A3(_0681_),
    .A4(_0702_),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2415_ (.A1(_0303_),
    .A2(_0671_),
    .A3(_0699_),
    .B(_0731_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2416_ (.A1(net136),
    .A2(_0637_),
    .B(_0291_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2417_ (.A1(_0606_),
    .A2(_0733_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2418_ (.A1(net152),
    .A2(_0734_),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2419_ (.A1(_0732_),
    .A2(_0735_),
    .Z(_1385_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2420_ (.I(_1254_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2421_ (.A1(\active_channel_count[2] ),
    .A2(\active_channel_count[3] ),
    .A3(_0736_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2422_ (.A1(net137),
    .A2(_0600_),
    .Z(_0737_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2423_ (.A1(_0919_),
    .A2(_0737_),
    .B1(_0710_),
    .B2(\channel_state[3][2] ),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2424_ (.A1(\channel_state[3][0] ),
    .A2(_0738_),
    .Z(_0739_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2425_ (.A1(net157),
    .A2(_0739_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2426_ (.A1(net4),
    .A2(_0638_),
    .A3(_0641_),
    .Z(_0740_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2427_ (.A1(\channel_state[2][2] ),
    .A2(_0643_),
    .Z(_0741_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2428_ (.A1(_0740_),
    .A2(_0741_),
    .B(_0283_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2429_ (.A1(net156),
    .A2(_0742_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2430_ (.A1(_0609_),
    .A2(_0292_),
    .B(_0732_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2431_ (.A1(_0828_),
    .A2(_0631_),
    .B1(_0632_),
    .B2(\channel_state[1][2] ),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2432_ (.A1(\channel_state[1][0] ),
    .A2(_0743_),
    .Z(_0744_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2433_ (.A1(net155),
    .A2(_0744_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2434_ (.I(net129),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2435_ (.I(net6),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2436_ (.A1(\transfer_count[2][30] ),
    .A2(_0399_),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2437_ (.A1(\transfer_count[2][26] ),
    .A2(_0385_),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2438_ (.I(net94),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2439_ (.I(net59),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2440_ (.A1(\transfer_count[1][8] ),
    .A2(_0434_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2441_ (.A1(\transfer_count[1][31] ),
    .A2(_0494_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2442_ (.A1(\transfer_count[1][30] ),
    .A2(_0491_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2443_ (.A1(\transfer_count[1][28] ),
    .A2(_0485_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2444_ (.A1(\transfer_count[1][27] ),
    .A2(_0481_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2445_ (.A1(\transfer_count[1][26] ),
    .A2(_0478_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2446_ (.A1(\transfer_count[1][24] ),
    .A2(_0473_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2447_ (.A1(\transfer_count[1][23] ),
    .A2(_0762_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2448_ (.A1(\transfer_count[1][22] ),
    .A2(_0468_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2449_ (.A1(\transfer_count[1][20] ),
    .A2(_0463_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2450_ (.A1(\transfer_count[1][19] ),
    .A2(_0460_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2451_ (.A1(\transfer_count[1][18] ),
    .A2(_0457_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2452_ (.A1(\transfer_count[1][16] ),
    .A2(_0451_),
    .Z(_1051_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2453_ (.A1(\transfer_count[3][31] ),
    .A2(_0280_),
    .Z(_1054_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2454_ (.A1(\transfer_count[3][30] ),
    .A2(_0276_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2455_ (.A1(\transfer_count[3][28] ),
    .A2(_0269_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2456_ (.A1(\transfer_count[3][26] ),
    .A2(_0263_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2457_ (.A1(\transfer_count[3][24] ),
    .A2(_0257_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2458_ (.A1(\transfer_count[3][22] ),
    .A2(_0251_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2459_ (.A1(\transfer_count[3][20] ),
    .A2(_0247_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2460_ (.A1(\transfer_count[3][18] ),
    .A2(_0243_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2461_ (.A1(\transfer_count[3][17] ),
    .A2(_0238_),
    .Z(_1096_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2462_ (.A1(\transfer_count[3][16] ),
    .A2(_0235_),
    .Z(_1099_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2463_ (.A1(\transfer_count[3][14] ),
    .A2(_0230_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2464_ (.A1(\transfer_count[3][6] ),
    .A2(_0210_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2465_ (.A1(\transfer_count[3][2] ),
    .A2(_1144_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2466_ (.A1(\transfer_count[0][3] ),
    .A2(_0928_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2467_ (.A1(\transfer_count[0][2] ),
    .A2(_1157_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2468_ (.A1(\transfer_count[0][7] ),
    .A2(_0935_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2469_ (.A1(\transfer_count[0][6] ),
    .A2(_0514_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2470_ (.A1(\transfer_count[0][15] ),
    .A2(_0537_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2471_ (.A1(\transfer_count[0][11] ),
    .A2(_0528_),
    .Z(_1192_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2472_ (.A1(\transfer_count[0][8] ),
    .A2(_0521_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2473_ (.A1(\transfer_count[0][31] ),
    .A2(_0584_),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2474_ (.A1(\transfer_count[0][30] ),
    .A2(_0581_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2475_ (.A1(\transfer_count[0][28] ),
    .A2(_0575_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2476_ (.A1(\transfer_count[0][27] ),
    .A2(_0572_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2477_ (.A1(\transfer_count[0][26] ),
    .A2(_0568_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2478_ (.A1(\transfer_count[0][24] ),
    .A2(_0563_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2479_ (.A1(\transfer_count[0][23] ),
    .A2(_0560_),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2480_ (.A1(\transfer_count[0][22] ),
    .A2(_0557_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2481_ (.A1(\transfer_count[0][20] ),
    .A2(_0551_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2482_ (.A1(\transfer_count[0][19] ),
    .A2(_0548_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2483_ (.A1(\transfer_count[0][18] ),
    .A2(_0545_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2484_ (.A1(\transfer_count[0][16] ),
    .A2(_0540_),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2485_ (.I(\active_channel_count[1] ),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2486_ (.A1(\transfer_count[2][31] ),
    .A2(_0403_),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2487_ (.A1(\transfer_count[2][28] ),
    .A2(_0392_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2488_ (.A1(\transfer_count[2][24] ),
    .A2(_0378_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2489_ (.A1(\transfer_count[2][22] ),
    .A2(_0370_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2490_ (.A1(\transfer_count[2][20] ),
    .A2(_0362_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2491_ (.A1(\transfer_count[2][18] ),
    .A2(_0356_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2492_ (.A1(\transfer_count[2][17] ),
    .A2(_0352_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2493_ (.A1(\transfer_count[2][16] ),
    .A2(_0349_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2494_ (.A1(\transfer_count[2][14] ),
    .A2(_0339_),
    .Z(_1309_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2495_ (.A1(\transfer_count[2][12] ),
    .A2(_0333_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2496_ (.A1(\transfer_count[2][10] ),
    .A2(_0326_),
    .ZN(_1321_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2497_ (.A1(\transfer_count[2][8] ),
    .A2(_0318_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2498_ (.A1(\transfer_count[2][6] ),
    .A2(_0311_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2499_ (.A1(\transfer_count[2][2] ),
    .A2(_1348_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2500_ (.A1(\transfer_count[1][3] ),
    .A2(_0418_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2501_ (.A1(_1361_),
    .A2(\transfer_count[1][2] ),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2502_ (.A1(\transfer_count[1][7] ),
    .A2(_0430_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2503_ (.A1(\transfer_count[1][6] ),
    .A2(_0427_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2504_ (.I(_1145_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2505_ (.I(_1158_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2506_ (.I(_1349_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2507_ (.I(_1362_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2508_ (.A1(\channel_state[0][2] ),
    .A2(_0950_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2509_ (.A1(\channel_state[0][2] ),
    .A2(_0618_),
    .B(_0745_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2510_ (.I0(_0766_),
    .I1(_0630_),
    .S(_0827_),
    .Z(_0142_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2511_ (.A1(_0285_),
    .A2(_0647_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2512_ (.A1(_0914_),
    .A2(_0712_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2513_ (.A1(net145),
    .A2(_0599_),
    .B(_0601_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2514_ (.A1(_0918_),
    .A2(_0746_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2515_ (.A(net75),
    .B(_0982_),
    .CO(_0983_),
    .S(_0984_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2516_ (.A(net74),
    .B(_0985_),
    .CO(_0986_),
    .S(_0987_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2517_ (.A(net73),
    .B(_0988_),
    .CO(_0989_),
    .S(_0990_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2518_ (.A(net72),
    .B(_0991_),
    .CO(_0992_),
    .S(_0993_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2519_ (.A(net71),
    .B(_0994_),
    .CO(_0995_),
    .S(_0996_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2520_ (.A(net70),
    .B(_0997_),
    .CO(_0998_),
    .S(_0999_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2521_ (.A(net69),
    .B(_1000_),
    .CO(_1001_),
    .S(_1002_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2522_ (.A(net68),
    .B(_1003_),
    .CO(_1004_),
    .S(_1005_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2523_ (.A(net93),
    .B(_1006_),
    .CO(_1007_),
    .S(_1008_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2524_ (.A(net92),
    .B(_1009_),
    .CO(_1010_),
    .S(_1011_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2525_ (.A(net91),
    .B(_1012_),
    .CO(_1013_),
    .S(_1014_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2526_ (.A(net90),
    .B(_1015_),
    .CO(_1016_),
    .S(_1017_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2527_ (.A(net88),
    .B(_1018_),
    .CO(_1019_),
    .S(_1020_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2528_ (.A(net87),
    .B(_1021_),
    .CO(_1022_),
    .S(_1023_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2529_ (.A(net86),
    .B(_1024_),
    .CO(_1025_),
    .S(_1026_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2530_ (.A(net85),
    .B(_1027_),
    .CO(_1028_),
    .S(_1029_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2531_ (.A(net84),
    .B(_1030_),
    .CO(_1031_),
    .S(_1032_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2532_ (.A(net83),
    .B(_1033_),
    .CO(_1034_),
    .S(_1035_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2533_ (.A(net82),
    .B(_1036_),
    .CO(_1037_),
    .S(_1038_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2534_ (.A(net81),
    .B(_1039_),
    .CO(_1040_),
    .S(_1041_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2535_ (.A(net80),
    .B(_1042_),
    .CO(_1043_),
    .S(_1044_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2536_ (.A(net79),
    .B(_1045_),
    .CO(_1046_),
    .S(_1047_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2537_ (.A(net77),
    .B(_1048_),
    .CO(_1049_),
    .S(_1050_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2538_ (.A(net76),
    .B(_1051_),
    .CO(_1052_),
    .S(_1053_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2539_ (.A(net36),
    .B(_1054_),
    .CO(_1055_),
    .S(_1056_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2540_ (.A(net35),
    .B(_1057_),
    .CO(_1058_),
    .S(_1059_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2541_ (.A(net34),
    .B(_1060_),
    .CO(_1061_),
    .S(_1062_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2542_ (.A(net33),
    .B(_1063_),
    .CO(_1064_),
    .S(_1065_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2543_ (.A(net32),
    .B(_1066_),
    .CO(_1067_),
    .S(_1068_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2544_ (.A(net31),
    .B(_1069_),
    .CO(_1070_),
    .S(_1071_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2545_ (.A(net30),
    .B(_1072_),
    .CO(_1073_),
    .S(_1074_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2546_ (.A(net29),
    .B(_1075_),
    .CO(_1076_),
    .S(_1077_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2547_ (.A(net27),
    .B(_1078_),
    .CO(_1079_),
    .S(_1080_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2548_ (.A(net26),
    .B(_1081_),
    .CO(_1082_),
    .S(_1083_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2549_ (.A(net25),
    .B(_1084_),
    .CO(_1085_),
    .S(_1086_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2550_ (.A(net24),
    .B(_1087_),
    .CO(_1088_),
    .S(_1089_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2551_ (.A(net23),
    .B(_1090_),
    .CO(_1091_),
    .S(_1092_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2552_ (.A(net22),
    .B(_1093_),
    .CO(_1094_),
    .S(_1095_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2553_ (.A(net21),
    .B(_1096_),
    .CO(_1097_),
    .S(_1098_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2554_ (.A(net20),
    .B(_1099_),
    .CO(_1100_),
    .S(_1101_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2555_ (.A(net19),
    .B(_1102_),
    .CO(_1103_),
    .S(_1104_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2556_ (.A(net18),
    .B(_1105_),
    .CO(_1106_),
    .S(_1107_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2557_ (.A(net16),
    .B(_1108_),
    .CO(_1109_),
    .S(_1110_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2558_ (.A(net15),
    .B(_1111_),
    .CO(_1112_),
    .S(_1113_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2559_ (.A(net14),
    .B(_1114_),
    .CO(_1115_),
    .S(_1116_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2560_ (.A(net13),
    .B(_1117_),
    .CO(_1118_),
    .S(_1119_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2561_ (.A(net12),
    .B(_1120_),
    .CO(_1121_),
    .S(_1122_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2562_ (.A(net11),
    .B(_1123_),
    .CO(_1124_),
    .S(_1125_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2563_ (.A(net10),
    .B(_1126_),
    .CO(_1127_),
    .S(_1128_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2564_ (.A(net9),
    .B(_1129_),
    .CO(_1130_),
    .S(_1131_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2565_ (.A(net8),
    .B(_1132_),
    .CO(_1133_),
    .S(_1134_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2566_ (.A(net7),
    .B(_1135_),
    .CO(_1136_),
    .S(_1137_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2567_ (.A(net132),
    .B(_1138_),
    .CO(_1139_),
    .S(_1140_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2568_ (.A(net131),
    .B(_1141_),
    .CO(_1142_),
    .S(_1143_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2569_ (.A(\transfer_count[3][0] ),
    .B(\transfer_count[3][1] ),
    .CO(_1144_),
    .S(_1145_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2570_ (.A(net130),
    .B(_1146_),
    .CO(_1147_),
    .S(_1148_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2571_ (.A(_1149_),
    .B(_1150_),
    .CO(_1151_),
    .S(_1152_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2572_ (.A(_1153_),
    .B(_1154_),
    .CO(_1155_),
    .S(_1156_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2573_ (.A(\transfer_count[0][0] ),
    .B(\transfer_count[0][1] ),
    .CO(_1157_),
    .S(_1158_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2574_ (.A(net45),
    .B(_1159_),
    .CO(_1160_),
    .S(_1161_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2575_ (.A(net67),
    .B(_1162_),
    .CO(_1163_),
    .S(_1164_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2576_ (.A(net56),
    .B(_1165_),
    .CO(_1166_),
    .S(_1167_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2577_ (.A(net111),
    .B(_1168_),
    .CO(_1169_),
    .S(_1170_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2578_ (.A(net100),
    .B(_1171_),
    .CO(_1172_),
    .S(_1173_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2579_ (.A(net89),
    .B(_1174_),
    .CO(_1175_),
    .S(_1176_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2580_ (.A(net78),
    .B(_1177_),
    .CO(_1178_),
    .S(_1179_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2581_ (.A(net40),
    .B(_1180_),
    .CO(_1181_),
    .S(_1182_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2582_ (.A(net39),
    .B(_1183_),
    .CO(_1184_),
    .S(_1185_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2583_ (.A(net38),
    .B(_1186_),
    .CO(_1187_),
    .S(_1188_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2584_ (.A(net37),
    .B(_1189_),
    .CO(_1190_),
    .S(_1191_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2585_ (.A(net28),
    .B(_1192_),
    .CO(_1193_),
    .S(_1194_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2586_ (.A(net17),
    .B(_1195_),
    .CO(_1196_),
    .S(_1197_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2587_ (.A(net133),
    .B(_1198_),
    .CO(_1199_),
    .S(_1200_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2588_ (.A(net122),
    .B(_1201_),
    .CO(_1202_),
    .S(_1203_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2589_ (.A(net58),
    .B(_1204_),
    .CO(_1205_),
    .S(_1206_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2590_ (.A(net57),
    .B(_1207_),
    .CO(_1208_),
    .S(_1209_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2591_ (.A(net55),
    .B(_1210_),
    .CO(_1211_),
    .S(_1212_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2592_ (.A(net54),
    .B(_1213_),
    .CO(_1214_),
    .S(_1215_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2593_ (.A(net53),
    .B(_1216_),
    .CO(_1217_),
    .S(_1218_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2594_ (.A(net52),
    .B(_1219_),
    .CO(_1220_),
    .S(_1221_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2595_ (.A(net51),
    .B(_1222_),
    .CO(_1223_),
    .S(_1224_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2596_ (.A(net50),
    .B(_1225_),
    .CO(_1226_),
    .S(_1227_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2597_ (.A(net49),
    .B(_1228_),
    .CO(_1229_),
    .S(_1230_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2598_ (.A(net48),
    .B(_1231_),
    .CO(_1232_),
    .S(_1233_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2599_ (.A(net47),
    .B(_1234_),
    .CO(_1235_),
    .S(_1236_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2600_ (.A(net46),
    .B(_1237_),
    .CO(_1238_),
    .S(_1239_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2601_ (.A(net44),
    .B(_1240_),
    .CO(_1241_),
    .S(_1242_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2602_ (.A(net43),
    .B(_1243_),
    .CO(_1244_),
    .S(_1245_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2603_ (.A(net42),
    .B(_1246_),
    .CO(_1247_),
    .S(_1248_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2604_ (.A(net41),
    .B(_1249_),
    .CO(_1250_),
    .S(_1251_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2605_ (.A(_1252_),
    .B(_1253_),
    .CO(_1254_),
    .S(_1255_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2606_ (.A(\active_channel_count[0] ),
    .B(\active_channel_count[1] ),
    .CO(_1256_),
    .S(_1257_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2607_ (.A(net128),
    .B(_1258_),
    .CO(_1259_),
    .S(_1260_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2608_ (.A(_1261_),
    .B(net127),
    .CO(_1262_),
    .S(_1263_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2609_ (.A(_1264_),
    .B(net126),
    .CO(_1265_),
    .S(_1266_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2610_ (.A(net125),
    .B(_1267_),
    .CO(_1268_),
    .S(_1269_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2611_ (.A(_1270_),
    .B(net124),
    .CO(_1271_),
    .S(_1272_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2612_ (.A(_1273_),
    .B(net123),
    .CO(_1274_),
    .S(_1275_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2613_ (.A(net121),
    .B(_1276_),
    .CO(_1277_),
    .S(_1278_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2614_ (.A(net120),
    .B(_1279_),
    .CO(_1280_),
    .S(_1281_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2615_ (.A(net119),
    .B(_1282_),
    .CO(_1283_),
    .S(_1284_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2616_ (.A(net118),
    .B(_1285_),
    .CO(_1286_),
    .S(_1287_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2617_ (.A(net117),
    .B(_1288_),
    .CO(_1289_),
    .S(_1290_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2618_ (.A(net116),
    .B(_1291_),
    .CO(_1292_),
    .S(_1293_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2619_ (.A(net115),
    .B(_1294_),
    .CO(_1295_),
    .S(_1296_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2620_ (.A(net114),
    .B(_1297_),
    .CO(_1298_),
    .S(_1299_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2621_ (.A(net113),
    .B(_1300_),
    .CO(_1301_),
    .S(_1302_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2622_ (.A(net112),
    .B(_1303_),
    .CO(_1304_),
    .S(_1305_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2623_ (.A(net110),
    .B(_1306_),
    .CO(_1307_),
    .S(_1308_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2624_ (.A(net109),
    .B(_1309_),
    .CO(_1310_),
    .S(_1311_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2625_ (.A(net108),
    .B(_1312_),
    .CO(_1313_),
    .S(_1314_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2626_ (.A(net107),
    .B(_1315_),
    .CO(_1316_),
    .S(_1317_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2627_ (.A(net106),
    .B(_1318_),
    .CO(_1319_),
    .S(_1320_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2628_ (.A(net105),
    .B(_1321_),
    .CO(_1322_),
    .S(_1323_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2629_ (.A(net104),
    .B(_1324_),
    .CO(_1325_),
    .S(_1326_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2630_ (.A(net103),
    .B(_1327_),
    .CO(_1328_),
    .S(_1329_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2631_ (.A(net102),
    .B(_1330_),
    .CO(_1331_),
    .S(_1332_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2632_ (.A(net101),
    .B(_1333_),
    .CO(_1334_),
    .S(_1335_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2633_ (.A(net99),
    .B(_1336_),
    .CO(_1337_),
    .S(_1338_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2634_ (.A(net98),
    .B(_1339_),
    .CO(_1340_),
    .S(_1341_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2635_ (.A(net97),
    .B(_1342_),
    .CO(_1343_),
    .S(_1344_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2636_ (.A(net96),
    .B(_1345_),
    .CO(_1346_),
    .S(_1347_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2637_ (.A(\transfer_count[2][0] ),
    .B(\transfer_count[2][1] ),
    .CO(_1348_),
    .S(_1349_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2638_ (.A(net95),
    .B(_1350_),
    .CO(_1351_),
    .S(_1352_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2639_ (.A(_1353_),
    .B(_1354_),
    .CO(_1355_),
    .S(_1356_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2640_ (.A(_1357_),
    .B(_1358_),
    .CO(_1359_),
    .S(_1360_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2641_ (.A(\transfer_count[1][0] ),
    .B(\transfer_count[1][1] ),
    .CO(_1361_),
    .S(_1362_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2642_ (.A(net60),
    .B(_1363_),
    .CO(_1364_),
    .S(_1365_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2643_ (.A(net62),
    .B(_1366_),
    .CO(_1367_),
    .S(_1368_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2644_ (.A(net61),
    .B(_1369_),
    .CO(_1370_),
    .S(_1371_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2645_ (.A(net66),
    .B(_1372_),
    .CO(_1373_),
    .S(_1374_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2646_ (.A(net65),
    .B(_1375_),
    .CO(_1376_),
    .S(_1377_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2647_ (.A(net64),
    .B(_1378_),
    .CO(_1379_),
    .S(_1380_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2648_ (.A(net63),
    .B(_1381_),
    .CO(_1382_),
    .S(_1383_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2650_ (.I(net175),
    .Z(debug_channel_state[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2651_ (.I(net176),
    .Z(debug_channel_state[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2652_ (.I(net177),
    .Z(debug_channel_state[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2653_ (.I(net178),
    .Z(debug_channel_state[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2654_ (.I(net179),
    .Z(debug_channel_state[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2655_ (.I(net180),
    .Z(debug_channel_state[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2656_ (.I(net181),
    .Z(debug_channel_state[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2657_ (.I(net182),
    .Z(debug_channel_state[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2658_ (.I(net183),
    .Z(debug_channel_state[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2659_ (.I(net184),
    .Z(debug_channel_state[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2660_ (.I(net185),
    .Z(debug_channel_state[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2661_ (.I(net186),
    .Z(debug_channel_state[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2662_ (.I(net187),
    .Z(debug_transfer_count[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2663_ (.I(net188),
    .Z(debug_transfer_count[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2664_ (.I(net189),
    .Z(debug_transfer_count[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2665_ (.I(net190),
    .Z(debug_transfer_count[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2666_ (.I(net191),
    .Z(debug_transfer_count[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2667_ (.I(net192),
    .Z(debug_transfer_count[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2668_ (.I(net193),
    .Z(debug_transfer_count[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2669_ (.I(net194),
    .Z(debug_transfer_count[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2670_ (.I(net195),
    .Z(debug_transfer_count[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2671_ (.I(net196),
    .Z(debug_transfer_count[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2672_ (.I(net197),
    .Z(debug_transfer_count[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2673_ (.I(net198),
    .Z(debug_transfer_count[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2674_ (.I(net199),
    .Z(debug_transfer_count[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2675_ (.I(net200),
    .Z(debug_transfer_count[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2676_ (.I(net201),
    .Z(debug_transfer_count[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2677_ (.I(net202),
    .Z(debug_transfer_count[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2678_ (.I(net203),
    .Z(debug_transfer_count[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2679_ (.I(net204),
    .Z(debug_transfer_count[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2680_ (.I(net205),
    .Z(debug_transfer_count[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2681_ (.I(net206),
    .Z(debug_transfer_count[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2682_ (.I(net207),
    .Z(debug_transfer_count[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2683_ (.I(net208),
    .Z(debug_transfer_count[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2684_ (.I(net209),
    .Z(debug_transfer_count[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2685_ (.I(net210),
    .Z(debug_transfer_count[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2686_ (.I(net211),
    .Z(debug_transfer_count[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2687_ (.I(net212),
    .Z(debug_transfer_count[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2688_ (.I(net213),
    .Z(debug_transfer_count[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2689_ (.I(net214),
    .Z(debug_transfer_count[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2690_ (.I(net215),
    .Z(debug_transfer_count[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2691_ (.I(net216),
    .Z(debug_transfer_count[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2692_ (.I(net217),
    .Z(debug_transfer_count[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2693_ (.I(net218),
    .Z(debug_transfer_count[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2694_ (.I(net219),
    .Z(debug_transfer_count[32]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2695_ (.I(net220),
    .Z(debug_transfer_count[33]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2696_ (.I(net221),
    .Z(debug_transfer_count[34]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2697_ (.I(net222),
    .Z(debug_transfer_count[35]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2698_ (.I(net223),
    .Z(debug_transfer_count[36]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2699_ (.I(net224),
    .Z(debug_transfer_count[37]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2700_ (.I(net225),
    .Z(debug_transfer_count[38]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2701_ (.I(net226),
    .Z(debug_transfer_count[39]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2702_ (.I(net227),
    .Z(debug_transfer_count[40]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2703_ (.I(net228),
    .Z(debug_transfer_count[41]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2704_ (.I(net229),
    .Z(debug_transfer_count[42]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2705_ (.I(net230),
    .Z(debug_transfer_count[43]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2706_ (.I(net231),
    .Z(debug_transfer_count[44]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2707_ (.I(net232),
    .Z(debug_transfer_count[45]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2708_ (.I(net233),
    .Z(debug_transfer_count[46]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2709_ (.I(net234),
    .Z(debug_transfer_count[47]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2710_ (.I(net235),
    .Z(debug_transfer_count[48]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2711_ (.I(net236),
    .Z(debug_transfer_count[49]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2712_ (.I(net237),
    .Z(debug_transfer_count[50]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2713_ (.I(net238),
    .Z(debug_transfer_count[51]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2714_ (.I(net239),
    .Z(debug_transfer_count[52]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2715_ (.I(net240),
    .Z(debug_transfer_count[53]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2716_ (.I(net241),
    .Z(debug_transfer_count[54]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2717_ (.I(net242),
    .Z(debug_transfer_count[55]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2718_ (.I(net243),
    .Z(debug_transfer_count[56]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2719_ (.I(net244),
    .Z(debug_transfer_count[57]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2720_ (.I(net245),
    .Z(debug_transfer_count[58]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2721_ (.I(net246),
    .Z(debug_transfer_count[59]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2722_ (.I(net247),
    .Z(debug_transfer_count[60]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2723_ (.I(net248),
    .Z(debug_transfer_count[61]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2724_ (.I(net249),
    .Z(debug_transfer_count[62]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2725_ (.I(net250),
    .Z(debug_transfer_count[63]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2726_ (.I(net251),
    .Z(debug_transfer_count[64]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2727_ (.I(net252),
    .Z(debug_transfer_count[65]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2728_ (.I(net253),
    .Z(debug_transfer_count[66]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2729_ (.I(net254),
    .Z(debug_transfer_count[67]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2730_ (.I(net255),
    .Z(debug_transfer_count[68]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2731_ (.I(net256),
    .Z(debug_transfer_count[69]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2732_ (.I(net257),
    .Z(debug_transfer_count[70]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2733_ (.I(net258),
    .Z(debug_transfer_count[71]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2734_ (.I(net259),
    .Z(debug_transfer_count[72]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2735_ (.I(net260),
    .Z(debug_transfer_count[73]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2736_ (.I(net261),
    .Z(debug_transfer_count[74]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2737_ (.I(net262),
    .Z(debug_transfer_count[75]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2738_ (.I(net263),
    .Z(debug_transfer_count[76]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2739_ (.I(net264),
    .Z(debug_transfer_count[77]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2740_ (.I(net265),
    .Z(debug_transfer_count[78]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2741_ (.I(net266),
    .Z(debug_transfer_count[79]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2742_ (.I(net267),
    .Z(debug_transfer_count[80]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2743_ (.I(net268),
    .Z(debug_transfer_count[81]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2744_ (.I(net269),
    .Z(debug_transfer_count[82]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2745_ (.I(net270),
    .Z(debug_transfer_count[83]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2746_ (.I(net271),
    .Z(debug_transfer_count[84]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2747_ (.I(net272),
    .Z(debug_transfer_count[85]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2748_ (.I(net273),
    .Z(debug_transfer_count[86]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2749_ (.I(net274),
    .Z(debug_transfer_count[87]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2750_ (.I(net275),
    .Z(debug_transfer_count[88]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2751_ (.I(net276),
    .Z(debug_transfer_count[89]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2752_ (.I(net277),
    .Z(debug_transfer_count[90]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2753_ (.I(net278),
    .Z(debug_transfer_count[91]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2754_ (.I(net279),
    .Z(debug_transfer_count[92]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2755_ (.I(net280),
    .Z(debug_transfer_count[93]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2756_ (.I(net281),
    .Z(debug_transfer_count[94]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2757_ (.I(net282),
    .Z(debug_transfer_count[95]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2758_ (.I(net283),
    .Z(debug_transfer_count[96]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2759_ (.I(net284),
    .Z(debug_transfer_count[97]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2760_ (.I(net285),
    .Z(debug_transfer_count[98]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2761_ (.I(net286),
    .Z(debug_transfer_count[99]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2762_ (.I(net287),
    .Z(debug_transfer_count[100]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2763_ (.I(net288),
    .Z(debug_transfer_count[101]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2764_ (.I(net289),
    .Z(debug_transfer_count[102]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2765_ (.I(net290),
    .Z(debug_transfer_count[103]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2766_ (.I(net291),
    .Z(debug_transfer_count[104]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2767_ (.I(net292),
    .Z(debug_transfer_count[105]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2768_ (.I(net293),
    .Z(debug_transfer_count[106]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2769_ (.I(net294),
    .Z(debug_transfer_count[107]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2770_ (.I(net295),
    .Z(debug_transfer_count[108]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2771_ (.I(net296),
    .Z(debug_transfer_count[109]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2772_ (.I(net297),
    .Z(debug_transfer_count[110]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2773_ (.I(net298),
    .Z(debug_transfer_count[111]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2774_ (.I(net299),
    .Z(debug_transfer_count[112]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2775_ (.I(net300),
    .Z(debug_transfer_count[113]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2776_ (.I(net301),
    .Z(debug_transfer_count[114]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2777_ (.I(net302),
    .Z(debug_transfer_count[115]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2778_ (.I(net303),
    .Z(debug_transfer_count[116]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2779_ (.I(net304),
    .Z(debug_transfer_count[117]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2780_ (.I(net305),
    .Z(debug_transfer_count[118]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2781_ (.I(net306),
    .Z(debug_transfer_count[119]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2782_ (.I(net307),
    .Z(debug_transfer_count[120]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2783_ (.I(net308),
    .Z(debug_transfer_count[121]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2784_ (.I(net309),
    .Z(debug_transfer_count[122]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2785_ (.I(net310),
    .Z(debug_transfer_count[123]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2786_ (.I(net311),
    .Z(debug_transfer_count[124]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2787_ (.I(net312),
    .Z(debug_transfer_count[125]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2788_ (.I(net313),
    .Z(debug_transfer_count[126]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2789_ (.I(net314),
    .Z(debug_transfer_count[127]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2790_ (.I(net315),
    .Z(dst_addr[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2791_ (.I(net316),
    .Z(dst_addr[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2792_ (.I(net317),
    .Z(dst_addr[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2793_ (.I(net318),
    .Z(dst_addr[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2794_ (.I(net319),
    .Z(dst_addr[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2795_ (.I(net320),
    .Z(dst_addr[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2796_ (.I(net321),
    .Z(dst_addr[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2797_ (.I(net322),
    .Z(dst_addr[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2798_ (.I(net323),
    .Z(dst_addr[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2799_ (.I(net324),
    .Z(dst_addr[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2800_ (.I(net325),
    .Z(dst_addr[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2801_ (.I(net326),
    .Z(dst_addr[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2802_ (.I(net327),
    .Z(dst_addr[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2803_ (.I(net328),
    .Z(dst_addr[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2804_ (.I(net329),
    .Z(dst_addr[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2805_ (.I(net330),
    .Z(dst_addr[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2806_ (.I(net331),
    .Z(dst_addr[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2807_ (.I(net332),
    .Z(dst_addr[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2808_ (.I(net333),
    .Z(dst_addr[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2809_ (.I(net334),
    .Z(dst_addr[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2810_ (.I(net335),
    .Z(dst_addr[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2811_ (.I(net336),
    .Z(dst_addr[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2812_ (.I(net337),
    .Z(dst_addr[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2813_ (.I(net338),
    .Z(dst_addr[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2814_ (.I(net339),
    .Z(dst_addr[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2815_ (.I(net340),
    .Z(dst_addr[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2816_ (.I(net341),
    .Z(dst_addr[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2817_ (.I(net342),
    .Z(dst_addr[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2818_ (.I(net343),
    .Z(dst_addr[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2819_ (.I(net344),
    .Z(dst_addr[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2820_ (.I(net345),
    .Z(dst_addr[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2821_ (.I(net346),
    .Z(dst_addr[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2822_ (.I(net347),
    .Z(dst_addr[32]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2823_ (.I(net348),
    .Z(dst_addr[33]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2824_ (.I(net349),
    .Z(dst_addr[34]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2825_ (.I(net350),
    .Z(dst_addr[35]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2826_ (.I(net351),
    .Z(dst_addr[36]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2827_ (.I(net352),
    .Z(dst_addr[37]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2828_ (.I(net353),
    .Z(dst_addr[38]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2829_ (.I(net354),
    .Z(dst_addr[39]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2830_ (.I(net355),
    .Z(dst_addr[40]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2831_ (.I(net356),
    .Z(dst_addr[41]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2832_ (.I(net357),
    .Z(dst_addr[42]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2833_ (.I(net358),
    .Z(dst_addr[43]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2834_ (.I(net359),
    .Z(dst_addr[44]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2835_ (.I(net360),
    .Z(dst_addr[45]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2836_ (.I(net361),
    .Z(dst_addr[46]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2837_ (.I(net362),
    .Z(dst_addr[47]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2838_ (.I(net363),
    .Z(dst_addr[48]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2839_ (.I(net364),
    .Z(dst_addr[49]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2840_ (.I(net365),
    .Z(dst_addr[50]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2841_ (.I(net366),
    .Z(dst_addr[51]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2842_ (.I(net367),
    .Z(dst_addr[52]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2843_ (.I(net368),
    .Z(dst_addr[53]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2844_ (.I(net369),
    .Z(dst_addr[54]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2845_ (.I(net370),
    .Z(dst_addr[55]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2846_ (.I(net371),
    .Z(dst_addr[56]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2847_ (.I(net372),
    .Z(dst_addr[57]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2848_ (.I(net373),
    .Z(dst_addr[58]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2849_ (.I(net374),
    .Z(dst_addr[59]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2850_ (.I(net375),
    .Z(dst_addr[60]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2851_ (.I(net376),
    .Z(dst_addr[61]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2852_ (.I(net377),
    .Z(dst_addr[62]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2853_ (.I(net378),
    .Z(dst_addr[63]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2854_ (.I(net379),
    .Z(dst_addr[64]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2855_ (.I(net380),
    .Z(dst_addr[65]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2856_ (.I(net381),
    .Z(dst_addr[66]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2857_ (.I(net382),
    .Z(dst_addr[67]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2858_ (.I(net383),
    .Z(dst_addr[68]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2859_ (.I(net384),
    .Z(dst_addr[69]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2860_ (.I(net385),
    .Z(dst_addr[70]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2861_ (.I(net386),
    .Z(dst_addr[71]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2862_ (.I(net387),
    .Z(dst_addr[72]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2863_ (.I(net388),
    .Z(dst_addr[73]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2864_ (.I(net389),
    .Z(dst_addr[74]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2865_ (.I(net390),
    .Z(dst_addr[75]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2866_ (.I(net391),
    .Z(dst_addr[76]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2867_ (.I(net392),
    .Z(dst_addr[77]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2868_ (.I(net393),
    .Z(dst_addr[78]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2869_ (.I(net394),
    .Z(dst_addr[79]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2870_ (.I(net395),
    .Z(dst_addr[80]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2871_ (.I(net396),
    .Z(dst_addr[81]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2872_ (.I(net397),
    .Z(dst_addr[82]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2873_ (.I(net398),
    .Z(dst_addr[83]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2874_ (.I(net399),
    .Z(dst_addr[84]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2875_ (.I(net400),
    .Z(dst_addr[85]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2876_ (.I(net401),
    .Z(dst_addr[86]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2877_ (.I(net402),
    .Z(dst_addr[87]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2878_ (.I(net403),
    .Z(dst_addr[88]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2879_ (.I(net404),
    .Z(dst_addr[89]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2880_ (.I(net405),
    .Z(dst_addr[90]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2881_ (.I(net406),
    .Z(dst_addr[91]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2882_ (.I(net407),
    .Z(dst_addr[92]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2883_ (.I(net408),
    .Z(dst_addr[93]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2884_ (.I(net409),
    .Z(dst_addr[94]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2885_ (.I(net410),
    .Z(dst_addr[95]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2886_ (.I(net411),
    .Z(dst_addr[96]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2887_ (.I(net412),
    .Z(dst_addr[97]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2888_ (.I(net413),
    .Z(dst_addr[98]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2889_ (.I(net414),
    .Z(dst_addr[99]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2890_ (.I(net415),
    .Z(dst_addr[100]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2891_ (.I(net416),
    .Z(dst_addr[101]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2892_ (.I(net417),
    .Z(dst_addr[102]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2893_ (.I(net418),
    .Z(dst_addr[103]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2894_ (.I(net419),
    .Z(dst_addr[104]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2895_ (.I(net420),
    .Z(dst_addr[105]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2896_ (.I(net421),
    .Z(dst_addr[106]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2897_ (.I(net422),
    .Z(dst_addr[107]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2898_ (.I(net423),
    .Z(dst_addr[108]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2899_ (.I(net424),
    .Z(dst_addr[109]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2900_ (.I(net425),
    .Z(dst_addr[110]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2901_ (.I(net426),
    .Z(dst_addr[111]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2902_ (.I(net427),
    .Z(dst_addr[112]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2903_ (.I(net428),
    .Z(dst_addr[113]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2904_ (.I(net429),
    .Z(dst_addr[114]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2905_ (.I(net430),
    .Z(dst_addr[115]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2906_ (.I(net431),
    .Z(dst_addr[116]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2907_ (.I(net432),
    .Z(dst_addr[117]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2908_ (.I(net433),
    .Z(dst_addr[118]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2909_ (.I(net434),
    .Z(dst_addr[119]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2910_ (.I(net435),
    .Z(dst_addr[120]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2911_ (.I(net436),
    .Z(dst_addr[121]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2912_ (.I(net437),
    .Z(dst_addr[122]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2913_ (.I(net438),
    .Z(dst_addr[123]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2914_ (.I(net439),
    .Z(dst_addr[124]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2915_ (.I(net440),
    .Z(dst_addr[125]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2916_ (.I(net441),
    .Z(dst_addr[126]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2917_ (.I(net442),
    .Z(dst_addr[127]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2918_ (.I(net443),
    .Z(dst_wdata[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2919_ (.I(net444),
    .Z(dst_wdata[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2920_ (.I(net445),
    .Z(dst_wdata[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2921_ (.I(net446),
    .Z(dst_wdata[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2922_ (.I(net447),
    .Z(dst_wdata[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2923_ (.I(net448),
    .Z(dst_wdata[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2924_ (.I(net449),
    .Z(dst_wdata[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2925_ (.I(net450),
    .Z(dst_wdata[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2926_ (.I(net451),
    .Z(dst_wdata[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2927_ (.I(net452),
    .Z(dst_wdata[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2928_ (.I(net453),
    .Z(dst_wdata[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2929_ (.I(net454),
    .Z(dst_wdata[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2930_ (.I(net455),
    .Z(dst_wdata[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2931_ (.I(net456),
    .Z(dst_wdata[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2932_ (.I(net457),
    .Z(dst_wdata[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2933_ (.I(net458),
    .Z(dst_wdata[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2934_ (.I(net459),
    .Z(dst_wdata[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2935_ (.I(net460),
    .Z(dst_wdata[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2936_ (.I(net461),
    .Z(dst_wdata[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2937_ (.I(net462),
    .Z(dst_wdata[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2938_ (.I(net463),
    .Z(dst_wdata[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2939_ (.I(net464),
    .Z(dst_wdata[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2940_ (.I(net465),
    .Z(dst_wdata[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2941_ (.I(net466),
    .Z(dst_wdata[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2942_ (.I(net467),
    .Z(dst_wdata[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2943_ (.I(net468),
    .Z(dst_wdata[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2944_ (.I(net469),
    .Z(dst_wdata[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2945_ (.I(net470),
    .Z(dst_wdata[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2946_ (.I(net471),
    .Z(dst_wdata[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2947_ (.I(net472),
    .Z(dst_wdata[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2948_ (.I(net473),
    .Z(dst_wdata[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2949_ (.I(net474),
    .Z(dst_wdata[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2950_ (.I(net475),
    .Z(dst_wdata[32]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2951_ (.I(net476),
    .Z(dst_wdata[33]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2952_ (.I(net477),
    .Z(dst_wdata[34]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2953_ (.I(net478),
    .Z(dst_wdata[35]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2954_ (.I(net479),
    .Z(dst_wdata[36]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2955_ (.I(net480),
    .Z(dst_wdata[37]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2956_ (.I(net481),
    .Z(dst_wdata[38]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2957_ (.I(net482),
    .Z(dst_wdata[39]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2958_ (.I(net483),
    .Z(dst_wdata[40]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2959_ (.I(net484),
    .Z(dst_wdata[41]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2960_ (.I(net485),
    .Z(dst_wdata[42]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2961_ (.I(net486),
    .Z(dst_wdata[43]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2962_ (.I(net487),
    .Z(dst_wdata[44]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2963_ (.I(net488),
    .Z(dst_wdata[45]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2964_ (.I(net489),
    .Z(dst_wdata[46]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2965_ (.I(net490),
    .Z(dst_wdata[47]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2966_ (.I(net491),
    .Z(dst_wdata[48]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2967_ (.I(net492),
    .Z(dst_wdata[49]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2968_ (.I(net493),
    .Z(dst_wdata[50]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2969_ (.I(net494),
    .Z(dst_wdata[51]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2970_ (.I(net495),
    .Z(dst_wdata[52]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2971_ (.I(net496),
    .Z(dst_wdata[53]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2972_ (.I(net497),
    .Z(dst_wdata[54]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2973_ (.I(net498),
    .Z(dst_wdata[55]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2974_ (.I(net499),
    .Z(dst_wdata[56]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2975_ (.I(net500),
    .Z(dst_wdata[57]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2976_ (.I(net501),
    .Z(dst_wdata[58]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2977_ (.I(net502),
    .Z(dst_wdata[59]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2978_ (.I(net503),
    .Z(dst_wdata[60]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2979_ (.I(net504),
    .Z(dst_wdata[61]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2980_ (.I(net505),
    .Z(dst_wdata[62]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2981_ (.I(net506),
    .Z(dst_wdata[63]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2982_ (.I(net507),
    .Z(dst_wdata[64]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2983_ (.I(net508),
    .Z(dst_wdata[65]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2984_ (.I(net509),
    .Z(dst_wdata[66]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2985_ (.I(net510),
    .Z(dst_wdata[67]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2986_ (.I(net511),
    .Z(dst_wdata[68]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2987_ (.I(net512),
    .Z(dst_wdata[69]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2988_ (.I(net513),
    .Z(dst_wdata[70]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2989_ (.I(net514),
    .Z(dst_wdata[71]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2990_ (.I(net515),
    .Z(dst_wdata[72]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2991_ (.I(net516),
    .Z(dst_wdata[73]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2992_ (.I(net517),
    .Z(dst_wdata[74]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2993_ (.I(net518),
    .Z(dst_wdata[75]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2994_ (.I(net519),
    .Z(dst_wdata[76]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2995_ (.I(net520),
    .Z(dst_wdata[77]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2996_ (.I(net521),
    .Z(dst_wdata[78]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2997_ (.I(net522),
    .Z(dst_wdata[79]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2998_ (.I(net523),
    .Z(dst_wdata[80]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _2999_ (.I(net524),
    .Z(dst_wdata[81]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3000_ (.I(net525),
    .Z(dst_wdata[82]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3001_ (.I(net526),
    .Z(dst_wdata[83]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3002_ (.I(net527),
    .Z(dst_wdata[84]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3003_ (.I(net528),
    .Z(dst_wdata[85]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3004_ (.I(net529),
    .Z(dst_wdata[86]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3005_ (.I(net530),
    .Z(dst_wdata[87]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3006_ (.I(net531),
    .Z(dst_wdata[88]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3007_ (.I(net532),
    .Z(dst_wdata[89]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3008_ (.I(net533),
    .Z(dst_wdata[90]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3009_ (.I(net534),
    .Z(dst_wdata[91]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3010_ (.I(net535),
    .Z(dst_wdata[92]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3011_ (.I(net536),
    .Z(dst_wdata[93]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3012_ (.I(net537),
    .Z(dst_wdata[94]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3013_ (.I(net538),
    .Z(dst_wdata[95]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3014_ (.I(net539),
    .Z(dst_wdata[96]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3015_ (.I(net540),
    .Z(dst_wdata[97]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3016_ (.I(net541),
    .Z(dst_wdata[98]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3017_ (.I(net542),
    .Z(dst_wdata[99]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3018_ (.I(net543),
    .Z(dst_wdata[100]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3019_ (.I(net544),
    .Z(dst_wdata[101]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3020_ (.I(net545),
    .Z(dst_wdata[102]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3021_ (.I(net546),
    .Z(dst_wdata[103]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3022_ (.I(net547),
    .Z(dst_wdata[104]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3023_ (.I(net548),
    .Z(dst_wdata[105]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3024_ (.I(net549),
    .Z(dst_wdata[106]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3025_ (.I(net550),
    .Z(dst_wdata[107]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3026_ (.I(net551),
    .Z(dst_wdata[108]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3027_ (.I(net552),
    .Z(dst_wdata[109]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3028_ (.I(net553),
    .Z(dst_wdata[110]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3029_ (.I(net554),
    .Z(dst_wdata[111]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3030_ (.I(net555),
    .Z(dst_wdata[112]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3031_ (.I(net556),
    .Z(dst_wdata[113]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3032_ (.I(net557),
    .Z(dst_wdata[114]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3033_ (.I(net558),
    .Z(dst_wdata[115]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3034_ (.I(net559),
    .Z(dst_wdata[116]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3035_ (.I(net560),
    .Z(dst_wdata[117]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3036_ (.I(net561),
    .Z(dst_wdata[118]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3037_ (.I(net562),
    .Z(dst_wdata[119]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3038_ (.I(net563),
    .Z(dst_wdata[120]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3039_ (.I(net564),
    .Z(dst_wdata[121]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3040_ (.I(net565),
    .Z(dst_wdata[122]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3041_ (.I(net566),
    .Z(dst_wdata[123]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3042_ (.I(net567),
    .Z(dst_wdata[124]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3043_ (.I(net568),
    .Z(dst_wdata[125]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3044_ (.I(net569),
    .Z(dst_wdata[126]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3045_ (.I(net570),
    .Z(dst_wdata[127]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3046_ (.I(net571),
    .Z(dst_wstrb[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3047_ (.I(net572),
    .Z(dst_wstrb[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3048_ (.I(net573),
    .Z(dst_wstrb[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3049_ (.I(net574),
    .Z(dst_wstrb[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3050_ (.I(net575),
    .Z(dst_wstrb[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3051_ (.I(net576),
    .Z(dst_wstrb[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3052_ (.I(net577),
    .Z(dst_wstrb[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3053_ (.I(net578),
    .Z(dst_wstrb[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3054_ (.I(net579),
    .Z(dst_wstrb[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3055_ (.I(net580),
    .Z(dst_wstrb[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3056_ (.I(net581),
    .Z(dst_wstrb[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3057_ (.I(net582),
    .Z(dst_wstrb[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3058_ (.I(net583),
    .Z(dst_wstrb[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3059_ (.I(net584),
    .Z(dst_wstrb[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3060_ (.I(net585),
    .Z(dst_wstrb[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3061_ (.I(net586),
    .Z(dst_wstrb[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3062_ (.I(net587),
    .Z(src_addr[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3063_ (.I(net588),
    .Z(src_addr[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3064_ (.I(net589),
    .Z(src_addr[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3065_ (.I(net590),
    .Z(src_addr[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3066_ (.I(net591),
    .Z(src_addr[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3067_ (.I(net592),
    .Z(src_addr[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3068_ (.I(net593),
    .Z(src_addr[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3069_ (.I(net594),
    .Z(src_addr[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3070_ (.I(net595),
    .Z(src_addr[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3071_ (.I(net596),
    .Z(src_addr[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3072_ (.I(net597),
    .Z(src_addr[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3073_ (.I(net598),
    .Z(src_addr[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3074_ (.I(net599),
    .Z(src_addr[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3075_ (.I(net600),
    .Z(src_addr[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3076_ (.I(net601),
    .Z(src_addr[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3077_ (.I(net602),
    .Z(src_addr[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3078_ (.I(net603),
    .Z(src_addr[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3079_ (.I(net604),
    .Z(src_addr[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3080_ (.I(net605),
    .Z(src_addr[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3081_ (.I(net606),
    .Z(src_addr[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3082_ (.I(net607),
    .Z(src_addr[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3083_ (.I(net608),
    .Z(src_addr[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3084_ (.I(net609),
    .Z(src_addr[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3085_ (.I(net610),
    .Z(src_addr[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3086_ (.I(net611),
    .Z(src_addr[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3087_ (.I(net612),
    .Z(src_addr[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3088_ (.I(net613),
    .Z(src_addr[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3089_ (.I(net614),
    .Z(src_addr[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3090_ (.I(net615),
    .Z(src_addr[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3091_ (.I(net616),
    .Z(src_addr[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3092_ (.I(net617),
    .Z(src_addr[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3093_ (.I(net618),
    .Z(src_addr[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3094_ (.I(net619),
    .Z(src_addr[32]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3095_ (.I(net620),
    .Z(src_addr[33]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3096_ (.I(net621),
    .Z(src_addr[34]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3097_ (.I(net622),
    .Z(src_addr[35]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3098_ (.I(net623),
    .Z(src_addr[36]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3099_ (.I(net624),
    .Z(src_addr[37]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3100_ (.I(net625),
    .Z(src_addr[38]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3101_ (.I(net626),
    .Z(src_addr[39]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3102_ (.I(net627),
    .Z(src_addr[40]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3103_ (.I(net628),
    .Z(src_addr[41]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3104_ (.I(net629),
    .Z(src_addr[42]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3105_ (.I(net630),
    .Z(src_addr[43]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3106_ (.I(net631),
    .Z(src_addr[44]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3107_ (.I(net632),
    .Z(src_addr[45]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3108_ (.I(net633),
    .Z(src_addr[46]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3109_ (.I(net634),
    .Z(src_addr[47]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3110_ (.I(net635),
    .Z(src_addr[48]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3111_ (.I(net636),
    .Z(src_addr[49]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3112_ (.I(net637),
    .Z(src_addr[50]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3113_ (.I(net638),
    .Z(src_addr[51]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3114_ (.I(net639),
    .Z(src_addr[52]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3115_ (.I(net640),
    .Z(src_addr[53]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3116_ (.I(net641),
    .Z(src_addr[54]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3117_ (.I(net642),
    .Z(src_addr[55]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3118_ (.I(net643),
    .Z(src_addr[56]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3119_ (.I(net644),
    .Z(src_addr[57]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3120_ (.I(net645),
    .Z(src_addr[58]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3121_ (.I(net646),
    .Z(src_addr[59]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3122_ (.I(net647),
    .Z(src_addr[60]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3123_ (.I(net648),
    .Z(src_addr[61]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3124_ (.I(net649),
    .Z(src_addr[62]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3125_ (.I(net650),
    .Z(src_addr[63]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3126_ (.I(net651),
    .Z(src_addr[64]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3127_ (.I(net652),
    .Z(src_addr[65]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3128_ (.I(net653),
    .Z(src_addr[66]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3129_ (.I(net654),
    .Z(src_addr[67]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3130_ (.I(net655),
    .Z(src_addr[68]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3131_ (.I(net656),
    .Z(src_addr[69]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3132_ (.I(net657),
    .Z(src_addr[70]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3133_ (.I(net658),
    .Z(src_addr[71]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3134_ (.I(net659),
    .Z(src_addr[72]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3135_ (.I(net660),
    .Z(src_addr[73]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3136_ (.I(net661),
    .Z(src_addr[74]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3137_ (.I(net662),
    .Z(src_addr[75]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3138_ (.I(net663),
    .Z(src_addr[76]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3139_ (.I(net664),
    .Z(src_addr[77]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3140_ (.I(net665),
    .Z(src_addr[78]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3141_ (.I(net666),
    .Z(src_addr[79]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3142_ (.I(net667),
    .Z(src_addr[80]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3143_ (.I(net668),
    .Z(src_addr[81]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3144_ (.I(net669),
    .Z(src_addr[82]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3145_ (.I(net670),
    .Z(src_addr[83]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3146_ (.I(net671),
    .Z(src_addr[84]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3147_ (.I(net672),
    .Z(src_addr[85]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3148_ (.I(net673),
    .Z(src_addr[86]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3149_ (.I(net674),
    .Z(src_addr[87]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3150_ (.I(net675),
    .Z(src_addr[88]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3151_ (.I(net676),
    .Z(src_addr[89]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3152_ (.I(net677),
    .Z(src_addr[90]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3153_ (.I(net678),
    .Z(src_addr[91]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3154_ (.I(net679),
    .Z(src_addr[92]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3155_ (.I(net680),
    .Z(src_addr[93]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3156_ (.I(net681),
    .Z(src_addr[94]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3157_ (.I(net682),
    .Z(src_addr[95]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3158_ (.I(net683),
    .Z(src_addr[96]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3159_ (.I(net684),
    .Z(src_addr[97]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3160_ (.I(net685),
    .Z(src_addr[98]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3161_ (.I(net686),
    .Z(src_addr[99]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3162_ (.I(net687),
    .Z(src_addr[100]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3163_ (.I(net688),
    .Z(src_addr[101]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3164_ (.I(net689),
    .Z(src_addr[102]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3165_ (.I(net690),
    .Z(src_addr[103]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3166_ (.I(net691),
    .Z(src_addr[104]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3167_ (.I(net692),
    .Z(src_addr[105]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3168_ (.I(net693),
    .Z(src_addr[106]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3169_ (.I(net694),
    .Z(src_addr[107]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3170_ (.I(net695),
    .Z(src_addr[108]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3171_ (.I(net696),
    .Z(src_addr[109]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3172_ (.I(net697),
    .Z(src_addr[110]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3173_ (.I(net698),
    .Z(src_addr[111]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3174_ (.I(net699),
    .Z(src_addr[112]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3175_ (.I(net700),
    .Z(src_addr[113]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3176_ (.I(net701),
    .Z(src_addr[114]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3177_ (.I(net702),
    .Z(src_addr[115]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3178_ (.I(net703),
    .Z(src_addr[116]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3179_ (.I(net704),
    .Z(src_addr[117]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3180_ (.I(net705),
    .Z(src_addr[118]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3181_ (.I(net706),
    .Z(src_addr[119]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3182_ (.I(net707),
    .Z(src_addr[120]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3183_ (.I(net708),
    .Z(src_addr[121]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3184_ (.I(net709),
    .Z(src_addr[122]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3185_ (.I(net710),
    .Z(src_addr[123]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3186_ (.I(net711),
    .Z(src_addr[124]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3187_ (.I(net712),
    .Z(src_addr[125]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3188_ (.I(net713),
    .Z(src_addr[126]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _3189_ (.I(net714),
    .Z(src_addr[127]));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \active_channel_count[0]$_DFF_PN0_  (.D(_0000_),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(\active_channel_count[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \active_channel_count[1]$_DFF_PN0_  (.D(_0001_),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(\active_channel_count[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \active_channel_count[2]$_DFF_PN0_  (.D(_0002_),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(\active_channel_count[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \active_channel_count[3]$_DFF_PN0_  (.D(_0003_),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(\active_channel_count[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \channel_busy[0]$_DFF_PN0_  (.D(_0004_),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(net146));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \channel_busy[1]$_DFF_PN0_  (.D(_0005_),
    .RN(net1),
    .CLK(clknet_4_12_0_clk),
    .Q(net147));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \channel_busy[2]$_DFF_PN0_  (.D(_0006_),
    .RN(net1),
    .CLK(clknet_4_6_0_clk),
    .Q(net148));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \channel_busy[3]$_DFF_PN0_  (.D(_0007_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(net149));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \channel_done[0]$_DFF_PN0_  (.D(_1390_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(net150));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \channel_done[1]$_DFF_PN0_  (.D(_1388_),
    .RN(net1),
    .CLK(clknet_4_12_0_clk),
    .Q(net151));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \channel_done[2]$_DFF_PN0_  (.D(_1385_),
    .RN(net1),
    .CLK(clknet_4_6_0_clk),
    .Q(net152));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \channel_done[3]$_DFF_PN0_  (.D(_1387_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(net153));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \channel_error[0]$_DFF_PN0_  (.D(_0008_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(net154));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \channel_error[1]$_DFF_PN0_  (.D(_0009_),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(net155));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \channel_error[2]$_DFF_PN0_  (.D(_0010_),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(net156));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \channel_error[3]$_DFF_PN0_  (.D(_0011_),
    .RN(net1),
    .CLK(clknet_4_12_0_clk),
    .Q(net157));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \channel_state[0][0]$_DFF_PN0_  (.D(_0979_),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(\channel_state[0][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \channel_state[0][1]$_DFF_PN0_  (.D(_0980_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(\channel_state[0][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \channel_state[0][2]$_DFF_PN0_  (.D(_0981_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(\channel_state[0][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \channel_state[1][0]$_DFF_PN0_  (.D(_0976_),
    .RN(net1),
    .CLK(clknet_4_12_0_clk),
    .Q(\channel_state[1][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \channel_state[1][1]$_DFF_PN0_  (.D(_0977_),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(\channel_state[1][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \channel_state[1][2]$_DFF_PN0_  (.D(_0978_),
    .RN(net1),
    .CLK(clknet_4_12_0_clk),
    .Q(\channel_state[1][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \channel_state[2][0]$_DFF_PN0_  (.D(_0973_),
    .RN(net1),
    .CLK(clknet_4_6_0_clk),
    .Q(\channel_state[2][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \channel_state[2][1]$_DFF_PN0_  (.D(_0974_),
    .RN(net1),
    .CLK(clknet_4_6_0_clk),
    .Q(\channel_state[2][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \channel_state[2][2]$_DFF_PN0_  (.D(_0975_),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\channel_state[2][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \channel_state[3][0]$_DFF_PN0_  (.D(_0970_),
    .RN(net1),
    .CLK(clknet_4_12_0_clk),
    .Q(\channel_state[3][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \channel_state[3][1]$_DFF_PN0_  (.D(_0971_),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(\channel_state[3][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \channel_state[3][2]$_DFF_PN0_  (.D(_0972_),
    .RN(net1),
    .CLK(clknet_4_14_0_clk),
    .Q(\channel_state[3][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \debug_active_channels[0]$_DFF_PN0_  (.D(\active_channel_count[0] ),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(net158));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \debug_active_channels[1]$_DFF_PN0_  (.D(\active_channel_count[1] ),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(net159));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \debug_active_channels[2]$_DFF_PN0_  (.D(\active_channel_count[2] ),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(net160));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \debug_active_channels[3]$_DFF_PN0_  (.D(\active_channel_count[3] ),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(net161));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \debug_has_active_channels$_DFF_PN0_  (.D(_0012_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(net162));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_write[0]$_DFFE_PN0P_  (.D(_0141_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(net163));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_write[1]$_DFFE_PN0P_  (.D(_0142_),
    .RN(net1),
    .CLK(clknet_4_12_0_clk),
    .Q(net164));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_write[2]$_DFFE_PN0P_  (.D(_0143_),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(net165));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_write[3]$_DFFE_PN0P_  (.D(_0144_),
    .RN(net1),
    .CLK(clknet_4_14_0_clk),
    .Q(net166));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_read[0]$_DFF_PN0_  (.D(_0968_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(net167));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_read[1]$_DFF_PN0_  (.D(_0967_),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(net168));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_read[2]$_DFF_PN0_  (.D(_0966_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(net169));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_read[3]$_DFF_PN0_  (.D(_0969_),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(net170));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_rready[0]$_DFF_PN0_  (.D(_1391_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(net171));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_rready[1]$_DFF_PN0_  (.D(_1389_),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(net172));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_rready[2]$_DFF_PN0_  (.D(_1386_),
    .RN(net1),
    .CLK(clknet_4_6_0_clk),
    .Q(net173));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_rready[3]$_DFFE_PN0P_  (.D(_0145_),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(net174));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][0]$_DFF_PN0_  (.D(_0013_),
    .RN(net1),
    .CLK(clknet_4_1_0_clk),
    .Q(\transfer_count[0][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][10]$_DFF_PN0_  (.D(_0014_),
    .RN(net1),
    .CLK(clknet_4_1_0_clk),
    .Q(\transfer_count[0][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][11]$_DFF_PN0_  (.D(_0015_),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\transfer_count[0][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][12]$_DFF_PN0_  (.D(_0016_),
    .RN(net1),
    .CLK(clknet_4_1_0_clk),
    .Q(\transfer_count[0][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][13]$_DFF_PN0_  (.D(_0017_),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\transfer_count[0][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][14]$_DFF_PN0_  (.D(_0018_),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\transfer_count[0][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][15]$_DFF_PN0_  (.D(_0019_),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\transfer_count[0][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][16]$_DFF_PN0_  (.D(_0020_),
    .RN(net1),
    .CLK(clknet_4_3_0_clk),
    .Q(\transfer_count[0][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][17]$_DFF_PN0_  (.D(_0021_),
    .RN(net1),
    .CLK(clknet_4_3_0_clk),
    .Q(\transfer_count[0][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][18]$_DFF_PN0_  (.D(_0022_),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(\transfer_count[0][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][19]$_DFF_PN0_  (.D(_0023_),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(\transfer_count[0][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][1]$_DFF_PN0_  (.D(_0024_),
    .RN(net1),
    .CLK(clknet_4_1_0_clk),
    .Q(\transfer_count[0][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][20]$_DFF_PN0_  (.D(_0025_),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\transfer_count[0][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][21]$_DFF_PN0_  (.D(_0026_),
    .RN(net1),
    .CLK(clknet_4_3_0_clk),
    .Q(\transfer_count[0][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][22]$_DFF_PN0_  (.D(_0027_),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\transfer_count[0][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][23]$_DFF_PN0_  (.D(_0028_),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\transfer_count[0][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][24]$_DFF_PN0_  (.D(_0029_),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\transfer_count[0][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][25]$_DFF_PN0_  (.D(_0030_),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\transfer_count[0][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][26]$_DFF_PN0_  (.D(_0031_),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\transfer_count[0][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][27]$_DFF_PN0_  (.D(_0032_),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\transfer_count[0][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][28]$_DFF_PN0_  (.D(_0033_),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\transfer_count[0][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][29]$_DFF_PN0_  (.D(_0034_),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\transfer_count[0][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][2]$_DFF_PN0_  (.D(_0035_),
    .RN(net1),
    .CLK(clknet_4_3_0_clk),
    .Q(\transfer_count[0][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][30]$_DFF_PN0_  (.D(_0036_),
    .RN(net1),
    .CLK(clknet_4_3_0_clk),
    .Q(\transfer_count[0][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][31]$_DFF_PN0_  (.D(_0037_),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\transfer_count[0][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][3]$_DFF_PN0_  (.D(_0038_),
    .RN(net1),
    .CLK(clknet_4_3_0_clk),
    .Q(\transfer_count[0][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][4]$_DFF_PN0_  (.D(_0039_),
    .RN(net1),
    .CLK(clknet_4_1_0_clk),
    .Q(\transfer_count[0][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][5]$_DFF_PN0_  (.D(_0040_),
    .RN(net1),
    .CLK(clknet_4_1_0_clk),
    .Q(\transfer_count[0][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][6]$_DFF_PN0_  (.D(_0041_),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\transfer_count[0][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][7]$_DFF_PN0_  (.D(_0042_),
    .RN(net1),
    .CLK(clknet_4_3_0_clk),
    .Q(\transfer_count[0][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][8]$_DFF_PN0_  (.D(_0043_),
    .RN(net1),
    .CLK(clknet_4_3_0_clk),
    .Q(\transfer_count[0][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[0][9]$_DFF_PN0_  (.D(_0044_),
    .RN(net1),
    .CLK(clknet_4_1_0_clk),
    .Q(\transfer_count[0][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][0]$_DFF_PN0_  (.D(_0045_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\transfer_count[1][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][10]$_DFF_PN0_  (.D(_0046_),
    .RN(net1),
    .CLK(clknet_4_14_0_clk),
    .Q(\transfer_count[1][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][11]$_DFF_PN0_  (.D(_0047_),
    .RN(net1),
    .CLK(clknet_4_14_0_clk),
    .Q(\transfer_count[1][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][12]$_DFF_PN0_  (.D(_0048_),
    .RN(net1),
    .CLK(clknet_4_14_0_clk),
    .Q(\transfer_count[1][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][13]$_DFF_PN0_  (.D(_0049_),
    .RN(net1),
    .CLK(clknet_4_14_0_clk),
    .Q(\transfer_count[1][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][14]$_DFF_PN0_  (.D(_0050_),
    .RN(net1),
    .CLK(clknet_4_14_0_clk),
    .Q(\transfer_count[1][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][15]$_DFF_PN0_  (.D(_0051_),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(\transfer_count[1][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][16]$_DFF_PN0_  (.D(_0052_),
    .RN(net1),
    .CLK(clknet_4_14_0_clk),
    .Q(\transfer_count[1][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][17]$_DFF_PN0_  (.D(_0053_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\transfer_count[1][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][18]$_DFF_PN0_  (.D(_0054_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\transfer_count[1][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][19]$_DFF_PN0_  (.D(_0055_),
    .RN(net1),
    .CLK(clknet_4_14_0_clk),
    .Q(\transfer_count[1][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][1]$_DFF_PN0_  (.D(_0056_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\transfer_count[1][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][20]$_DFF_PN0_  (.D(_0057_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\transfer_count[1][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][21]$_DFF_PN0_  (.D(_0058_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\transfer_count[1][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][22]$_DFF_PN0_  (.D(_0059_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\transfer_count[1][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][23]$_DFF_PN0_  (.D(_0060_),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(\transfer_count[1][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][24]$_DFF_PN0_  (.D(_0061_),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(\transfer_count[1][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][25]$_DFF_PN0_  (.D(_0062_),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(\transfer_count[1][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][26]$_DFF_PN0_  (.D(_0063_),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(\transfer_count[1][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][27]$_DFF_PN0_  (.D(_0064_),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(\transfer_count[1][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][28]$_DFF_PN0_  (.D(_0065_),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(\transfer_count[1][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][29]$_DFF_PN0_  (.D(_0066_),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(\transfer_count[1][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][2]$_DFF_PN0_  (.D(_0067_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\transfer_count[1][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][30]$_DFF_PN0_  (.D(_0068_),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(\transfer_count[1][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][31]$_DFF_PN0_  (.D(_0069_),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(\transfer_count[1][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][3]$_DFF_PN0_  (.D(_0070_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\transfer_count[1][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][4]$_DFF_PN0_  (.D(_0071_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\transfer_count[1][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][5]$_DFF_PN0_  (.D(_0072_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\transfer_count[1][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][6]$_DFF_PN0_  (.D(_0073_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\transfer_count[1][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][7]$_DFF_PN0_  (.D(_0074_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\transfer_count[1][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][8]$_DFF_PN0_  (.D(_0075_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\transfer_count[1][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[1][9]$_DFF_PN0_  (.D(_0076_),
    .RN(net1),
    .CLK(clknet_4_14_0_clk),
    .Q(\transfer_count[1][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][0]$_DFF_PN0_  (.D(_0077_),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(\transfer_count[2][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][10]$_DFF_PN0_  (.D(_0078_),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\transfer_count[2][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][11]$_DFF_PN0_  (.D(_0079_),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\transfer_count[2][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][12]$_DFF_PN0_  (.D(_0080_),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\transfer_count[2][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][13]$_DFF_PN0_  (.D(_0081_),
    .RN(net1),
    .CLK(clknet_4_6_0_clk),
    .Q(\transfer_count[2][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][14]$_DFF_PN0_  (.D(_0082_),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(\transfer_count[2][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][15]$_DFF_PN0_  (.D(_0083_),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\transfer_count[2][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][16]$_DFF_PN0_  (.D(_0084_),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\transfer_count[2][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][17]$_DFF_PN0_  (.D(_0085_),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\transfer_count[2][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][18]$_DFF_PN0_  (.D(_0086_),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\transfer_count[2][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][19]$_DFF_PN0_  (.D(_0087_),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\transfer_count[2][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][1]$_DFF_PN0_  (.D(_0088_),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(\transfer_count[2][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][20]$_DFF_PN0_  (.D(_0089_),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\transfer_count[2][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][21]$_DFF_PN0_  (.D(_0090_),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\transfer_count[2][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][22]$_DFF_PN0_  (.D(_0091_),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\transfer_count[2][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][23]$_DFF_PN0_  (.D(_0092_),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(\transfer_count[2][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][24]$_DFF_PN0_  (.D(_0093_),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(\transfer_count[2][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][25]$_DFF_PN0_  (.D(_0094_),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(\transfer_count[2][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][26]$_DFF_PN0_  (.D(_0095_),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(\transfer_count[2][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][27]$_DFF_PN0_  (.D(_0096_),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(\transfer_count[2][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][28]$_DFF_PN0_  (.D(_0097_),
    .RN(net1),
    .CLK(clknet_4_6_0_clk),
    .Q(\transfer_count[2][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][29]$_DFF_PN0_  (.D(_0098_),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(\transfer_count[2][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][2]$_DFF_PN0_  (.D(_0099_),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(\transfer_count[2][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][30]$_DFF_PN0_  (.D(_0100_),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(\transfer_count[2][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][31]$_DFF_PN0_  (.D(_0101_),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(\transfer_count[2][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][3]$_DFF_PN0_  (.D(_0102_),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(\transfer_count[2][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][4]$_DFF_PN0_  (.D(_0103_),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(\transfer_count[2][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][5]$_DFF_PN0_  (.D(_0104_),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(\transfer_count[2][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][6]$_DFF_PN0_  (.D(_0105_),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(\transfer_count[2][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][7]$_DFF_PN0_  (.D(_0106_),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(\transfer_count[2][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][8]$_DFF_PN0_  (.D(_0107_),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(\transfer_count[2][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[2][9]$_DFF_PN0_  (.D(_0108_),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\transfer_count[2][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][0]$_DFF_PN0_  (.D(_0109_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][10]$_DFF_PN0_  (.D(_0110_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(\transfer_count[3][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][11]$_DFF_PN0_  (.D(_0111_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][12]$_DFF_PN0_  (.D(_0112_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(\transfer_count[3][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][13]$_DFF_PN0_  (.D(_0113_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\transfer_count[3][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][14]$_DFF_PN0_  (.D(_0114_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\transfer_count[3][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][15]$_DFF_PN0_  (.D(_0115_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][16]$_DFF_PN0_  (.D(_0116_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\transfer_count[3][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][17]$_DFF_PN0_  (.D(_0117_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\transfer_count[3][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][18]$_DFF_PN0_  (.D(_0118_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\transfer_count[3][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][19]$_DFF_PN0_  (.D(_0119_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\transfer_count[3][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][1]$_DFF_PN0_  (.D(_0120_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][20]$_DFF_PN0_  (.D(_0121_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\transfer_count[3][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][21]$_DFF_PN0_  (.D(_0122_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\transfer_count[3][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][22]$_DFF_PN0_  (.D(_0123_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][23]$_DFF_PN0_  (.D(_0124_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][24]$_DFF_PN0_  (.D(_0125_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][25]$_DFF_PN0_  (.D(_0126_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][26]$_DFF_PN0_  (.D(_0127_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][27]$_DFF_PN0_  (.D(_0128_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][28]$_DFF_PN0_  (.D(_0129_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][29]$_DFF_PN0_  (.D(_0130_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\transfer_count[3][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][2]$_DFF_PN0_  (.D(_0131_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][30]$_DFF_PN0_  (.D(_0132_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\transfer_count[3][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][31]$_DFF_PN0_  (.D(_0133_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\transfer_count[3][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][3]$_DFF_PN0_  (.D(_0134_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][4]$_DFF_PN0_  (.D(_0135_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][5]$_DFF_PN0_  (.D(_0136_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][6]$_DFF_PN0_  (.D(_0137_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][7]$_DFF_PN0_  (.D(_0138_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(\transfer_count[3][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][8]$_DFF_PN0_  (.D(_0139_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(\transfer_count[3][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \transfer_count[3][9]$_DFF_PN0_  (.D(_0140_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(\transfer_count[3][9] ));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 hold1 (.I(net715),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Right_145 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Right_146 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Right_147 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Right_148 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Right_149 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Right_150 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Right_151 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Right_152 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Right_153 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Right_154 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Right_155 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Right_156 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Right_157 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Right_158 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_159_Right_159 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_160_Right_160 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_161_Right_161 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_162_Right_162 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_163_Right_163 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_164_Right_164 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_165_Right_165 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_166_Right_166 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_167_Right_167 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_168_Right_168 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_169_Right_169 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_170_Right_170 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_171_Right_171 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_172_Right_172 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_173_Right_173 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_174_Right_174 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_175_Right_175 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_176_Right_176 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_177_Right_177 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_178_Right_178 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_179_Right_179 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_180_Right_180 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_181_Right_181 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_182_Right_182 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_183_Right_183 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_184_Right_184 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_185_Right_185 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_186 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_187 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_188 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_189 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_190 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_191 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_192 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_193 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_194 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_195 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_196 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_197 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_198 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_199 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_200 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_201 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_202 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_203 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_204 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_205 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_206 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_207 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_208 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_209 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_210 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_211 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_212 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_213 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_214 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_215 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_216 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_217 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_218 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_219 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_220 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_221 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_222 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_223 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_224 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_225 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_226 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_227 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_228 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Left_229 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Left_230 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Left_231 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Left_232 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Left_233 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Left_234 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Left_235 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Left_236 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Left_237 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Left_238 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Left_239 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Left_240 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Left_241 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Left_242 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Left_243 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Left_244 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Left_245 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Left_246 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Left_247 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Left_248 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Left_249 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Left_250 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Left_251 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Left_252 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Left_253 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Left_254 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Left_255 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Left_256 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Left_257 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Left_258 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Left_259 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Left_260 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Left_261 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Left_262 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Left_263 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Left_264 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Left_265 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Left_266 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Left_267 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Left_268 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Left_269 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Left_270 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Left_271 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Left_272 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Left_273 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Left_274 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Left_275 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Left_276 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Left_277 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Left_278 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Left_279 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Left_280 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Left_281 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Left_282 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Left_283 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Left_284 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Left_285 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Left_286 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Left_287 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Left_288 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Left_289 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Left_290 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Left_291 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Left_292 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Left_293 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Left_294 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Left_295 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Left_296 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Left_297 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Left_298 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Left_299 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Left_300 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Left_301 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Left_302 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Left_303 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Left_304 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Left_305 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Left_306 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Left_307 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Left_308 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Left_309 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Left_310 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Left_311 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Left_312 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Left_313 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Left_314 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Left_315 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Left_316 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Left_317 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Left_318 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Left_319 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Left_320 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Left_321 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Left_322 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Left_323 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Left_324 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Left_325 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Left_326 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Left_327 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Left_328 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Left_329 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Left_330 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Left_331 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Left_332 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Left_333 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Left_334 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Left_335 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Left_336 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Left_337 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Left_338 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Left_339 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Left_340 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Left_341 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Left_342 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Left_343 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Left_344 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_159_Left_345 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_160_Left_346 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_161_Left_347 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_162_Left_348 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_163_Left_349 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_164_Left_350 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_165_Left_351 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_166_Left_352 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_167_Left_353 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_168_Left_354 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_169_Left_355 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_170_Left_356 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_171_Left_357 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_172_Left_358 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_173_Left_359 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_174_Left_360 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_175_Left_361 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_176_Left_362 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_177_Left_363 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_178_Left_364 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_179_Left_365 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_180_Left_366 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_181_Left_367 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_182_Left_368 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_183_Left_369 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_184_Left_370 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_185_Left_371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_375 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_376 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_377 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_378 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_379 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_380 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_381 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_382 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_383 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_384 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_385 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_386 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_387 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_388 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_467 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_468 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_961 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_962 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_963 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_964 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_965 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_966 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_967 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_968 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_969 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_970 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_971 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_972 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_973 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_974 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_975 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_976 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_977 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_978 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_979 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_980 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_981 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_982 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_983 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_984 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_985 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_986 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_987 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_988 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_989 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_990 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_991 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_992 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_993 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_994 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_995 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_996 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_997 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_998 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_999 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input1 (.I(channel_enable[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(channel_enable[1]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input3 (.I(channel_enable[2]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(channel_enable[3]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(channel_length[0]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(channel_length[100]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(channel_length[101]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(channel_length[102]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(channel_length[103]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(channel_length[104]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input11 (.I(channel_length[105]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input12 (.I(channel_length[106]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input13 (.I(channel_length[107]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input14 (.I(channel_length[108]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input15 (.I(channel_length[109]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input16 (.I(channel_length[10]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input17 (.I(channel_length[110]),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input18 (.I(channel_length[111]),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input19 (.I(channel_length[112]),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input20 (.I(channel_length[113]),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input21 (.I(channel_length[114]),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input22 (.I(channel_length[115]),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input23 (.I(channel_length[116]),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input24 (.I(channel_length[117]),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input25 (.I(channel_length[118]),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input26 (.I(channel_length[119]),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input27 (.I(channel_length[11]),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input28 (.I(channel_length[120]),
    .Z(net29));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input29 (.I(channel_length[121]),
    .Z(net30));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input30 (.I(channel_length[122]),
    .Z(net31));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input31 (.I(channel_length[123]),
    .Z(net32));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input32 (.I(channel_length[124]),
    .Z(net33));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input33 (.I(channel_length[125]),
    .Z(net34));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input34 (.I(channel_length[126]),
    .Z(net35));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input35 (.I(channel_length[127]),
    .Z(net36));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input36 (.I(channel_length[12]),
    .Z(net37));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input37 (.I(channel_length[13]),
    .Z(net38));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input38 (.I(channel_length[14]),
    .Z(net39));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input39 (.I(channel_length[15]),
    .Z(net40));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input40 (.I(channel_length[16]),
    .Z(net41));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input41 (.I(channel_length[17]),
    .Z(net42));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input42 (.I(channel_length[18]),
    .Z(net43));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input43 (.I(channel_length[19]),
    .Z(net44));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input44 (.I(channel_length[1]),
    .Z(net45));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input45 (.I(channel_length[20]),
    .Z(net46));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input46 (.I(channel_length[21]),
    .Z(net47));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input47 (.I(channel_length[22]),
    .Z(net48));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input48 (.I(channel_length[23]),
    .Z(net49));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input49 (.I(channel_length[24]),
    .Z(net50));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input50 (.I(channel_length[25]),
    .Z(net51));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input51 (.I(channel_length[26]),
    .Z(net52));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input52 (.I(channel_length[27]),
    .Z(net53));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input53 (.I(channel_length[28]),
    .Z(net54));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input54 (.I(channel_length[29]),
    .Z(net55));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input55 (.I(channel_length[2]),
    .Z(net56));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input56 (.I(channel_length[30]),
    .Z(net57));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input57 (.I(channel_length[31]),
    .Z(net58));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input58 (.I(channel_length[32]),
    .Z(net59));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input59 (.I(channel_length[33]),
    .Z(net60));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input60 (.I(channel_length[34]),
    .Z(net61));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input61 (.I(channel_length[35]),
    .Z(net62));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input62 (.I(channel_length[36]),
    .Z(net63));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input63 (.I(channel_length[37]),
    .Z(net64));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input64 (.I(channel_length[38]),
    .Z(net65));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input65 (.I(channel_length[39]),
    .Z(net66));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input66 (.I(channel_length[3]),
    .Z(net67));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input67 (.I(channel_length[40]),
    .Z(net68));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input68 (.I(channel_length[41]),
    .Z(net69));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input69 (.I(channel_length[42]),
    .Z(net70));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input70 (.I(channel_length[43]),
    .Z(net71));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input71 (.I(channel_length[44]),
    .Z(net72));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input72 (.I(channel_length[45]),
    .Z(net73));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input73 (.I(channel_length[46]),
    .Z(net74));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input74 (.I(channel_length[47]),
    .Z(net75));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input75 (.I(channel_length[48]),
    .Z(net76));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input76 (.I(channel_length[49]),
    .Z(net77));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input77 (.I(channel_length[4]),
    .Z(net78));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input78 (.I(channel_length[50]),
    .Z(net79));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input79 (.I(channel_length[51]),
    .Z(net80));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input80 (.I(channel_length[52]),
    .Z(net81));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input81 (.I(channel_length[53]),
    .Z(net82));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input82 (.I(channel_length[54]),
    .Z(net83));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input83 (.I(channel_length[55]),
    .Z(net84));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input84 (.I(channel_length[56]),
    .Z(net85));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input85 (.I(channel_length[57]),
    .Z(net86));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input86 (.I(channel_length[58]),
    .Z(net87));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input87 (.I(channel_length[59]),
    .Z(net88));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input88 (.I(channel_length[5]),
    .Z(net89));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input89 (.I(channel_length[60]),
    .Z(net90));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input90 (.I(channel_length[61]),
    .Z(net91));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input91 (.I(channel_length[62]),
    .Z(net92));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input92 (.I(channel_length[63]),
    .Z(net93));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input93 (.I(channel_length[64]),
    .Z(net94));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input94 (.I(channel_length[65]),
    .Z(net95));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input95 (.I(channel_length[66]),
    .Z(net96));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input96 (.I(channel_length[67]),
    .Z(net97));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input97 (.I(channel_length[68]),
    .Z(net98));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input98 (.I(channel_length[69]),
    .Z(net99));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input99 (.I(channel_length[6]),
    .Z(net100));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input100 (.I(channel_length[70]),
    .Z(net101));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input101 (.I(channel_length[71]),
    .Z(net102));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input102 (.I(channel_length[72]),
    .Z(net103));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input103 (.I(channel_length[73]),
    .Z(net104));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input104 (.I(channel_length[74]),
    .Z(net105));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input105 (.I(channel_length[75]),
    .Z(net106));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input106 (.I(channel_length[76]),
    .Z(net107));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input107 (.I(channel_length[77]),
    .Z(net108));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input108 (.I(channel_length[78]),
    .Z(net109));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input109 (.I(channel_length[79]),
    .Z(net110));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input110 (.I(channel_length[7]),
    .Z(net111));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input111 (.I(channel_length[80]),
    .Z(net112));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input112 (.I(channel_length[81]),
    .Z(net113));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input113 (.I(channel_length[82]),
    .Z(net114));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input114 (.I(channel_length[83]),
    .Z(net115));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input115 (.I(channel_length[84]),
    .Z(net116));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input116 (.I(channel_length[85]),
    .Z(net117));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input117 (.I(channel_length[86]),
    .Z(net118));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input118 (.I(channel_length[87]),
    .Z(net119));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input119 (.I(channel_length[88]),
    .Z(net120));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input120 (.I(channel_length[89]),
    .Z(net121));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input121 (.I(channel_length[8]),
    .Z(net122));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input122 (.I(channel_length[90]),
    .Z(net123));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input123 (.I(channel_length[91]),
    .Z(net124));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input124 (.I(channel_length[92]),
    .Z(net125));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input125 (.I(channel_length[93]),
    .Z(net126));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input126 (.I(channel_length[94]),
    .Z(net127));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input127 (.I(channel_length[95]),
    .Z(net128));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input128 (.I(channel_length[96]),
    .Z(net129));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input129 (.I(channel_length[97]),
    .Z(net130));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input130 (.I(channel_length[98]),
    .Z(net131));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input131 (.I(channel_length[99]),
    .Z(net132));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input132 (.I(channel_length[9]),
    .Z(net133));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input133 (.I(channel_start[0]),
    .Z(net134));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input134 (.I(channel_start[1]),
    .Z(net135));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input135 (.I(net716),
    .Z(net136));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input136 (.I(net717),
    .Z(net137));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input137 (.I(dst_wready[0]),
    .Z(net138));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input138 (.I(dst_wready[1]),
    .Z(net139));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input139 (.I(dst_wready[2]),
    .Z(net140));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input140 (.I(dst_wready[3]),
    .Z(net141));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input141 (.I(src_rvalid[0]),
    .Z(net142));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input142 (.I(src_rvalid[1]),
    .Z(net143));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input143 (.I(src_rvalid[2]),
    .Z(net144));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input144 (.I(src_rvalid[3]),
    .Z(net145));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output145 (.I(net146),
    .Z(channel_busy[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output146 (.I(net147),
    .Z(channel_busy[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output147 (.I(net148),
    .Z(channel_busy[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output148 (.I(net149),
    .Z(channel_busy[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output149 (.I(net150),
    .Z(channel_done[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output150 (.I(net151),
    .Z(channel_done[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output151 (.I(net152),
    .Z(channel_done[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output152 (.I(net153),
    .Z(channel_done[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output153 (.I(net154),
    .Z(channel_error[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output154 (.I(net155),
    .Z(channel_error[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output155 (.I(net156),
    .Z(channel_error[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output156 (.I(net157),
    .Z(channel_error[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output157 (.I(net158),
    .Z(debug_active_channels[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output158 (.I(net159),
    .Z(debug_active_channels[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output159 (.I(net160),
    .Z(debug_active_channels[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output160 (.I(net161),
    .Z(debug_active_channels[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output161 (.I(net162),
    .Z(debug_has_active_channels));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output162 (.I(net163),
    .Z(dst_write[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output163 (.I(net164),
    .Z(dst_write[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output164 (.I(net165),
    .Z(dst_write[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output165 (.I(net166),
    .Z(dst_write[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output166 (.I(net167),
    .Z(src_read[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output167 (.I(net168),
    .Z(src_read[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output168 (.I(net169),
    .Z(src_read[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output169 (.I(net170),
    .Z(src_read[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output170 (.I(net171),
    .Z(src_rready[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output171 (.I(net172),
    .Z(src_rready[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output172 (.I(net173),
    .Z(src_rready[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output173 (.I(net174),
    .Z(src_rready[3]));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2650__174 (.ZN(net175));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2651__175 (.ZN(net176));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2652__176 (.ZN(net177));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2653__177 (.ZN(net178));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2654__178 (.ZN(net179));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2655__179 (.ZN(net180));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2656__180 (.ZN(net181));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2657__181 (.ZN(net182));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2658__182 (.ZN(net183));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2659__183 (.ZN(net184));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2660__184 (.ZN(net185));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2661__185 (.ZN(net186));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2662__186 (.ZN(net187));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2663__187 (.ZN(net188));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2664__188 (.ZN(net189));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2665__189 (.ZN(net190));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2666__190 (.ZN(net191));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2667__191 (.ZN(net192));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2668__192 (.ZN(net193));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2669__193 (.ZN(net194));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2670__194 (.ZN(net195));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2671__195 (.ZN(net196));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2672__196 (.ZN(net197));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2673__197 (.ZN(net198));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2674__198 (.ZN(net199));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2675__199 (.ZN(net200));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2676__200 (.ZN(net201));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2677__201 (.ZN(net202));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2678__202 (.ZN(net203));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2679__203 (.ZN(net204));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2680__204 (.ZN(net205));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2681__205 (.ZN(net206));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2682__206 (.ZN(net207));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2683__207 (.ZN(net208));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2684__208 (.ZN(net209));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2685__209 (.ZN(net210));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2686__210 (.ZN(net211));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2687__211 (.ZN(net212));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2688__212 (.ZN(net213));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2689__213 (.ZN(net214));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2690__214 (.ZN(net215));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2691__215 (.ZN(net216));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2692__216 (.ZN(net217));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2693__217 (.ZN(net218));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2694__218 (.ZN(net219));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2695__219 (.ZN(net220));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2696__220 (.ZN(net221));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2697__221 (.ZN(net222));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2698__222 (.ZN(net223));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2699__223 (.ZN(net224));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2700__224 (.ZN(net225));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2701__225 (.ZN(net226));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2702__226 (.ZN(net227));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2703__227 (.ZN(net228));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2704__228 (.ZN(net229));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2705__229 (.ZN(net230));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2706__230 (.ZN(net231));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2707__231 (.ZN(net232));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2708__232 (.ZN(net233));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2709__233 (.ZN(net234));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2710__234 (.ZN(net235));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2711__235 (.ZN(net236));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2712__236 (.ZN(net237));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2713__237 (.ZN(net238));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2714__238 (.ZN(net239));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2715__239 (.ZN(net240));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2716__240 (.ZN(net241));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2717__241 (.ZN(net242));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2718__242 (.ZN(net243));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2719__243 (.ZN(net244));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2720__244 (.ZN(net245));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2721__245 (.ZN(net246));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2722__246 (.ZN(net247));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2723__247 (.ZN(net248));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2724__248 (.ZN(net249));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2725__249 (.ZN(net250));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2726__250 (.ZN(net251));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2727__251 (.ZN(net252));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2728__252 (.ZN(net253));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2729__253 (.ZN(net254));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2730__254 (.ZN(net255));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2731__255 (.ZN(net256));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2732__256 (.ZN(net257));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2733__257 (.ZN(net258));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2734__258 (.ZN(net259));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2735__259 (.ZN(net260));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2736__260 (.ZN(net261));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2737__261 (.ZN(net262));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2738__262 (.ZN(net263));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2739__263 (.ZN(net264));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2740__264 (.ZN(net265));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2741__265 (.ZN(net266));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2742__266 (.ZN(net267));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2743__267 (.ZN(net268));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2744__268 (.ZN(net269));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2745__269 (.ZN(net270));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2746__270 (.ZN(net271));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2747__271 (.ZN(net272));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2748__272 (.ZN(net273));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2749__273 (.ZN(net274));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2750__274 (.ZN(net275));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2751__275 (.ZN(net276));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2752__276 (.ZN(net277));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2753__277 (.ZN(net278));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2754__278 (.ZN(net279));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2755__279 (.ZN(net280));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2756__280 (.ZN(net281));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2757__281 (.ZN(net282));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2758__282 (.ZN(net283));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2759__283 (.ZN(net284));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2760__284 (.ZN(net285));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2761__285 (.ZN(net286));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2762__286 (.ZN(net287));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2763__287 (.ZN(net288));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2764__288 (.ZN(net289));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2765__289 (.ZN(net290));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2766__290 (.ZN(net291));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2767__291 (.ZN(net292));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2768__292 (.ZN(net293));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2769__293 (.ZN(net294));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2770__294 (.ZN(net295));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2771__295 (.ZN(net296));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2772__296 (.ZN(net297));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2773__297 (.ZN(net298));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2774__298 (.ZN(net299));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2775__299 (.ZN(net300));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2776__300 (.ZN(net301));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2777__301 (.ZN(net302));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2778__302 (.ZN(net303));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2779__303 (.ZN(net304));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2780__304 (.ZN(net305));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2781__305 (.ZN(net306));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2782__306 (.ZN(net307));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2783__307 (.ZN(net308));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2784__308 (.ZN(net309));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2785__309 (.ZN(net310));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2786__310 (.ZN(net311));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2787__311 (.ZN(net312));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2788__312 (.ZN(net313));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2789__313 (.ZN(net314));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2790__314 (.ZN(net315));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2791__315 (.ZN(net316));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2792__316 (.ZN(net317));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2793__317 (.ZN(net318));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2794__318 (.ZN(net319));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2795__319 (.ZN(net320));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2796__320 (.ZN(net321));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2797__321 (.ZN(net322));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2798__322 (.ZN(net323));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2799__323 (.ZN(net324));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2800__324 (.ZN(net325));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2801__325 (.ZN(net326));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2802__326 (.ZN(net327));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2803__327 (.ZN(net328));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2804__328 (.ZN(net329));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2805__329 (.ZN(net330));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2806__330 (.ZN(net331));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2807__331 (.ZN(net332));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2808__332 (.ZN(net333));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2809__333 (.ZN(net334));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2810__334 (.ZN(net335));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2811__335 (.ZN(net336));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2812__336 (.ZN(net337));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2813__337 (.ZN(net338));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2814__338 (.ZN(net339));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2815__339 (.ZN(net340));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2816__340 (.ZN(net341));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2817__341 (.ZN(net342));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2818__342 (.ZN(net343));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2819__343 (.ZN(net344));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2820__344 (.ZN(net345));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2821__345 (.ZN(net346));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2822__346 (.ZN(net347));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2823__347 (.ZN(net348));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2824__348 (.ZN(net349));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2825__349 (.ZN(net350));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2826__350 (.ZN(net351));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2827__351 (.ZN(net352));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2828__352 (.ZN(net353));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2829__353 (.ZN(net354));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2830__354 (.ZN(net355));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2831__355 (.ZN(net356));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2832__356 (.ZN(net357));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2833__357 (.ZN(net358));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2834__358 (.ZN(net359));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2835__359 (.ZN(net360));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2836__360 (.ZN(net361));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2837__361 (.ZN(net362));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2838__362 (.ZN(net363));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2839__363 (.ZN(net364));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2840__364 (.ZN(net365));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2841__365 (.ZN(net366));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2842__366 (.ZN(net367));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2843__367 (.ZN(net368));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2844__368 (.ZN(net369));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2845__369 (.ZN(net370));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2846__370 (.ZN(net371));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2847__371 (.ZN(net372));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2848__372 (.ZN(net373));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2849__373 (.ZN(net374));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2850__374 (.ZN(net375));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2851__375 (.ZN(net376));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2852__376 (.ZN(net377));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2853__377 (.ZN(net378));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2854__378 (.ZN(net379));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2855__379 (.ZN(net380));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2856__380 (.ZN(net381));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2857__381 (.ZN(net382));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2858__382 (.ZN(net383));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2859__383 (.ZN(net384));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2860__384 (.ZN(net385));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2861__385 (.ZN(net386));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2862__386 (.ZN(net387));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2863__387 (.ZN(net388));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2864__388 (.ZN(net389));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2865__389 (.ZN(net390));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2866__390 (.ZN(net391));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2867__391 (.ZN(net392));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2868__392 (.ZN(net393));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2869__393 (.ZN(net394));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2870__394 (.ZN(net395));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2871__395 (.ZN(net396));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2872__396 (.ZN(net397));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2873__397 (.ZN(net398));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2874__398 (.ZN(net399));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2875__399 (.ZN(net400));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2876__400 (.ZN(net401));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2877__401 (.ZN(net402));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2878__402 (.ZN(net403));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2879__403 (.ZN(net404));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2880__404 (.ZN(net405));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2881__405 (.ZN(net406));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2882__406 (.ZN(net407));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2883__407 (.ZN(net408));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2884__408 (.ZN(net409));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2885__409 (.ZN(net410));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2886__410 (.ZN(net411));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2887__411 (.ZN(net412));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2888__412 (.ZN(net413));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2889__413 (.ZN(net414));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2890__414 (.ZN(net415));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2891__415 (.ZN(net416));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2892__416 (.ZN(net417));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2893__417 (.ZN(net418));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2894__418 (.ZN(net419));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2895__419 (.ZN(net420));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2896__420 (.ZN(net421));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2897__421 (.ZN(net422));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2898__422 (.ZN(net423));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2899__423 (.ZN(net424));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2900__424 (.ZN(net425));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2901__425 (.ZN(net426));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2902__426 (.ZN(net427));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2903__427 (.ZN(net428));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2904__428 (.ZN(net429));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2905__429 (.ZN(net430));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2906__430 (.ZN(net431));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2907__431 (.ZN(net432));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2908__432 (.ZN(net433));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2909__433 (.ZN(net434));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2910__434 (.ZN(net435));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2911__435 (.ZN(net436));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2912__436 (.ZN(net437));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2913__437 (.ZN(net438));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2914__438 (.ZN(net439));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2915__439 (.ZN(net440));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2916__440 (.ZN(net441));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2917__441 (.ZN(net442));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2918__442 (.ZN(net443));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2919__443 (.ZN(net444));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2920__444 (.ZN(net445));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2921__445 (.ZN(net446));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2922__446 (.ZN(net447));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2923__447 (.ZN(net448));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2924__448 (.ZN(net449));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2925__449 (.ZN(net450));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2926__450 (.ZN(net451));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2927__451 (.ZN(net452));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2928__452 (.ZN(net453));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2929__453 (.ZN(net454));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2930__454 (.ZN(net455));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2931__455 (.ZN(net456));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2932__456 (.ZN(net457));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2933__457 (.ZN(net458));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2934__458 (.ZN(net459));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2935__459 (.ZN(net460));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2936__460 (.ZN(net461));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2937__461 (.ZN(net462));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2938__462 (.ZN(net463));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2939__463 (.ZN(net464));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2940__464 (.ZN(net465));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2941__465 (.ZN(net466));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2942__466 (.ZN(net467));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2943__467 (.ZN(net468));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2944__468 (.ZN(net469));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2945__469 (.ZN(net470));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2946__470 (.ZN(net471));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2947__471 (.ZN(net472));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2948__472 (.ZN(net473));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2949__473 (.ZN(net474));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2950__474 (.ZN(net475));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2951__475 (.ZN(net476));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2952__476 (.ZN(net477));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2953__477 (.ZN(net478));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2954__478 (.ZN(net479));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2955__479 (.ZN(net480));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2956__480 (.ZN(net481));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2957__481 (.ZN(net482));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2958__482 (.ZN(net483));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2959__483 (.ZN(net484));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2960__484 (.ZN(net485));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2961__485 (.ZN(net486));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2962__486 (.ZN(net487));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2963__487 (.ZN(net488));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2964__488 (.ZN(net489));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2965__489 (.ZN(net490));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2966__490 (.ZN(net491));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2967__491 (.ZN(net492));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2968__492 (.ZN(net493));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2969__493 (.ZN(net494));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2970__494 (.ZN(net495));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2971__495 (.ZN(net496));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2972__496 (.ZN(net497));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2973__497 (.ZN(net498));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2974__498 (.ZN(net499));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2975__499 (.ZN(net500));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2976__500 (.ZN(net501));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2977__501 (.ZN(net502));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2978__502 (.ZN(net503));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2979__503 (.ZN(net504));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2980__504 (.ZN(net505));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2981__505 (.ZN(net506));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2982__506 (.ZN(net507));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2983__507 (.ZN(net508));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2984__508 (.ZN(net509));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2985__509 (.ZN(net510));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2986__510 (.ZN(net511));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2987__511 (.ZN(net512));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2988__512 (.ZN(net513));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2989__513 (.ZN(net514));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2990__514 (.ZN(net515));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2991__515 (.ZN(net516));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2992__516 (.ZN(net517));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2993__517 (.ZN(net518));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2994__518 (.ZN(net519));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2995__519 (.ZN(net520));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2996__520 (.ZN(net521));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2997__521 (.ZN(net522));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2998__522 (.ZN(net523));
 gf180mcu_fd_sc_mcu9t5v0__tiel _2999__523 (.ZN(net524));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3000__524 (.ZN(net525));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3001__525 (.ZN(net526));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3002__526 (.ZN(net527));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3003__527 (.ZN(net528));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3004__528 (.ZN(net529));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3005__529 (.ZN(net530));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3006__530 (.ZN(net531));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3007__531 (.ZN(net532));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3008__532 (.ZN(net533));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3009__533 (.ZN(net534));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3010__534 (.ZN(net535));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3011__535 (.ZN(net536));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3012__536 (.ZN(net537));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3013__537 (.ZN(net538));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3014__538 (.ZN(net539));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3015__539 (.ZN(net540));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3016__540 (.ZN(net541));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3017__541 (.ZN(net542));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3018__542 (.ZN(net543));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3019__543 (.ZN(net544));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3020__544 (.ZN(net545));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3021__545 (.ZN(net546));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3022__546 (.ZN(net547));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3023__547 (.ZN(net548));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3024__548 (.ZN(net549));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3025__549 (.ZN(net550));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3026__550 (.ZN(net551));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3027__551 (.ZN(net552));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3028__552 (.ZN(net553));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3029__553 (.ZN(net554));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3030__554 (.ZN(net555));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3031__555 (.ZN(net556));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3032__556 (.ZN(net557));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3033__557 (.ZN(net558));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3034__558 (.ZN(net559));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3035__559 (.ZN(net560));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3036__560 (.ZN(net561));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3037__561 (.ZN(net562));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3038__562 (.ZN(net563));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3039__563 (.ZN(net564));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3040__564 (.ZN(net565));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3041__565 (.ZN(net566));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3042__566 (.ZN(net567));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3043__567 (.ZN(net568));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3044__568 (.ZN(net569));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3045__569 (.ZN(net570));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3046__570 (.ZN(net571));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3047__571 (.ZN(net572));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3048__572 (.ZN(net573));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3049__573 (.ZN(net574));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3050__574 (.ZN(net575));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3051__575 (.ZN(net576));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3052__576 (.ZN(net577));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3053__577 (.ZN(net578));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3054__578 (.ZN(net579));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3055__579 (.ZN(net580));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3056__580 (.ZN(net581));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3057__581 (.ZN(net582));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3058__582 (.ZN(net583));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3059__583 (.ZN(net584));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3060__584 (.ZN(net585));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3061__585 (.ZN(net586));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3062__586 (.ZN(net587));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3063__587 (.ZN(net588));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3064__588 (.ZN(net589));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3065__589 (.ZN(net590));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3066__590 (.ZN(net591));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3067__591 (.ZN(net592));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3068__592 (.ZN(net593));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3069__593 (.ZN(net594));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3070__594 (.ZN(net595));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3071__595 (.ZN(net596));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3072__596 (.ZN(net597));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3073__597 (.ZN(net598));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3074__598 (.ZN(net599));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3075__599 (.ZN(net600));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3076__600 (.ZN(net601));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3077__601 (.ZN(net602));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3078__602 (.ZN(net603));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3079__603 (.ZN(net604));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3080__604 (.ZN(net605));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3081__605 (.ZN(net606));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3082__606 (.ZN(net607));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3083__607 (.ZN(net608));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3084__608 (.ZN(net609));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3085__609 (.ZN(net610));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3086__610 (.ZN(net611));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3087__611 (.ZN(net612));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3088__612 (.ZN(net613));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3089__613 (.ZN(net614));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3090__614 (.ZN(net615));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3091__615 (.ZN(net616));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3092__616 (.ZN(net617));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3093__617 (.ZN(net618));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3094__618 (.ZN(net619));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3095__619 (.ZN(net620));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3096__620 (.ZN(net621));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3097__621 (.ZN(net622));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3098__622 (.ZN(net623));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3099__623 (.ZN(net624));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3100__624 (.ZN(net625));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3101__625 (.ZN(net626));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3102__626 (.ZN(net627));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3103__627 (.ZN(net628));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3104__628 (.ZN(net629));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3105__629 (.ZN(net630));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3106__630 (.ZN(net631));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3107__631 (.ZN(net632));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3108__632 (.ZN(net633));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3109__633 (.ZN(net634));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3110__634 (.ZN(net635));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3111__635 (.ZN(net636));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3112__636 (.ZN(net637));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3113__637 (.ZN(net638));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3114__638 (.ZN(net639));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3115__639 (.ZN(net640));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3116__640 (.ZN(net641));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3117__641 (.ZN(net642));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3118__642 (.ZN(net643));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3119__643 (.ZN(net644));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3120__644 (.ZN(net645));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3121__645 (.ZN(net646));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3122__646 (.ZN(net647));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3123__647 (.ZN(net648));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3124__648 (.ZN(net649));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3125__649 (.ZN(net650));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3126__650 (.ZN(net651));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3127__651 (.ZN(net652));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3128__652 (.ZN(net653));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3129__653 (.ZN(net654));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3130__654 (.ZN(net655));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3131__655 (.ZN(net656));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3132__656 (.ZN(net657));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3133__657 (.ZN(net658));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3134__658 (.ZN(net659));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3135__659 (.ZN(net660));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3136__660 (.ZN(net661));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3137__661 (.ZN(net662));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3138__662 (.ZN(net663));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3139__663 (.ZN(net664));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3140__664 (.ZN(net665));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3141__665 (.ZN(net666));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3142__666 (.ZN(net667));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3143__667 (.ZN(net668));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3144__668 (.ZN(net669));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3145__669 (.ZN(net670));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3146__670 (.ZN(net671));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3147__671 (.ZN(net672));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3148__672 (.ZN(net673));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3149__673 (.ZN(net674));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3150__674 (.ZN(net675));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3151__675 (.ZN(net676));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3152__676 (.ZN(net677));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3153__677 (.ZN(net678));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3154__678 (.ZN(net679));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3155__679 (.ZN(net680));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3156__680 (.ZN(net681));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3157__681 (.ZN(net682));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3158__682 (.ZN(net683));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3159__683 (.ZN(net684));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3160__684 (.ZN(net685));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3161__685 (.ZN(net686));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3162__686 (.ZN(net687));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3163__687 (.ZN(net688));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3164__688 (.ZN(net689));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3165__689 (.ZN(net690));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3166__690 (.ZN(net691));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3167__691 (.ZN(net692));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3168__692 (.ZN(net693));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3169__693 (.ZN(net694));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3170__694 (.ZN(net695));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3171__695 (.ZN(net696));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3172__696 (.ZN(net697));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3173__697 (.ZN(net698));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3174__698 (.ZN(net699));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3175__699 (.ZN(net700));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3176__700 (.ZN(net701));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3177__701 (.ZN(net702));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3178__702 (.ZN(net703));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3179__703 (.ZN(net704));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3180__704 (.ZN(net705));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3181__705 (.ZN(net706));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3182__706 (.ZN(net707));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3183__707 (.ZN(net708));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3184__708 (.ZN(net709));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3185__709 (.ZN(net710));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3186__710 (.ZN(net711));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3187__711 (.ZN(net712));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3188__712 (.ZN(net713));
 gf180mcu_fd_sc_mcu9t5v0__tiel _3189__713 (.ZN(net714));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_0_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_1_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_2_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_3_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_4_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_5_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_6_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_7_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_8_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_9_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_10_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_11_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_12_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_13_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_14_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_15_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 clkload0 (.I(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 clkload1 (.I(clknet_4_1_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload2 (.I(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkload3 (.I(clknet_4_3_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload4 (.I(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload5 (.I(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 clkload6 (.I(clknet_4_6_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 clkload7 (.I(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload8 (.I(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload9 (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload10 (.I(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 clkload11 (.I(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload12 (.I(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload13 (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload14 (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net715));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold3 (.I(channel_start[2]),
    .Z(net716));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold4 (.I(channel_start[3]),
    .Z(net717));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_1 (.I(net149));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_2 (.I(net153));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_3 (.I(net157));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_4 (.I(net157));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_5 (.I(net166));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_27 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1675 ();
endmodule
