module bsg_async_credit_counter (r_clk_i,
    r_credits_avail_o,
    r_dec_credit_i,
    r_infinite_credits_i,
    r_reset_i,
    w_clk_i,
    w_inc_token_i,
    w_reset_i);
 input r_clk_i;
 output r_credits_avail_o;
 input r_dec_credit_i;
 input r_infinite_credits_i;
 input r_reset_i;
 input w_clk_i;
 input w_inc_token_i;
 input w_reset_i;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire \bapg.w_ptr_binary_r_o[0] ;
 wire \bapg.w_ptr_binary_r_o[1] ;
 wire \bapg.w_ptr_binary_r_o[2] ;
 wire \bapg.w_ptr_gray_r[0] ;
 wire \bapg.w_ptr_gray_r[1] ;
 wire \bapg.w_ptr_gray_r_rsync_o[0] ;
 wire \bapg.w_ptr_gray_r_rsync_o[1] ;
 wire \bapg.w_ptr_gray_r_rsync_o[2] ;
 wire \bapg.w_ptr_gray_r_rsync_r[0][0] ;
 wire \bapg.w_ptr_gray_r_rsync_r[0][1] ;
 wire \bapg.w_ptr_gray_r_rsync_r[0][2] ;
 wire \bapg.w_ptr_n[0] ;
 wire \bapg.w_ptr_n[1] ;
 wire \r_counter_r[0] ;
 wire \r_counter_r[1] ;
 wire \r_counter_r[2] ;
 wire \r_counter_r_hi_bits_gray[0] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire clknet_0_w_clk_i;
 wire clknet_1_0__leaf_w_clk_i;
 wire clknet_1_1__leaf_w_clk_i;

 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30_ (.I(net6),
    .ZN(_08_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31_ (.A1(\bapg.w_ptr_n[0] ),
    .A2(\bapg.w_ptr_n[1] ),
    .Z(_09_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _32_ (.I0(\bapg.w_ptr_gray_r[0] ),
    .I1(_09_),
    .S(net5),
    .Z(_10_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _33_ (.A1(_08_),
    .A2(_10_),
    .Z(_00_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _34_ (.A1(\bapg.w_ptr_binary_r_o[2] ),
    .A2(\bapg.w_ptr_n[1] ),
    .A3(_28_),
    .Z(_11_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _35_ (.I0(\bapg.w_ptr_gray_r[1] ),
    .I1(_11_),
    .S(net5),
    .Z(_12_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _36_ (.A1(_08_),
    .A2(_12_),
    .Z(_01_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _37_ (.A1(net5),
    .A2(_28_),
    .ZN(_13_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _38_ (.A1(\bapg.w_ptr_binary_r_o[2] ),
    .A2(_13_),
    .ZN(_14_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _39_ (.A1(_08_),
    .A2(_14_),
    .Z(_02_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _40_ (.I0(\bapg.w_ptr_binary_r_o[0] ),
    .I1(\bapg.w_ptr_n[0] ),
    .S(net5),
    .Z(_15_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _41_ (.A1(_08_),
    .A2(_15_),
    .Z(_03_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _42_ (.I0(\bapg.w_ptr_binary_r_o[1] ),
    .I1(\bapg.w_ptr_n[1] ),
    .S(net5),
    .Z(_16_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _43_ (.A1(_08_),
    .A2(_16_),
    .Z(_04_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _44_ (.I(net4),
    .ZN(_17_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _45_ (.A1(\r_counter_r[0] ),
    .A2(net2),
    .Z(_18_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _46_ (.A1(_17_),
    .A2(_18_),
    .Z(_05_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _47_ (.I0(\r_counter_r[1] ),
    .I1(\r_counter_r_hi_bits_gray[0] ),
    .S(net2),
    .Z(_19_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _48_ (.A1(_17_),
    .A2(_19_),
    .Z(_06_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _49_ (.A1(_29_),
    .A2(net2),
    .Z(_20_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _50_ (.A1(\r_counter_r[2] ),
    .A2(_20_),
    .ZN(_21_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _51_ (.A1(_17_),
    .A2(_21_),
    .ZN(_07_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _52_ (.A1(\r_counter_r[2] ),
    .A2(\bapg.w_ptr_gray_r_rsync_o[2] ),
    .ZN(_22_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _53_ (.A1(\r_counter_r[2] ),
    .A2(\bapg.w_ptr_gray_r_rsync_o[2] ),
    .Z(_23_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _54_ (.A1(\r_counter_r[1] ),
    .A2(\bapg.w_ptr_gray_r_rsync_o[1] ),
    .ZN(_24_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _55_ (.I0(_22_),
    .I1(_23_),
    .S(_24_),
    .Z(_25_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _56_ (.A1(\r_counter_r_hi_bits_gray[0] ),
    .A2(\bapg.w_ptr_gray_r_rsync_o[0] ),
    .Z(_26_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _57_ (.A1(net3),
    .A2(_25_),
    .A3(_26_),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _58_ (.A(net5),
    .B(\bapg.w_ptr_binary_r_o[0] ),
    .CO(_27_),
    .S(\bapg.w_ptr_n[0] ));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _59_ (.A(\bapg.w_ptr_binary_r_o[1] ),
    .B(_27_),
    .CO(_28_),
    .S(\bapg.w_ptr_n[1] ));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _60_ (.A(\r_counter_r[0] ),
    .B(\r_counter_r[1] ),
    .CO(_29_),
    .S(\r_counter_r_hi_bits_gray[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \bapg.w_ptr_gray_r[0]$_SDFFE_PP0P_  (.D(_00_),
    .CLK(clknet_1_1__leaf_w_clk_i),
    .Q(\bapg.w_ptr_gray_r[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \bapg.w_ptr_gray_r[1]$_SDFFE_PP0P_  (.D(_01_),
    .CLK(clknet_1_1__leaf_w_clk_i),
    .Q(\bapg.w_ptr_gray_r[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \bapg.w_ptr_gray_r[2]$_SDFFE_PP0P_  (.D(_02_),
    .CLK(clknet_1_1__leaf_w_clk_i),
    .Q(\bapg.w_ptr_binary_r_o[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \bapg.w_ptr_gray_r_rsync_r[0][0]$_DFF_P_  (.D(\bapg.w_ptr_gray_r[0] ),
    .CLK(net1),
    .Q(\bapg.w_ptr_gray_r_rsync_r[0][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \bapg.w_ptr_gray_r_rsync_r[0][1]$_DFF_P_  (.D(\bapg.w_ptr_gray_r[1] ),
    .CLK(net1),
    .Q(\bapg.w_ptr_gray_r_rsync_r[0][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \bapg.w_ptr_gray_r_rsync_r[0][2]$_DFF_P_  (.D(\bapg.w_ptr_binary_r_o[2] ),
    .CLK(net1),
    .Q(\bapg.w_ptr_gray_r_rsync_r[0][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \bapg.w_ptr_gray_r_rsync_r[1][0]$_DFF_P_  (.D(\bapg.w_ptr_gray_r_rsync_r[0][0] ),
    .CLK(net1),
    .Q(\bapg.w_ptr_gray_r_rsync_o[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \bapg.w_ptr_gray_r_rsync_r[1][1]$_DFF_P_  (.D(\bapg.w_ptr_gray_r_rsync_r[0][1] ),
    .CLK(net1),
    .Q(\bapg.w_ptr_gray_r_rsync_o[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \bapg.w_ptr_gray_r_rsync_r[1][2]$_DFF_P_  (.D(\bapg.w_ptr_gray_r_rsync_r[0][2] ),
    .CLK(net1),
    .Q(\bapg.w_ptr_gray_r_rsync_o[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \bapg.w_ptr_r[0]$_SDFFE_PP0P_  (.D(_03_),
    .CLK(clknet_1_0__leaf_w_clk_i),
    .Q(\bapg.w_ptr_binary_r_o[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \bapg.w_ptr_r[1]$_SDFFE_PP0P_  (.D(_04_),
    .CLK(clknet_1_0__leaf_w_clk_i),
    .Q(\bapg.w_ptr_binary_r_o[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \r_counter_r[0]$_SDFFE_PP0P_  (.D(_05_),
    .CLK(net1),
    .Q(\r_counter_r[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \r_counter_r[1]$_SDFFE_PP0P_  (.D(_06_),
    .CLK(net1),
    .Q(\r_counter_r[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \r_counter_r[2]$_SDFFE_PP1P_  (.D(_07_),
    .CLK(net1),
    .Q(\r_counter_r[2] ));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_46 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_47 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_48 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_49 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_50 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_51 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_52 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_53 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_54 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_55 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_56 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_57 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input1 (.I(r_clk_i),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(r_dec_credit_i),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(r_infinite_credits_i),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(r_reset_i),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input5 (.I(w_inc_token_i),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(w_reset_i),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output7 (.I(net7),
    .Z(r_credits_avail_o));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_0_w_clk_i (.I(w_clk_i),
    .Z(clknet_0_w_clk_i));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_0__f_w_clk_i (.I(clknet_0_w_clk_i),
    .Z(clknet_1_0__leaf_w_clk_i));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_1__f_w_clk_i (.I(clknet_0_w_clk_i),
    .Z(clknet_1_1__leaf_w_clk_i));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload0 (.I(clknet_1_0__leaf_w_clk_i));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_23 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_7 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_212 ();
endmodule
