module fixed_spi_master (clk,
    rst_n,
    rx_valid,
    spi_clk,
    spi_cs_n,
    spi_miso,
    spi_mosi,
    tx_ready,
    tx_valid,
    rx_data,
    tx_data);
 input clk;
 input rst_n;
 output rx_valid;
 output spi_clk;
 output spi_cs_n;
 input spi_miso;
 output spi_mosi;
 output tx_ready;
 input tx_valid;
 output [7:0] rx_data;
 input [7:0] tx_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire \bit_counter[0] ;
 wire \bit_counter[1] ;
 wire \bit_counter[2] ;
 wire \bit_counter[3] ;
 wire \rx_shift_reg[0] ;
 wire \rx_shift_reg[1] ;
 wire \rx_shift_reg[2] ;
 wire \rx_shift_reg[3] ;
 wire \rx_shift_reg[4] ;
 wire \rx_shift_reg[5] ;
 wire \rx_shift_reg[6] ;
 wire \rx_shift_reg[7] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \tx_shift_reg[0] ;
 wire \tx_shift_reg[1] ;
 wire \tx_shift_reg[2] ;
 wire \tx_shift_reg[3] ;
 wire \tx_shift_reg[4] ;
 wire \tx_shift_reg[5] ;
 wire \tx_shift_reg[6] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 BUF_X4 _210_ (.A(\bit_counter[2] ),
    .Z(_156_));
 BUF_X4 _211_ (.A(_191_),
    .Z(_157_));
 NAND2_X1 _212_ (.A1(_156_),
    .A2(_157_),
    .ZN(_158_));
 OR2_X2 _213_ (.A1(\bit_counter[3] ),
    .A2(_158_),
    .ZN(_197_));
 INV_X1 _214_ (.A(_197_),
    .ZN(_204_));
 CLKBUF_X2 _215_ (.A(rst_n),
    .Z(_037_));
 INV_X1 _216_ (.A(_037_),
    .ZN(_038_));
 CLKBUF_X3 _217_ (.A(_038_),
    .Z(_039_));
 BUF_X4 _218_ (.A(\state[2] ),
    .Z(_040_));
 CLKBUF_X3 _219_ (.A(_040_),
    .Z(_041_));
 NOR3_X1 _220_ (.A1(\bit_counter[3] ),
    .A2(_200_),
    .A3(_158_),
    .ZN(_042_));
 BUF_X2 _221_ (.A(net20),
    .Z(_043_));
 INV_X1 _222_ (.A(_200_),
    .ZN(_044_));
 OAI21_X1 _223_ (.A(_043_),
    .B1(_004_),
    .B2(_044_),
    .ZN(_045_));
 OAI21_X1 _224_ (.A(_041_),
    .B1(_042_),
    .B2(_045_),
    .ZN(_046_));
 BUF_X2 _225_ (.A(\state[0] ),
    .Z(_047_));
 NAND2_X1 _226_ (.A1(net10),
    .A2(_047_),
    .ZN(_048_));
 AOI21_X1 _227_ (.A(_039_),
    .B1(_046_),
    .B2(_048_),
    .ZN(_002_));
 BUF_X2 _228_ (.A(_037_),
    .Z(_049_));
 BUF_X2 _229_ (.A(\state[1] ),
    .Z(_050_));
 INV_X1 _230_ (.A(_050_),
    .ZN(_051_));
 CLKBUF_X3 _231_ (.A(_051_),
    .Z(_052_));
 INV_X1 _232_ (.A(net10),
    .ZN(_053_));
 NAND2_X1 _233_ (.A1(_053_),
    .A2(_047_),
    .ZN(_054_));
 NAND3_X1 _234_ (.A1(_049_),
    .A2(_052_),
    .A3(_054_),
    .ZN(_001_));
 BUF_X2 _235_ (.A(_202_),
    .Z(_055_));
 AND4_X1 _236_ (.A1(_049_),
    .A2(_043_),
    .A3(_041_),
    .A4(_055_),
    .ZN(_000_));
 BUF_X2 _237_ (.A(\bit_counter[0] ),
    .Z(_056_));
 NAND3_X1 _238_ (.A1(_156_),
    .A2(_056_),
    .A3(\bit_counter[1] ),
    .ZN(_194_));
 OR2_X1 _239_ (.A1(\bit_counter[3] ),
    .A2(_194_),
    .ZN(_207_));
 INV_X2 _240_ (.A(_040_),
    .ZN(_057_));
 NOR2_X1 _241_ (.A1(_057_),
    .A2(_056_),
    .ZN(_058_));
 INV_X2 _242_ (.A(_047_),
    .ZN(_059_));
 NAND2_X1 _243_ (.A1(_043_),
    .A2(_040_),
    .ZN(_060_));
 OAI22_X4 _244_ (.A1(_059_),
    .A2(_040_),
    .B1(_055_),
    .B2(_060_),
    .ZN(_061_));
 MUX2_X1 _245_ (.A(_056_),
    .B(_058_),
    .S(_061_),
    .Z(_062_));
 AND2_X1 _246_ (.A1(_049_),
    .A2(_062_),
    .ZN(_005_));
 INV_X1 _247_ (.A(_192_),
    .ZN(_063_));
 NOR2_X1 _248_ (.A1(_057_),
    .A2(_063_),
    .ZN(_064_));
 MUX2_X1 _249_ (.A(\bit_counter[1] ),
    .B(_064_),
    .S(_061_),
    .Z(_065_));
 AND2_X1 _250_ (.A1(_049_),
    .A2(_065_),
    .ZN(_006_));
 INV_X1 _251_ (.A(_055_),
    .ZN(_066_));
 AND2_X1 _252_ (.A1(_043_),
    .A2(_041_),
    .ZN(_067_));
 AOI22_X1 _253_ (.A1(_047_),
    .A2(_057_),
    .B1(_066_),
    .B2(_067_),
    .ZN(_068_));
 NOR2_X1 _254_ (.A1(_157_),
    .A2(_057_),
    .ZN(_069_));
 OAI21_X1 _255_ (.A(_156_),
    .B1(_068_),
    .B2(_069_),
    .ZN(_070_));
 NOR2_X1 _256_ (.A1(_156_),
    .A2(_057_),
    .ZN(_071_));
 NAND3_X1 _257_ (.A1(_157_),
    .A2(_061_),
    .A3(_071_),
    .ZN(_072_));
 AOI21_X1 _258_ (.A(_039_),
    .B1(_070_),
    .B2(_072_),
    .ZN(_007_));
 INV_X1 _259_ (.A(_196_),
    .ZN(_073_));
 NOR2_X1 _260_ (.A1(_057_),
    .A2(_073_),
    .ZN(_074_));
 MUX2_X1 _261_ (.A(\bit_counter[3] ),
    .B(_074_),
    .S(_061_),
    .Z(_075_));
 AND2_X1 _262_ (.A1(_049_),
    .A2(_075_),
    .ZN(_008_));
 CLKBUF_X3 _263_ (.A(_038_),
    .Z(_076_));
 NAND2_X1 _264_ (.A1(_050_),
    .A2(\rx_shift_reg[0] ),
    .ZN(_077_));
 NAND2_X1 _265_ (.A1(_052_),
    .A2(net11),
    .ZN(_078_));
 AOI21_X1 _266_ (.A(_076_),
    .B1(_077_),
    .B2(_078_),
    .ZN(_009_));
 NAND2_X1 _267_ (.A1(_050_),
    .A2(\rx_shift_reg[1] ),
    .ZN(_079_));
 NAND2_X1 _268_ (.A1(_052_),
    .A2(net12),
    .ZN(_080_));
 AOI21_X1 _269_ (.A(_076_),
    .B1(_079_),
    .B2(_080_),
    .ZN(_010_));
 NAND2_X1 _270_ (.A1(_050_),
    .A2(\rx_shift_reg[2] ),
    .ZN(_081_));
 NAND2_X1 _271_ (.A1(_052_),
    .A2(net13),
    .ZN(_082_));
 AOI21_X1 _272_ (.A(_076_),
    .B1(_081_),
    .B2(_082_),
    .ZN(_011_));
 NAND2_X1 _273_ (.A1(_050_),
    .A2(\rx_shift_reg[3] ),
    .ZN(_083_));
 NAND2_X1 _274_ (.A1(_052_),
    .A2(net14),
    .ZN(_084_));
 AOI21_X1 _275_ (.A(_076_),
    .B1(_083_),
    .B2(_084_),
    .ZN(_012_));
 NAND2_X1 _276_ (.A1(_050_),
    .A2(\rx_shift_reg[4] ),
    .ZN(_085_));
 NAND2_X1 _277_ (.A1(_052_),
    .A2(net15),
    .ZN(_086_));
 AOI21_X1 _278_ (.A(_076_),
    .B1(_085_),
    .B2(_086_),
    .ZN(_013_));
 NAND2_X1 _279_ (.A1(_050_),
    .A2(\rx_shift_reg[5] ),
    .ZN(_087_));
 NAND2_X1 _280_ (.A1(_052_),
    .A2(net16),
    .ZN(_088_));
 AOI21_X1 _281_ (.A(_076_),
    .B1(_087_),
    .B2(_088_),
    .ZN(_014_));
 NAND2_X1 _282_ (.A1(_050_),
    .A2(\rx_shift_reg[6] ),
    .ZN(_089_));
 NAND2_X1 _283_ (.A1(_052_),
    .A2(net17),
    .ZN(_090_));
 AOI21_X1 _284_ (.A(_076_),
    .B1(_089_),
    .B2(_090_),
    .ZN(_015_));
 NAND2_X1 _285_ (.A1(_050_),
    .A2(\rx_shift_reg[7] ),
    .ZN(_091_));
 NAND2_X1 _286_ (.A1(_051_),
    .A2(net18),
    .ZN(_092_));
 AOI21_X1 _287_ (.A(_076_),
    .B1(_091_),
    .B2(_092_),
    .ZN(_016_));
 AND2_X1 _288_ (.A1(_049_),
    .A2(\rx_shift_reg[0] ),
    .ZN(_093_));
 AND2_X1 _289_ (.A1(_037_),
    .A2(net1),
    .ZN(_094_));
 OR2_X1 _290_ (.A1(_043_),
    .A2(_055_),
    .ZN(_095_));
 OR4_X1 _291_ (.A1(_057_),
    .A2(_003_),
    .A3(_192_),
    .A4(_095_),
    .ZN(_096_));
 XNOR2_X2 _292_ (.A(_156_),
    .B(_157_),
    .ZN(_097_));
 NOR2_X1 _293_ (.A1(_055_),
    .A2(_205_),
    .ZN(_098_));
 NAND4_X1 _294_ (.A1(_199_),
    .A2(_196_),
    .A3(_097_),
    .A4(_098_),
    .ZN(_099_));
 NOR2_X1 _295_ (.A1(_195_),
    .A2(_208_),
    .ZN(_100_));
 AND2_X1 _296_ (.A1(_199_),
    .A2(_209_),
    .ZN(_101_));
 AND2_X1 _297_ (.A1(_195_),
    .A2(_208_),
    .ZN(_102_));
 NOR2_X1 _298_ (.A1(_199_),
    .A2(_209_),
    .ZN(_103_));
 AOI22_X1 _299_ (.A1(_100_),
    .A2(_101_),
    .B1(_102_),
    .B2(_103_),
    .ZN(_104_));
 NOR3_X1 _300_ (.A1(_096_),
    .A2(_099_),
    .A3(_104_),
    .ZN(_105_));
 MUX2_X1 _301_ (.A(_093_),
    .B(_094_),
    .S(_105_),
    .Z(_017_));
 AND2_X1 _302_ (.A1(_049_),
    .A2(\rx_shift_reg[1] ),
    .ZN(_106_));
 OR4_X1 _303_ (.A1(_057_),
    .A2(_196_),
    .A3(_095_),
    .A4(_097_),
    .ZN(_107_));
 NAND3_X2 _304_ (.A1(_098_),
    .A2(_102_),
    .A3(_103_),
    .ZN(_108_));
 NOR4_X1 _305_ (.A1(_056_),
    .A2(_063_),
    .A3(_107_),
    .A4(_108_),
    .ZN(_109_));
 MUX2_X1 _306_ (.A(_106_),
    .B(_094_),
    .S(_109_),
    .Z(_018_));
 AND2_X1 _307_ (.A1(_049_),
    .A2(\rx_shift_reg[2] ),
    .ZN(_110_));
 NOR4_X1 _308_ (.A1(_003_),
    .A2(_063_),
    .A3(_107_),
    .A4(_108_),
    .ZN(_111_));
 MUX2_X1 _309_ (.A(_110_),
    .B(_094_),
    .S(_111_),
    .Z(_019_));
 AND2_X1 _310_ (.A1(_037_),
    .A2(\rx_shift_reg[3] ),
    .ZN(_112_));
 NOR4_X1 _311_ (.A1(_056_),
    .A2(_192_),
    .A3(_107_),
    .A4(_108_),
    .ZN(_113_));
 MUX2_X1 _312_ (.A(_112_),
    .B(_094_),
    .S(_113_),
    .Z(_020_));
 AND2_X1 _313_ (.A1(_037_),
    .A2(\rx_shift_reg[4] ),
    .ZN(_114_));
 NOR4_X1 _314_ (.A1(_196_),
    .A2(_096_),
    .A3(_097_),
    .A4(_108_),
    .ZN(_115_));
 MUX2_X1 _315_ (.A(_114_),
    .B(_094_),
    .S(_115_),
    .Z(_021_));
 AND2_X1 _316_ (.A1(_037_),
    .A2(\rx_shift_reg[5] ),
    .ZN(_116_));
 NOR2_X1 _317_ (.A1(_043_),
    .A2(_055_),
    .ZN(_117_));
 NAND4_X2 _318_ (.A1(_040_),
    .A2(_073_),
    .A3(_117_),
    .A4(_097_),
    .ZN(_118_));
 NOR4_X1 _319_ (.A1(_056_),
    .A2(_063_),
    .A3(_108_),
    .A4(_118_),
    .ZN(_119_));
 MUX2_X1 _320_ (.A(_116_),
    .B(_094_),
    .S(_119_),
    .Z(_022_));
 AND2_X1 _321_ (.A1(_037_),
    .A2(\rx_shift_reg[6] ),
    .ZN(_120_));
 NOR4_X1 _322_ (.A1(_003_),
    .A2(_063_),
    .A3(_108_),
    .A4(_118_),
    .ZN(_121_));
 MUX2_X1 _323_ (.A(_120_),
    .B(_094_),
    .S(_121_),
    .Z(_023_));
 AND2_X1 _324_ (.A1(_037_),
    .A2(\rx_shift_reg[7] ),
    .ZN(_122_));
 NOR4_X1 _325_ (.A1(_056_),
    .A2(_192_),
    .A3(_108_),
    .A4(_118_),
    .ZN(_123_));
 MUX2_X1 _326_ (.A(_122_),
    .B(_094_),
    .S(_123_),
    .Z(_024_));
 NOR2_X1 _327_ (.A1(_039_),
    .A2(_052_),
    .ZN(_025_));
 MUX2_X1 _328_ (.A(_043_),
    .B(_004_),
    .S(_041_),
    .Z(_124_));
 AND4_X1 _329_ (.A1(_049_),
    .A2(_059_),
    .A3(_051_),
    .A4(_124_),
    .ZN(_026_));
 NAND2_X1 _330_ (.A1(_059_),
    .A2(net21),
    .ZN(_125_));
 NAND4_X1 _331_ (.A1(_049_),
    .A2(_052_),
    .A3(_054_),
    .A4(_125_),
    .ZN(_027_));
 OAI21_X1 _332_ (.A(_043_),
    .B1(_004_),
    .B2(_200_),
    .ZN(_126_));
 NAND2_X2 _333_ (.A1(_041_),
    .A2(_126_),
    .ZN(_127_));
 MUX2_X2 _334_ (.A(_041_),
    .B(net10),
    .S(_047_),
    .Z(_128_));
 AOI21_X1 _335_ (.A(net22),
    .B1(_127_),
    .B2(_128_),
    .ZN(_129_));
 AND2_X1 _336_ (.A1(_040_),
    .A2(_126_),
    .ZN(_130_));
 BUF_X2 _337_ (.A(_130_),
    .Z(_131_));
 MUX2_X2 _338_ (.A(_053_),
    .B(_057_),
    .S(_059_),
    .Z(_132_));
 MUX2_X1 _339_ (.A(net9),
    .B(\tx_shift_reg[6] ),
    .S(_041_),
    .Z(_133_));
 NOR3_X1 _340_ (.A1(_131_),
    .A2(_132_),
    .A3(_133_),
    .ZN(_134_));
 NOR3_X1 _341_ (.A1(_039_),
    .A2(_129_),
    .A3(_134_),
    .ZN(_028_));
 AOI21_X1 _342_ (.A(_076_),
    .B1(_059_),
    .B2(net23),
    .ZN(_135_));
 NAND2_X1 _343_ (.A1(_054_),
    .A2(_135_),
    .ZN(_029_));
 OAI21_X1 _344_ (.A(\tx_shift_reg[0] ),
    .B1(_131_),
    .B2(_132_),
    .ZN(_136_));
 NAND3_X1 _345_ (.A1(_057_),
    .A2(net2),
    .A3(_128_),
    .ZN(_137_));
 AOI21_X1 _346_ (.A(_076_),
    .B1(_136_),
    .B2(_137_),
    .ZN(_030_));
 AOI21_X1 _347_ (.A(\tx_shift_reg[1] ),
    .B1(_127_),
    .B2(_128_),
    .ZN(_138_));
 MUX2_X1 _348_ (.A(net3),
    .B(\tx_shift_reg[0] ),
    .S(_041_),
    .Z(_139_));
 NOR3_X1 _349_ (.A1(_131_),
    .A2(_132_),
    .A3(_139_),
    .ZN(_140_));
 NOR3_X1 _350_ (.A1(_039_),
    .A2(_138_),
    .A3(_140_),
    .ZN(_031_));
 AOI21_X1 _351_ (.A(\tx_shift_reg[2] ),
    .B1(_127_),
    .B2(_128_),
    .ZN(_141_));
 MUX2_X1 _352_ (.A(net4),
    .B(\tx_shift_reg[1] ),
    .S(_041_),
    .Z(_142_));
 NOR3_X1 _353_ (.A1(_131_),
    .A2(_132_),
    .A3(_142_),
    .ZN(_143_));
 NOR3_X1 _354_ (.A1(_039_),
    .A2(_141_),
    .A3(_143_),
    .ZN(_032_));
 AOI21_X1 _355_ (.A(\tx_shift_reg[3] ),
    .B1(_127_),
    .B2(_128_),
    .ZN(_144_));
 MUX2_X1 _356_ (.A(net5),
    .B(\tx_shift_reg[2] ),
    .S(_041_),
    .Z(_145_));
 NOR3_X1 _357_ (.A1(_131_),
    .A2(_132_),
    .A3(_145_),
    .ZN(_146_));
 NOR3_X1 _358_ (.A1(_039_),
    .A2(_144_),
    .A3(_146_),
    .ZN(_033_));
 AOI21_X1 _359_ (.A(\tx_shift_reg[4] ),
    .B1(_127_),
    .B2(_128_),
    .ZN(_147_));
 MUX2_X1 _360_ (.A(net6),
    .B(\tx_shift_reg[3] ),
    .S(_040_),
    .Z(_148_));
 NOR3_X1 _361_ (.A1(_131_),
    .A2(_132_),
    .A3(_148_),
    .ZN(_149_));
 NOR3_X1 _362_ (.A1(_039_),
    .A2(_147_),
    .A3(_149_),
    .ZN(_034_));
 AOI21_X1 _363_ (.A(\tx_shift_reg[5] ),
    .B1(_127_),
    .B2(_128_),
    .ZN(_150_));
 MUX2_X1 _364_ (.A(net7),
    .B(\tx_shift_reg[4] ),
    .S(_040_),
    .Z(_151_));
 NOR3_X1 _365_ (.A1(_131_),
    .A2(_132_),
    .A3(_151_),
    .ZN(_152_));
 NOR3_X1 _366_ (.A1(_039_),
    .A2(_150_),
    .A3(_152_),
    .ZN(_035_));
 AOI21_X1 _367_ (.A(\tx_shift_reg[6] ),
    .B1(_127_),
    .B2(_128_),
    .ZN(_153_));
 MUX2_X1 _368_ (.A(net8),
    .B(\tx_shift_reg[5] ),
    .S(_040_),
    .Z(_154_));
 NOR3_X1 _369_ (.A1(_131_),
    .A2(_132_),
    .A3(_154_),
    .ZN(_155_));
 NOR3_X1 _370_ (.A1(_039_),
    .A2(_153_),
    .A3(_155_),
    .ZN(_036_));
 HA_X1 _371_ (.A(\bit_counter[0] ),
    .B(\bit_counter[1] ),
    .CO(_191_),
    .S(_192_));
 HA_X1 _372_ (.A(_193_),
    .B(_194_),
    .CO(_195_),
    .S(_196_));
 HA_X1 _373_ (.A(_193_),
    .B(_197_),
    .CO(_198_),
    .S(_199_));
 HA_X1 _374_ (.A(_193_),
    .B(_197_),
    .CO(_200_),
    .S(_201_));
 HA_X1 _375_ (.A(\bit_counter[3] ),
    .B(_197_),
    .CO(_202_),
    .S(_203_));
 HA_X1 _376_ (.A(\bit_counter[3] ),
    .B(_204_),
    .CO(_205_),
    .S(_206_));
 HA_X1 _377_ (.A(_193_),
    .B(_207_),
    .CO(_208_),
    .S(_209_));
 DFF_X1 \bit_counter[0]$_SDFFE_PN0P_  (.D(_005_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\bit_counter[0] ),
    .QN(_003_));
 DFF_X1 \bit_counter[1]$_SDFFE_PN0P_  (.D(_006_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\bit_counter[1] ),
    .QN(_187_));
 DFF_X1 \bit_counter[2]$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\bit_counter[2] ),
    .QN(_186_));
 DFF_X2 \bit_counter[3]$_SDFFE_PN0P_  (.D(_008_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\bit_counter[3] ),
    .QN(_193_));
 DFF_X1 \rx_data[0]$_SDFFE_PN0P_  (.D(_009_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net11),
    .QN(_185_));
 DFF_X1 \rx_data[1]$_SDFFE_PN0P_  (.D(_010_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net12),
    .QN(_184_));
 DFF_X1 \rx_data[2]$_SDFFE_PN0P_  (.D(_011_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net13),
    .QN(_183_));
 DFF_X1 \rx_data[3]$_SDFFE_PN0P_  (.D(_012_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net14),
    .QN(_182_));
 DFF_X1 \rx_data[4]$_SDFFE_PN0P_  (.D(_013_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net15),
    .QN(_181_));
 DFF_X1 \rx_data[5]$_SDFFE_PN0P_  (.D(_014_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net16),
    .QN(_180_));
 DFF_X1 \rx_data[6]$_SDFFE_PN0P_  (.D(_015_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net17),
    .QN(_179_));
 DFF_X1 \rx_data[7]$_SDFFE_PN0P_  (.D(_016_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net18),
    .QN(_178_));
 DFF_X1 \rx_shift_reg[0]$_SDFFE_PN0P_  (.D(_017_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\rx_shift_reg[0] ),
    .QN(_177_));
 DFF_X1 \rx_shift_reg[1]$_SDFFE_PN0P_  (.D(_018_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\rx_shift_reg[1] ),
    .QN(_176_));
 DFF_X1 \rx_shift_reg[2]$_SDFFE_PN0P_  (.D(_019_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\rx_shift_reg[2] ),
    .QN(_175_));
 DFF_X1 \rx_shift_reg[3]$_SDFFE_PN0P_  (.D(_020_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\rx_shift_reg[3] ),
    .QN(_174_));
 DFF_X1 \rx_shift_reg[4]$_SDFFE_PN0P_  (.D(_021_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\rx_shift_reg[4] ),
    .QN(_173_));
 DFF_X1 \rx_shift_reg[5]$_SDFFE_PN0P_  (.D(_022_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\rx_shift_reg[5] ),
    .QN(_172_));
 DFF_X1 \rx_shift_reg[6]$_SDFFE_PN0P_  (.D(_023_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\rx_shift_reg[6] ),
    .QN(_171_));
 DFF_X1 \rx_shift_reg[7]$_SDFFE_PN0P_  (.D(_024_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\rx_shift_reg[7] ),
    .QN(_170_));
 DFF_X1 \rx_valid$_SDFF_PN0_  (.D(_025_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net19),
    .QN(_169_));
 DFF_X1 \spi_clk$_SDFFE_PN0P_  (.D(_026_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net20),
    .QN(_004_));
 DFF_X1 \spi_cs_n$_SDFFE_PN1P_  (.D(_027_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net21),
    .QN(_168_));
 DFF_X1 \spi_mosi$_SDFFE_PN0P_  (.D(_028_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net22),
    .QN(_188_));
 DFF_X1 \state[0]$_DFF_P_  (.D(_001_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\state[0] ),
    .QN(_189_));
 DFF_X1 \state[1]$_DFF_P_  (.D(_000_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\state[1] ),
    .QN(_190_));
 DFF_X1 \state[2]$_DFF_P_  (.D(_002_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\state[2] ),
    .QN(_167_));
 DFF_X1 \tx_ready$_SDFFE_PN1P_  (.D(_029_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net23),
    .QN(_166_));
 DFF_X1 \tx_shift_reg[0]$_SDFFE_PN0P_  (.D(_030_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\tx_shift_reg[0] ),
    .QN(_165_));
 DFF_X1 \tx_shift_reg[1]$_SDFFE_PN0P_  (.D(_031_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\tx_shift_reg[1] ),
    .QN(_164_));
 DFF_X1 \tx_shift_reg[2]$_SDFFE_PN0P_  (.D(_032_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\tx_shift_reg[2] ),
    .QN(_163_));
 DFF_X1 \tx_shift_reg[3]$_SDFFE_PN0P_  (.D(_033_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\tx_shift_reg[3] ),
    .QN(_162_));
 DFF_X1 \tx_shift_reg[4]$_SDFFE_PN0P_  (.D(_034_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\tx_shift_reg[4] ),
    .QN(_161_));
 DFF_X1 \tx_shift_reg[5]$_SDFFE_PN0P_  (.D(_035_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\tx_shift_reg[5] ),
    .QN(_160_));
 DFF_X1 \tx_shift_reg[6]$_SDFFE_PN0P_  (.D(_036_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\tx_shift_reg[6] ),
    .QN(_159_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_47 ();
 BUF_X1 input1 (.A(spi_miso),
    .Z(net1));
 BUF_X1 input2 (.A(tx_data[0]),
    .Z(net2));
 BUF_X1 input3 (.A(tx_data[1]),
    .Z(net3));
 BUF_X1 input4 (.A(tx_data[2]),
    .Z(net4));
 BUF_X1 input5 (.A(tx_data[3]),
    .Z(net5));
 BUF_X1 input6 (.A(tx_data[4]),
    .Z(net6));
 BUF_X1 input7 (.A(tx_data[5]),
    .Z(net7));
 BUF_X1 input8 (.A(tx_data[6]),
    .Z(net8));
 BUF_X1 input9 (.A(tx_data[7]),
    .Z(net9));
 BUF_X1 input10 (.A(tx_valid),
    .Z(net10));
 BUF_X1 output11 (.A(net11),
    .Z(rx_data[0]));
 BUF_X1 output12 (.A(net12),
    .Z(rx_data[1]));
 BUF_X1 output13 (.A(net13),
    .Z(rx_data[2]));
 BUF_X1 output14 (.A(net14),
    .Z(rx_data[3]));
 BUF_X1 output15 (.A(net15),
    .Z(rx_data[4]));
 BUF_X1 output16 (.A(net16),
    .Z(rx_data[5]));
 BUF_X1 output17 (.A(net17),
    .Z(rx_data[6]));
 BUF_X1 output18 (.A(net18),
    .Z(rx_data[7]));
 BUF_X1 output19 (.A(net19),
    .Z(rx_valid));
 BUF_X1 output20 (.A(net20),
    .Z(spi_clk));
 BUF_X1 output21 (.A(net21),
    .Z(spi_cs_n));
 BUF_X1 output22 (.A(net22),
    .Z(spi_mosi));
 BUF_X1 output23 (.A(net23),
    .Z(tx_ready));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 CLKBUF_X3 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 CLKBUF_X3 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 CLKBUF_X3 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 INV_X2 clkload0 (.A(clknet_2_0__leaf_clk));
 INV_X1 clkload1 (.A(clknet_2_2__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X16 FILLER_0_33 ();
 FILLCELL_X8 FILLER_0_49 ();
 FILLCELL_X2 FILLER_0_57 ();
 FILLCELL_X1 FILLER_0_59 ();
 FILLCELL_X2 FILLER_0_63 ();
 FILLCELL_X2 FILLER_0_68 ();
 FILLCELL_X1 FILLER_0_116 ();
 FILLCELL_X4 FILLER_0_125 ();
 FILLCELL_X1 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_147 ();
 FILLCELL_X1 FILLER_0_179 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X2 FILLER_1_76 ();
 FILLCELL_X1 FILLER_1_78 ();
 FILLCELL_X1 FILLER_1_107 ();
 FILLCELL_X1 FILLER_1_112 ();
 FILLCELL_X32 FILLER_1_138 ();
 FILLCELL_X8 FILLER_1_170 ();
 FILLCELL_X2 FILLER_1_178 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X16 FILLER_2_33 ();
 FILLCELL_X4 FILLER_2_49 ();
 FILLCELL_X2 FILLER_2_53 ();
 FILLCELL_X1 FILLER_2_55 ();
 FILLCELL_X4 FILLER_2_81 ();
 FILLCELL_X2 FILLER_2_85 ();
 FILLCELL_X1 FILLER_2_87 ();
 FILLCELL_X8 FILLER_2_92 ();
 FILLCELL_X4 FILLER_2_100 ();
 FILLCELL_X2 FILLER_2_104 ();
 FILLCELL_X1 FILLER_2_106 ();
 FILLCELL_X2 FILLER_2_110 ();
 FILLCELL_X1 FILLER_2_112 ();
 FILLCELL_X32 FILLER_2_124 ();
 FILLCELL_X16 FILLER_2_156 ();
 FILLCELL_X8 FILLER_2_172 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X16 FILLER_3_33 ();
 FILLCELL_X8 FILLER_3_49 ();
 FILLCELL_X2 FILLER_3_57 ();
 FILLCELL_X16 FILLER_3_84 ();
 FILLCELL_X2 FILLER_3_100 ();
 FILLCELL_X1 FILLER_3_102 ();
 FILLCELL_X32 FILLER_3_144 ();
 FILLCELL_X4 FILLER_3_176 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X16 FILLER_4_33 ();
 FILLCELL_X2 FILLER_4_49 ();
 FILLCELL_X1 FILLER_4_51 ();
 FILLCELL_X1 FILLER_4_80 ();
 FILLCELL_X1 FILLER_4_89 ();
 FILLCELL_X2 FILLER_4_103 ();
 FILLCELL_X32 FILLER_4_130 ();
 FILLCELL_X16 FILLER_4_162 ();
 FILLCELL_X2 FILLER_4_178 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X8 FILLER_5_65 ();
 FILLCELL_X4 FILLER_5_73 ();
 FILLCELL_X2 FILLER_5_77 ();
 FILLCELL_X1 FILLER_5_79 ();
 FILLCELL_X1 FILLER_5_105 ();
 FILLCELL_X2 FILLER_5_119 ();
 FILLCELL_X16 FILLER_5_124 ();
 FILLCELL_X8 FILLER_5_140 ();
 FILLCELL_X4 FILLER_5_148 ();
 FILLCELL_X1 FILLER_5_152 ();
 FILLCELL_X8 FILLER_5_170 ();
 FILLCELL_X2 FILLER_5_178 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X2 FILLER_6_86 ();
 FILLCELL_X1 FILLER_6_88 ();
 FILLCELL_X1 FILLER_6_93 ();
 FILLCELL_X2 FILLER_6_115 ();
 FILLCELL_X8 FILLER_6_120 ();
 FILLCELL_X1 FILLER_6_128 ();
 FILLCELL_X1 FILLER_6_146 ();
 FILLCELL_X8 FILLER_6_160 ();
 FILLCELL_X2 FILLER_6_168 ();
 FILLCELL_X4 FILLER_6_173 ();
 FILLCELL_X2 FILLER_6_177 ();
 FILLCELL_X1 FILLER_6_179 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X8 FILLER_7_65 ();
 FILLCELL_X2 FILLER_7_73 ();
 FILLCELL_X1 FILLER_7_75 ();
 FILLCELL_X2 FILLER_7_83 ();
 FILLCELL_X1 FILLER_7_87 ();
 FILLCELL_X2 FILLER_7_113 ();
 FILLCELL_X1 FILLER_7_115 ();
 FILLCELL_X8 FILLER_7_122 ();
 FILLCELL_X2 FILLER_7_130 ();
 FILLCELL_X1 FILLER_7_132 ();
 FILLCELL_X8 FILLER_7_137 ();
 FILLCELL_X1 FILLER_7_145 ();
 FILLCELL_X16 FILLER_7_157 ();
 FILLCELL_X4 FILLER_7_173 ();
 FILLCELL_X2 FILLER_7_177 ();
 FILLCELL_X1 FILLER_7_179 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X8 FILLER_8_65 ();
 FILLCELL_X1 FILLER_8_73 ();
 FILLCELL_X1 FILLER_8_92 ();
 FILLCELL_X2 FILLER_8_114 ();
 FILLCELL_X8 FILLER_8_122 ();
 FILLCELL_X8 FILLER_8_135 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X16 FILLER_9_33 ();
 FILLCELL_X8 FILLER_9_49 ();
 FILLCELL_X4 FILLER_9_57 ();
 FILLCELL_X2 FILLER_9_61 ();
 FILLCELL_X1 FILLER_9_63 ();
 FILLCELL_X8 FILLER_9_68 ();
 FILLCELL_X4 FILLER_9_76 ();
 FILLCELL_X2 FILLER_9_90 ();
 FILLCELL_X4 FILLER_9_107 ();
 FILLCELL_X2 FILLER_9_114 ();
 FILLCELL_X1 FILLER_9_116 ();
 FILLCELL_X1 FILLER_9_121 ();
 FILLCELL_X8 FILLER_9_143 ();
 FILLCELL_X4 FILLER_9_151 ();
 FILLCELL_X2 FILLER_9_155 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X16 FILLER_10_33 ();
 FILLCELL_X4 FILLER_10_49 ();
 FILLCELL_X2 FILLER_10_53 ();
 FILLCELL_X1 FILLER_10_55 ();
 FILLCELL_X8 FILLER_10_75 ();
 FILLCELL_X1 FILLER_10_83 ();
 FILLCELL_X1 FILLER_10_89 ();
 FILLCELL_X1 FILLER_10_100 ();
 FILLCELL_X2 FILLER_10_114 ();
 FILLCELL_X2 FILLER_10_119 ();
 FILLCELL_X2 FILLER_10_128 ();
 FILLCELL_X2 FILLER_10_156 ();
 FILLCELL_X4 FILLER_10_162 ();
 FILLCELL_X1 FILLER_10_166 ();
 FILLCELL_X4 FILLER_10_170 ();
 FILLCELL_X1 FILLER_10_174 ();
 FILLCELL_X2 FILLER_10_178 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X8 FILLER_11_65 ();
 FILLCELL_X2 FILLER_11_73 ();
 FILLCELL_X1 FILLER_11_75 ();
 FILLCELL_X2 FILLER_11_83 ();
 FILLCELL_X1 FILLER_11_85 ();
 FILLCELL_X4 FILLER_11_89 ();
 FILLCELL_X2 FILLER_11_93 ();
 FILLCELL_X1 FILLER_11_95 ();
 FILLCELL_X1 FILLER_11_130 ();
 FILLCELL_X16 FILLER_11_138 ();
 FILLCELL_X2 FILLER_11_154 ();
 FILLCELL_X8 FILLER_11_159 ();
 FILLCELL_X4 FILLER_11_167 ();
 FILLCELL_X2 FILLER_11_171 ();
 FILLCELL_X1 FILLER_11_173 ();
 FILLCELL_X2 FILLER_11_177 ();
 FILLCELL_X1 FILLER_11_179 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X16 FILLER_12_33 ();
 FILLCELL_X8 FILLER_12_49 ();
 FILLCELL_X4 FILLER_12_57 ();
 FILLCELL_X2 FILLER_12_61 ();
 FILLCELL_X2 FILLER_12_87 ();
 FILLCELL_X4 FILLER_12_96 ();
 FILLCELL_X2 FILLER_12_100 ();
 FILLCELL_X8 FILLER_12_104 ();
 FILLCELL_X2 FILLER_12_112 ();
 FILLCELL_X4 FILLER_12_130 ();
 FILLCELL_X8 FILLER_12_146 ();
 FILLCELL_X2 FILLER_12_178 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X4 FILLER_13_65 ();
 FILLCELL_X2 FILLER_13_69 ();
 FILLCELL_X1 FILLER_13_71 ();
 FILLCELL_X2 FILLER_13_79 ();
 FILLCELL_X8 FILLER_13_98 ();
 FILLCELL_X4 FILLER_13_106 ();
 FILLCELL_X2 FILLER_13_110 ();
 FILLCELL_X1 FILLER_13_112 ();
 FILLCELL_X1 FILLER_13_119 ();
 FILLCELL_X8 FILLER_13_125 ();
 FILLCELL_X2 FILLER_13_133 ();
 FILLCELL_X1 FILLER_13_139 ();
 FILLCELL_X1 FILLER_13_157 ();
 FILLCELL_X2 FILLER_13_175 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X16 FILLER_14_33 ();
 FILLCELL_X8 FILLER_14_49 ();
 FILLCELL_X4 FILLER_14_57 ();
 FILLCELL_X2 FILLER_14_61 ();
 FILLCELL_X1 FILLER_14_63 ();
 FILLCELL_X4 FILLER_14_68 ();
 FILLCELL_X1 FILLER_14_72 ();
 FILLCELL_X2 FILLER_14_80 ();
 FILLCELL_X1 FILLER_14_82 ();
 FILLCELL_X2 FILLER_14_86 ();
 FILLCELL_X1 FILLER_14_88 ();
 FILLCELL_X1 FILLER_14_93 ();
 FILLCELL_X4 FILLER_14_104 ();
 FILLCELL_X2 FILLER_14_108 ();
 FILLCELL_X1 FILLER_14_110 ();
 FILLCELL_X8 FILLER_14_122 ();
 FILLCELL_X1 FILLER_14_130 ();
 FILLCELL_X8 FILLER_14_146 ();
 FILLCELL_X2 FILLER_14_154 ();
 FILLCELL_X2 FILLER_14_163 ();
 FILLCELL_X8 FILLER_14_168 ();
 FILLCELL_X4 FILLER_14_176 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X16 FILLER_15_33 ();
 FILLCELL_X8 FILLER_15_49 ();
 FILLCELL_X1 FILLER_15_57 ();
 FILLCELL_X2 FILLER_15_86 ();
 FILLCELL_X1 FILLER_15_88 ();
 FILLCELL_X8 FILLER_15_103 ();
 FILLCELL_X4 FILLER_15_111 ();
 FILLCELL_X2 FILLER_15_115 ();
 FILLCELL_X1 FILLER_15_119 ();
 FILLCELL_X2 FILLER_15_125 ();
 FILLCELL_X1 FILLER_15_127 ();
 FILLCELL_X2 FILLER_15_152 ();
 FILLCELL_X1 FILLER_15_161 ();
 FILLCELL_X2 FILLER_15_166 ();
 FILLCELL_X4 FILLER_15_171 ();
 FILLCELL_X2 FILLER_15_175 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X16 FILLER_16_65 ();
 FILLCELL_X8 FILLER_16_98 ();
 FILLCELL_X2 FILLER_16_106 ();
 FILLCELL_X1 FILLER_16_108 ();
 FILLCELL_X2 FILLER_16_129 ();
 FILLCELL_X2 FILLER_16_155 ();
 FILLCELL_X1 FILLER_16_157 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X8 FILLER_17_97 ();
 FILLCELL_X1 FILLER_17_105 ();
 FILLCELL_X4 FILLER_17_108 ();
 FILLCELL_X1 FILLER_17_112 ();
 FILLCELL_X8 FILLER_17_120 ();
 FILLCELL_X2 FILLER_17_128 ();
 FILLCELL_X8 FILLER_17_137 ();
 FILLCELL_X4 FILLER_17_145 ();
 FILLCELL_X8 FILLER_17_172 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X4 FILLER_18_123 ();
 FILLCELL_X2 FILLER_18_127 ();
 FILLCELL_X2 FILLER_18_153 ();
 FILLCELL_X1 FILLER_18_155 ();
 FILLCELL_X16 FILLER_18_160 ();
 FILLCELL_X4 FILLER_18_176 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X8 FILLER_19_97 ();
 FILLCELL_X2 FILLER_19_105 ();
 FILLCELL_X4 FILLER_19_117 ();
 FILLCELL_X1 FILLER_19_121 ();
 FILLCELL_X32 FILLER_19_133 ();
 FILLCELL_X8 FILLER_19_165 ();
 FILLCELL_X4 FILLER_19_173 ();
 FILLCELL_X2 FILLER_19_177 ();
 FILLCELL_X1 FILLER_19_179 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X16 FILLER_20_65 ();
 FILLCELL_X8 FILLER_20_81 ();
 FILLCELL_X4 FILLER_20_89 ();
 FILLCELL_X2 FILLER_20_93 ();
 FILLCELL_X1 FILLER_20_95 ();
 FILLCELL_X2 FILLER_20_120 ();
 FILLCELL_X1 FILLER_20_122 ();
 FILLCELL_X32 FILLER_20_143 ();
 FILLCELL_X4 FILLER_20_175 ();
 FILLCELL_X1 FILLER_20_179 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X8 FILLER_21_97 ();
 FILLCELL_X4 FILLER_21_105 ();
 FILLCELL_X2 FILLER_21_109 ();
 FILLCELL_X1 FILLER_21_111 ();
 FILLCELL_X2 FILLER_21_116 ();
 FILLCELL_X1 FILLER_21_118 ();
 FILLCELL_X8 FILLER_21_126 ();
 FILLCELL_X4 FILLER_21_134 ();
 FILLCELL_X2 FILLER_21_138 ();
 FILLCELL_X32 FILLER_21_147 ();
 FILLCELL_X1 FILLER_21_179 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X16 FILLER_22_65 ();
 FILLCELL_X8 FILLER_22_81 ();
 FILLCELL_X4 FILLER_22_89 ();
 FILLCELL_X1 FILLER_22_93 ();
 FILLCELL_X1 FILLER_22_114 ();
 FILLCELL_X2 FILLER_22_132 ();
 FILLCELL_X16 FILLER_22_151 ();
 FILLCELL_X8 FILLER_22_167 ();
 FILLCELL_X4 FILLER_22_175 ();
 FILLCELL_X1 FILLER_22_179 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X2 FILLER_23_97 ();
 FILLCELL_X1 FILLER_23_99 ();
 FILLCELL_X2 FILLER_23_104 ();
 FILLCELL_X1 FILLER_23_106 ();
 FILLCELL_X1 FILLER_23_113 ();
 FILLCELL_X4 FILLER_23_118 ();
 FILLCELL_X2 FILLER_23_122 ();
 FILLCELL_X16 FILLER_23_127 ();
 FILLCELL_X2 FILLER_23_143 ();
 FILLCELL_X32 FILLER_23_148 ();
endmodule
