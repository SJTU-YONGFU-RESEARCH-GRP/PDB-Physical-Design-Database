module parameterized_cam (clk,
    compare_enable,
    match,
    rst_n,
    valid,
    write_enable,
    compare_data,
    match_addr,
    write_addr,
    write_data);
 input clk;
 input compare_enable;
 output match;
 input rst_n;
 output valid;
 input write_enable;
 input [7:0] compare_data;
 output [3:0] match_addr;
 input [3:0] write_addr;
 input [7:0] write_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire _433_;
 wire _434_;
 wire _435_;
 wire _436_;
 wire _437_;
 wire _438_;
 wire _439_;
 wire _440_;
 wire _441_;
 wire _442_;
 wire _443_;
 wire _444_;
 wire _445_;
 wire _446_;
 wire _447_;
 wire _448_;
 wire _449_;
 wire _450_;
 wire _451_;
 wire _452_;
 wire _453_;
 wire _454_;
 wire _455_;
 wire _456_;
 wire _457_;
 wire _458_;
 wire _459_;
 wire _460_;
 wire _461_;
 wire _462_;
 wire _463_;
 wire _464_;
 wire _465_;
 wire _466_;
 wire _467_;
 wire _468_;
 wire _469_;
 wire _470_;
 wire \cam_memory[0][0] ;
 wire \cam_memory[0][1] ;
 wire \cam_memory[0][2] ;
 wire \cam_memory[0][3] ;
 wire \cam_memory[0][4] ;
 wire \cam_memory[0][5] ;
 wire \cam_memory[0][6] ;
 wire \cam_memory[0][7] ;
 wire \cam_memory[10][0] ;
 wire \cam_memory[10][1] ;
 wire \cam_memory[10][2] ;
 wire \cam_memory[10][3] ;
 wire \cam_memory[10][4] ;
 wire \cam_memory[10][5] ;
 wire \cam_memory[10][6] ;
 wire \cam_memory[10][7] ;
 wire \cam_memory[11][0] ;
 wire \cam_memory[11][1] ;
 wire \cam_memory[11][2] ;
 wire \cam_memory[11][3] ;
 wire \cam_memory[11][4] ;
 wire \cam_memory[11][5] ;
 wire \cam_memory[11][6] ;
 wire \cam_memory[11][7] ;
 wire \cam_memory[12][0] ;
 wire \cam_memory[12][1] ;
 wire \cam_memory[12][2] ;
 wire \cam_memory[12][3] ;
 wire \cam_memory[12][4] ;
 wire \cam_memory[12][5] ;
 wire \cam_memory[12][6] ;
 wire \cam_memory[12][7] ;
 wire \cam_memory[13][0] ;
 wire \cam_memory[13][1] ;
 wire \cam_memory[13][2] ;
 wire \cam_memory[13][3] ;
 wire \cam_memory[13][4] ;
 wire \cam_memory[13][5] ;
 wire \cam_memory[13][6] ;
 wire \cam_memory[13][7] ;
 wire \cam_memory[14][0] ;
 wire \cam_memory[14][1] ;
 wire \cam_memory[14][2] ;
 wire \cam_memory[14][3] ;
 wire \cam_memory[14][4] ;
 wire \cam_memory[14][5] ;
 wire \cam_memory[14][6] ;
 wire \cam_memory[14][7] ;
 wire \cam_memory[15][0] ;
 wire \cam_memory[15][1] ;
 wire \cam_memory[15][2] ;
 wire \cam_memory[15][3] ;
 wire \cam_memory[15][4] ;
 wire \cam_memory[15][5] ;
 wire \cam_memory[15][6] ;
 wire \cam_memory[15][7] ;
 wire \cam_memory[1][0] ;
 wire \cam_memory[1][1] ;
 wire \cam_memory[1][2] ;
 wire \cam_memory[1][3] ;
 wire \cam_memory[1][4] ;
 wire \cam_memory[1][5] ;
 wire \cam_memory[1][6] ;
 wire \cam_memory[1][7] ;
 wire \cam_memory[2][0] ;
 wire \cam_memory[2][1] ;
 wire \cam_memory[2][2] ;
 wire \cam_memory[2][3] ;
 wire \cam_memory[2][4] ;
 wire \cam_memory[2][5] ;
 wire \cam_memory[2][6] ;
 wire \cam_memory[2][7] ;
 wire \cam_memory[3][0] ;
 wire \cam_memory[3][1] ;
 wire \cam_memory[3][2] ;
 wire \cam_memory[3][3] ;
 wire \cam_memory[3][4] ;
 wire \cam_memory[3][5] ;
 wire \cam_memory[3][6] ;
 wire \cam_memory[3][7] ;
 wire \cam_memory[4][0] ;
 wire \cam_memory[4][1] ;
 wire \cam_memory[4][2] ;
 wire \cam_memory[4][3] ;
 wire \cam_memory[4][4] ;
 wire \cam_memory[4][5] ;
 wire \cam_memory[4][6] ;
 wire \cam_memory[4][7] ;
 wire \cam_memory[5][0] ;
 wire \cam_memory[5][1] ;
 wire \cam_memory[5][2] ;
 wire \cam_memory[5][3] ;
 wire \cam_memory[5][4] ;
 wire \cam_memory[5][5] ;
 wire \cam_memory[5][6] ;
 wire \cam_memory[5][7] ;
 wire \cam_memory[6][0] ;
 wire \cam_memory[6][1] ;
 wire \cam_memory[6][2] ;
 wire \cam_memory[6][3] ;
 wire \cam_memory[6][4] ;
 wire \cam_memory[6][5] ;
 wire \cam_memory[6][6] ;
 wire \cam_memory[6][7] ;
 wire \cam_memory[7][0] ;
 wire \cam_memory[7][1] ;
 wire \cam_memory[7][2] ;
 wire \cam_memory[7][3] ;
 wire \cam_memory[7][4] ;
 wire \cam_memory[7][5] ;
 wire \cam_memory[7][6] ;
 wire \cam_memory[7][7] ;
 wire \cam_memory[8][0] ;
 wire \cam_memory[8][1] ;
 wire \cam_memory[8][2] ;
 wire \cam_memory[8][3] ;
 wire \cam_memory[8][4] ;
 wire \cam_memory[8][5] ;
 wire \cam_memory[8][6] ;
 wire \cam_memory[8][7] ;
 wire \cam_memory[9][0] ;
 wire \cam_memory[9][1] ;
 wire \cam_memory[9][2] ;
 wire \cam_memory[9][3] ;
 wire \cam_memory[9][4] ;
 wire \cam_memory[9][5] ;
 wire \cam_memory[9][6] ;
 wire \cam_memory[9][7] ;
 wire \valid_bits[0] ;
 wire \valid_bits[10] ;
 wire \valid_bits[11] ;
 wire \valid_bits[12] ;
 wire \valid_bits[13] ;
 wire \valid_bits[14] ;
 wire \valid_bits[15] ;
 wire \valid_bits[1] ;
 wire \valid_bits[2] ;
 wire \valid_bits[3] ;
 wire \valid_bits[4] ;
 wire \valid_bits[5] ;
 wire \valid_bits[6] ;
 wire \valid_bits[7] ;
 wire \valid_bits[8] ;
 wire \valid_bits[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net20;
 wire net21;

 sky130_fd_sc_hd__buf_6 _471_ (.A(compare_data[1]),
    .X(_149_));
 sky130_fd_sc_hd__xnor2_1 _472_ (.A(_149_),
    .B(\cam_memory[14][1] ),
    .Y(_150_));
 sky130_fd_sc_hd__nand2_1 _473_ (.A(\valid_bits[14] ),
    .B(_150_),
    .Y(_151_));
 sky130_fd_sc_hd__buf_6 _474_ (.A(compare_data[6]),
    .X(_152_));
 sky130_fd_sc_hd__xnor2_1 _475_ (.A(_152_),
    .B(\cam_memory[14][6] ),
    .Y(_153_));
 sky130_fd_sc_hd__buf_6 _476_ (.A(compare_data[5]),
    .X(_154_));
 sky130_fd_sc_hd__xnor2_1 _477_ (.A(_154_),
    .B(\cam_memory[14][5] ),
    .Y(_155_));
 sky130_fd_sc_hd__buf_6 _478_ (.A(compare_data[7]),
    .X(_156_));
 sky130_fd_sc_hd__xnor2_1 _479_ (.A(_156_),
    .B(\cam_memory[14][7] ),
    .Y(_157_));
 sky130_fd_sc_hd__nand3_1 _480_ (.A(_153_),
    .B(_155_),
    .C(_157_),
    .Y(_158_));
 sky130_fd_sc_hd__buf_6 _481_ (.A(compare_data[4]),
    .X(_159_));
 sky130_fd_sc_hd__xnor2_1 _482_ (.A(_159_),
    .B(\cam_memory[14][4] ),
    .Y(_160_));
 sky130_fd_sc_hd__buf_6 _483_ (.A(compare_data[2]),
    .X(_161_));
 sky130_fd_sc_hd__xnor2_1 _484_ (.A(_161_),
    .B(\cam_memory[14][2] ),
    .Y(_162_));
 sky130_fd_sc_hd__buf_6 _485_ (.A(compare_data[3]),
    .X(_163_));
 sky130_fd_sc_hd__xnor2_1 _486_ (.A(_163_),
    .B(\cam_memory[14][3] ),
    .Y(_164_));
 sky130_fd_sc_hd__buf_6 _487_ (.A(compare_data[0]),
    .X(_165_));
 sky130_fd_sc_hd__xnor2_1 _488_ (.A(_165_),
    .B(\cam_memory[14][0] ),
    .Y(_166_));
 sky130_fd_sc_hd__nand4_1 _489_ (.A(_160_),
    .B(_162_),
    .C(_164_),
    .D(_166_),
    .Y(_167_));
 sky130_fd_sc_hd__nor3_2 _490_ (.A(_151_),
    .B(_158_),
    .C(_167_),
    .Y(_168_));
 sky130_fd_sc_hd__buf_16 _491_ (.A(_165_),
    .X(_169_));
 sky130_fd_sc_hd__xnor2_1 _492_ (.A(_169_),
    .B(\cam_memory[15][0] ),
    .Y(_170_));
 sky130_fd_sc_hd__nand2_1 _493_ (.A(\valid_bits[15] ),
    .B(_170_),
    .Y(_171_));
 sky130_fd_sc_hd__buf_8 _494_ (.A(_154_),
    .X(_172_));
 sky130_fd_sc_hd__xnor2_1 _495_ (.A(_172_),
    .B(\cam_memory[15][5] ),
    .Y(_173_));
 sky130_fd_sc_hd__buf_8 _496_ (.A(_152_),
    .X(_174_));
 sky130_fd_sc_hd__xnor2_1 _497_ (.A(_174_),
    .B(\cam_memory[15][6] ),
    .Y(_175_));
 sky130_fd_sc_hd__buf_16 _498_ (.A(_156_),
    .X(_176_));
 sky130_fd_sc_hd__xnor2_1 _499_ (.A(_176_),
    .B(\cam_memory[15][7] ),
    .Y(_177_));
 sky130_fd_sc_hd__nand3_1 _500_ (.A(_173_),
    .B(_175_),
    .C(_177_),
    .Y(_178_));
 sky130_fd_sc_hd__buf_6 _501_ (.A(_159_),
    .X(_179_));
 sky130_fd_sc_hd__xnor2_1 _502_ (.A(_179_),
    .B(\cam_memory[15][4] ),
    .Y(_180_));
 sky130_fd_sc_hd__buf_6 _503_ (.A(_161_),
    .X(_181_));
 sky130_fd_sc_hd__xnor2_1 _504_ (.A(_181_),
    .B(\cam_memory[15][2] ),
    .Y(_182_));
 sky130_fd_sc_hd__buf_6 _505_ (.A(_149_),
    .X(_183_));
 sky130_fd_sc_hd__xnor2_1 _506_ (.A(_183_),
    .B(\cam_memory[15][1] ),
    .Y(_184_));
 sky130_fd_sc_hd__buf_6 _507_ (.A(_163_),
    .X(_185_));
 sky130_fd_sc_hd__xnor2_1 _508_ (.A(_185_),
    .B(\cam_memory[15][3] ),
    .Y(_186_));
 sky130_fd_sc_hd__nand4_1 _509_ (.A(_180_),
    .B(_182_),
    .C(_184_),
    .D(_186_),
    .Y(_187_));
 sky130_fd_sc_hd__nor3_1 _510_ (.A(_171_),
    .B(_178_),
    .C(_187_),
    .Y(_188_));
 sky130_fd_sc_hd__xnor2_1 _511_ (.A(_183_),
    .B(\cam_memory[12][1] ),
    .Y(_189_));
 sky130_fd_sc_hd__nand2_1 _512_ (.A(\valid_bits[12] ),
    .B(_189_),
    .Y(_190_));
 sky130_fd_sc_hd__xnor2_1 _513_ (.A(_176_),
    .B(\cam_memory[12][7] ),
    .Y(_191_));
 sky130_fd_sc_hd__xnor2_1 _514_ (.A(_181_),
    .B(\cam_memory[12][2] ),
    .Y(_192_));
 sky130_fd_sc_hd__xnor2_1 _515_ (.A(_174_),
    .B(\cam_memory[12][6] ),
    .Y(_193_));
 sky130_fd_sc_hd__nand3_1 _516_ (.A(_191_),
    .B(_192_),
    .C(_193_),
    .Y(_194_));
 sky130_fd_sc_hd__xnor2_1 _517_ (.A(_172_),
    .B(\cam_memory[12][5] ),
    .Y(_195_));
 sky130_fd_sc_hd__xnor2_1 _518_ (.A(_185_),
    .B(\cam_memory[12][3] ),
    .Y(_196_));
 sky130_fd_sc_hd__xnor2_1 _519_ (.A(_169_),
    .B(\cam_memory[12][0] ),
    .Y(_197_));
 sky130_fd_sc_hd__xnor2_1 _520_ (.A(_179_),
    .B(\cam_memory[12][4] ),
    .Y(_198_));
 sky130_fd_sc_hd__nand4_1 _521_ (.A(_195_),
    .B(_196_),
    .C(_197_),
    .D(_198_),
    .Y(_199_));
 sky130_fd_sc_hd__nor3_2 _522_ (.A(_190_),
    .B(_194_),
    .C(_199_),
    .Y(_200_));
 sky130_fd_sc_hd__xnor2_1 _523_ (.A(_183_),
    .B(\cam_memory[13][1] ),
    .Y(_201_));
 sky130_fd_sc_hd__xor2_1 _524_ (.A(_152_),
    .B(\cam_memory[13][6] ),
    .X(_202_));
 sky130_fd_sc_hd__xor2_1 _525_ (.A(_159_),
    .B(\cam_memory[13][4] ),
    .X(_203_));
 sky130_fd_sc_hd__xor2_1 _526_ (.A(_176_),
    .B(\cam_memory[13][7] ),
    .X(_204_));
 sky130_fd_sc_hd__nor3_1 _527_ (.A(_202_),
    .B(_203_),
    .C(_204_),
    .Y(_205_));
 sky130_fd_sc_hd__xor2_1 _528_ (.A(_163_),
    .B(\cam_memory[13][3] ),
    .X(_206_));
 sky130_fd_sc_hd__xor2_1 _529_ (.A(_154_),
    .B(\cam_memory[13][5] ),
    .X(_207_));
 sky130_fd_sc_hd__xor2_1 _530_ (.A(_161_),
    .B(\cam_memory[13][2] ),
    .X(_208_));
 sky130_fd_sc_hd__xor2_1 _531_ (.A(_165_),
    .B(\cam_memory[13][0] ),
    .X(_209_));
 sky130_fd_sc_hd__nor4_1 _532_ (.A(_206_),
    .B(_207_),
    .C(_208_),
    .D(_209_),
    .Y(_210_));
 sky130_fd_sc_hd__nand4_1 _533_ (.A(\valid_bits[13] ),
    .B(_201_),
    .C(_205_),
    .D(_210_),
    .Y(_211_));
 sky130_fd_sc_hd__nor4b_2 _534_ (.A(_168_),
    .B(_188_),
    .C(_200_),
    .D_N(_211_),
    .Y(_212_));
 sky130_fd_sc_hd__xnor2_1 _535_ (.A(_165_),
    .B(\cam_memory[9][0] ),
    .Y(_213_));
 sky130_fd_sc_hd__nand2_1 _536_ (.A(\valid_bits[9] ),
    .B(_213_),
    .Y(_214_));
 sky130_fd_sc_hd__xnor2_1 _537_ (.A(_152_),
    .B(\cam_memory[9][6] ),
    .Y(_215_));
 sky130_fd_sc_hd__xnor2_1 _538_ (.A(_154_),
    .B(\cam_memory[9][5] ),
    .Y(_216_));
 sky130_fd_sc_hd__xnor2_1 _539_ (.A(_156_),
    .B(\cam_memory[9][7] ),
    .Y(_217_));
 sky130_fd_sc_hd__nand3_1 _540_ (.A(_215_),
    .B(_216_),
    .C(_217_),
    .Y(_218_));
 sky130_fd_sc_hd__xnor2_1 _541_ (.A(_163_),
    .B(\cam_memory[9][3] ),
    .Y(_219_));
 sky130_fd_sc_hd__xnor2_1 _542_ (.A(_161_),
    .B(\cam_memory[9][2] ),
    .Y(_220_));
 sky130_fd_sc_hd__xnor2_1 _543_ (.A(_149_),
    .B(\cam_memory[9][1] ),
    .Y(_221_));
 sky130_fd_sc_hd__xnor2_1 _544_ (.A(_159_),
    .B(\cam_memory[9][4] ),
    .Y(_222_));
 sky130_fd_sc_hd__nand4_2 _545_ (.A(_219_),
    .B(_220_),
    .C(_221_),
    .D(_222_),
    .Y(_223_));
 sky130_fd_sc_hd__nor3_4 _546_ (.A(_214_),
    .B(_218_),
    .C(_223_),
    .Y(_224_));
 sky130_fd_sc_hd__xnor2_1 _547_ (.A(_183_),
    .B(\cam_memory[11][1] ),
    .Y(_225_));
 sky130_fd_sc_hd__nand2_1 _548_ (.A(\valid_bits[11] ),
    .B(_225_),
    .Y(_226_));
 sky130_fd_sc_hd__xnor2_1 _549_ (.A(_174_),
    .B(\cam_memory[11][6] ),
    .Y(_227_));
 sky130_fd_sc_hd__xnor2_1 _550_ (.A(_172_),
    .B(\cam_memory[11][5] ),
    .Y(_228_));
 sky130_fd_sc_hd__xnor2_1 _551_ (.A(_176_),
    .B(\cam_memory[11][7] ),
    .Y(_229_));
 sky130_fd_sc_hd__nand3_1 _552_ (.A(_227_),
    .B(_228_),
    .C(_229_),
    .Y(_230_));
 sky130_fd_sc_hd__xnor2_1 _553_ (.A(_185_),
    .B(\cam_memory[11][3] ),
    .Y(_231_));
 sky130_fd_sc_hd__xnor2_1 _554_ (.A(_179_),
    .B(\cam_memory[11][4] ),
    .Y(_232_));
 sky130_fd_sc_hd__xnor2_1 _555_ (.A(_181_),
    .B(\cam_memory[11][2] ),
    .Y(_233_));
 sky130_fd_sc_hd__xnor2_1 _556_ (.A(_169_),
    .B(\cam_memory[11][0] ),
    .Y(_234_));
 sky130_fd_sc_hd__nand4_1 _557_ (.A(_231_),
    .B(_232_),
    .C(_233_),
    .D(_234_),
    .Y(_235_));
 sky130_fd_sc_hd__nor3_1 _558_ (.A(_226_),
    .B(_230_),
    .C(_235_),
    .Y(_236_));
 sky130_fd_sc_hd__xnor2_1 _559_ (.A(_149_),
    .B(\cam_memory[8][1] ),
    .Y(_237_));
 sky130_fd_sc_hd__nand2_1 _560_ (.A(\valid_bits[8] ),
    .B(_237_),
    .Y(_238_));
 sky130_fd_sc_hd__xnor2_1 _561_ (.A(_174_),
    .B(\cam_memory[8][6] ),
    .Y(_239_));
 sky130_fd_sc_hd__xnor2_1 _562_ (.A(_156_),
    .B(\cam_memory[8][7] ),
    .Y(_240_));
 sky130_fd_sc_hd__xnor2_1 _563_ (.A(_161_),
    .B(\cam_memory[8][2] ),
    .Y(_241_));
 sky130_fd_sc_hd__nand3_1 _564_ (.A(_239_),
    .B(_240_),
    .C(_241_),
    .Y(_242_));
 sky130_fd_sc_hd__xnor2_1 _565_ (.A(_172_),
    .B(\cam_memory[8][5] ),
    .Y(_243_));
 sky130_fd_sc_hd__xnor2_1 _566_ (.A(_163_),
    .B(\cam_memory[8][3] ),
    .Y(_244_));
 sky130_fd_sc_hd__xnor2_1 _567_ (.A(_179_),
    .B(\cam_memory[8][4] ),
    .Y(_245_));
 sky130_fd_sc_hd__xnor2_1 _568_ (.A(_165_),
    .B(\cam_memory[8][0] ),
    .Y(_246_));
 sky130_fd_sc_hd__nand4_2 _569_ (.A(_243_),
    .B(_244_),
    .C(_245_),
    .D(_246_),
    .Y(_247_));
 sky130_fd_sc_hd__nor3_4 _570_ (.A(_238_),
    .B(_242_),
    .C(_247_),
    .Y(_248_));
 sky130_fd_sc_hd__xnor2_1 _571_ (.A(_165_),
    .B(\cam_memory[10][0] ),
    .Y(_249_));
 sky130_fd_sc_hd__nand2_1 _572_ (.A(\valid_bits[10] ),
    .B(_249_),
    .Y(_250_));
 sky130_fd_sc_hd__xnor2_1 _573_ (.A(_152_),
    .B(\cam_memory[10][6] ),
    .Y(_251_));
 sky130_fd_sc_hd__xnor2_1 _574_ (.A(_154_),
    .B(\cam_memory[10][5] ),
    .Y(_252_));
 sky130_fd_sc_hd__xnor2_1 _575_ (.A(_156_),
    .B(\cam_memory[10][7] ),
    .Y(_253_));
 sky130_fd_sc_hd__nand3_1 _576_ (.A(_251_),
    .B(_252_),
    .C(_253_),
    .Y(_254_));
 sky130_fd_sc_hd__xnor2_1 _577_ (.A(_163_),
    .B(\cam_memory[10][3] ),
    .Y(_255_));
 sky130_fd_sc_hd__xnor2_1 _578_ (.A(_149_),
    .B(\cam_memory[10][1] ),
    .Y(_256_));
 sky130_fd_sc_hd__xnor2_1 _579_ (.A(_161_),
    .B(\cam_memory[10][2] ),
    .Y(_257_));
 sky130_fd_sc_hd__xnor2_1 _580_ (.A(_159_),
    .B(\cam_memory[10][4] ),
    .Y(_258_));
 sky130_fd_sc_hd__nand4_1 _581_ (.A(_255_),
    .B(_256_),
    .C(_257_),
    .D(_258_),
    .Y(_259_));
 sky130_fd_sc_hd__nor3_1 _582_ (.A(_250_),
    .B(_254_),
    .C(_259_),
    .Y(_260_));
 sky130_fd_sc_hd__nor4_2 _583_ (.A(_224_),
    .B(_236_),
    .C(_248_),
    .D(_260_),
    .Y(_261_));
 sky130_fd_sc_hd__xnor2_1 _584_ (.A(_149_),
    .B(\cam_memory[7][1] ),
    .Y(_262_));
 sky130_fd_sc_hd__nand2_1 _585_ (.A(\valid_bits[7] ),
    .B(_262_),
    .Y(_263_));
 sky130_fd_sc_hd__xnor2_1 _586_ (.A(_152_),
    .B(\cam_memory[7][6] ),
    .Y(_264_));
 sky130_fd_sc_hd__xnor2_1 _587_ (.A(_154_),
    .B(\cam_memory[7][5] ),
    .Y(_265_));
 sky130_fd_sc_hd__xnor2_1 _588_ (.A(_156_),
    .B(\cam_memory[7][7] ),
    .Y(_266_));
 sky130_fd_sc_hd__nand3_1 _589_ (.A(_264_),
    .B(_265_),
    .C(_266_),
    .Y(_267_));
 sky130_fd_sc_hd__xnor2_1 _590_ (.A(_185_),
    .B(\cam_memory[7][3] ),
    .Y(_268_));
 sky130_fd_sc_hd__xnor2_1 _591_ (.A(_169_),
    .B(\cam_memory[7][0] ),
    .Y(_269_));
 sky130_fd_sc_hd__xnor2_1 _592_ (.A(_181_),
    .B(\cam_memory[7][2] ),
    .Y(_270_));
 sky130_fd_sc_hd__xnor2_1 _593_ (.A(_159_),
    .B(\cam_memory[7][4] ),
    .Y(_271_));
 sky130_fd_sc_hd__nand4_1 _594_ (.A(_268_),
    .B(_269_),
    .C(_270_),
    .D(_271_),
    .Y(_272_));
 sky130_fd_sc_hd__nor3_2 _595_ (.A(_263_),
    .B(_267_),
    .C(_272_),
    .Y(_273_));
 sky130_fd_sc_hd__xnor2_1 _596_ (.A(_169_),
    .B(\cam_memory[5][0] ),
    .Y(_274_));
 sky130_fd_sc_hd__nand2_1 _597_ (.A(\valid_bits[5] ),
    .B(_274_),
    .Y(_275_));
 sky130_fd_sc_hd__xnor2_1 _598_ (.A(_176_),
    .B(\cam_memory[5][7] ),
    .Y(_276_));
 sky130_fd_sc_hd__xnor2_1 _599_ (.A(_181_),
    .B(\cam_memory[5][2] ),
    .Y(_277_));
 sky130_fd_sc_hd__xnor2_1 _600_ (.A(_174_),
    .B(\cam_memory[5][6] ),
    .Y(_278_));
 sky130_fd_sc_hd__nand3_1 _601_ (.A(_276_),
    .B(_277_),
    .C(_278_),
    .Y(_279_));
 sky130_fd_sc_hd__xnor2_1 _602_ (.A(_179_),
    .B(\cam_memory[5][4] ),
    .Y(_280_));
 sky130_fd_sc_hd__xnor2_1 _603_ (.A(_183_),
    .B(\cam_memory[5][1] ),
    .Y(_281_));
 sky130_fd_sc_hd__xnor2_1 _604_ (.A(_185_),
    .B(\cam_memory[5][3] ),
    .Y(_282_));
 sky130_fd_sc_hd__xnor2_1 _605_ (.A(_172_),
    .B(\cam_memory[5][5] ),
    .Y(_283_));
 sky130_fd_sc_hd__nand4_1 _606_ (.A(_280_),
    .B(_281_),
    .C(_282_),
    .D(_283_),
    .Y(_284_));
 sky130_fd_sc_hd__nor3_1 _607_ (.A(_275_),
    .B(_279_),
    .C(_284_),
    .Y(_285_));
 sky130_fd_sc_hd__xnor2_1 _608_ (.A(_169_),
    .B(\cam_memory[6][0] ),
    .Y(_286_));
 sky130_fd_sc_hd__nand2_1 _609_ (.A(\valid_bits[6] ),
    .B(_286_),
    .Y(_287_));
 sky130_fd_sc_hd__xnor2_1 _610_ (.A(_174_),
    .B(\cam_memory[6][6] ),
    .Y(_288_));
 sky130_fd_sc_hd__xnor2_1 _611_ (.A(_172_),
    .B(\cam_memory[6][5] ),
    .Y(_289_));
 sky130_fd_sc_hd__xnor2_1 _612_ (.A(_176_),
    .B(\cam_memory[6][7] ),
    .Y(_290_));
 sky130_fd_sc_hd__nand3_1 _613_ (.A(_288_),
    .B(_289_),
    .C(_290_),
    .Y(_291_));
 sky130_fd_sc_hd__xnor2_1 _614_ (.A(_181_),
    .B(\cam_memory[6][2] ),
    .Y(_292_));
 sky130_fd_sc_hd__xnor2_1 _615_ (.A(_183_),
    .B(\cam_memory[6][1] ),
    .Y(_293_));
 sky130_fd_sc_hd__xnor2_1 _616_ (.A(_185_),
    .B(\cam_memory[6][3] ),
    .Y(_294_));
 sky130_fd_sc_hd__xnor2_1 _617_ (.A(_179_),
    .B(\cam_memory[6][4] ),
    .Y(_295_));
 sky130_fd_sc_hd__nand4_1 _618_ (.A(_292_),
    .B(_293_),
    .C(_294_),
    .D(_295_),
    .Y(_296_));
 sky130_fd_sc_hd__nor3_2 _619_ (.A(_287_),
    .B(_291_),
    .C(_296_),
    .Y(_297_));
 sky130_fd_sc_hd__xnor2_1 _620_ (.A(_165_),
    .B(\cam_memory[4][0] ),
    .Y(_298_));
 sky130_fd_sc_hd__nand2_1 _621_ (.A(\valid_bits[4] ),
    .B(_298_),
    .Y(_299_));
 sky130_fd_sc_hd__xnor2_1 _622_ (.A(_154_),
    .B(\cam_memory[4][5] ),
    .Y(_300_));
 sky130_fd_sc_hd__xnor2_1 _623_ (.A(_159_),
    .B(\cam_memory[4][4] ),
    .Y(_301_));
 sky130_fd_sc_hd__xnor2_1 _624_ (.A(_156_),
    .B(\cam_memory[4][7] ),
    .Y(_302_));
 sky130_fd_sc_hd__nand3_1 _625_ (.A(_300_),
    .B(_301_),
    .C(_302_),
    .Y(_303_));
 sky130_fd_sc_hd__xnor2_1 _626_ (.A(_163_),
    .B(\cam_memory[4][3] ),
    .Y(_304_));
 sky130_fd_sc_hd__xnor2_1 _627_ (.A(_149_),
    .B(\cam_memory[4][1] ),
    .Y(_305_));
 sky130_fd_sc_hd__xnor2_1 _628_ (.A(_161_),
    .B(\cam_memory[4][2] ),
    .Y(_306_));
 sky130_fd_sc_hd__xnor2_1 _629_ (.A(_152_),
    .B(\cam_memory[4][6] ),
    .Y(_307_));
 sky130_fd_sc_hd__nand4_1 _630_ (.A(_304_),
    .B(_305_),
    .C(_306_),
    .D(_307_),
    .Y(_308_));
 sky130_fd_sc_hd__or3_2 _631_ (.A(_299_),
    .B(_303_),
    .C(_308_),
    .X(_309_));
 sky130_fd_sc_hd__nor4b_1 _632_ (.A(_273_),
    .B(_285_),
    .C(_297_),
    .D_N(_309_),
    .Y(_310_));
 sky130_fd_sc_hd__xnor2_1 _633_ (.A(_183_),
    .B(\cam_memory[3][1] ),
    .Y(_311_));
 sky130_fd_sc_hd__nand2_1 _634_ (.A(\valid_bits[3] ),
    .B(_311_),
    .Y(_312_));
 sky130_fd_sc_hd__xnor2_1 _635_ (.A(_174_),
    .B(\cam_memory[3][6] ),
    .Y(_313_));
 sky130_fd_sc_hd__xnor2_1 _636_ (.A(_179_),
    .B(\cam_memory[3][4] ),
    .Y(_314_));
 sky130_fd_sc_hd__xnor2_1 _637_ (.A(_176_),
    .B(\cam_memory[3][7] ),
    .Y(_315_));
 sky130_fd_sc_hd__nand3_1 _638_ (.A(_313_),
    .B(_314_),
    .C(_315_),
    .Y(_316_));
 sky130_fd_sc_hd__xnor2_1 _639_ (.A(_181_),
    .B(\cam_memory[3][2] ),
    .Y(_317_));
 sky130_fd_sc_hd__xnor2_1 _640_ (.A(_169_),
    .B(\cam_memory[3][0] ),
    .Y(_318_));
 sky130_fd_sc_hd__xnor2_1 _641_ (.A(_185_),
    .B(\cam_memory[3][3] ),
    .Y(_319_));
 sky130_fd_sc_hd__xnor2_1 _642_ (.A(_172_),
    .B(\cam_memory[3][5] ),
    .Y(_320_));
 sky130_fd_sc_hd__nand4_1 _643_ (.A(_317_),
    .B(_318_),
    .C(_319_),
    .D(_320_),
    .Y(_321_));
 sky130_fd_sc_hd__nor3_1 _644_ (.A(_312_),
    .B(_316_),
    .C(_321_),
    .Y(_322_));
 sky130_fd_sc_hd__xnor2_1 _645_ (.A(_169_),
    .B(\cam_memory[2][0] ),
    .Y(_323_));
 sky130_fd_sc_hd__nand2_1 _646_ (.A(\valid_bits[2] ),
    .B(_323_),
    .Y(_324_));
 sky130_fd_sc_hd__xnor2_1 _647_ (.A(_174_),
    .B(\cam_memory[2][6] ),
    .Y(_325_));
 sky130_fd_sc_hd__xnor2_1 _648_ (.A(_172_),
    .B(\cam_memory[2][5] ),
    .Y(_326_));
 sky130_fd_sc_hd__xnor2_1 _649_ (.A(_176_),
    .B(\cam_memory[2][7] ),
    .Y(_327_));
 sky130_fd_sc_hd__nand3_1 _650_ (.A(_325_),
    .B(_326_),
    .C(_327_),
    .Y(_328_));
 sky130_fd_sc_hd__xnor2_1 _651_ (.A(_185_),
    .B(\cam_memory[2][3] ),
    .Y(_329_));
 sky130_fd_sc_hd__xnor2_1 _652_ (.A(_183_),
    .B(\cam_memory[2][1] ),
    .Y(_330_));
 sky130_fd_sc_hd__xnor2_1 _653_ (.A(_181_),
    .B(\cam_memory[2][2] ),
    .Y(_331_));
 sky130_fd_sc_hd__xnor2_1 _654_ (.A(_179_),
    .B(\cam_memory[2][4] ),
    .Y(_332_));
 sky130_fd_sc_hd__nand4_1 _655_ (.A(_329_),
    .B(_330_),
    .C(_331_),
    .D(_332_),
    .Y(_333_));
 sky130_fd_sc_hd__nor3_2 _656_ (.A(_324_),
    .B(_328_),
    .C(_333_),
    .Y(_334_));
 sky130_fd_sc_hd__xnor2_1 _657_ (.A(_183_),
    .B(\cam_memory[0][1] ),
    .Y(_335_));
 sky130_fd_sc_hd__nand2_1 _658_ (.A(\valid_bits[0] ),
    .B(_335_),
    .Y(_336_));
 sky130_fd_sc_hd__xnor2_1 _659_ (.A(_174_),
    .B(\cam_memory[0][6] ),
    .Y(_337_));
 sky130_fd_sc_hd__xnor2_1 _660_ (.A(_179_),
    .B(\cam_memory[0][4] ),
    .Y(_338_));
 sky130_fd_sc_hd__xnor2_1 _661_ (.A(_176_),
    .B(\cam_memory[0][7] ),
    .Y(_339_));
 sky130_fd_sc_hd__nand3_1 _662_ (.A(_337_),
    .B(_338_),
    .C(_339_),
    .Y(_340_));
 sky130_fd_sc_hd__xnor2_1 _663_ (.A(_185_),
    .B(\cam_memory[0][3] ),
    .Y(_341_));
 sky130_fd_sc_hd__xnor2_1 _664_ (.A(_172_),
    .B(\cam_memory[0][5] ),
    .Y(_342_));
 sky130_fd_sc_hd__xnor2_1 _665_ (.A(_169_),
    .B(\cam_memory[0][0] ),
    .Y(_343_));
 sky130_fd_sc_hd__xnor2_1 _666_ (.A(_181_),
    .B(\cam_memory[0][2] ),
    .Y(_344_));
 sky130_fd_sc_hd__nand4_1 _667_ (.A(_341_),
    .B(_342_),
    .C(_343_),
    .D(_344_),
    .Y(_345_));
 sky130_fd_sc_hd__nor3_1 _668_ (.A(_336_),
    .B(_340_),
    .C(_345_),
    .Y(_346_));
 sky130_fd_sc_hd__xnor2_1 _669_ (.A(_169_),
    .B(\cam_memory[1][0] ),
    .Y(_347_));
 sky130_fd_sc_hd__nand2_1 _670_ (.A(\valid_bits[1] ),
    .B(_347_),
    .Y(_348_));
 sky130_fd_sc_hd__xnor2_1 _671_ (.A(_174_),
    .B(\cam_memory[1][6] ),
    .Y(_349_));
 sky130_fd_sc_hd__xnor2_1 _672_ (.A(_172_),
    .B(\cam_memory[1][5] ),
    .Y(_350_));
 sky130_fd_sc_hd__xnor2_1 _673_ (.A(_176_),
    .B(\cam_memory[1][7] ),
    .Y(_351_));
 sky130_fd_sc_hd__nand3_1 _674_ (.A(_349_),
    .B(_350_),
    .C(_351_),
    .Y(_352_));
 sky130_fd_sc_hd__xnor2_1 _675_ (.A(_179_),
    .B(\cam_memory[1][4] ),
    .Y(_353_));
 sky130_fd_sc_hd__xnor2_1 _676_ (.A(_185_),
    .B(\cam_memory[1][3] ),
    .Y(_354_));
 sky130_fd_sc_hd__xnor2_1 _677_ (.A(_183_),
    .B(\cam_memory[1][1] ),
    .Y(_355_));
 sky130_fd_sc_hd__xnor2_1 _678_ (.A(_181_),
    .B(\cam_memory[1][2] ),
    .Y(_356_));
 sky130_fd_sc_hd__nand4_1 _679_ (.A(_353_),
    .B(_354_),
    .C(_355_),
    .D(_356_),
    .Y(_357_));
 sky130_fd_sc_hd__nor3_1 _680_ (.A(_348_),
    .B(_352_),
    .C(_357_),
    .Y(_358_));
 sky130_fd_sc_hd__nor4_1 _681_ (.A(_322_),
    .B(_334_),
    .C(_346_),
    .D(_358_),
    .Y(_359_));
 sky130_fd_sc_hd__inv_1 _682_ (.A(net2),
    .Y(_360_));
 sky130_fd_sc_hd__a41oi_2 _683_ (.A1(_212_),
    .A2(_261_),
    .A3(_310_),
    .A4(_359_),
    .B1(_360_),
    .Y(_000_));
 sky130_fd_sc_hd__inv_1 _684_ (.A(net3),
    .Y(_461_));
 sky130_fd_sc_hd__inv_1 _685_ (.A(net4),
    .Y(_462_));
 sky130_fd_sc_hd__buf_4 _686_ (.A(net13),
    .X(_361_));
 sky130_fd_sc_hd__clkbuf_4 _687_ (.A(_463_),
    .X(_362_));
 sky130_fd_sc_hd__buf_4 _688_ (.A(write_addr[3]),
    .X(_363_));
 sky130_fd_sc_hd__buf_4 _689_ (.A(write_addr[2]),
    .X(_364_));
 sky130_fd_sc_hd__nor2_1 _690_ (.A(_363_),
    .B(_364_),
    .Y(_365_));
 sky130_fd_sc_hd__and3_1 _691_ (.A(_361_),
    .B(_362_),
    .C(_365_),
    .X(_366_));
 sky130_fd_sc_hd__clkbuf_4 _692_ (.A(_366_),
    .X(_367_));
 sky130_fd_sc_hd__mux2_1 _693_ (.A0(\cam_memory[0][0] ),
    .A1(net5),
    .S(_367_),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _694_ (.A0(\cam_memory[0][1] ),
    .A1(net6),
    .S(_367_),
    .X(_002_));
 sky130_fd_sc_hd__mux2_1 _695_ (.A0(\cam_memory[0][2] ),
    .A1(net7),
    .S(_367_),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _696_ (.A0(\cam_memory[0][3] ),
    .A1(net8),
    .S(_367_),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _697_ (.A0(\cam_memory[0][4] ),
    .A1(net9),
    .S(_367_),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _698_ (.A0(\cam_memory[0][5] ),
    .A1(net10),
    .S(_367_),
    .X(_006_));
 sky130_fd_sc_hd__mux2_1 _699_ (.A0(\cam_memory[0][6] ),
    .A1(net11),
    .S(_367_),
    .X(_007_));
 sky130_fd_sc_hd__mux2_1 _700_ (.A0(\cam_memory[0][7] ),
    .A1(net12),
    .S(_367_),
    .X(_008_));
 sky130_fd_sc_hd__buf_4 _701_ (.A(net5),
    .X(_368_));
 sky130_fd_sc_hd__buf_6 _702_ (.A(_361_),
    .X(_369_));
 sky130_fd_sc_hd__clkbuf_4 _703_ (.A(_465_),
    .X(_370_));
 sky130_fd_sc_hd__nor2b_1 _704_ (.A(_364_),
    .B_N(_363_),
    .Y(_371_));
 sky130_fd_sc_hd__clkbuf_4 _705_ (.A(_371_),
    .X(_372_));
 sky130_fd_sc_hd__nand3_4 _706_ (.A(_369_),
    .B(_370_),
    .C(_372_),
    .Y(_373_));
 sky130_fd_sc_hd__mux2_1 _707_ (.A0(_368_),
    .A1(\cam_memory[10][0] ),
    .S(_373_),
    .X(_009_));
 sky130_fd_sc_hd__clkbuf_4 _708_ (.A(net6),
    .X(_374_));
 sky130_fd_sc_hd__mux2_1 _709_ (.A0(_374_),
    .A1(\cam_memory[10][1] ),
    .S(_373_),
    .X(_010_));
 sky130_fd_sc_hd__buf_4 _710_ (.A(net7),
    .X(_375_));
 sky130_fd_sc_hd__mux2_1 _711_ (.A0(_375_),
    .A1(\cam_memory[10][2] ),
    .S(_373_),
    .X(_011_));
 sky130_fd_sc_hd__buf_4 _712_ (.A(net8),
    .X(_376_));
 sky130_fd_sc_hd__mux2_1 _713_ (.A0(_376_),
    .A1(\cam_memory[10][3] ),
    .S(_373_),
    .X(_012_));
 sky130_fd_sc_hd__buf_4 _714_ (.A(net9),
    .X(_377_));
 sky130_fd_sc_hd__mux2_1 _715_ (.A0(_377_),
    .A1(\cam_memory[10][4] ),
    .S(_373_),
    .X(_013_));
 sky130_fd_sc_hd__buf_4 _716_ (.A(net10),
    .X(_378_));
 sky130_fd_sc_hd__mux2_1 _717_ (.A0(_378_),
    .A1(\cam_memory[10][5] ),
    .S(_373_),
    .X(_014_));
 sky130_fd_sc_hd__buf_4 _718_ (.A(net11),
    .X(_379_));
 sky130_fd_sc_hd__mux2_1 _719_ (.A0(_379_),
    .A1(\cam_memory[10][6] ),
    .S(_373_),
    .X(_015_));
 sky130_fd_sc_hd__buf_4 _720_ (.A(net12),
    .X(_380_));
 sky130_fd_sc_hd__mux2_1 _721_ (.A0(_380_),
    .A1(\cam_memory[10][7] ),
    .S(_373_),
    .X(_016_));
 sky130_fd_sc_hd__buf_4 _722_ (.A(_469_),
    .X(_381_));
 sky130_fd_sc_hd__nand3_4 _723_ (.A(_369_),
    .B(_381_),
    .C(_372_),
    .Y(_382_));
 sky130_fd_sc_hd__mux2_1 _724_ (.A0(_368_),
    .A1(\cam_memory[11][0] ),
    .S(_382_),
    .X(_017_));
 sky130_fd_sc_hd__mux2_1 _725_ (.A0(_374_),
    .A1(\cam_memory[11][1] ),
    .S(_382_),
    .X(_018_));
 sky130_fd_sc_hd__mux2_1 _726_ (.A0(_375_),
    .A1(\cam_memory[11][2] ),
    .S(_382_),
    .X(_019_));
 sky130_fd_sc_hd__mux2_1 _727_ (.A0(_376_),
    .A1(\cam_memory[11][3] ),
    .S(_382_),
    .X(_020_));
 sky130_fd_sc_hd__mux2_1 _728_ (.A0(_377_),
    .A1(\cam_memory[11][4] ),
    .S(_382_),
    .X(_021_));
 sky130_fd_sc_hd__mux2_1 _729_ (.A0(_378_),
    .A1(\cam_memory[11][5] ),
    .S(_382_),
    .X(_022_));
 sky130_fd_sc_hd__mux2_1 _730_ (.A0(_379_),
    .A1(\cam_memory[11][6] ),
    .S(_382_),
    .X(_023_));
 sky130_fd_sc_hd__mux2_1 _731_ (.A0(_380_),
    .A1(\cam_memory[11][7] ),
    .S(_382_),
    .X(_024_));
 sky130_fd_sc_hd__nand4_4 _732_ (.A(_363_),
    .B(_364_),
    .C(_361_),
    .D(_362_),
    .Y(_383_));
 sky130_fd_sc_hd__mux2_1 _733_ (.A0(_368_),
    .A1(\cam_memory[12][0] ),
    .S(_383_),
    .X(_025_));
 sky130_fd_sc_hd__mux2_1 _734_ (.A0(_374_),
    .A1(\cam_memory[12][1] ),
    .S(_383_),
    .X(_026_));
 sky130_fd_sc_hd__mux2_1 _735_ (.A0(_375_),
    .A1(\cam_memory[12][2] ),
    .S(_383_),
    .X(_027_));
 sky130_fd_sc_hd__mux2_1 _736_ (.A0(_376_),
    .A1(\cam_memory[12][3] ),
    .S(_383_),
    .X(_028_));
 sky130_fd_sc_hd__mux2_1 _737_ (.A0(_377_),
    .A1(\cam_memory[12][4] ),
    .S(_383_),
    .X(_029_));
 sky130_fd_sc_hd__mux2_1 _738_ (.A0(_378_),
    .A1(\cam_memory[12][5] ),
    .S(_383_),
    .X(_030_));
 sky130_fd_sc_hd__mux2_1 _739_ (.A0(_379_),
    .A1(\cam_memory[12][6] ),
    .S(_383_),
    .X(_031_));
 sky130_fd_sc_hd__mux2_1 _740_ (.A0(_380_),
    .A1(\cam_memory[12][7] ),
    .S(_383_),
    .X(_032_));
 sky130_fd_sc_hd__clkbuf_4 _741_ (.A(_467_),
    .X(_384_));
 sky130_fd_sc_hd__nand4_4 _742_ (.A(_363_),
    .B(_364_),
    .C(_361_),
    .D(_384_),
    .Y(_385_));
 sky130_fd_sc_hd__mux2_1 _743_ (.A0(_368_),
    .A1(\cam_memory[13][0] ),
    .S(_385_),
    .X(_033_));
 sky130_fd_sc_hd__mux2_1 _744_ (.A0(_374_),
    .A1(\cam_memory[13][1] ),
    .S(_385_),
    .X(_034_));
 sky130_fd_sc_hd__mux2_1 _745_ (.A0(_375_),
    .A1(\cam_memory[13][2] ),
    .S(_385_),
    .X(_035_));
 sky130_fd_sc_hd__mux2_1 _746_ (.A0(_376_),
    .A1(\cam_memory[13][3] ),
    .S(_385_),
    .X(_036_));
 sky130_fd_sc_hd__mux2_1 _747_ (.A0(_377_),
    .A1(\cam_memory[13][4] ),
    .S(_385_),
    .X(_037_));
 sky130_fd_sc_hd__mux2_1 _748_ (.A0(_378_),
    .A1(\cam_memory[13][5] ),
    .S(_385_),
    .X(_038_));
 sky130_fd_sc_hd__mux2_1 _749_ (.A0(_379_),
    .A1(\cam_memory[13][6] ),
    .S(_385_),
    .X(_039_));
 sky130_fd_sc_hd__mux2_1 _750_ (.A0(_380_),
    .A1(\cam_memory[13][7] ),
    .S(_385_),
    .X(_040_));
 sky130_fd_sc_hd__nand4_4 _751_ (.A(_363_),
    .B(_364_),
    .C(_361_),
    .D(_370_),
    .Y(_386_));
 sky130_fd_sc_hd__mux2_1 _752_ (.A0(_368_),
    .A1(\cam_memory[14][0] ),
    .S(_386_),
    .X(_041_));
 sky130_fd_sc_hd__mux2_1 _753_ (.A0(_374_),
    .A1(\cam_memory[14][1] ),
    .S(_386_),
    .X(_042_));
 sky130_fd_sc_hd__mux2_1 _754_ (.A0(_375_),
    .A1(\cam_memory[14][2] ),
    .S(_386_),
    .X(_043_));
 sky130_fd_sc_hd__mux2_1 _755_ (.A0(_376_),
    .A1(\cam_memory[14][3] ),
    .S(_386_),
    .X(_044_));
 sky130_fd_sc_hd__mux2_1 _756_ (.A0(_377_),
    .A1(\cam_memory[14][4] ),
    .S(_386_),
    .X(_045_));
 sky130_fd_sc_hd__mux2_1 _757_ (.A0(_378_),
    .A1(\cam_memory[14][5] ),
    .S(_386_),
    .X(_046_));
 sky130_fd_sc_hd__mux2_1 _758_ (.A0(_379_),
    .A1(\cam_memory[14][6] ),
    .S(_386_),
    .X(_047_));
 sky130_fd_sc_hd__mux2_1 _759_ (.A0(_380_),
    .A1(\cam_memory[14][7] ),
    .S(_386_),
    .X(_048_));
 sky130_fd_sc_hd__nand4_4 _760_ (.A(_363_),
    .B(_364_),
    .C(_361_),
    .D(_381_),
    .Y(_387_));
 sky130_fd_sc_hd__mux2_1 _761_ (.A0(_368_),
    .A1(\cam_memory[15][0] ),
    .S(_387_),
    .X(_049_));
 sky130_fd_sc_hd__mux2_1 _762_ (.A0(_374_),
    .A1(\cam_memory[15][1] ),
    .S(_387_),
    .X(_050_));
 sky130_fd_sc_hd__mux2_1 _763_ (.A0(_375_),
    .A1(\cam_memory[15][2] ),
    .S(_387_),
    .X(_051_));
 sky130_fd_sc_hd__mux2_1 _764_ (.A0(_376_),
    .A1(\cam_memory[15][3] ),
    .S(_387_),
    .X(_052_));
 sky130_fd_sc_hd__mux2_1 _765_ (.A0(_377_),
    .A1(\cam_memory[15][4] ),
    .S(_387_),
    .X(_053_));
 sky130_fd_sc_hd__mux2_1 _766_ (.A0(_378_),
    .A1(\cam_memory[15][5] ),
    .S(_387_),
    .X(_054_));
 sky130_fd_sc_hd__mux2_1 _767_ (.A0(_379_),
    .A1(\cam_memory[15][6] ),
    .S(_387_),
    .X(_055_));
 sky130_fd_sc_hd__mux2_1 _768_ (.A0(_380_),
    .A1(\cam_memory[15][7] ),
    .S(_387_),
    .X(_056_));
 sky130_fd_sc_hd__and3_1 _769_ (.A(_361_),
    .B(_384_),
    .C(_365_),
    .X(_388_));
 sky130_fd_sc_hd__clkbuf_4 _770_ (.A(_388_),
    .X(_389_));
 sky130_fd_sc_hd__mux2_1 _771_ (.A0(\cam_memory[1][0] ),
    .A1(net5),
    .S(_389_),
    .X(_057_));
 sky130_fd_sc_hd__mux2_1 _772_ (.A0(\cam_memory[1][1] ),
    .A1(net6),
    .S(_389_),
    .X(_058_));
 sky130_fd_sc_hd__mux2_1 _773_ (.A0(\cam_memory[1][2] ),
    .A1(net7),
    .S(_389_),
    .X(_059_));
 sky130_fd_sc_hd__mux2_1 _774_ (.A0(\cam_memory[1][3] ),
    .A1(net8),
    .S(_389_),
    .X(_060_));
 sky130_fd_sc_hd__mux2_1 _775_ (.A0(\cam_memory[1][4] ),
    .A1(net9),
    .S(_389_),
    .X(_061_));
 sky130_fd_sc_hd__mux2_1 _776_ (.A0(\cam_memory[1][5] ),
    .A1(net10),
    .S(_389_),
    .X(_062_));
 sky130_fd_sc_hd__mux2_1 _777_ (.A0(\cam_memory[1][6] ),
    .A1(net11),
    .S(_389_),
    .X(_063_));
 sky130_fd_sc_hd__mux2_1 _778_ (.A0(\cam_memory[1][7] ),
    .A1(net12),
    .S(_389_),
    .X(_064_));
 sky130_fd_sc_hd__and3_1 _779_ (.A(_361_),
    .B(_370_),
    .C(_365_),
    .X(_390_));
 sky130_fd_sc_hd__buf_2 _780_ (.A(_390_),
    .X(_391_));
 sky130_fd_sc_hd__mux2_1 _781_ (.A0(\cam_memory[2][0] ),
    .A1(net5),
    .S(_391_),
    .X(_065_));
 sky130_fd_sc_hd__mux2_1 _782_ (.A0(\cam_memory[2][1] ),
    .A1(net6),
    .S(_391_),
    .X(_066_));
 sky130_fd_sc_hd__mux2_1 _783_ (.A0(\cam_memory[2][2] ),
    .A1(net7),
    .S(_391_),
    .X(_067_));
 sky130_fd_sc_hd__mux2_1 _784_ (.A0(\cam_memory[2][3] ),
    .A1(net8),
    .S(_391_),
    .X(_068_));
 sky130_fd_sc_hd__mux2_1 _785_ (.A0(\cam_memory[2][4] ),
    .A1(net9),
    .S(_391_),
    .X(_069_));
 sky130_fd_sc_hd__mux2_1 _786_ (.A0(\cam_memory[2][5] ),
    .A1(net10),
    .S(_391_),
    .X(_070_));
 sky130_fd_sc_hd__mux2_1 _787_ (.A0(\cam_memory[2][6] ),
    .A1(net11),
    .S(_391_),
    .X(_071_));
 sky130_fd_sc_hd__mux2_1 _788_ (.A0(\cam_memory[2][7] ),
    .A1(net12),
    .S(_391_),
    .X(_072_));
 sky130_fd_sc_hd__and3_1 _789_ (.A(_361_),
    .B(_381_),
    .C(_365_),
    .X(_392_));
 sky130_fd_sc_hd__clkbuf_4 _790_ (.A(_392_),
    .X(_393_));
 sky130_fd_sc_hd__mux2_1 _791_ (.A0(\cam_memory[3][0] ),
    .A1(net5),
    .S(_393_),
    .X(_073_));
 sky130_fd_sc_hd__mux2_1 _792_ (.A0(\cam_memory[3][1] ),
    .A1(net6),
    .S(_393_),
    .X(_074_));
 sky130_fd_sc_hd__mux2_1 _793_ (.A0(\cam_memory[3][2] ),
    .A1(net7),
    .S(_393_),
    .X(_075_));
 sky130_fd_sc_hd__mux2_1 _794_ (.A0(\cam_memory[3][3] ),
    .A1(net8),
    .S(_393_),
    .X(_076_));
 sky130_fd_sc_hd__mux2_1 _795_ (.A0(\cam_memory[3][4] ),
    .A1(net9),
    .S(_393_),
    .X(_077_));
 sky130_fd_sc_hd__mux2_1 _796_ (.A0(\cam_memory[3][5] ),
    .A1(net10),
    .S(_393_),
    .X(_078_));
 sky130_fd_sc_hd__mux2_1 _797_ (.A0(\cam_memory[3][6] ),
    .A1(net11),
    .S(_393_),
    .X(_079_));
 sky130_fd_sc_hd__mux2_1 _798_ (.A0(\cam_memory[3][7] ),
    .A1(net12),
    .S(_393_),
    .X(_080_));
 sky130_fd_sc_hd__nor2b_1 _799_ (.A(_363_),
    .B_N(_364_),
    .Y(_394_));
 sky130_fd_sc_hd__clkbuf_4 _800_ (.A(_394_),
    .X(_395_));
 sky130_fd_sc_hd__nand3_4 _801_ (.A(_369_),
    .B(_362_),
    .C(_395_),
    .Y(_396_));
 sky130_fd_sc_hd__mux2_1 _802_ (.A0(_368_),
    .A1(\cam_memory[4][0] ),
    .S(_396_),
    .X(_081_));
 sky130_fd_sc_hd__mux2_1 _803_ (.A0(_374_),
    .A1(\cam_memory[4][1] ),
    .S(_396_),
    .X(_082_));
 sky130_fd_sc_hd__mux2_1 _804_ (.A0(_375_),
    .A1(\cam_memory[4][2] ),
    .S(_396_),
    .X(_083_));
 sky130_fd_sc_hd__mux2_1 _805_ (.A0(_376_),
    .A1(\cam_memory[4][3] ),
    .S(_396_),
    .X(_084_));
 sky130_fd_sc_hd__mux2_1 _806_ (.A0(_377_),
    .A1(\cam_memory[4][4] ),
    .S(_396_),
    .X(_085_));
 sky130_fd_sc_hd__mux2_1 _807_ (.A0(_378_),
    .A1(\cam_memory[4][5] ),
    .S(_396_),
    .X(_086_));
 sky130_fd_sc_hd__mux2_1 _808_ (.A0(_379_),
    .A1(\cam_memory[4][6] ),
    .S(_396_),
    .X(_087_));
 sky130_fd_sc_hd__mux2_1 _809_ (.A0(_380_),
    .A1(\cam_memory[4][7] ),
    .S(_396_),
    .X(_088_));
 sky130_fd_sc_hd__nand3_4 _810_ (.A(_369_),
    .B(_384_),
    .C(_395_),
    .Y(_397_));
 sky130_fd_sc_hd__mux2_1 _811_ (.A0(_368_),
    .A1(\cam_memory[5][0] ),
    .S(_397_),
    .X(_089_));
 sky130_fd_sc_hd__mux2_1 _812_ (.A0(_374_),
    .A1(\cam_memory[5][1] ),
    .S(_397_),
    .X(_090_));
 sky130_fd_sc_hd__mux2_1 _813_ (.A0(_375_),
    .A1(\cam_memory[5][2] ),
    .S(_397_),
    .X(_091_));
 sky130_fd_sc_hd__mux2_1 _814_ (.A0(_376_),
    .A1(\cam_memory[5][3] ),
    .S(_397_),
    .X(_092_));
 sky130_fd_sc_hd__mux2_1 _815_ (.A0(_377_),
    .A1(\cam_memory[5][4] ),
    .S(_397_),
    .X(_093_));
 sky130_fd_sc_hd__mux2_1 _816_ (.A0(_378_),
    .A1(\cam_memory[5][5] ),
    .S(_397_),
    .X(_094_));
 sky130_fd_sc_hd__mux2_1 _817_ (.A0(_379_),
    .A1(\cam_memory[5][6] ),
    .S(_397_),
    .X(_095_));
 sky130_fd_sc_hd__mux2_1 _818_ (.A0(_380_),
    .A1(\cam_memory[5][7] ),
    .S(_397_),
    .X(_096_));
 sky130_fd_sc_hd__nand3_4 _819_ (.A(_369_),
    .B(_370_),
    .C(_395_),
    .Y(_398_));
 sky130_fd_sc_hd__mux2_1 _820_ (.A0(_368_),
    .A1(\cam_memory[6][0] ),
    .S(_398_),
    .X(_097_));
 sky130_fd_sc_hd__mux2_1 _821_ (.A0(_374_),
    .A1(\cam_memory[6][1] ),
    .S(_398_),
    .X(_098_));
 sky130_fd_sc_hd__mux2_1 _822_ (.A0(_375_),
    .A1(\cam_memory[6][2] ),
    .S(_398_),
    .X(_099_));
 sky130_fd_sc_hd__mux2_1 _823_ (.A0(_376_),
    .A1(\cam_memory[6][3] ),
    .S(_398_),
    .X(_100_));
 sky130_fd_sc_hd__mux2_1 _824_ (.A0(_377_),
    .A1(\cam_memory[6][4] ),
    .S(_398_),
    .X(_101_));
 sky130_fd_sc_hd__mux2_1 _825_ (.A0(_378_),
    .A1(\cam_memory[6][5] ),
    .S(_398_),
    .X(_102_));
 sky130_fd_sc_hd__mux2_1 _826_ (.A0(_379_),
    .A1(\cam_memory[6][6] ),
    .S(_398_),
    .X(_103_));
 sky130_fd_sc_hd__mux2_1 _827_ (.A0(_380_),
    .A1(\cam_memory[6][7] ),
    .S(_398_),
    .X(_104_));
 sky130_fd_sc_hd__nand3_4 _828_ (.A(_369_),
    .B(_381_),
    .C(_395_),
    .Y(_399_));
 sky130_fd_sc_hd__mux2_1 _829_ (.A0(_368_),
    .A1(\cam_memory[7][0] ),
    .S(_399_),
    .X(_105_));
 sky130_fd_sc_hd__mux2_1 _830_ (.A0(_374_),
    .A1(\cam_memory[7][1] ),
    .S(_399_),
    .X(_106_));
 sky130_fd_sc_hd__mux2_1 _831_ (.A0(_375_),
    .A1(\cam_memory[7][2] ),
    .S(_399_),
    .X(_107_));
 sky130_fd_sc_hd__mux2_1 _832_ (.A0(_376_),
    .A1(\cam_memory[7][3] ),
    .S(_399_),
    .X(_108_));
 sky130_fd_sc_hd__mux2_1 _833_ (.A0(_377_),
    .A1(\cam_memory[7][4] ),
    .S(_399_),
    .X(_109_));
 sky130_fd_sc_hd__mux2_1 _834_ (.A0(_378_),
    .A1(\cam_memory[7][5] ),
    .S(_399_),
    .X(_110_));
 sky130_fd_sc_hd__mux2_1 _835_ (.A0(_379_),
    .A1(\cam_memory[7][6] ),
    .S(_399_),
    .X(_111_));
 sky130_fd_sc_hd__mux2_1 _836_ (.A0(_380_),
    .A1(\cam_memory[7][7] ),
    .S(_399_),
    .X(_112_));
 sky130_fd_sc_hd__nand3_4 _837_ (.A(_369_),
    .B(_362_),
    .C(_372_),
    .Y(_400_));
 sky130_fd_sc_hd__mux2_1 _838_ (.A0(net5),
    .A1(\cam_memory[8][0] ),
    .S(_400_),
    .X(_113_));
 sky130_fd_sc_hd__mux2_1 _839_ (.A0(net6),
    .A1(\cam_memory[8][1] ),
    .S(_400_),
    .X(_114_));
 sky130_fd_sc_hd__mux2_1 _840_ (.A0(net7),
    .A1(\cam_memory[8][2] ),
    .S(_400_),
    .X(_115_));
 sky130_fd_sc_hd__mux2_1 _841_ (.A0(net8),
    .A1(\cam_memory[8][3] ),
    .S(_400_),
    .X(_116_));
 sky130_fd_sc_hd__mux2_1 _842_ (.A0(net9),
    .A1(\cam_memory[8][4] ),
    .S(_400_),
    .X(_117_));
 sky130_fd_sc_hd__mux2_1 _843_ (.A0(net10),
    .A1(\cam_memory[8][5] ),
    .S(_400_),
    .X(_118_));
 sky130_fd_sc_hd__mux2_1 _844_ (.A0(net11),
    .A1(\cam_memory[8][6] ),
    .S(_400_),
    .X(_119_));
 sky130_fd_sc_hd__mux2_1 _845_ (.A0(net12),
    .A1(\cam_memory[8][7] ),
    .S(_400_),
    .X(_120_));
 sky130_fd_sc_hd__nand3_4 _846_ (.A(_369_),
    .B(_384_),
    .C(_372_),
    .Y(_401_));
 sky130_fd_sc_hd__mux2_1 _847_ (.A0(net5),
    .A1(\cam_memory[9][0] ),
    .S(_401_),
    .X(_121_));
 sky130_fd_sc_hd__mux2_1 _848_ (.A0(net6),
    .A1(\cam_memory[9][1] ),
    .S(_401_),
    .X(_122_));
 sky130_fd_sc_hd__mux2_1 _849_ (.A0(net7),
    .A1(\cam_memory[9][2] ),
    .S(_401_),
    .X(_123_));
 sky130_fd_sc_hd__mux2_1 _850_ (.A0(net8),
    .A1(\cam_memory[9][3] ),
    .S(_401_),
    .X(_124_));
 sky130_fd_sc_hd__mux2_1 _851_ (.A0(net9),
    .A1(\cam_memory[9][4] ),
    .S(_401_),
    .X(_125_));
 sky130_fd_sc_hd__mux2_1 _852_ (.A0(net10),
    .A1(\cam_memory[9][5] ),
    .S(_401_),
    .X(_126_));
 sky130_fd_sc_hd__mux2_1 _853_ (.A0(net11),
    .A1(\cam_memory[9][6] ),
    .S(_401_),
    .X(_127_));
 sky130_fd_sc_hd__mux2_1 _854_ (.A0(net12),
    .A1(\cam_memory[9][7] ),
    .S(_401_),
    .X(_128_));
 sky130_fd_sc_hd__nor2_1 _855_ (.A(_273_),
    .B(_285_),
    .Y(_402_));
 sky130_fd_sc_hd__or3_1 _856_ (.A(_348_),
    .B(_352_),
    .C(_357_),
    .X(_403_));
 sky130_fd_sc_hd__a21oi_1 _857_ (.A1(_346_),
    .A2(_403_),
    .B1(_334_),
    .Y(_404_));
 sky130_fd_sc_hd__o21ai_0 _858_ (.A1(_322_),
    .A2(_404_),
    .B1(_309_),
    .Y(_405_));
 sky130_fd_sc_hd__nand2b_1 _859_ (.A_N(_273_),
    .B(_297_),
    .Y(_406_));
 sky130_fd_sc_hd__nor4_1 _860_ (.A(_168_),
    .B(_200_),
    .C(_248_),
    .D(_260_),
    .Y(_407_));
 sky130_fd_sc_hd__nand2_1 _861_ (.A(_406_),
    .B(_407_),
    .Y(_408_));
 sky130_fd_sc_hd__a21o_1 _862_ (.A1(_402_),
    .A2(_405_),
    .B1(_408_),
    .X(_409_));
 sky130_fd_sc_hd__or3_1 _863_ (.A(_250_),
    .B(_254_),
    .C(_259_),
    .X(_410_));
 sky130_fd_sc_hd__a21oi_1 _864_ (.A1(_224_),
    .A2(_410_),
    .B1(_236_),
    .Y(_411_));
 sky130_fd_sc_hd__o21ai_0 _865_ (.A1(_200_),
    .A2(_411_),
    .B1(_211_),
    .Y(_412_));
 sky130_fd_sc_hd__nand2b_1 _866_ (.A_N(_168_),
    .B(_412_),
    .Y(_413_));
 sky130_fd_sc_hd__nand3_1 _867_ (.A(_170_),
    .B(_173_),
    .C(_175_),
    .Y(_414_));
 sky130_fd_sc_hd__nand4_1 _868_ (.A(_177_),
    .B(_180_),
    .C(_182_),
    .D(_184_),
    .Y(_415_));
 sky130_fd_sc_hd__nor2_1 _869_ (.A(_414_),
    .B(_415_),
    .Y(_416_));
 sky130_fd_sc_hd__nor2b_1 _870_ (.A(net2),
    .B_N(net15),
    .Y(_417_));
 sky130_fd_sc_hd__a31oi_1 _871_ (.A1(\valid_bits[15] ),
    .A2(_186_),
    .A3(_416_),
    .B1(_417_),
    .Y(_418_));
 sky130_fd_sc_hd__nor2_1 _872_ (.A(_000_),
    .B(_417_),
    .Y(_419_));
 sky130_fd_sc_hd__a31oi_1 _873_ (.A1(_409_),
    .A2(_413_),
    .A3(_418_),
    .B1(_419_),
    .Y(_129_));
 sky130_fd_sc_hd__nor2_1 _874_ (.A(_346_),
    .B(_358_),
    .Y(_420_));
 sky130_fd_sc_hd__nand3_1 _875_ (.A(_274_),
    .B(_276_),
    .C(_277_),
    .Y(_421_));
 sky130_fd_sc_hd__nand4_1 _876_ (.A(_278_),
    .B(_280_),
    .C(_281_),
    .D(_282_),
    .Y(_422_));
 sky130_fd_sc_hd__nand2_1 _877_ (.A(\valid_bits[5] ),
    .B(_283_),
    .Y(_423_));
 sky130_fd_sc_hd__nor3_1 _878_ (.A(_421_),
    .B(_422_),
    .C(_423_),
    .Y(_424_));
 sky130_fd_sc_hd__nand3_1 _879_ (.A(_298_),
    .B(_300_),
    .C(_301_),
    .Y(_425_));
 sky130_fd_sc_hd__nand4_1 _880_ (.A(_302_),
    .B(_304_),
    .C(_305_),
    .D(_306_),
    .Y(_426_));
 sky130_fd_sc_hd__nand2_1 _881_ (.A(\valid_bits[4] ),
    .B(_307_),
    .Y(_427_));
 sky130_fd_sc_hd__nor3_1 _882_ (.A(_425_),
    .B(_426_),
    .C(_427_),
    .Y(_428_));
 sky130_fd_sc_hd__nor4_1 _883_ (.A(_224_),
    .B(_248_),
    .C(_424_),
    .D(_428_),
    .Y(_429_));
 sky130_fd_sc_hd__o31a_1 _884_ (.A1(_322_),
    .A2(_334_),
    .A3(_420_),
    .B1(_429_),
    .X(_430_));
 sky130_fd_sc_hd__nor2_1 _885_ (.A(_273_),
    .B(_297_),
    .Y(_431_));
 sky130_fd_sc_hd__nand3_1 _886_ (.A(_249_),
    .B(_251_),
    .C(_252_),
    .Y(_432_));
 sky130_fd_sc_hd__nand4_1 _887_ (.A(_253_),
    .B(_255_),
    .C(_256_),
    .D(_257_),
    .Y(_433_));
 sky130_fd_sc_hd__nor2_1 _888_ (.A(_432_),
    .B(_433_),
    .Y(_434_));
 sky130_fd_sc_hd__nand3_1 _889_ (.A(_225_),
    .B(_227_),
    .C(_228_),
    .Y(_435_));
 sky130_fd_sc_hd__nand4_1 _890_ (.A(_229_),
    .B(_231_),
    .C(_232_),
    .D(_233_),
    .Y(_436_));
 sky130_fd_sc_hd__nand2_1 _891_ (.A(\valid_bits[11] ),
    .B(_234_),
    .Y(_437_));
 sky130_fd_sc_hd__nor3_1 _892_ (.A(_435_),
    .B(_436_),
    .C(_437_),
    .Y(_438_));
 sky130_fd_sc_hd__a31oi_1 _893_ (.A1(\valid_bits[10] ),
    .A2(_258_),
    .A3(_434_),
    .B1(_438_),
    .Y(_439_));
 sky130_fd_sc_hd__o31ai_1 _894_ (.A1(_224_),
    .A2(_248_),
    .A3(_431_),
    .B1(_439_),
    .Y(_440_));
 sky130_fd_sc_hd__nor2b_1 _895_ (.A(_200_),
    .B_N(_211_),
    .Y(_441_));
 sky130_fd_sc_hd__o21ai_0 _896_ (.A1(_430_),
    .A2(_440_),
    .B1(_441_),
    .Y(_442_));
 sky130_fd_sc_hd__nor2b_1 _897_ (.A(net2),
    .B_N(net16),
    .Y(_443_));
 sky130_fd_sc_hd__nor3_1 _898_ (.A(_168_),
    .B(_188_),
    .C(_443_),
    .Y(_444_));
 sky130_fd_sc_hd__nor2_1 _899_ (.A(_000_),
    .B(_443_),
    .Y(_445_));
 sky130_fd_sc_hd__a21oi_1 _900_ (.A1(_442_),
    .A2(_444_),
    .B1(_445_),
    .Y(_130_));
 sky130_fd_sc_hd__nand2b_1 _901_ (.A_N(_310_),
    .B(_261_),
    .Y(_446_));
 sky130_fd_sc_hd__nor2_1 _902_ (.A(net2),
    .B(net17),
    .Y(_447_));
 sky130_fd_sc_hd__a31oi_1 _903_ (.A1(net2),
    .A2(_212_),
    .A3(_446_),
    .B1(_447_),
    .Y(_131_));
 sky130_fd_sc_hd__nor2_1 _904_ (.A(net2),
    .B(net18),
    .Y(_448_));
 sky130_fd_sc_hd__a31oi_1 _905_ (.A1(net2),
    .A2(_212_),
    .A3(_261_),
    .B1(_448_),
    .Y(_132_));
 sky130_fd_sc_hd__nor3_2 _906_ (.A(_364_),
    .B(net3),
    .C(net4),
    .Y(_449_));
 sky130_fd_sc_hd__xor2_4 _907_ (.A(_363_),
    .B(_449_),
    .X(_450_));
 sky130_fd_sc_hd__nor2_2 _908_ (.A(net3),
    .B(_464_),
    .Y(_451_));
 sky130_fd_sc_hd__a31o_1 _909_ (.A1(_367_),
    .A2(_450_),
    .A3(_451_),
    .B1(\valid_bits[0] ),
    .X(_133_));
 sky130_fd_sc_hd__xnor2_1 _910_ (.A(_364_),
    .B(_362_),
    .Y(_452_));
 sky130_fd_sc_hd__nand2_1 _911_ (.A(_361_),
    .B(_452_),
    .Y(_453_));
 sky130_fd_sc_hd__nor2b_1 _912_ (.A(_453_),
    .B_N(_450_),
    .Y(_454_));
 sky130_fd_sc_hd__a21o_1 _913_ (.A1(_370_),
    .A2(_454_),
    .B1(\valid_bits[10] ),
    .X(_134_));
 sky130_fd_sc_hd__a21o_1 _914_ (.A1(_381_),
    .A2(_454_),
    .B1(\valid_bits[11] ),
    .X(_135_));
 sky130_fd_sc_hd__a21o_1 _915_ (.A1(_451_),
    .A2(_454_),
    .B1(\valid_bits[12] ),
    .X(_136_));
 sky130_fd_sc_hd__nand2b_1 _916_ (.A_N(_452_),
    .B(net13),
    .Y(_455_));
 sky130_fd_sc_hd__nor2b_1 _917_ (.A(_455_),
    .B_N(_450_),
    .Y(_456_));
 sky130_fd_sc_hd__a21o_1 _918_ (.A1(_384_),
    .A2(_456_),
    .B1(\valid_bits[13] ),
    .X(_137_));
 sky130_fd_sc_hd__a21o_1 _919_ (.A1(_370_),
    .A2(_456_),
    .B1(\valid_bits[14] ),
    .X(_138_));
 sky130_fd_sc_hd__a21o_1 _920_ (.A1(_381_),
    .A2(_456_),
    .B1(\valid_bits[15] ),
    .X(_139_));
 sky130_fd_sc_hd__nand3_1 _921_ (.A(_369_),
    .B(_384_),
    .C(_452_),
    .Y(_457_));
 sky130_fd_sc_hd__o21bai_1 _922_ (.A1(_450_),
    .A2(_457_),
    .B1_N(\valid_bits[1] ),
    .Y(_140_));
 sky130_fd_sc_hd__nor2_1 _923_ (.A(_450_),
    .B(_453_),
    .Y(_458_));
 sky130_fd_sc_hd__a21o_1 _924_ (.A1(_370_),
    .A2(_458_),
    .B1(\valid_bits[2] ),
    .X(_141_));
 sky130_fd_sc_hd__a21o_1 _925_ (.A1(_381_),
    .A2(_458_),
    .B1(\valid_bits[3] ),
    .X(_142_));
 sky130_fd_sc_hd__a21o_1 _926_ (.A1(_451_),
    .A2(_458_),
    .B1(\valid_bits[4] ),
    .X(_143_));
 sky130_fd_sc_hd__nor2_2 _927_ (.A(_450_),
    .B(_455_),
    .Y(_459_));
 sky130_fd_sc_hd__a21o_1 _928_ (.A1(_384_),
    .A2(_459_),
    .B1(\valid_bits[5] ),
    .X(_144_));
 sky130_fd_sc_hd__a21o_1 _929_ (.A1(_370_),
    .A2(_459_),
    .B1(\valid_bits[6] ),
    .X(_145_));
 sky130_fd_sc_hd__a21o_1 _930_ (.A1(_381_),
    .A2(_459_),
    .B1(\valid_bits[7] ),
    .X(_146_));
 sky130_fd_sc_hd__nand2_1 _931_ (.A(_362_),
    .B(_365_),
    .Y(_460_));
 sky130_fd_sc_hd__a31o_1 _932_ (.A1(_451_),
    .A2(_459_),
    .A3(_460_),
    .B1(\valid_bits[8] ),
    .X(_147_));
 sky130_fd_sc_hd__a41o_1 _933_ (.A1(_369_),
    .A2(_384_),
    .A3(_450_),
    .A4(_452_),
    .B1(\valid_bits[9] ),
    .X(_148_));
 sky130_fd_sc_hd__ha_1 _934_ (.A(_461_),
    .B(_462_),
    .COUT(_463_),
    .SUM(_464_));
 sky130_fd_sc_hd__ha_1 _935_ (.A(_461_),
    .B(net4),
    .COUT(_465_),
    .SUM(_466_));
 sky130_fd_sc_hd__ha_1 _936_ (.A(net3),
    .B(_462_),
    .COUT(_467_),
    .SUM(_468_));
 sky130_fd_sc_hd__ha_1 _937_ (.A(net3),
    .B(net4),
    .COUT(_469_),
    .SUM(_470_));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[0][0]$_DFFE_PN0P_  (.D(_001_),
    .Q(\cam_memory[0][0] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[0][1]$_DFFE_PN0P_  (.D(_002_),
    .Q(\cam_memory[0][1] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[0][2]$_DFFE_PN0P_  (.D(_003_),
    .Q(\cam_memory[0][2] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[0][3]$_DFFE_PN0P_  (.D(_004_),
    .Q(\cam_memory[0][3] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[0][4]$_DFFE_PN0P_  (.D(_005_),
    .Q(\cam_memory[0][4] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[0][5]$_DFFE_PN0P_  (.D(_006_),
    .Q(\cam_memory[0][5] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[0][6]$_DFFE_PN0P_  (.D(_007_),
    .Q(\cam_memory[0][6] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[0][7]$_DFFE_PN0P_  (.D(_008_),
    .Q(\cam_memory[0][7] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[10][0]$_DFFE_PN0P_  (.D(_009_),
    .Q(\cam_memory[10][0] ),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[10][1]$_DFFE_PN0P_  (.D(_010_),
    .Q(\cam_memory[10][1] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[10][2]$_DFFE_PN0P_  (.D(_011_),
    .Q(\cam_memory[10][2] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[10][3]$_DFFE_PN0P_  (.D(_012_),
    .Q(\cam_memory[10][3] ),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[10][4]$_DFFE_PN0P_  (.D(_013_),
    .Q(\cam_memory[10][4] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[10][5]$_DFFE_PN0P_  (.D(_014_),
    .Q(\cam_memory[10][5] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[10][6]$_DFFE_PN0P_  (.D(_015_),
    .Q(\cam_memory[10][6] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[10][7]$_DFFE_PN0P_  (.D(_016_),
    .Q(\cam_memory[10][7] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[11][0]$_DFFE_PN0P_  (.D(_017_),
    .Q(\cam_memory[11][0] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[11][1]$_DFFE_PN0P_  (.D(_018_),
    .Q(\cam_memory[11][1] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[11][2]$_DFFE_PN0P_  (.D(_019_),
    .Q(\cam_memory[11][2] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[11][3]$_DFFE_PN0P_  (.D(_020_),
    .Q(\cam_memory[11][3] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[11][4]$_DFFE_PN0P_  (.D(_021_),
    .Q(\cam_memory[11][4] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[11][5]$_DFFE_PN0P_  (.D(_022_),
    .Q(\cam_memory[11][5] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[11][6]$_DFFE_PN0P_  (.D(_023_),
    .Q(\cam_memory[11][6] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[11][7]$_DFFE_PN0P_  (.D(_024_),
    .Q(\cam_memory[11][7] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[12][0]$_DFFE_PN0P_  (.D(_025_),
    .Q(\cam_memory[12][0] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[12][1]$_DFFE_PN0P_  (.D(_026_),
    .Q(\cam_memory[12][1] ),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[12][2]$_DFFE_PN0P_  (.D(_027_),
    .Q(\cam_memory[12][2] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[12][3]$_DFFE_PN0P_  (.D(_028_),
    .Q(\cam_memory[12][3] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[12][4]$_DFFE_PN0P_  (.D(_029_),
    .Q(\cam_memory[12][4] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[12][5]$_DFFE_PN0P_  (.D(_030_),
    .Q(\cam_memory[12][5] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[12][6]$_DFFE_PN0P_  (.D(_031_),
    .Q(\cam_memory[12][6] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[12][7]$_DFFE_PN0P_  (.D(_032_),
    .Q(\cam_memory[12][7] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[13][0]$_DFFE_PN0P_  (.D(_033_),
    .Q(\cam_memory[13][0] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[13][1]$_DFFE_PN0P_  (.D(_034_),
    .Q(\cam_memory[13][1] ),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[13][2]$_DFFE_PN0P_  (.D(_035_),
    .Q(\cam_memory[13][2] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[13][3]$_DFFE_PN0P_  (.D(_036_),
    .Q(\cam_memory[13][3] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[13][4]$_DFFE_PN0P_  (.D(_037_),
    .Q(\cam_memory[13][4] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[13][5]$_DFFE_PN0P_  (.D(_038_),
    .Q(\cam_memory[13][5] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[13][6]$_DFFE_PN0P_  (.D(_039_),
    .Q(\cam_memory[13][6] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[13][7]$_DFFE_PN0P_  (.D(_040_),
    .Q(\cam_memory[13][7] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[14][0]$_DFFE_PN0P_  (.D(_041_),
    .Q(\cam_memory[14][0] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[14][1]$_DFFE_PN0P_  (.D(_042_),
    .Q(\cam_memory[14][1] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[14][2]$_DFFE_PN0P_  (.D(_043_),
    .Q(\cam_memory[14][2] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[14][3]$_DFFE_PN0P_  (.D(_044_),
    .Q(\cam_memory[14][3] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[14][4]$_DFFE_PN0P_  (.D(_045_),
    .Q(\cam_memory[14][4] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[14][5]$_DFFE_PN0P_  (.D(_046_),
    .Q(\cam_memory[14][5] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[14][6]$_DFFE_PN0P_  (.D(_047_),
    .Q(\cam_memory[14][6] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[14][7]$_DFFE_PN0P_  (.D(_048_),
    .Q(\cam_memory[14][7] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[15][0]$_DFFE_PN0P_  (.D(_049_),
    .Q(\cam_memory[15][0] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[15][1]$_DFFE_PN0P_  (.D(_050_),
    .Q(\cam_memory[15][1] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[15][2]$_DFFE_PN0P_  (.D(_051_),
    .Q(\cam_memory[15][2] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[15][3]$_DFFE_PN0P_  (.D(_052_),
    .Q(\cam_memory[15][3] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[15][4]$_DFFE_PN0P_  (.D(_053_),
    .Q(\cam_memory[15][4] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[15][5]$_DFFE_PN0P_  (.D(_054_),
    .Q(\cam_memory[15][5] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[15][6]$_DFFE_PN0P_  (.D(_055_),
    .Q(\cam_memory[15][6] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[15][7]$_DFFE_PN0P_  (.D(_056_),
    .Q(\cam_memory[15][7] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[1][0]$_DFFE_PN0P_  (.D(_057_),
    .Q(\cam_memory[1][0] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[1][1]$_DFFE_PN0P_  (.D(_058_),
    .Q(\cam_memory[1][1] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[1][2]$_DFFE_PN0P_  (.D(_059_),
    .Q(\cam_memory[1][2] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[1][3]$_DFFE_PN0P_  (.D(_060_),
    .Q(\cam_memory[1][3] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[1][4]$_DFFE_PN0P_  (.D(_061_),
    .Q(\cam_memory[1][4] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[1][5]$_DFFE_PN0P_  (.D(_062_),
    .Q(\cam_memory[1][5] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[1][6]$_DFFE_PN0P_  (.D(_063_),
    .Q(\cam_memory[1][6] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[1][7]$_DFFE_PN0P_  (.D(_064_),
    .Q(\cam_memory[1][7] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[2][0]$_DFFE_PN0P_  (.D(_065_),
    .Q(\cam_memory[2][0] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[2][1]$_DFFE_PN0P_  (.D(_066_),
    .Q(\cam_memory[2][1] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[2][2]$_DFFE_PN0P_  (.D(_067_),
    .Q(\cam_memory[2][2] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[2][3]$_DFFE_PN0P_  (.D(_068_),
    .Q(\cam_memory[2][3] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[2][4]$_DFFE_PN0P_  (.D(_069_),
    .Q(\cam_memory[2][4] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[2][5]$_DFFE_PN0P_  (.D(_070_),
    .Q(\cam_memory[2][5] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[2][6]$_DFFE_PN0P_  (.D(_071_),
    .Q(\cam_memory[2][6] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[2][7]$_DFFE_PN0P_  (.D(_072_),
    .Q(\cam_memory[2][7] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[3][0]$_DFFE_PN0P_  (.D(_073_),
    .Q(\cam_memory[3][0] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[3][1]$_DFFE_PN0P_  (.D(_074_),
    .Q(\cam_memory[3][1] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[3][2]$_DFFE_PN0P_  (.D(_075_),
    .Q(\cam_memory[3][2] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[3][3]$_DFFE_PN0P_  (.D(_076_),
    .Q(\cam_memory[3][3] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[3][4]$_DFFE_PN0P_  (.D(_077_),
    .Q(\cam_memory[3][4] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[3][5]$_DFFE_PN0P_  (.D(_078_),
    .Q(\cam_memory[3][5] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[3][6]$_DFFE_PN0P_  (.D(_079_),
    .Q(\cam_memory[3][6] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[3][7]$_DFFE_PN0P_  (.D(_080_),
    .Q(\cam_memory[3][7] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[4][0]$_DFFE_PN0P_  (.D(_081_),
    .Q(\cam_memory[4][0] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[4][1]$_DFFE_PN0P_  (.D(_082_),
    .Q(\cam_memory[4][1] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[4][2]$_DFFE_PN0P_  (.D(_083_),
    .Q(\cam_memory[4][2] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[4][3]$_DFFE_PN0P_  (.D(_084_),
    .Q(\cam_memory[4][3] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[4][4]$_DFFE_PN0P_  (.D(_085_),
    .Q(\cam_memory[4][4] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[4][5]$_DFFE_PN0P_  (.D(_086_),
    .Q(\cam_memory[4][5] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[4][6]$_DFFE_PN0P_  (.D(_087_),
    .Q(\cam_memory[4][6] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[4][7]$_DFFE_PN0P_  (.D(_088_),
    .Q(\cam_memory[4][7] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[5][0]$_DFFE_PN0P_  (.D(_089_),
    .Q(\cam_memory[5][0] ),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[5][1]$_DFFE_PN0P_  (.D(_090_),
    .Q(\cam_memory[5][1] ),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[5][2]$_DFFE_PN0P_  (.D(_091_),
    .Q(\cam_memory[5][2] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[5][3]$_DFFE_PN0P_  (.D(_092_),
    .Q(\cam_memory[5][3] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[5][4]$_DFFE_PN0P_  (.D(_093_),
    .Q(\cam_memory[5][4] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[5][5]$_DFFE_PN0P_  (.D(_094_),
    .Q(\cam_memory[5][5] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[5][6]$_DFFE_PN0P_  (.D(_095_),
    .Q(\cam_memory[5][6] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[5][7]$_DFFE_PN0P_  (.D(_096_),
    .Q(\cam_memory[5][7] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[6][0]$_DFFE_PN0P_  (.D(_097_),
    .Q(\cam_memory[6][0] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[6][1]$_DFFE_PN0P_  (.D(_098_),
    .Q(\cam_memory[6][1] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[6][2]$_DFFE_PN0P_  (.D(_099_),
    .Q(\cam_memory[6][2] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[6][3]$_DFFE_PN0P_  (.D(_100_),
    .Q(\cam_memory[6][3] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[6][4]$_DFFE_PN0P_  (.D(_101_),
    .Q(\cam_memory[6][4] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[6][5]$_DFFE_PN0P_  (.D(_102_),
    .Q(\cam_memory[6][5] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[6][6]$_DFFE_PN0P_  (.D(_103_),
    .Q(\cam_memory[6][6] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[6][7]$_DFFE_PN0P_  (.D(_104_),
    .Q(\cam_memory[6][7] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[7][0]$_DFFE_PN0P_  (.D(_105_),
    .Q(\cam_memory[7][0] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[7][1]$_DFFE_PN0P_  (.D(_106_),
    .Q(\cam_memory[7][1] ),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[7][2]$_DFFE_PN0P_  (.D(_107_),
    .Q(\cam_memory[7][2] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[7][3]$_DFFE_PN0P_  (.D(_108_),
    .Q(\cam_memory[7][3] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[7][4]$_DFFE_PN0P_  (.D(_109_),
    .Q(\cam_memory[7][4] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[7][5]$_DFFE_PN0P_  (.D(_110_),
    .Q(\cam_memory[7][5] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[7][6]$_DFFE_PN0P_  (.D(_111_),
    .Q(\cam_memory[7][6] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[7][7]$_DFFE_PN0P_  (.D(_112_),
    .Q(\cam_memory[7][7] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[8][0]$_DFFE_PN0P_  (.D(_113_),
    .Q(\cam_memory[8][0] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[8][1]$_DFFE_PN0P_  (.D(_114_),
    .Q(\cam_memory[8][1] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[8][2]$_DFFE_PN0P_  (.D(_115_),
    .Q(\cam_memory[8][2] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[8][3]$_DFFE_PN0P_  (.D(_116_),
    .Q(\cam_memory[8][3] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[8][4]$_DFFE_PN0P_  (.D(_117_),
    .Q(\cam_memory[8][4] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[8][5]$_DFFE_PN0P_  (.D(_118_),
    .Q(\cam_memory[8][5] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[8][6]$_DFFE_PN0P_  (.D(_119_),
    .Q(\cam_memory[8][6] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[8][7]$_DFFE_PN0P_  (.D(_120_),
    .Q(\cam_memory[8][7] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[9][0]$_DFFE_PN0P_  (.D(_121_),
    .Q(\cam_memory[9][0] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[9][1]$_DFFE_PN0P_  (.D(_122_),
    .Q(\cam_memory[9][1] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[9][2]$_DFFE_PN0P_  (.D(_123_),
    .Q(\cam_memory[9][2] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[9][3]$_DFFE_PN0P_  (.D(_124_),
    .Q(\cam_memory[9][3] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[9][4]$_DFFE_PN0P_  (.D(_125_),
    .Q(\cam_memory[9][4] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[9][5]$_DFFE_PN0P_  (.D(_126_),
    .Q(\cam_memory[9][5] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[9][6]$_DFFE_PN0P_  (.D(_127_),
    .Q(\cam_memory[9][6] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cam_memory[9][7]$_DFFE_PN0P_  (.D(_128_),
    .Q(\cam_memory[9][7] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \match$_DFF_PN0_  (.D(_000_),
    .Q(net14),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \match_addr[0]$_DFFE_PN0P_  (.D(_129_),
    .Q(net15),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \match_addr[1]$_DFFE_PN0P_  (.D(_130_),
    .Q(net16),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \match_addr[2]$_DFFE_PN0P_  (.D(_131_),
    .Q(net17),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \match_addr[3]$_DFFE_PN0P_  (.D(_132_),
    .Q(net18),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid$_DFF_PN0_  (.D(net2),
    .Q(net19),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid_bits[0]$_DFFE_PN0P_  (.D(_133_),
    .Q(\valid_bits[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid_bits[10]$_DFFE_PN0P_  (.D(_134_),
    .Q(\valid_bits[10] ),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid_bits[11]$_DFFE_PN0P_  (.D(_135_),
    .Q(\valid_bits[11] ),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid_bits[12]$_DFFE_PN0P_  (.D(_136_),
    .Q(\valid_bits[12] ),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid_bits[13]$_DFFE_PN0P_  (.D(_137_),
    .Q(\valid_bits[13] ),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid_bits[14]$_DFFE_PN0P_  (.D(_138_),
    .Q(\valid_bits[14] ),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid_bits[15]$_DFFE_PN0P_  (.D(_139_),
    .Q(\valid_bits[15] ),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid_bits[1]$_DFFE_PN0P_  (.D(_140_),
    .Q(\valid_bits[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid_bits[2]$_DFFE_PN0P_  (.D(_141_),
    .Q(\valid_bits[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid_bits[3]$_DFFE_PN0P_  (.D(_142_),
    .Q(\valid_bits[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid_bits[4]$_DFFE_PN0P_  (.D(_143_),
    .Q(\valid_bits[4] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid_bits[5]$_DFFE_PN0P_  (.D(_144_),
    .Q(\valid_bits[5] ),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid_bits[6]$_DFFE_PN0P_  (.D(_145_),
    .Q(\valid_bits[6] ),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid_bits[7]$_DFFE_PN0P_  (.D(_146_),
    .Q(\valid_bits[7] ),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid_bits[8]$_DFFE_PN0P_  (.D(_147_),
    .Q(\valid_bits[8] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid_bits[9]$_DFFE_PN0P_  (.D(_148_),
    .Q(\valid_bits[9] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__buf_16 hold1 (.A(net20),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_175 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(net21),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(write_addr[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(write_addr[1]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input4 (.A(write_data[0]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(write_data[1]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input6 (.A(write_data[2]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input7 (.A(write_data[3]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(write_data[4]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(write_data[5]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input10 (.A(write_data[6]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input11 (.A(write_data[7]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(write_enable),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 output13 (.A(net14),
    .X(match));
 sky130_fd_sc_hd__clkbuf_1 output14 (.A(net15),
    .X(match_addr[0]));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net16),
    .X(match_addr[1]));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net17),
    .X(match_addr[2]));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net18),
    .X(match_addr[3]));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net19),
    .X(valid));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload0 (.A(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload1 (.A(clknet_4_2_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload2 (.A(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload3 (.A(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload4 (.A(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload5 (.A(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload6 (.A(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload7 (.A(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload8 (.A(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload9 (.A(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload10 (.A(clknet_4_11_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload11 (.A(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload12 (.A(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload13 (.A(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload14 (.A(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net20));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(compare_enable),
    .X(net21));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_182 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_126 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_122 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_76 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_94 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_162 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_150 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_174 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_90 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_249 ();
endmodule
